��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\����q�?��e�I8�b�Ǽ$��"����ׯ1�V0���'�#����'����iX���R,4�	�W�bn���.�Ss�mY���dA]�����{mJ�4h86���q��tW��&�i�ܙ����0v����i�o�B`rR�}&��X�H&`͐]�������&�mzA�׉+Wş�ɮͳ�P6�Ȣ���'ď�4�%͂��J�%߽����
�1`b ��u����|��&7񟵒�������q�P4��'���Yt�(e���tJ�T�Z�>�~�=���̵|y�r����f��P��U�h~/� ���H8$
.QP�i������F�e
�#�?�6��Q6h:*�����х`PAl�[.�oؒ���_r�.4�'��s@��
���� ��;�<�J�m�{n��+�N"�F�J��ۯ��U�t�����C"�}��Sd�Q��I �}��s�\�x'Z��L��z]�4댱�`a��N��Zk9j�h�9�QƠC��u��7�;!b��ŉvX���ej1�`>Cm1o�^\��B�=0��]H���JH��0�/��v�����C��3Ã���.Y x���hvS�@b��1��0��4ΙV��3�=��e�D2�$����N�*�v�wi�1ީ\�Y�P� �ћ�0F��kOG3?�Lp,��8��#�U�*�~��X���,n�a~m���d���B4���H�zTq4ύؓ����:�����|Z	-���(6wE����
dI��Y�PС����$ҧ��+�HeT���_/�Ý8�
��M�^��)2��P���a{��p�3Hh�[�9t�\�C/O���vҙ��V6�jE��16K��E��".�oiUQGZj!�����Q1q��C�|>|K�"\b��e6^�߶+���s�TCգ��!r�a��.�w;�h�����%bF�E�P �j��8�Zԟ~�u��a���.c���@�r��CU��,��*	7��{9�+02��s'���x8�gRl�N���p��0c
�#��Gm���)↨
���JP�(�(�,4͍�خC�����2@P��A��br�q�ҒS�k�rʶ6m��WsR�`{���m�����yYp�U�Z��O��=�0Y�r!���u�Q���L���ڍ]�Q^�:LBh]����|I8����	tN�* ����k��Ƶ�P��d��[��ʎ��)f��ݯ�Wa��J�!�u���S�+f�P�YU��4���Q�~��OQC8�M՞��1��B��Gd3�_�
>B������M�d�Ay��D�Ӗ��@e�0bH=�d�xM,f�"=�.|���=O�kcX��Q�g$��P�T�Ts�M�rW8De�5+"��B9�I�iԈuh�x�h;�Ӏz-���.L�=^��m�G�-=�#^��\5�^�t .���Ww��~�Z������R���Z"�C�#y��r���P�� 
��v���q��%sp{W|Ƶ���/of���9�~��xL�kY=�	�U�� �sA�d����u`�Y	��W6���4r����O��C�o?ZM�z��p!���ګ���b/�k�X����ԲD�N�>�vt_m�I����"�g�s~HE�*H��@+������"HU�-ե_�K����c ��.a�!�z����F0W��u�dĘ�i8���Α�L�1�M��3z�=zW{����[�\mh4qt(����5��X[�手�c�}JNe�����:L`���?��hC
����h�#ߋ�ߜng׽;��ՙ��S��Q����|�%��D��:&��2q̟�~�S��IT��`�-�v����!���[�Xn�Ӹ�xк���X��	�B����!��*�᭚���&0ی����M?%+¡M��zt#��2r�"�vYC|��F��;���A�ה-��oo��@�J��4:_	��ťs-����p!WLj*,��E�M T�{���:�aU�����.liܫ�'sIJb#\P7W�uj���σ����΁n����`���Ү1]��-��2P�α���� ����L0�KW��
߬�ڿvհN�h�%����6�����B[z�b�ۍ�T}�q@q������o���(0�#��W�q�P{���Rf�(F�Ӡ��q�m��+_�Y�n�!L��}M��W��J��Ҕ=�,T��}�V��-,x���=;d�X� �qߎ�1ct׮�D)�����2Txl\&$,u�I�n��ҳ^�נ"��O����=�8cԯ�L���Vc�a�dt���\���Ka�5@L�`�җh�L�62�{����\N��e�&7J?Շٳl�8�Qa6-��%�Lˆ��q�6_�y���|�,8J���.�C}'! ,6��Z���b�q�^�;L>�W�t�	����{+{l�x�����F��~�U�A��Eԡ4�6BA�%w^�H����(�O�'r0惣���f�T�hA�{D�+����v*N��2�0�����%O~[��j%;�-c�q����A��r8R�r�����B���?>�@���k�j�~�g�x�=eGO�9�Rв�aXce�x0T�G����c8䴑�I�:��;	ŀ��*u��S�b�^��_#V� ��÷gՇ�w%�%�s�P���$6�@����m�O~���~Vz��s��֡�Mμ�ǝ^6r?o �}�:����A���?��r�K��}Jl�g���%`��QG7���A�'��O�ޟk\~���«��#nI"zv�o�N0��+���ը����qT�s��	�2��g��:�)�Azr���o{ӟ.�a@>�Vq���A�n�
�]��P"u.0���	v�˞�n0�+�ml�G���^Z��U�ɷ���ߧiD��7�uw�v�u�n09���༡���y���G��:���r	ϟ*Ƙ~w�� l��w#EG���Y���j�b���X*>�"%9���w䊄�y�<-u{�) ���Ǧ��u��֎sH����e.$�ãz#_g�	t4��R�M�Vo���py;ݨ�r��P<�b��er�
��»%��Ǿr�s��0d��|B�Yt!�QQ!G�}�-���7'�����5�J��!k��GI�c��M���xye��'�z���~�:v�#C�u�e�w��]�6w����1�w���O�dYyEg^��g�]@'����
�*GϹ+ښlE��	�`�1'���;�ܾ�R�!��pqQ�)���'�YY�د��K�iZ�-k��􏚩O*�0�[��Ѯ��M�g"���Us��./��Z/41�'�f�&��;��P����HON<G�k�_�穈4�_:hB3g��'=q'�햀�%��{U�L��yg}��h�P���:��uԯ�zb�>��X���$}c56��-�tg���"���� �������L�
�^�7qz�^z��k�R�xex����L���7ˣ�#N��?=p9IF���N��j���Y�C>$;,��`v�H�q[�1�`�x��@��_�X�4h9R�kD٢6�O�G��̤��gn�krC΍{NV�Ld�Jx�ܻa�]��dX��TBT��1h��O�C�v,wk�%���N_wݬԗ	�rt��"�Ǔ��6�����&�Ə�^q9���k����;����� ί�+�d���P$E�m�Y2Xs+���a{���{�2:D�͗�1�/y���ӝ+�V��GtWMtϸ�<��sV����=Cs�xl!ҝ�b����aT��<�h�*�z�Me�Cٽ��3Fg[�4Ճ�= ���L+��m\;���NO�Ñ6�J8������*�m�,ೄ���5�ey�5��J��-�0��̚�HI�|���k^+1�4(���=���!��&�e/��\e�l։�ݛ~��NI-C'�;z��0�TR�g��J�1�1;��r}���z;o�8�~f��?��V1�m�zzAęy1(�����%�H9�������CyA����TI�� �(b\�*?V�M/
�"M�6��lu��i^������DhU�%y���	�]�˰~�/ 2?$*���,���GnNwѯܠ{���Gи�s���`��":|Q�x�q�j��Y�3ˤEa滑-K�,�Ȍ5��[���j0���H\�ji �Ƶ�*����R�W��o�&(�j���N���r�o���-*����V?�~�ӿ�XII*�_,c���ċ~5=���1M\�f����0�Ο�B/��_�V�#V��mR)n	�
�n�y���������ь��
g��I|p���`�)��wPa@���ԑ��i�yO5pg��_C!��C8���;E�7�ѭ�,����J�譞gr��
�� 0鼨�"����5U��ɵ����Dt�%:����'a1������}�/��-���\�;�-�x]_@ͻ��)���D�F(���*X[��ZNN��R�5.̚��T�("=��49�<�L��k�T���}�m	z�]Z��^�����C��o�5J��k��#����&����=��O!�1J#u@!{���rVw׍����JΔ���IۮTEe �9��]5��a��Cid��,x�$�_0
���F'�������
���9���׺�c�ś%u��6O�k#�=�1�5�M���b���)�A/�(���k� ���[�ޗ�E_k��S���O0���d$�,O'Ix_�d\����K��+��p0���OX���y�/"
��K1�o#�#1��M[g��$���X���} ��\)z������&x�{n��F������섙����oDW�,3vAKV�S	���N[��E ���,��[ᛵ�*+�h�������Qۗ ���-��Id�=ˋH�XS��!��(��n�S-��3��(g��5h�A���\�2���O��Ѐ����!����R�p���i5V�����+���
w����K�����͜��*�D�.iҼ$|�/u�ۨ��M5���]@�~A�&��>%�n������\���d4_:fkT�y�}NY����_��e�x[��
��X�<ln_�;�W�r����s�R�P�΂G$z�F2�))�p��K�R섢��	��G,�g��E_�Ơ��k��aI���׈�r�̇���xB�+��tm�@;J����TU�k���!^g�5��&c�:w;��\��\$��=���WF�"k?/X�9%n,o�������jv�NSfz��_�0F�3§L�L�L���iv�������� >���㸖��]_)8�ՌYDX���\��6Sl=%�٬�`K�?��O�&��k�O:Y��w���v%(Y.�2�j}!� ly�T�ywUJ�*�x�t����F�������?Ra��p�ƲI<��A�/S�xE=�S�1$��$�X+W�a��I�ʍb��|'om�w������e�^o�����J�R�1��ț��� ��ڵF�I-�^T�0䣺h��B��w$W��`��L/��2Ey2�R2,$}������c;:��s{�nV�	[���g��-�`$���+�	�9B!�G}���y��Z��߈�W��n�I�Pu-%��\� ����=o'M �Jl��7ם!�����?n�"��D�a<��j�2�b�����;��ϑӫ�g��L�Qj[r���Ԅxrk�}����$�]:V*5�FC�t�Ϥ蟢M���7sv������2 �_�,��>ivU�MHM�x$�|���(UEtm(���x��Ӌ�v��(�j��Đ�j�h�<"��N�k΢H'���m��� ����^'ˢ��ճ&{x�)�y6)��N�P�$;� �8��K��[��O�����/$�"lG�� �g�S@�П/�v�j��ֳ6�B��F��{�0��lhQ4¼v��،R7�O��L9"��i��_M:�F��I�>`5N������s3K~Pɛ��6	��;;���F��OFȊa��P�4�H�p�܌�����3Ɉ:�È���r��ڷS�$*�y8���R~�z�S8�4cZLr,
�xi�s�2�����ڑ��OB=�x�`����~�S�������OٰV�]"8lt諭��SHֺ�?�e�X�̽!LW/;Z6��=�h��y�Y�n^h!ѴN�t�����emk���@\�6:
�[4�[e�+F��ፈ�
�tβ':�n�M1lM�X�i�s�{co��=���5PX�����2y����ef�3x�גӇ�f`B����y�������3f�-0o6�_CgkW;�B�J�nY�[���m�ʪ�N(�w	��F����s<�Q�������3�%>౧����q�y������21G����/E]b�b׍���I��{�y<��V�T����nxqMԚ�Dc}���W/X��tt�
��b���MHw��A�K�݄��>����<3S�h���0�X�_)��KI��c��|r�;2��H̄n #�=z�d�:�"|g��8����(�m!N[N�%���x*>51ڴ��I���4��\��.�_w5�K�|��̅m���E}���N�|��;#9�A�"�*��l��Z)�rF\�Z���0)�Xw��ϟ�i�7���{=�e���E�RPT�\.�Q��+���2Z��R���v,.}
4f0�2�l��Q�1[��+e&Do����O��m���<�HV㛬C�R����=�1��vN^�'����1=��+��B�"�ڰ�V�\8Cz&β������M��	Ey]��ɭI怍:�J�W�Al�w��CC]�ht-	V�ӪÂ�j�j�=0q"�W!�YLR/7a�$.���7P?����3�S�]�y��'���D���ᙻ��j��Ĭ�������!>uN�w���}���+�ƻ������� ���>J�F]��dO�����Ŭ�hfR{g��|ֿ���[��; �t,�OrTHȖJYd5�� Ҕ(nv}��{����PG�']F�X �m~LBD�z��[�D�#���|C7�#Oo����m9BY��D`:$�U�E�̺6¹4�_R݀�P���qNC�%
b��<E���b�:��DW����y��#z���7x~�����?�PV��9 ?����$��@���E2��D��ȸ����@���V|}f�M�G!�0�r������8krF�)*��q��tE���w~�Âxv�~ff��~X5�$�G�[�Ѳ�a0�B�k������zgiq��|G��Z�ӓ{��L!8⓲m��K^?���'���<�������������^�Ғ���m��F�����a�0zQv��L\*_�1���~f�t�p\�`��3S�"�]� ����O� �F��&s�#��H�k+	��6���B��S�0�!B?���Nf��+P�{�/���T-�1_�rls7[�k�-9���u�	�o�x{U�H�)i`V����F�|8&miȥ���&Gܗ.1B��=@B��A��+�a�(�H�BuO�+V������b�{b�:ܲ�^uȜ��ǹU�J���5���s���)�(~.tJ�R��%mU���穋&ކ�:<�]e�F^�`v��4�=s�.�0�UQ�ΤQ�A����T�Q<��+<��=�`ky:�Հ�Y��O�u�fa�A&,�D���$�A	����� ���Ɖ蘅PvV��?q$�rb���������'�NjA�LM���S�W|A�7�s=%{M�.}}���Ԧh!���e�u���zԣ��YB?-dؖ;��%Pv �A���ހ� *z̠[����3{�8�S(�#���e벬��:g����q��#�x�����Oz%�{47��B�`��$���:�&ە�K�1�~|)M��#��sÂ�Z�H��aV��fz�;1�E@%=�k�v�{-�;�4Of/��CZƫ%I�����r�#W�P��v����/K��jz����UT��,�B�r��{^yRg�=�ژ/%$q��*4�i�l�j�9�tmm�)�{R�ѰI:��DeY���h3ڻS�æ?��9�_ �?�o�G�BnJ�)�8�4��dTrIYX�.�M��`Kݨ��hB%�jcws��L���,˶v9~�g�d���> (��%w͑�BOy�����g}K�L���gm$�D�e���71�e� �ZR��5���ȼΚT!DW��%��*Ln%�O����kV��6�3I��ՃcQ���..�Y�����ñ���-������ךiv͗=}�ņS�w&�~����u�B���6�+�~@����.4�²���'0�#d��HG����A��(0���#��l%B�]���d�c���P��_U���k1��P.��dL��l�c�=j�Ad���e)k��Ek�N��Iޠ�S���m���9I1t�F���f�i,V�y��|S騫̶x@۫iA��d%j+��cRF��b�a�4���8�>��.S^��o��q�����?�f�Qn �ˤCC� ���r�㰺��>��?ޏBϚ ��2ޡ��KޒJ=��స�Bf�kN.b��ȩ���LWӸ=����6�]����Ҡ�Y�9����7[��WV]�B�4����u^��Ȇ&lS�z����8kA�e�6yڰNN<�S��g�[m�愗�pg�0Y��1��.��6�n�K�z���\QT�`��A�ϮVjC�	�.�L.跟�L�4��eC��Ǥ�T���I|
̓>���N�4�V�ק�9����7�1���V�n�6{�f��Aa���4�4@��mH�nQ?S��r�V�K�F�3}P�Ú�pF_.��3�AvD�m֥�}��o�i��#z�� �mb.���i�������Ӭ�HOK�V�O�+H�[�f��