��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\����q�?��e�I8�b�Ǽ$��"����ׯ1�V0�����v��"�F$�|��a2��|mP��� Εi��$�q$ � �?�kZ��
R�Q\��f���Z$��c5B�v�S� ���y�aV��խzg�_�*X5|G�}�	@f��l��&R����A,��)���X�rk�V�ˀ ��d78�6a��yǰ�[鐗�K�M���,+f<��skq}��S�Z. �yne����Pp�Gp��In�6%��.(i��WN�I���G��2f�|v�;�w�¾g��B�f?1<٧l��Z��I��uƭ����{����Zt���LM��0K��A�X��~֞7�f� �N��i6>:���In��R�Fʍs�F^���^�ve�qd����~7�eoD�n'�r �T�xRW��?]m�i$���
u ����g{� ]����mI+�D���]σ}��ZhM1B�������n���_����R�"�XDb��6$b�"�IwU��͇,�A�u���O	�c�l�<�%`p�"T��"Kb�A����%o����4��O�5��M[;!}��g�'��B\2g��r~�d%�5����3�s��Pz�lӤY�'2��Hjre�W+�d?vZ�?Cid�'qlm�A黍O%��2�v""VA�S=t^��w��S�t�4�yêb'�-��^�\�mǒ�0�+	�f�"��o��yG��^�.�"�j���i-8l���p��X`�|6� �.EK%�(t�rL�{�ٖ�A�: ܐ7�DuZ��T��k���b�/�v�-�"[���O�9�r�yz$> �nx��XM�Y��E�i)\)�v���B�Hc1c5�û�R��Y�A�;Pv�  /]�M��B�❁���g��Nk��A9������֌�v����p�>@|�:wh��c�5ר��4z��t�ׇ]���<	���_P\�y۲�{QMk�P'�U�c��	�҇H�,�3�K�����*W�A�%����R]DC0��`�w��=��[��F[��v�}�Ӧ��y�#�&{q�߫f���DxL�z��O���fA�)L����G��x��~�LYA��xㄨ��� ~0k��AJ�p��P�)2Q2D{2���|�Y@��H"g��!ʋ�o��L��		v3��?�������
Ǥj�/l.�!�ܭ����Y�.*��3\D��3ۃ��S�[���ڧ;��~;��X�{��|�!�����a-�����	^��,���_ɉ
>�u�Ea6��'�@»L��^�3�7[�y�`k��X�u���[x��24�lH��X�S� k ���.��]齪8)$g �Ӯ����4(�X/{�#��Q�����=�`Kc!�t q��~ɛ�Iɝ�#۱����r��#.J2�j���wj�h�<6_�<��v�*��8�>xO�CE�!�1E疪�վ�s17�-9���9o�����tR�#0��h}��뮀�+E�[���&� ���C��I�ey~\|K�K�c��D�c�|�.�ׇ�s�=�5����GE����Q�ݢ���0��H9P�e�_�]P��o_C�v�:X͆��j�s|�5���t2��t'��k��z*��Txb�д��f��y/�)ǽ�<f��V���}����1nI� jl-]td�O��wL�m��4r���.�D�����L6�(�ڀ�h�\#ܙ���ѹE�*Cx�w� n�s���$b>d�w��O�.M���0��b�:���\W����@�A��@W�	�Bu�e�SC�$f�{.n�(��3^���)�#kj��N{L���fG/�4G��f�4 \ѐ������?./�L.�>�4|��]�o�_`o�(>y'�~�����|Lг�a��*qL1�&��kk��ʔ��4���z�E�}ƾ��k�H�On{Jd���I�1���.	x�%��[8�J!��kԟҤ��\����&�N7+��n�}�f����d� +LAp�f�����rYZ�.�:�D&kH��sOs�P"b`���ζ���=���'�묱���q/��]k�7I��:aeEZ����5�"Gy���!�pޛ�%If�H��WD�~t��8���/&�!�V�~7�Rh��0��9��2��Vt�����
�;�|!��G��>�S��NHyTV��[LIC9��/8-a#Iw�?�Z�_�]��r�:����MH�O1��~���V�1�tj���ah��� �2/�XN�R�����1�����wg���H�/��|��-��}�#N@��<7ȋxF�D�36��ݨ���5��`wZJOo>�ZmO�JYz��rn��R��vt�s��������h�ëtz�C�m��Ŕ�.��ݬ���I�K�j�$��!�dQPR_�'���������i-�dl���sV�x�ֿ5��+�絯�#�*����W��V�5�~�z�)�I(U&-�;N����dh��e1)6��XB&d�``XX��/��)�zp}�}c{���2�ޗ��,�ù�y�}�gZ0����]��MQ�b,&�r����.D2�"a|�/e�������m��o��]g���볠{�r��/,�r���z����v2b[������q&$sL��!�a<� N�g���0����$�~�r���J������QK�}�D����h���Zy��	�a@���X+��u!|V���]��QT��)W�Q����|�p��:�����cj-8�e��g���8F��V/�z��LD�
!�R���^
�]�&mTS����P�u˴G�����X@p��5�c�n�K?̹�K����-�Y$4y�� �+��`��<�J�����hÊ�I�c>TV"�����![�
��}������(,,_�S�!g�W`�g�)��h��uSx'�w�ĸ=���0��W�z�U:ep�C�&�SHT�H��[�)"M��\+��W5�%y>���|eBj��g�>b�Q~;�E�j��y����ܯ�$��51`o0�oc��ˊn -�r�M��"�t�q��w-�v+��)����e����M;��ZM6��3��\@g�h�>qJ�gM\ܴsh�ZQ�j!	��ؿh���ɂs;����g
�z��T����k0 qs�ݶ(��j`��#8�sGS>��a�`VFg���N
t�˩�F��a'�n�S�7{� �i+�K�g>�A:���;
���� �D��z���<;չ4�!�62g�3>�}f!z�P���e�"�n)��[^�h���%�Q$�K6&eK<p�5�Ս#�U7iD�����b�
��5����%k���)"`�W��b\��4�w��t�{LX�7��s��P�D�VP�K��A*���P��(���������[i�_��Zە/���덵�"���M�r4���o�`�m���j��^�vE���Eyŝ�@s���ʈS�oF2��<�	*�|���w�$Y�g����&��mH�=����z�PJ��XN��p�!1Y[w������ C�SՉx��0C�w�]�l20��,��qWT��&,h��L��g���P���v%D^�2�O���qT��r'��n��/5�k	WX�p" ��J��.�sF��{K�;�hϑea���R[�c(�� �D���M� ��S�$4���^a#�z�"Zr�����N��H���o${IR�r�����w�A�VHY��#�%2�o�L�!.�RD~�Μ���S�pW��t���V���u`m����r������' 2����
|��<j���e�k��"���2�ٖ�֧U���/�pfmu۲��Z�Lx1�y�M�).[��Z��\t�����0<,s��)�EB�#s�y\ͤ?��+QHhW����9���as#x||�E"��*�	�I�=������;�_����٪�i?�̡Pn�!��֕P����O$M�Qu��@%���%Y�k�S�Y/��iz��&��٫ =�*1;Y2��K�������]��dw�����IIJ��816D��s4>�9��d;�\��������"�\j,.)��h���ӯ�b�Nabo{#�3v���=�)e8���(v	��}3'��Or����Mr=��Vl`n������thV;a����z�<���>�-���ن'n���~�m�ˎ 8�	"*���V��2�� b1�{4����9:�Y�i ���z�l���9��{�c�f!��x���D+�[���{��QWr%��Z4�P|��_�?Xg�uNC�A�~[B&G�u�}Rp��;���1���.��0��
0�l߾i��#JK�A"�"9���Ĉ������\�p����mR�NRf��ҧo��\�:��;��W�K��(l*��1]>��pl[u��L�x���� J}�zT�1���6���R�df��+���/��!@?RU��3ma��c�<I�P�?�Y����r�4��߇x��O-f=J��������Յ�S�2�N�3,�k��`��rH'&�`Q��*k2W>G�}�Ԙ1����'���֔���y��1�
�#�����5���M���Y��4I�"|<��	u���E3�2߮A�ˮ���ro��� ��=@K��q����}��D�8x�k��BA�^*�����!���J&�ٯ��A�]��b̝�h�̱@���
�y��rpx���"'9���P���c���̓���-��6����F&u^�r�jT� ����u���{��D�սF���0K�+�|��;�0)��253�-9�"|���G��O��\�i����%�,'P6��C`p��n��x��~}��n����B)o�ֽ��X�8B�8��ȋ{t�n��o>/1��Y�d�|���!&�P�j��{�V8Tz�~+=�/[����wa�T��FC/�۸��7����T�a���k鷱J�̲e�fՇ��gXf��FljQ�1�%�Jj�v.�X1.�|��y#�����t�X��r�����S�����7�o���������bpߓ�C,�v��`�f�a�7WjQ}�ZLz�Ҳ#ڥ]�#�M��^�$��A(�+�|����rE�Wk�.�����K3\�@'��Í8�{�mf~�<�9��������|��\�X�O�}��r� �tg�Z���0,Re1����k��aNN�~��	@�1�<\r�nIJ���DE��U��W����>����1��޹�n�Rb�z�W=̦+Uf`��z9����sJ�����U��E� ;!cG��p8����#�qx��P����{(#$j6�������/˵�]i�d����왗�M���W����O�,��j��ũ^�/�*)6!,��辏�C��,Ʊ*u���q�"��v;n�0�ш�M���0�۠��መ�HRFfƹ��Z��D*����Bɶ�,R�岅^P�q��34a�f|N�>\[hv��h���1w��0G�Y���\�Z�ވX�d�m,�j�4I����7�0Wɘ!T��1���]U?9L�^MSw	�;9����(�/�BT _ڵ,[����Fl?��:����[#��@���慏:4x����]K�п�E{%����Z�N>����ܶtO�2'��.z�Wb�cto�\R�:k4 ��	Er������D��܍�\~�5���5��g��ߔz���"H�v}~�ӱuL�6�
��Dv�<R�V\�qUGb�.���������T�è�.��Lp�<P=���Rgˑ�Zz늩��+����`�j����<^,��g ��$8���q?�GS&*$�RX4C�r����a�F�n�ѡ}T�7��aE�D����-�����Zԋ<��Hs��俛�)Y�����ug+~���ｋ�oA ��j��pT��;��4��(�@��g���}6��ANɲ�B�t8���O1���,Qo( ��N��G=��tԄ�_\��d��/�6�~5�t�+[��Yۙ]/�.�T���=��N�a�"�:ZkMJ�}�x�!X��F8-�j��L���f��cX�����:&:�yPe��opT�Ty�>"ܷx���{\+N��@�d�"2��_�p��<b^����^�G�>�ʴ<;\_N`����>z������A�@*rP!��Zg@��	�B��7p��s-�� 3aJ���/�O��3ω���1�箱OT�3��U�k�����z�7.��.'9��w��.f�W�͓ ����=�>�����!�]�}J-�E���u<`,��[���^%CW�Pӱ�3���'�҃�$���3�Qx+���L�a����Y�^�BFzϯ,��M5�� ����	1Y���{�� ������Ŏт	7��a�����<�hL����Z��~l���Hc�O�Y��<T��c�j�����5�7�NS� x_�Ϥ�k�B�тG����X���zD�}�JU��y��-i#�!��О��
�ٌ��!���(JT���B�P�e�;P�\B��:�A��d>�ma��̿�.m�! 0	��<s�x�l3z���4B�k��g�_��eԛ���S����|�l}��;l,�\�O�o,�«k��Vh����=�V#���|�v��!WY�(�jÁ�w�{Ym��1��w�~Oe}���tu�J�Vc^.?�'.J繡o�5�\����ǃ�� �|��"v�Y���j\�զ�Ѹ(~��<������\���3�뛻��y5A41���Pڟ	�Y�e�NK�B5U�p���nѨ�YR� ��8scӥ���Iv�,�EQ,���8Ѱ��p��ː�z,�xF5nͥ���R�o��-�|T&�6�8�B�k$��x?h�w��D���~����جS�oowoM��&b�M�x���~���U�r|X�Z�zU�僳����m����l�{�%7�3�2ߋ��ы�+-sykG��#'�{p0e�=���