��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@���$U[H_#�/8�y��,��F��`G�m6f�f�aiI`������tC����dl���=eZ��^�٭����B�FYĸX�G�����݁�]}~�s�cC�_ �c��2)����$�a<��d�6�q��tӏ�ˡ\s�$�L���Ÿ|^*��g�@U�*2�X���2��^�:9��D<��;�h��É}����a$;��몬g��>��W��iv���o�ăN�G\\�[�4�������W4xl��0�;O���V^��@��l5f+��\�&�7F�CqϮ�Y"�� C�T���/��Ƹg"���l ����~G�_y�kIe�+E�9�>Ǹ=�oWS�|���WV��P����������L��΋I2�G�r	y�i&�l��vЦ5�o�#����T�WrkV#��+�ڛ����C��ɀeG31>�����k�\�%�̶�@J�%A-�@�'2�}�0�΋ha���RN;zy�Q}N��5Z��}L���Z��¼�1<}M�����g�) $�8��Ρ�g���}E����G�@).�b���L��<�1�~:�~"�S��Y�p*-��^(Yj�����k��=98VK�ϲ�=�Zhy��� �#��_���c���~���YƯXrh"� Sao�%��Ƭ�;���cE��:�<:���6��E����Mr`2C���L�g.�T�"/)(dAX �B\\�xG�� ����	��r=�ى��x�⿐�z{�&��!�$�ȠC���}���?pEp�����p���р�e��Tu�M�@(���v6�ɥ.D�{(��Ķ)B0�h.ˢ�ا--��I�OtQ��I�ǧ�b:�ot����'�� �AvY��ɲ��c�Q��h�v�z�Fo�6$�ǧA��h�;�X��?F�4�E���j���X�Qd�i�� �C���¤T&=Ò�z#������z?��:�]q���� ���O��]*�h<�w2���9h}�{�/��Ԡ��vg��ӱ�Fι�\7���0�>�^�{�,�Xm�+�~��	��=}J
�J̜�zAH�e$z�b�����ֆ�`Pթ]��^�	]�~4�
��q�N���2�F���9,~�c8@?W�\��}���u3^D�l"����J�g��Ї�@G��ݻtq��Ҿ�	A�R�S��&)?f(��G��`��^X��_>=s+}ƹ՜ ��qgU�),��LЫ�&F�6�h?hy@��2�XL3-mV�O��p�w�s��>P{'��3N��x�Ŏ����er�i�k��&�%�����8�Wֻ�0��q4�no�{ۦRk"�32o(B�'f��	��r�s{)7���x]ۨ��s/[����IόM`�ԍ��X���F���(�����ti��S��B��q�B�ٟ�E �y���Ϫ�f3�¨qf�ލÉZla��}����*���ӛx��)����I)+�}��QM���*�jb��%qv����CR����.�?e�Y�E���F���}���5���U��}�)~����-�I�0�\w��i��\�6#�HB�^�`���y�/�/4��cZ|l���C�p)
��%BepZ[�Fطzup�
i��!>��M |Y��7�Y�;�V��M�� �rC��Cj���m�aϺeI_�����`&�l�$*ߊ�d���E�Y���U�8���b2FUjϟ�QG����n)�'���L�I��Ai�ȁ1���� �z˂�M*�b�>jtU�ҳ%�J���ia̍}ь4��`�\!��e�����rU�n��*�K_Fo=�N�m���35���=
a�6K�G�Hi9C7�+ �x{<�}B��72��o�Zo�q7n,�M��L��fA�������@G�a�����lP[f����R�V������P?v'6}PeɥN٣�F��;V�%$\s40�4���R����/+��,<^���`�Ѐ�� ;�ʹ-�\~J�e����w�q�t������M����F����4e])w<0���#�����'�t�+ ��$��L����z��m��l5�6F����4JvƠ��*�)H
��m:��j�J��St�~��6=v�>��f�پvyt��:D�Б��]�dP/$��k;���z*�"t{�G��ۧڶ�r�/a�k�P�X�7���Ս�?���M�m�����\ ��7Ad�qq7�N(��5w�v=ݴ�u#�0�%h�2���}��2޲O�ܻ�q�PV'��J�[ڑR��Ũ�":�O�6�	���m��1S�$���j�nLca�c<�����x]�e�ܝ\��ge��r/@�w�t��l�H�r�~��:�7(�Ϯ��p������ L��7!�.�L2B ��@��ڐ��6��,������i�m��w+���P��D?x��Ř������>��E�`&���p!���볝�S�vu[�f�j���80m4�èL�Ԕ���YMZO�h�`G::�dL]:4i�g�2�����*K��e%3��봩8���WԎ���kF���_QM(��9�\��\jP��=-�oI��F�W�<��t�,��-3?1q|4�`y�6|@(��ӹ�=o�A�-���Z�,.�*Q������
E��L�R'�dJ<M���O�s�X�X�"3����'c��ZXTU���7(�ݐ�ͦ1��YǪ#s���|ޜ���O����/-l�.��^�\���1x:����z�x҉?�R�ysqܬ���F��j��[�[��޽��P���Gk�s�����$��Auuz�X�,+<�,BȂ� ~�y��ҁ�x�w�D�l�݌)��X��\�!khg)�wדX��0��7ü�8���T|�����iR��N��M��/��hb�G���s�4>��Fz�����ңluOc?8�l��q��W�c�"���$�;�������wd��j���y<�y��<N�������A�,=[˧�����n��8�f�̸��ʂ����l�}O�ʖU�O��rFM��g�ZĘXkG02�c*�td�;�6����+�F\�(F,z	�_��|��#�ȹu�;�����������7�w@��Q�F���p�(��W�p
J��`��hA�7Kn�E��^̼���\��-t]�d�j*��4���{��%#�39QK�q�m=�@�N8����S�֥�9iZ��]7Zt�Sy����s��a�(��tgKW��W���u}O�r���t([����I��N B]�T��c� T4議$
��Zk3�k�N���h��ו�,�G�m+:��;��i��E�1!dރ���]�7�s,Q�${OV�6j��z�&��A�/��	��B�[�[�c]����5)�na��v�'?��h�$��(X@zLߔD�@�VO���6�[�W����O�4m���#t���kB�����O�������6Z�����H?'��lo��jב�IU���@�e?"�(�Ј�]T�d�?���x��6t#P�o.�p3��%0:�H\�^�UO���*�{���7"=:���1�>1�rRb�>dz��cj�iRϮ��ͧpƧZ҉�(g�Oʕc=�^"T��o+RH2A;vǒ|�Ռ����\�)�qp����'Z�(�~�&�9�_S�&�4&�*M 5:E�`�,���F�s�,1�+6!�bv\:�B��xd�<��׾`1��L���D附?������bO����q�JXF:.�h�3Qik;)Oa��b=$u0@��)Nd������1�[Cczq�g�p��D�~#D�(���r���w�S���6�x���c[�]���]�����ԔzrE��D�O6��7�{�����·��e�j���O��edѳ��:��Q����p��·wo�>�U�Z��z��:��#��	\b�7Kè�"�
X�t��9W$���+A�@��ٚ�8�ǭ�]ML+j�}�1OK�^�sPRv�v�\�e�5�=��Ôޯ�"�z?7/}H۠v�|Z2��X)rj����G)C/�`������1�YՉ`( ��Jr�Vb�WB"!ɕ2[���󾃵�}*1��,q��(�7zJ_
q���#��L�G����@T`2�C��^p5����^�G�+� �m���#Z5��zfd�T_7D���F�4���?�т^�틈�cu����s;J8d��}�a��b�5w����k�Cݴ�	�����n_����~��~�^�����,IT ͽY��n���]����l5_W�fbG��XH>�&r%?}N�
)�)�޴����T�O�Ca����ǭz�K¶�����T����cxii^F�:�l�Ab<"s(z���:$�K�na;�6�(	pS)��Y�D�໸O�?e��67�+_��Ӵ�mmdnȧ�c-�iw���h�M���&�}�oN����[����Ghb=����ɋ���ob!��\��؏���Kfi������;0��*Ét��as��!K��6K7<d{v�l�c�<� /b����=Iu
�֎��J�F�_����1���ۛ�3n��9��B�����YF?E0���D�M�D8j���6�bi��+	�v�����	8�[KR�7�F_�&m�i�ws��U~�������\ɖ��1U*v��0�N��֑������=����SQGj���Ĕ��Ǣv��&=R�;jӽ�YT=��١R�	"�&���k�S(u��7$���J�F��A�9� �h���}9(��+�>?ש��� Ӡ�i-m֪������ļ����q��qx�O���k.`���;&:�Ip����q۩A��hs�LH�j����&gU��ɰ֊^� z:z|�u-���k��^��z��V+GeF�ڬ[�)�����Ù1��� �8�T�p��)�P����|����F�/�l}2?�V*ƪ$�%��rSQRi�#�+�5�Xk�� �?2����$]RA���&��l��%B�w�E�+�|�T��K���`��2E�Bs
����A��Ԓ�v͊n�2��,�s���	x�����̣��t�9�u5_�K�`�[讆�\H�6��y��{�q�[���i�$낣Vo�Ae� ��#���YP��bK�V7-A2bk3 �!�EV%L��獱�䇪����9���i�#�D2A
�wǗ�kJ<����8Ԇ�</@B��8R9I��p��V=3]qߥ:�#�����
�,��^�I��������L��z���~��JӁi��J	�X��B�L��C2�k������t��D�?�6�Y'䋉mP��~�1�,WGA<��!������%��Ug�1@���VB�1@�  �������yQ�|�B.]cL�83���v���<�	Kk{w������j���屸p
�I��@�7�~�U���I�q��W�;4��|CX�����^WmR4�1;nZ�h�S����/�ǰ�[�j,���)��(�2^���� Cv���x��n���Y*眮����JrW��l(�J�ܓ�m沿ǛK�� 	�)h�*>l,��oj��T���)�I�9���=���*|��ͭ�H�-��(�oh�kL��}��M�k�*����3FJ�p0�?G#co&1�9dV�o=�W}ˀ��>qK`|xX�7�@c����^,T�b��KJiYمH/)�9�)�V0pA��J���F��.^��}�f=�L��`k�6Y�����F�`@/,���Nz��i��h���#D��N��b�w˥�HU�8���W�.oj򉉁�Q�o���������M�q�m�\p���]߿��k���;/9��-�