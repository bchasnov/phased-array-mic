��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|��I�ɖ�<���/������
����V|Z�y�l��%�0B���1���|"|{��s��i�˫�Ol$�&��P��]P�����\����~�
-Qh�Z�}��7hs��1��s��1C��� r�0')���}QPT�wSG�){���ǕG�Cj�T~7���y�4��ZSVd��n<��4��d��/��~�������Z5�C��A�?ff/ �K��|�g�܃����hw��l��rѵ���"��@��G�/+(�ڦ��wQ���i���D&�&Y��2U�o���H�D�,�!q6���TD.�f��V�����<5*���1Δ�ੴ�]^b�/�̈�O%��xގ��Xi�+�M,��Ğ��1���;�4���jb���K)i��.�]D��L1w��1ɿ�B��P��dB:C�^�����sI��&W|�wR_}��v�����*�b��|& �[���&=5XD�����5M'k��&�U�����+$�b��: �j*�C��*Z�x�~�{�� �eEF)�۬���s�R_gmS��T�pԖc�0��fK����R��6)��L��*�zoZڟo36�Q�ҝ�~x��*N���R{���(��BM)��_.���%�E)6���C�`A��nyW.y���8c���s���t�O�s�Y��!�:��X�>���2�\+�C�8�͎H��U���r�.
�����tf���p̖HH��Jm�`��$ �����i��2�H��L1���r�<�.�3Q����'��Z�/ف�V(x�5B2��|�_��Of��-���N�s��"�m��(2;q=�*$M8�����(<��y3{���.N�Н8o^Sذ�iB\�_#D�̠�_1?��A�|܋0޺6�`��.���LL0=Wx�.��#	]�&wP���w�<J�p�?;ن%�'J<ג=�wD�GH ޞ�r��q!��-�6-�2�[��V)ӯ�����:8��o�Uz�ҒJ7[��H������L*`ӛ�X2�02�ǈ�xR�d��**�i�w�q��y_���K@�\؆c��/����x^��c�,��dʃ��sv,�୩���JIx#�>�g�k�㈅w����2�X9ji��Rqǁ��M�5g/.�EYd:r�^�^!b2���f�}I��b1R�,��Dp��0&�D�ǆPP
���L����y���͚w�4�F��6�%T�.EF��d�K3e�:/I��a*^�ݧ�;���,����΀���>��~��s����.-Y˜�i�[�V�4~�',ln�S�$���>8���u쌐�͚S�0&��V�Έ:-�B��qL�+�c�JA���/i�>�8"ۦS
�B?�8���T"u)#�c_�sچg��{�e��UI�N�S��=�~�r��������6�rBܣܿ��B��IW�c Mޞ��Y�$%gO��.6�QcP��M-�"qZ��l���s�/�!X�g��U�V�\��@S��d��܀"����U����J�к1K��6*�֦�˩Zo��w�j���b�޷���Ã�cF�E*���P`��.���"���v����_�`��1"��V�e���ͬ�g�Hϑ(���\g���qm}�8�����}��,����^vYNYb#��Wa0u[&r��w��|�mЎo��onE��g5Dm��ܗ��ߠ-rWE��c��-��_GϮg���4�jF���~���rK ��\(M>y�%z'���XQ��-4���h,(�+jF�ީ�|�5V��i0�u�,�q�wW����,쮅,��H����2���	�I����ah�j�B:��.R{�=,�Ggoߔ��  �^%`�]a$]����ߩ��4H���S��I��!���������a���9:l��4N��PB�O����t�O%��X3�>�i/1qA7Y����l�� n����p�����$��9�����j�a^~%�����J� Mkw�rb2�t�^O,��������cÝ���[:�kZ��u����vn�FD_�Q�lc�~�������K�r���Kd��EΚ�L@Di�y3x���z?7��I��ԗ�
�΍���'�J�e=W'�e�����B�s�h�O#/��*�O�J��LP\�_���p��4I�j���+%��Ŏ�����^��9���`�G�S��K��W��8p^��܈����ms�M}H��w;pn΀�����-�{ :�lR��qQ|��Qx�RT|���R�"��ι���m�$/���������wQ�z]�e�)��jM������#\��gvJ=���n�������6���'� ?
�Q���	�i�톐1�#5W2��S��趌��D��U��������
���+=��ߝ���[�6�v�db�h������w��I��*o���-�*G'kSkب��Rc���; ��#^P	3����}�Ǳ�'��G�2:��f�����4�y�}q��ۏ������>=�
��W=|����"80^d�ݏ¢���W[���C��)�)�|0�ew��Z��L�Ӳ�,��5W5L�hv(G;�O�`��M�A�q��7�^�&�ѹ2:�O~��b�5�%����E�#���e���n(�x,"�3���r*�Y�>�u���(˝v[��؜5I&��u2�΍d�SM4.b^�:���'\VnK[���,�Q���[b�n�eFp����m�W�E��(���!LJ,�X��1▩�_`��|�:�@�dVr� ��(b@��͊�1����=M��vMD��v�*>˷��X��=w���T�t%сM���|N��$X������ж�H.�9��6(��Zj%�;�ɈFd�=ܺ���V/�ө�ISᎱB�ʾ*j���gw�<���7����h�^V០�xB�!cyu��gi��`�x�|o/�^�V0�o�7�X�c�����2��NnY�qf��]�3��}�zۨB�5�����=by���e �t,��@|
�0���6�C��#�ǧ�&n�i����J���!�Y跎nD<Ӷy�g%7�=6���P��ͽ��x��Z(�9x�a�ֆ*r>�<K�5=?K�6λH�
dei�>#S`�Z�`�hyƷ̈ ^�y�0�6=JNY�D�A��k�����0oe́,aQ$�z�)R0O�����q�{ٌ�hhWPf��2S#\VH�載��c,�8��O�ߣZ�l�����M,¾�\7��4Lμ���`�\q�����>9��_(@p����|�pb���б��I@����b/��.�C�"�B��?���Kr���PJ�������f�w�ش����U�rL7���6�Vʋk������kH����#���˯�B��dz��g�$��� �51%��y�dv[�@]ֿ��p[B���7��������j8��U	�) g����
D���E)k��� �4���B�ZZ�*O0�W=��ղ������g����N�pJX�vw�d��;$����kn���ᩁ�]� >�t�Ŗw���O���K�0�.W���(���=O�Z�fr��?���|�1H�U(�P3�E6V�A��T�;M^�R"ݱÕ)e�L�7çï���ӆ���7)Oz鐟�X_�ӹ�T�����C�d��bN���?�����;ɞP!�AR ��i��+�PW4�ZP�8��?��x�1�m����&+��o.�E�T&g�T\�����w��f��������-yڬ�fK8&��}Qs�58R�;�����7S9�~!�@�VǵI���