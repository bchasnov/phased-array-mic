��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1���e}ʲ��cg�t�ϙ�a�:�KR�%���ݧw���ȼ���E��� �(�����q�֭}s�j�O�%)�Q�����^$���[bqbٍ���f�?� ����v�Ϡ�Adز*���{J!�pC�lL-��N��2�)�	�o�A����WǍd�L ��C�,<<%���I�QB�M-"k
���H��M�6��.�s=
���@1V1�x�e�X�Ӂ��&��}�7m��$�*O���2�"��(Ojd�C7�8��L��r_X��ƛ����3_	A�(���'���ԧ��V.�$��)3�;�>�Vx�g�Ӂ�-E�}�)c�4����s��j���GWZ�����C�
���g=�_����!�PF�@n�	+�E��a�fJ�G���8"p]��ES�怙��`p*W�X��3-�7͹A�JѸ")[�T��w������<~>�;DC�bu�\ C�n@w��L#����[o��儶�@!����
{-~y�K7�a�P�÷.�᣻{b����l�^
!�"$�<K�h�'�ٴ�V������vI_1:;:
Z`iC����*��$Y �����5>����a�Uz37�'�P��Mj���HB�$VhF��N����W	��Aj������a{�-������x0 PEsr��"j��&L��Q��KN��?�����4��g�躙����Vo����)8%�I��:����_`r�QY4��N��V;��y ��M�V���ظɌ�T�:MY-vQ�P�7��y�%q1:x���cW�l��";�oo���DE�H��Rl;Dl���~���\��~G���-��
���d�A� �mV�STD�\�1�m��l�{���&�M����c�I��Qj� ��7=oL�JT��%� ��pU��;�[��΋m��F���LR���؛N#V��3�C�c#4|hF�{�[׉��@�m�^���OVP��I�g}�y�b����'�m��a�)Od�C�/�b1>��V��$���m�R���j��d�����o�t�~gY_����xj;(t�����߀�$а�|����F��tP�j��b;�ۗM_-B4�qO��4�������eO���J�Mj�Fi�g�������XA��۠B�)RtTg ~=.!�A�r�Ƃbs�SV%�Ր2�;
�I����7.��( N�x�)�6���.��T=8b���V1��#����h��յ�:��9��*m�FB�:�������d.Ja�f/��m����{n�,�&��koj�VEj~cއ�P�,�K(�J��2�:�D1�*�G�F�P��eȟ��E9rD�/h]d�g�uv�v�9)&?��֭7�r{Ps[}%*��~SB��l_30���~�iX��Z'_c�:=�]2�.�:��[���c}��Td��^���H�D����\ƫa��V��Z� �����c��ρǄi���߅��W�n7ȷ!���O[u%���`:O�_�ϥn�����"�ޒ��*��Ҙ�D\�#[&)����i��8���#ޕ{��8�^�"c�U�!�E��E����.\�
�]���W7�+0��xsQu3��ӱ*=�W1��'��ta0>ϐ'n9ct.���9bl(t����ѥ
��fH┻�Nw�����Ei<�0�̚8�Jpb9� \��NT)�`Er�~S�v�5���R����@f�c����F.�9"%���Gڥ�ߍ�h��lY�D^-'��?���op3I>W�d)I�Y�{#r�N3����݁�t�|icn�6KEȦ���r���E�9~���X)�ɻ��<c޵jW���~��P����(�$��P��+%�C�{ؖ�!�"�&�6L?L`�*%�WqU�Wn�[�#w(��&�D�̝N��� ��^I�H�>,�����ƪl�Iu�߰�%��H���㏢]q��$����'n�e�Q/�ÿu��C Jʅ�v��
7��,p�MPKp��y��J�h-.Ѯb��L���a��eb�����,<�
���� �?�����.�<��
����V�����ӕ��=i�s0���1�C[1�*���"o�*d䪥�� Y�rwuƻ}RA�n��hv�ch8P���a���P�3���=�V�<��K�;�Y�����ly�;AV���y�T�����Ĭ�{Ίm�P�b�(�+�s�X6��QQqِ���u^9�~ F�@;�ws9�:u�L>���n\�,��0$\�(��6~�K�	����ȪG)B_#�����Ѕ{UTM+�k�rꕦ�Ճ�T^L<|I���իS�� ��y���0�Q=lC*Լ�M܁HblM���+l;�͙��<��>y��*~�4���BRL6ߖ�H}4�)��b���ڢ�8g<}+;�L_�X�dE��6���%���y���h��w2�����:7��'Q�6(�wd��>F7n&���t�'����ق�s�?�q	.,I��?:��G:XR/		(�ˁ�Ƃ���P�u+�C�sq1$[sq򖋴����	Gi"J"; �`���PE��eo�h+��g$�U�E?{6�{Dp{eMؕK�>��'��Eȗ�<tʢ>X�å�Gv��:%�'Ȏ{U	�/�;+PF�C����o~_�i>�M�^����7D����
����v�Oj��"�q���	E�J��K��Yl�֖���7r�Z�/�ܫ1s?M�U�YV9��=�,D��B��=��j��˓(I�����\�3S]���
Õ�2�#��y�j�.�5��d�4l�
O�^�3+�,E=��7��W���*.�f}�ԕ�v�W��D"�'�����q���I����.�L4��Y|����?:a��k<Rϫ������M_�c�e=b	�����ta< `7AX�F�3�\³ׯ�wn��V}KR|�����T��������P�ӡiy�XJkx��c�'���W$����]���w#���a��М���i��"�T�h5��:���E�����X��ӻO��!���-�b�8PN�%�Ƨ��Q�4z�gٜ�P�{�ES�'�~���`�s6K9�n��b�B�E�4��a1�bs���<5΋6
w:�U+��r��?K�Ω�p6��0���25��![9�*�3V��E`�H�G��:q];'���N��Zo?��K?z����`���q���!ԁ��Z/�s��4���� ��%b�h��R�	)��R:�����<}i�����s.����T�f���~�W:��b�3H<�m�	�y���pc�czW62�
�����+����c���.�	�(��r^���$�d<1�V�q?��Y�M�¬��'�""���?�sS���<=yT6������p���U:�%��՚�G\:;��8'e�/��7<��d��nWsX�c׌��֛�l�e�����G�IR��~V@(�hW&�?]V|�'*!�)�x�ǀ�Y�<�Z�6ň�;O���U��� c�-}������(I�?bLiר�����`]�HM�����)*�h̾Ø!�Z���)	!��98���^��(���+ѽ��@��r-2]'�D�գ��� |���_4d�uPg����_p��6�O�(��/
h��hTH�N�bTm��Е�hK�-��^+��۞�c�>[�; ���_^�@���;�Q� ,�el�X{Z���Y��/6�4��C������re��.��LE����Z��#P���+���WX�>��{��Ǒ�s�*҇�]QHM�G��~դ}�Ux��!��2Ðי�G��6N�y�O��R�#~�Y4:��?�yE?�C;m��;%����BHHj2��uJ��!f�#\�ڋ%<t1�񅸩zc��� y��r�{���j���������=�Px��k¾�3�\O�3���P�q��I��ꆽAC�Jw5�`�0lݷ͏�����R�����za.�G�&�ʑ�
��ŗT^����~���H|ύ$	���"b�];�>�K�G��o�Qr��W�b�.�JL�`xp@v�cTV�X�!�V��V�4���Q��_����A;�OY�q�Y͡��Tv�C������*��Y÷����آQʥ��[{������a�Զ�)�����(�y��������˼�^Tq��G�o��	�z��q�vrK�	�\=�c&��_yf^�:RTW�x��r_g��k�^�L:֢qi(����q����DuGXO�z���X�b �=��=-�'�=[�.��$�򴙗��E���t��eg��$�#�,A��\//%�b��%��x�1b�Mf���Y����{qK-m����Oָ)��G#�0$�I�_�f~:�H��d^4�k�@i��+��$oޣ���4��r��ql#��]�&��\2s.ôMȢ��9��K+n��>5m�ӯ�J����_��p�U�V������g����_ۃU�<@DD|�O�(��N�	8�����w^2�p�0�?1l�#���H\��ń�\u�a	TO�M�.�|}{�(��Jy8-��C�Y��AK����vX�7�Z���$�4�p�����Тg�u����܈���	R���lǝ�|~�@b�o�8���g��4���#��	�Z�q����
�I�^� ?a��ñ�H|�b�`�I����߀_X�^C�Y�b���F?�� 빗Єl�PO1�#�������R8NY�\���Р��f'1�Y��͈��l��zL1?�����U�����2��0�7��J��zA0h����o=��n��i�a[79K�sP��̀ji�C��j�)wQ����H^���߽��q�T���r\
d��Z�6�	�=�1�{ۿ.�|�Y��\�HP� O��̀����U_)M���c&W�H�[��WXV}�~r��>ߵ�����y�Wz� �S�W����s=! `\=G9|F}�D�Z���'�@p��6�YY\vg���@>��]�y�{�V�tQ�x%� F�e��>���V'���P �=,���׃����w�L�˫���4)��W�ߺ�����}�˦6� �Ø��Y��zd_�g|�=mɧ332�[�,�q<w���G�O���Ơxބ�V�Rep��%�\e�
u�E���l����DNV�j6h�*��+�<�$D�	:|�}u�a �^�����pC��bH�P�<���Y�����؞R�z��N���>�!���V��1�褟�@yN�i�z���_�-d���Xٷ��̥"�n����)����'3*�Ś�DY!���f��My����B,<���d.ɠߤދ�@�A+����s}rGy,.�.��z���m_�<�VQ��E�Ғ�KBe"�۸���I�l��c�����֪�^x}%�|S��R��b���ZJC��ZR5)��v�����n	g�p��҃	Wu:��[�A�)��
�,���t8(�� +#��4Ks��QEK���["��[*����(��td���mR0����A����B�>���"�v�Ց�� {�9�V�����c��#�栄�	֣�m�������ngίmtIKlq��тz�xO�o���a`� .&IcZ
�e:�u%�`��}dR�6�����y�m�û,s���{����=]���  ��fƽ>F�/�2NQ���#�u�9:�^B4�������i��`���7��hcL&��'`�)�"x­���П�Wmnuy��ҽ��]�kNkhKDpy�^!�!�,x����\�TF��m�Y�uG�j��8V8�A�L���j�M�Js�
��@"c���}�kh�O�W��)�u[t����W_|��-��+��2R�-3YX� �2#P�8p	��	}puq�C�jg��<߉3���Ԟ�5�ې_bTG=� ���P�G�@��7���GB@�w�
�)���[�/2��<��(i{�\r�758���dN�����gtݶ9��g�]�P6�#� dо[��?(rri�!���*�즮6�:�<�]
���tp��z�uy4OӅ��Ɛ���ez�C)�d��6����
*J���y���ȣ41^����o��C:�#<�.*�Ι��vQ/����X��h�[w���:�>`��[�� �˰�img� ����R*�oE���~�<�A͂���0"�p��g^/���?m�����s�'�t��5L�"���i�=e_��ri�S�M��E��e�9����9��Z��
�O%p(s��l-���b�fS����u�+
��7MZ	 ��}�M�;`�+/��n��R��0����_U���QYRT��u����\�<��ܽ�ug��h�zP�w�f��o�F[i4E�%ktc%���A �����ˉ|%�6�qAy����;oh�W�cG/��������Ѭ��
5�������?�W��^by�^R���Y�b�(i��>7W{x��="Bw3�<�-�T6*l��vnG�~6��}Hȿd/I;��?O��ύi��N��/�懀A�A@a��+0���c�R\�3�������
v��$��0�궨H�e�#)�Ь��JlC�{�W�<֟H+x���w�R�������ѿ��{a��r���9�#��zMGo�-�Rs1��;iWA.V�Ӌ�tJ�6 �7�+8^pS���e�k�qWZ���Kb4�x��4��}� �Rm`��(��[��N�^��𝄙��|��	>~�� 
�]	�)TZ��4���}����Q�L'Ĕ ��Bt��/8�(�!Nm���ǋP�ǪV�
,����r�_�\g^�9�T79ٛi���(������r��<+D���m0A4�";�ڄX9���i�u�NuM�u���ہ-�c�v0�L�TU~�h�bAq�f>_��"��5+���K��og����Ⱥ��w��%�+M��ZqG#�4F쭽fF�v�o�۳�P�H�d�T�K�5C�:I�k���[ᓐH�����0�N���n0��.HH�IkA 3�Y��!����
��L��D�~�q>ڨ�	����=&�9A���i3inh��|���0ax'�ƹ�O�GW�@{�����T+L���zw)�c�n��Qx/���.�F���>�[��ݦ,B >��֚+s�&)��³��\�+�"aID�z��7��p�Uq|˧�;J���Sb�F��-����:��j���������AG��w�#-�0z�h�ƥs'�M�^�f} ?�K��*����sU�_��
�'L�g ��w�d�����^ ���Y4�D��qo�{��-7쀥��	m376ƁlA�6j�Ю��R6P%t:��Z���9�~)o����������(�G�K-\ 4(�*��j�$QC��`�<R/]ʹ��D��ڹ�K��+��G�U��2mR��"����9j�6:zrk����U�}k�T��aݾ�1T�^�DTAY�y�eWA<X��W�FN�7�[�e�[���s�@��(θ�s4��u��Z�(<�wس$_O�,�ؑ[�^��!}������B�P��p����� ~�rG���dK�[��N''
Q�OR�}+����-����b��yoH�<�w��П�OK��a�sN���wf^,�y	�$4t8e����
Y�>���GS�f?��#��=)1
��Rky����ԹE�q��ĉJ�Vf����"t���@J���|�4}�����C� }���g��u���$��.>d����ǂ@�fp���_�g6OC�Il���z�ހ�]w��U�����#PT8���e��^����8	�/{�-�|��G5��5v��٘_���e��\��
�-'���Z�i�۾"��	�IPj���$�3c�.���v��TQ����hY����Oy���B��r�1L�V.8Ϳ	�.7a���Dm��.�~r���r�<�ă�x��rh�e�N��q�"B���B�N�R
���?���\b���-qK$�l-�g���=�F�-%��~`ו	q0hk�rm�\��sL���p���1������¤.�+�N�'O�w)��u5�٭{[��;Q`�c�=����������fs�Cit-�m1Y���i�ֽK5���Z?g���q�{ݤ�Ǐ9��3�dXn�nT�����.��8��`�Zk@х�ZH@r�YV?�%�M�z��+����T��<��ٛN������u���q�?��sR��!/���b\$��I��{�ivn�vv �l��t���\h~9>jqH��B��D�|��
�9�%O1�.�T�e��&�;Pny��ӣnZ�"�FˈR�,��
d+���R��*٫��OÎ�HCrG��R�%��<T�A��%F�IŚ��#��[�L��i�\C���72�{�7�gu|�E6{{eO�*xb�C)�w'�;�GY�+d�.\���V�3��"q#B�I,��?� &�3A�)|���\ ��$G�E����]�́	��(�$�lW-l���Ѓ�ե�pV���<tr	�|ܕF�G3�0���?2):|~�C�ׄ�@�-���u�E��Kި��V�d�:�C4(pyB�����
br�wa��o1\��i9ѐ>5��{I3$��AL�9�����).�68�onJ�8Jy�vɢ�K���C�����@~�n�F�t@$y�A3����'oU����À�����b�t����XACA,�G����+aI6���	��鐫8t~�ûH��0o���,2���>�x��y~�n�ZF'��.��%�ÌRQSI��9�%n6��V�Q;v�J=(�/fX�>��AI�Ή��:����V�W�$�X�}'I�=�}�?��Vǽ"ʀ����8����8-765�:_s�S}�Ԓ�:��:�}��o��Z���}��f�nW�#j��,��p��t�8 o�g�(=�=[璋�Xp�m�JIY�q��^�f'G�<p#�9���X,F��Ax]�A�i�t`��'+��ʏƾ߹�p�X��{'7�$��VG�H��Q��A�Y��%1A���)���'�6�u�;�6KԨ�?�pO�8�s��
��<=��
ǯww��^�㴦��|�宆�h�fxl�^|/�1���2�;x��9�"��`E��Qt���%A�g���� ��d
}�g
�hB9Ϊ2r����~�>�LF��g	H����^��5�����6�lg��a0���*�^�k\�Ѐ�	� C�	�I�-��g]vJz/n�r�ˊ?�w����h愄]D��Ω���#lj�a�՛�l�~8�Sl�i�(��nw]ή�O-��FH2�� z�p)��P��6��5���T9���rL"��,��|��p*a������/�I�n.�1�h��$�js$'�K�a��xҰ-��ݵM�)�z��L:�sǆ��RKuV>���w��{Si���� Da���O���]�[����:�*�nZ�� Y���aۋ\��	�Tp3�V3�hr$�%h�t��Nq��HVz�}*w#���qg*o8e�-i+�ӕ�LJrL!Q{�`C<�?.�F����(B7�5��F}�
��4w<.��ؾ�6����T�D�}_K�����q*&h��}�4�v���9�B���H�P[�k-v�G�{kH$s*-�ˡ<��ba��t� �:�O#�Z�҉��i��K�.v#��&��7[tџ���(^�g�v����uJ5!S^�����Z�v3
�ԣ%o���'>Ct"�Nq��^�����S7��t5���re��+W��Wɠ>/z�NpC�衤Z�S�fȭ�r�` fϸ��r�,�\/�+�K2�#8K~�@��E�k���	�������xl� �G�s��%/�G{d"����[[�BI���-��Çxo�j>��on�wJHS�ɏDmU�أwXe�启S��l>ૃ?���t�e��wD�V�y�C���"��C��y�-�p��'�&r$���l�/��QWM3�5Y�2
9��X�8P�A���Mmoq�����,0�$DW���X�����i�lm�@Łq.:����B���V����p)f���h�N��sQ�=֤jr��mO��9�Q{c��R��e�n���nI������NV
���v��a�5�^5��*����NB�)&��=!�'y՗׸�S�Q���B���xט7��COC�l���#�NI3Y�}hb��w������b��8L�ff�z1��D���/�H�x
�e�2B�2z�7ni���В+&�wn�������ܟH,q	��1�J�J���:�Je'E~B�ȬP�U�Cw�j��3%���h"I�7j�+�=�P��0���o��/�Z��7TD�4�M���HKBt�6�6�4K��	_��8����W��g����Q�nE�"o���~��w9Zdfb���/��0�	��X��� ����Qly�\�$��̉>UOk�����(��Ώ�og�*�X��v��IS�Lu���U}�KZ�ם�j���1�]�D>���_:�p�3��)X�������֍�����ʓa��B+�f�3&�j����I�$� ��h�6�-)�{��˜*��˯��R��4��mg	[�}�}J��'K�� z� T�o�( �j�-�j��i�mi����v�ԢBF�ѴGm�x������B�y�a�}u�wm�u���N*>] �+�Z#�9g����+����Ǉ�02k��|+�p ��%ǀo��=<H�؈4�`�+Eێx��ܙS����d���kN�贀~��D��pTY7�̎�*|"M�/����L�T��\UT}��o�΀R�2��O��Fl��I��X��D�m�s����7����4,�̀R�G�L`~Z�[vLV̑� ڀ�n�!���o��I&�c@-���"�WY��\���š�|��Q4q���-��^P�}����o�~��|L���=�u����/���ߒ��I�iI�Z�������&)��ͻ��2��|��-�l���u�!Y�g̭����*��!YO1n+W"���,*˛�(��YK�íQ����RO�y!��x�^��ϜyD��)M���-�>B��zw��	�.�d����㸃L�0�ᤜ�S��9m��9��Ϲ>?�VDb�[�L��t=�L����K�]�~�l4���jΧ�������X"�.헜��	����Y�x�@/|�jR�����	=I#����0�ӑ���@� ��Ķ�C�ųsi#��M
C3RO�9"���/f�0�}� ���^nD�$��d��|\&�|ҟA���*���!�80������D�}�D9�����~����ҙ[
:1~�=��_BAUi3��������,�{���ޅ����P�O��T�$2{_M�@#����+;�/���f��'p-��u7�j�8G�Y�j$���̧�A1-M���c�i�����mņI��e����"�	���ķ��A���7TTm�j�ww��
��h�����3���o�>�P���ʣ`���X�DC��������>�4(�7�F:��h�W�}4	Q#Ym[W@Cs�-[�/������:��`͏�2�"�N/����u��)���g5��&�|�g�j�.]o��X��]e��s�}����u��H�Z�?85�Ix��k �ڃ�y��N�c�z��0��E0�{���(4��J���k�R(�%C��J����З�'Xu��:�X����X�/,р2�?*����c��h�V���ñ��D�4T9���X�+}�{�ǘ��g��,:��2k\P*<�����O��K�dNȘ�N��|u�M�?��9/�"��6�:P��Ĕ!?�w�%��-��b��~Zɴ�AC͏���1:�B�� �BX�m�1���B䋘|YU�"��V���@�X5A�ٴ/�fw�>��c`G�b�#���ц�zR�����͆;,|�!L�O;�0��o:-OD	����t�r���rx �w�_�μ��7 #�t������f:�~�y΁�53n,ϡ��4���[z�x�.���K�R��,8����3�P����C��o�fvR]x����;Hג4(�:!�zYH31}�L�0�,��p��{\zۇ�@%M��m�b|�/����?��mA��Jf"^��sҬ�t2
��`�$�J\+��DI{�/�!����H��Ґ@pi�\�b�uk8t���<Du|*/�;Ĕ�/q�1�h]��d��L�q	C�J?uE*���@?If=%��G ��fG2|7����i�"�ܮ�&C8�z�_ݕ9Ĺd�[��R��˹�~�w������IQQ��w�DZ6lc���-A���-b�P�]�U�������>�1���Q���q�w�cY����KX9k��LXަ'��l�b}�CY:���v��*���0��#� m:�k�o��a�Kxt�@ٻ�:�Q�=�]�Y�BhE!�m���uCIݦߪ	�ʻ۴ �}0{�9x�qg��6���BGR�,�D���A�w�q,i�U�HMux��V�!x�юP�r[iZV�Sw2K[u��hx9_e���9��8��*�P���6s,��Vڂ]��4.F��,~�`�}kW�_�㯸�r֙^�SF�A盙���H�n�$˒�+��]��8�����pW�2D�y�.{�y��C-Ip�J'	Ԫ�j��V{���J��xz�g�{���Wx�04,Aշ��FOFMOh��s�6�A-�M��X�Ĕ(f��"�JzT��!R���pxv��t�\DC2G���h����s6i�N��0���f]�}}��Vg1���68�ZYj#��|m��l���ֶ+��)�J2:�%|��9Kl�1��.��)6�P_Aq�,��U
/�q���4�<��78�m.�I��^���c��Z����ҟ=��*�`�- ��Ia�n��3@�eCUH�`��y�f�+�ߖ	����K2���V�Y��|�hF�E�J���S�p�H^l�3.�=*@L���/��4��:���x�"#�Ӣ�58�|P�������*L�1�=x6����u�#��ȶ:$k�l>�l䳛!����2��H��ƪ�(6�j�|���6��u(V�N��M�a���R�!w��z�_SkxǹΜ��Ǫs��pTۡ!e;r	���]�*�8� G�3W�|�d��5h@:Gq.�GIM���[��yЌP��\�J�U(�����x?�M4}�ΎlM?2ߠ2:�=}Z�m<��*���ȪX�'�6
�O�����ϥ�m�Kx�, �|����Ag#IX�@�>ɘ������;.)5t���.:�O��\jK
�7Qý6��]B:�Hr���omY�>-�A�(�׻E��E��~�(�CGZ�w���N�-{��A�*���b����P��G��
���*x���Y�Q�kL�"��R�Kp+�5,lކ�al�7���{r4�>*	nԵ."�ڼ��Y��&lU��Z��
���	]pDy"g�w��C����V��p��H�|���*A�}x孧לW2<��zO�R�t�˹��4�H�l��{o��v��X��/���7�/�R��usR��R�����&���Q�+��ʳ�΃��vF��x��\�w�{��©Ei�R^��[�f[�~�Z#�z�\H|�h	$��W7Z�3�$�E3�s��&�vǭ�r��������$�}��)����L�~qS�'ZާW�f��f��'�N�t���FpbS�?_$A�7Er��Ω�-B�� {��<y"fNJ��fj�}!�U/f�6{0�Fv�t�ɡg�R�"c�J1Z@s�T�s����o��/��%A-��\sn��\�o��1;v?7�]���@5á8�8m/�ϥ�����q8�٫[���ge��c������%�ܷw�;v��U��MH"�b@�ۯl�#�ZOz�b��]o�sȒy:��^x�g��_0WB����δ5HEA*�����"1<�R� �r�W�A�� L��`����9�c��>���.��(J�5iV�������ŀ����C|^�oY�ОHaS�\���� S��5�&�"����J�q��PxEյ���H��9���p�N���k��3��+�z$�*�뺺�YZ�e�ʽ�+oԥ�����/�ޮ��B.�	�����X�w����9�SNboAW��8ԡV���_�K&=�=�o��� �q �����@v�tt��;���Nt�ʹ����5���bsնD�O"�R)�;�3�`��r.Q�<F��f�:�Ơ<��{C1�?��%��{��p�� �
<H��4�m,)�:9=�N�=[�	*��'2cΤG�磺a�W1H,�Xpۙ���?�I I��I"1vg�6��ԡ +��0�,%Y35�eE'�g�pؤ1���
 �����?)DF�Af]@..@�]����yp:O[�-�@�Y 4��0�_� �J3��N�t���K�gm�M����ֱ	s�W�|�'4b�_f[pS����2��A���I"��1��K<>S��O��ŽH�oJ2�D���(�̞�w7��'��*���� s5�
�*��{,'�E� w
i/M%*mT$�kFH�	!��!V���\׷�n~�.J�S�u	Ǔ;ˎR��F���䩢g��RUq4��0�8��5=��_�T��Fj�����ei�OC
4� �;�'`�\�%���RB�+O,�4!`4���_B����4��O@wU+w֩e��H��ea����z�z������N�A�?�sq��9BȾ�j��`	
����8߱@D��-�DY!&m����rw[�"h� T�&p�����2����0�8w*��W�Gxw˜^Sc��Q�1�q��I������y6�0WG
�b�+����w�CF�pd-Ś��Q/�3�><XZ\-Ye�`KX�X7V��"R�C�E�MUnl� ?C8��M���s���ēoM�>���/�B����N��Ϯ>�qnZ��ջo�Y��o��hrJ�;�6f_�0���z	^��ᛣ�pȓePa���b�8�6<��p^@AX��?.I��ؔ��rx߃c�>�h�lH���1�
k����#8$5�f��9��y	���L��(��1b��d��Lq`AW�'����d0>�����l�s;%�����e����}�p���G�0��p�jև�/�3��"��v�+�zE��n�6�`�;v�c�͟���ݬ����1�=e�J�w��`0��!]GL�`Ҧ�k_��X�a���䙽ˬ�N��)��ߏ�a�3�l4U�����5�MA��!*�UڥY*t�ϥ����R���D�a�E��FF2��3�scl��,��x�Hٙ�`���:�� �;C���M�vW�13�W7y�d����զ�9�����p�0�f]%��?z�!�nN=i�/X��CS���I��gN���C��4������H�ͳ}����.�Q(���w'Cxap<�8�"�t��b,�����I�������M���e�D�L������a�����4>](�Cfd�q
����U�v���pe��3����:?�]y˱S7W<�XG��6-��k�����*~5�}TL1ڧH�`fS%A��ۼL�q�Q\l������P�y�,o��eVi��Bq�E6�o��l���W�����ݟ��=�ip�l�M��߬!�����r�*.y#�\U�V��6�H�k���=A~5He���H�V S�����D�(+�=�ʲ�`:��C���'�F�WyŢ��)!e��A[xG�E]Y�5�H��^�>�9U=琯l��)��hB�	K{$3�
2�����2���b���<�����E�i�ܿh�(�~���#�^#yC�D�\�wn�:T�ם�د�e|��C�B�N����~i�!W������$.��e(�磝�O���Y�Tw.�?u�~'1L���[�E&����]4�y�dd$��,w�O��0$1!MW����ˈ�O{�>���?aFց�ј�ӭ��[�л���T�ђ1$��q��TjW�bIs	3<�ڝ���6�r4����[h�)�EEn���}��Hڹ����p����3aP&m�u�m ���/�aW��3e�ځwB��y��hiyA����Խ5��H��[u�/#y>�������s��UT*���n��~"*��jM�'�u�5���
��&�S}܉��Tټ�>OC��{2a����8������x9�w�]��B������RXР�'��~b�n���(]H5����D��Z�{��:���N�]��v
M��b��1�l����R�ڂPM�,v����2�X�Ä���[�4��v�{�����8v�v�08s�����	��g����R�LxU�Rj���o'�EXx���-����3���������&��!�c�ܰqM��5,B���6��;/Q8@�rsҀ�C,�<Sz\T *m&�t5����?��2Ct��Kn�xɔ}M���s,Ꮪ�G�w�[�X���d�b�89�,������$Y�im����&�f)91����|2�IH�wL��-���]�&��@�����[`G�E���$������;�j&� g,��j圃g{�V��	��*�URW1��N+�}1�D$�v�P�{���5Ah|Hڮ��r$�Q���/�?hٙ((��Pě|�V�n�Tt�E��G�	�;V�D�L�.� ���.��Hn��f��?x��m�$l�V~Bv��#���H�-�Tiea`�Sg2�M�a4QA9�c.�o��7������6\���	"��hbNn `Pc���WT�uqR�QS6��`�V~���\UNb�z�
3��n~Sqr���")�z�7*<$m{��	�9_&b|�7n��=&kN4N��FH �YG}%�m����U����S%�JwK��

CU;�aQ�	��϶��V"TQX�#�sK������F�R�肋Lp�3 #�unov01�� y��+Է�ĳw,�Z'j��(���ɰEO�m�vF}�W��"�e�eS�-O�$20�g O�)�$ �1������V�02�<&���F0����;p-�'�-Q4���z�Z�Qh�Eu�D|�X�``dH�B�Y�`8�H ����}�V�q���1��'�yW�t�����*��]g���
��a$Gs.�.Z�UI�����B��_��mң�Q�gRm`�]���:�JV��������$DrR8�4�R��`dL�v�N�$����y��)9kHc���F�|v�ǎ�e�ؤB��Ι��@�'��IT�X����M�&Bo��e��_����,�'��m������<6t���k��%�$$ʥ��s�7��U����ԇ��F(����x��f:�:�N�c�2n�B��x��er*~��ҡ����J��hX�ul���?'�&T2>���0�j+�"��A�Z/PR���� NWP�z�����"��ʟl�|c&p�&�D<�s�!��aiHHz��y�����鹡a{K�GH��&��=�)��g�]�+�nM4�$s�u�G��Zs+�˅�G��[4��±����O�~�ޟ���$��0gn���Ԟ�KJ��*#(�h��щ*a������&�B��/�p��=0���_y���ú�'���U����U�Ku�߷BH�m�`V����x�>��b�ZcڲO�UI9[o&,3}�����w$y��:�nxZ,M58�(J��=8�ݎ�^V�d�J��@<	+rB]���y?�S��q���ŵw����˭G���@Ӵl
� (���φʿem��YÁ�J"�j��/��Q�G5��@�,�B�6B����[��z?�q(��E����P���F�|�C�9pşfxkL�^%7x6w/��c�g�� �ZƽD���������,�l�JP�}�71�GP�1�����">΋$&����9�ߦ[	zΜ>��-�N*ܚl����{0�5�~�i�f)���[V>�@O�9>�\��{��R�Ҥ5�3�`��x������&L�`+�r��8I�Ha���@㎃Y(��z29"T�A >�?�]5�%��������v���Z6:Mrܴ%	Ww8�
���#����͂�K����Mb���;��n(_��o����E���)8J1��I���n;�Ӫs6쳄� ��^��ML]����d�xFj=D�!�9��JS�R�������y��!�k3ў8�������H&�v"Dӌo��F�?z����֏rY�L�M.T�Q��}?�'��E����/gόX!J�����|�v]�	IX���+��i��H�g-�a�b��Ȏ{	H���7�����@/��L-⍀N�3S�J� ���:�UC�M�|ĝK�%�:�u�#�U���Vb/XZ}�8�#
h{)�Iw����Cb��ɦ����i�u�	&-[f�L��&��-R����At�e*���m�����.��I�	ڕM��,,6�&�px5	����4��.� b��"�M.!򆌮��̞����㭎+|���=s��hAM�rXR5g���Ko���E�
�e{�����q�����iH�� �
��G�K�*ք9����es|ڤ������$�f!�]-}u��&�{���;��Z{���3]��0ն�G�yHU|���m��̲����vl�Q�9@�T���V�����,�}>�����(S ����^��