��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1���e}ʲ��cg�t�ϙ�a�:�KR�%���ݧw���ȼ�L�����Q ��UB�j7�o����fٟ8�1�X�:p����U�PQ��B�˞"u��d]�6V ή;��ӯ���V��� �-�Af�hL=%>���؄��Rވ�$S��m3�"������D��|�X������F�'�/��0�%�j�0�?g�!2Ńq,���5K���
[!��ډY�@|��]CD��F2��(�r�4�������mr�j⋆�^e�~� ��# ��yI^cV�hH�f �� �- -�����@�0*��h�[*��\�6�o�7�R����d3���%�fA'=������D��G�Zu7#��h�_��������ɜ����\r�����ѱ�zW��?p�0��=�$$B�2�����+p���
�� �]��2��{�.�P:-���7�xO.����T�9�r]sl"��U��=�����/�/x�*+�IG0��?�Z`7�_O)�t�F�t��T2�NݜjB�L�T^�n
��g��[�ᯡe�󳶤;wK�`=���z'C�7���{�ό��"���m5=���7��g���ED�Y��� Ki�����.�U�k��82.dO��U��[y��otx�Ǻ�"��n���;4f.Pp��X^ֳ�0>�ʥ���k�6�}@����f6A��R��� /��C�F��
gՙ�������ך� us���1��A�7�G�D� ^;�1xrVy6�c��v_X�p�0�M�;��"}�u�3�3���K	�_��j��WA��3���nK�x�|.��dWu(��6rR"@���j=�[��*L��j�?�:��Tm��B5����
���x�gu���]�jl��q���[=3Q�9�-�l�C>�]%k.fs��Z>�y�koQ���hA�S�O&|ZH��!�(�i��5����4h�BH]��9���� �8��Cuϯd�mc��mu���Q~k���d_�ŧw�������a�|el��q��
��V|�-�j�Zs\:�t� ̃4Du���x��������YE$~`7�K�Yf(� ��J "�Gc���Q�_�ڜc��,Uҥ_bG���%7�ߚk�WC�6��G`�Q��W�
�"|D�gk<���cq K�v�Į"��J����B�#��������YNE��r�&V�y,�,ߚ����Ը>�CP�	Ĉ���_��.YU�r�bE�< �6��A�5�y�I�D���0��58������y��H��aĎ2;$������8�Y���Ey��K��0 *r���Y������I0�p�E�#`���7�C�i�Vj�)��M��<���uh��:�lO���Q�-=��O���{��$'�(�5�IK"[�N��.����?u��NfX�$��
�IP�9�t)K����-� �}W��AfA6�Yk?�+Bb�|X�Ů@�Op�D�O?�fk��)���3q+
Q��a���J��mF�2}�`EℐbB��(��T�x��Pf��ā\�=_.�W7�ԩ���2W�C,9�K��Da�^E��
>����srk�`�y¼Mг{ʥ�&���Ub�c�yt ���V[j�^��^.�h���!"T�Q�bn�>p��wv�\@79b	�4���-�;��_iȎX��צC˸�@��|D ����z���{D��ߑ�DZ2��N���Z�`î�T��0L"�G!�����g@j��W����$�o�OR���E������mE�������.$������hj��N;a9},�j�J�w2���S��ƕ�����_�q���h���f�Z�����f���p@��9UM��E�	�`ͳ��Y�����=g�Ը�'������u�7����v�z�րiqkkT�1�HJ���([M��(+E�������h���Z0o>�Zv,�������fR�I!_���FR�a��6����G�E��
��y8a%'� �%mKr;S��|)�}���#'�O<��v�#�f�Ç��O�.ſ~�V��ŋ���pd>
>^�O_]��-�N�{Ƨ��/N�̔��Wk��l H��F��:>G������9qߖ�h��<���h6���i �;[1@62~��K�G5���tf%a5D1�H�X
gZn8����?6��?�e4�_[SXۇɲo�q@���m�˵䝣qE_�'2I(��y���pO=���5�h֠��.����\I�T�~^)�ʷ<}�~�ѩPQ�������A��7�  �ό�+Z{\�����{N�:�K�a�E^����d���Z+�RYŒ34e�T1,�%��M���ڃ��.���*K��^Jr6�#�^"b��n���"�+"4
~�����^4�AO���"V�!uiћ�BM&���*!�	�����ga�!F�������>���R���]��ˣ��pk;p�����}��	f��-��� w���%��\
������#��pՋ������TX+��X����Cz(��^`O'�4r����d�!z�aH�;>q�b�J�x��������\m�����u��>�����;�������৴2���>08��W������)��M	
�eh��S�<�]��Z�Ē�ۍ��#|�JGZ�$D�먧����x�N�]:SM[)6��,�h)�xk�/�!v�ԙڙ톍��?a�'�=������(�N'��7b{/�B��
������S�[B)��
u7��5^���E�?`�<@S`�T�ެR�A�k�#7��[K�)��4��(NZu�R��Aw�9����v�Et9aQ�;'F�R�qk��Y/yC>��V��6��w�#m�������5���{U�bp�=�!�d*e��Iq�y��������iI��4Tp�!j� �ndP)���+�tf?�2�dK^���ܜ�>��X �������5�`ua[y�������=�M fb���T���_ܣ�n��!���YwK���[��SGՕS�F~����vk�Q��@L�Y�^K��@p੽8\�2�T]N"/rHc����()�gnNj0dPJׅi�Ͳڏ����閒���+wP��{�\}8���#�([\B���*���&��4 ���c�g�JȬ�4uG�������PN���e��59��yQQ�؋�å<���|��v$��=�y�L:A���r�O�k��0ṃ#��A�p���K�l��N!��y����Cڢ�$��.����	��1goܑǞ�]�_*?)�~�X��t<�U*�K�!Mg�n��;��^n����Z�\�x���k8��{y�B9�	%3�Nr0��[�*���Y(A� k��=�#,6±���C��[�8]��-8!�Ŕ���[��ɥ\�����X��K(30���������F?a�1ۍ����� ��^TC�7g�����UO��8x�Yd&��L��5�V�br����NȽ ר��E+�.����U��~�-��������Y$乮�[�>E&�Ҿ<��E�����:T�#!�U	0����w�\Ѿ� ���]�zՈH#�)^�]ք/EU]�������ؖ�ހ;��% �&�Ј1�^9����]��
�'�/EIT�:8�9L+B����$�F�{biwo��W#"9#�M��V�n2`��dL$r�C($�c�7�CB��,h�
�|�?�(�f�thʝ粲[�|j�C>K�}MmL�|�q�3L�Wu�90��3h�|���3=˴�y��E�i��{�-團�u�QQf�%�z����V+B͙�N�9*L�y�������x�KR�� �����f�ä���aO�������y�\��H�����p�QO�b�w���xI^rP�L:)��G#c�6�\���6,α�D�R;4[ċ�F7+�:L�����^k���=qj�A���4��Oo���H�od<��},�,���l�c˓cn�L��?�����H6Z�<�֖���ù�qi�AHTc��)>���-)���u��\�� ����z���,�c�q�V�-d[��^zQ��f�m���� �Y9�b���f֐U��[��%��'\z٤��b�0�E��d�q�T\�G=L�����w�t�Hҝ�. �8"�[u>~�3��F!�h�K
�����k��t`���N�ʄ����~4:�"���FͮZ�������.��Y��sėI��BU��8����2�־�H�5�;3Q�B/�>�	���lo�LvV^��8�נ���x�7�W�vN� m�Ԁ����O3�-�9�C��<�B9�e5M	+�?�Q�
�"�˕�=�G7�����|�Z�r�,�{��>�X�@�o˷ld�Y��2��^Xf#8���G���򾣵���Ri�WNE{���E4#���A�I�)��֭�măj.�*�X?(t�S�c���z��⒌�н�-=��]��qsJ�q[�f��5�dش&�{�+�BO�E�e�x��~%]���֟B
�u�`T��"3�ݨ_ve8{@髀��@�
s7��$NOnNn%��f�NZ�"w��i�b(Yߑ�; v;�mV�~����Ib*aӀ1e*�u��l�<D��N�C:g����t�7�vtw��~�TaY�w���(��u1�C�������_���n8��l��\	޴k
|�b�Y� �re��h��<ZÏS@Fו���1`�e,m���ҏ�)�Jb�0V�h<�k�gV�7� �����~���F�y���>#J�`��1�Y9�v·t��
��U_����l��` �-J�+�����7�V��"�n�����?�n��2�o�ˋ��ȳt��YhĲ�����/�!U�����l�W1mVhR�_~�)�����j����~����#P�K�4�u�ʏИ��{�����3�W�$Av���4]*x�z͵>� ��^�FX����r(�?�b\�<|(��H���R+��X8�CK�M�)q��*����F�Vq�gk��,���S)62O$5�X栚؍@<���^Rq7E�?��J;z��S%s���c�s�q@���ռLQ@Q��oR�t���6��Yѣ�F@��j��`�@�q��I���h��R��:k
��(�j�ft>j��6�3�a�M�ʈ�m#g��e�V�*RWk�i���Qc�(n'��Gx%�`m8i7�s��RS�~��(?E��⡻�g�Kͨ�4�u.���Y�(r�=,v��U�`j^���R����>��{��Qr���ū�ɠR�<�rB\p²����v��k՛��y�[zo�3O��������	� Ŕx��.��3�C���4#Ӱ�^`����O��ԪF��9=%tu�j)e��nl&��&����?�~g��Y�w��#����a��3��o���* �����'������L�7ߺ!]c�ah�-9	┘���fN�N{�����-��a����f����`A�jn��d8C������n���yFOy+8�����!�F�tb"@�9M6��\��0��V[X�< >Q���
�n6BEl��b� ��V4Km,E��Ø�����1-Ѣ_#&s?��%�e�r�ۣ ��˕�ap3�)���0�d��5GZo��hz�ێ��
��g���-ɞF%W<��A��ְ"�\���������kyVX�������ۍ��{_��{��X	&G�'"��u��dR�k�K�����,.@�̓�<phi��s������3l�c�kr^�C&��7X`k������V�,#0��x�q���U�q��h�Z�4E�i
�k!��>���Luv��~�ݔ���n�@1~�W,]�&���9������9P(�]�����^���uiAyb���������&G��;P`���ɒj�㧡@`Lu���>ྯ��m�	��k���JX�1^Vf|��
���W��A]�Dy3��la����{��Q6�ە�e��#/���Kr ��|����#Q<�0���Z*��F)ǣu��AlX�&&�.�N���� �}ަ,(�7����W�:Y#�S��6OcT�wԛG���Z&D�ɹ�� �Ph4�-�����@��b�N�Ӟŗ�>)���g�bu�u�yi�%2��#�$j��˯�b]�n�ݿ%"4�Hq˘ד�\e����g ��f��H��Ǭ#�Ӣ��w]*���a�Fӭ�H�uh�w��Q���+ʍG�|�F�ʋ��6\WdFL�gb�r�B.t��F��ag�p���zmdO6.S
?D���@�� ���t��h� 9N��E`KN|��������u�fy�ς�_�x�x�y�V���8ݖ�	�M lߘ�z�4옣C��OGo1)����4m�!�;��@�ͣ��Y�H��Q�qX�,�Ϊ��ž	���n��o%��:r/���P�����>���|Ct���q�s&7Ɂy��p�yz�Ԓ�·��MR}�ٮF���+*|d�#����:n����ȏV͜Pl�'����y}��]dք�gꞨ'�5]�9�K��)']y�	�!���į�c�oY��^���#�7��=¨����I%�8]�d2��!&�:ku �!$��g�����ˏl2(�+TIr�%�:��RN@t�i��l�Q�҃���jtŅ'�c��8*G)����,��S�{*�̛�Ճ%��m��
^��@�z4\c�󀍧�CdK��/&u8!�i5�U�+��c����3������EK�ڈ�����lDap�R9�Wڶ�I�8A� /���r��B���@@B�Q�a�V�U��&�R��oN�iO�9δH���ˣ�2��1s?���y;�?PX�#�=��*]O�D���F������}�C���
�S����8��P�Z�e���MP{N���f.��e�Ř�AD���T�3\ݹ�q,���q>Rՠ�6�(g6&,/I�����t��A��
�R�Pg�����q��#�;�W��c�oٳ�����]A�b/~R� �>���Z��3��0�?���v���I��I|vLZ;U��J�Odg=�|XuZ����[�]�4s��I� �[�e7@��_��Z�pF������?��e�0��ڥv1|5ތ�?fe�l���2��qu�t�L|劾�_��l��[[�dDؿ\Q՟ps\A=��$��u�'���W^��ǭ��d��2O������㸈3d
��d9��ζ,-\�^�#�Ea�K��N�g���]��b��c��,��D�V��g;�j!��j�A�&�+�R��2ŷ���z���I`^?���N���E	����Q3H��I�7�����ug�!wy���q��̾�q��|�<�ǿ{V��Cs����#��-��.��o�Wk�ߊA2$W��AJ��=q_I�!�ﺡ�G	+2?�{�_�N�G
�LF�	&�:�SS�\�r�ސAv��n��zmB����X��FF%�ʫ��������?�A�8כȟ&Iʙ9��{��١�������+u��k��Rx�^'0Tp�1w��[����I�tt�}�7�*�8uQ��� ��z�E�C"�����XH�opK��+��N% *D�_a� ��1�J]i�
���w(�6�p�zV[w�,�����@Й�����M��/��ͳsu�FP�J�T�S����t}&բ6�"T��������<t qS��X�Y� y�F�Oe��y_�lU�gF=�B����;���8̬Aq�P̯�M��R(Xa���Y�thx/�%�P�������sgg�vV�L=�>.�����~l�]m�z
����`0��cfRR��dd"�t�L�08�Y���K%����n��� �/q�l�~Z��;Nܫ�,�h.�6{�KmɠP�M��10r7�A��s[8���e�ʻ.�m����Z�9;�]C-���ЖvCty�q$�V��ň̜%'8i���K���-'x��P�s�j:���P���f�0ĆP@M�X�'Vʫ�ۜ���2���Y�b��F��O}*�c$�n�),��G��k��^��?��
��1WQ�W�Sg�a���E�˙�$	��q�zOC�;��x^����@p Dn����e��������(�-����8��ç�Fu��-f��J/����Tr2�^*ּ�aW ��������e�'��4����r-*z)�J�j�:ܰN��n��Į�¿¦�_�ii?��o�/�VO 8�3��L�]�M�z�`���@��Y��f�~k���3�<�l/G��聉�6��v�]�z;�?j�hhR.�p��#����P[2 �念����m]����IC��h��ۨS��GH�:4��\x5�O�B�y��o�r�⠛:k���~7��kyK�q�W�^t��U-��u���5Bh��zu7T���i�ѩ��rӰ�Q���~@��ٺ��.��Ek�wg'b	lL:��d�}�&�dUYB� ��y;�mJi��d��d��#"��H��F��M������"���;�ka�_^C2�g��6�g��ф���ބ�Z̀�� ��l}Ƕ�q�	h����S�B ސ
AcP�X��a�1�8�;IL7JN�r��M�}�����w�v�V UC~gW�I�T�OF��`W�$���-.f�:��%��δK��f+"�)#8Ƞ	Pl1C
` �@I/��wG(�������ޥ2A>S?&� /��z{ؔ捻�[�Yp��Si�!d�w�"�%Y�Ye��ۚ�<�������a{�)�S��2`@��&���3@������H�ѕy�:�ygޘ���(�O�r���ZߕzeR$��������o�Šd/��v_dh���H��� �ڡ���~0��>Q_1R�E�#w�R��E��������TT#�sy~�M"!Ս��1���H��M=��,jɛy�Ay�@V�	�,��Īj�V1�Z%��M̒T]
��HR��}U{b�?�3��`�t;��,�|H{g�j��(�b�������|��Wqb�ے}������p3]hͰ�����֠Mӓzk2L����a,��R�dإ�Ax�5����<]8i��
��T�����PgnG�9H~��w�>�)�>I8�g3u� ���[�͗W��%- >,w����_&̔3�M76�S) %4Ð<��g��Ț�
�PM����Hۜ���"�sȩ�y8����Av�r��B�ӷ4�)h%�����>�P<�]�a�@;v~��#����"*����
z=O��C$�h菧m�$v�j>��ÍP(�t�~�$+Ȧ6(�^�vO<g�>��u(�i��wGe�<T�epYT���>84�Y�Ң�Ik3o���w��z8��6���H۬�9Z>r���_�@!̉�QM/��B%&��;M�Cڠ��C��t�Ӊ��Rdԩ�A��u�zi"�`r:q<�F���daܨc�o��v$�ڍ:��o'�T��̆[�����-�ל����`P������u���3�0�Z����I��<;ȭE� y��-	�wU&�v!J�uF�_��Oo�̏�:z����u«��~v3��W��]9� o8��l��N[���1di���c#��[��RNK��
��4��M�̆�H4���mI��_��d;� �	 ���Z��}0�P�I�^��r+�[E���o<�]7-�(��Z�nV�^����3!�׫z��C��8�v��M��ʤ�85���e�#.s����h3'D�+���e�E`/uO���f�V=̇�rq���>W`�;��yg���5���QOY�<�(n��ı�Ϛs���I�;�-�r������W�A��AT��K���A���3c�9��L��(���<��ӎV��� ���_�)�f��wQ�6<�]��=�鑸���Ԉ����mԸ���p=By2�5�S�I]�M��`�E����~܋�A���;{�����;З����-	i	{��ԣ�?+���M]0,	d�^�ⷁкc�	�-	6���ߩ��CJ�O�6~��o#���u���yd�i��E՚��7$t��dm�Lul�!�����v0YF?#���Z 4���~�(gv�0fߤ5]��H9�Vg@zii�����鸘�)K�
����8�D�3�}$G����{E�&�d�/k���J�Ĩؽ�ߟHt�#����7fi�ڷ���l��r���á�I@�9�%`��h�~TV��[��%�I5��Kx�}�T ]f��x7l��ؒ�+�<� h%�)�!��-��{A�����t��z�]����W\��3Q�)�.J��@U�+��~=煍g� K����(ۈ����������P�"�O� �H?��B�;�G|��g�>�Dp��8�?�.�x��Sj5����3������]�Ά 7�Tm�}[�Sr���괮��T���A�Uz������<f��p�璑�L��5�΍�*���'o��Z#�aoL+ �
�
[���V��G��0��zi'�"�Y��[�;g7_]��;I�Q�D_�D|J��ǘ�u���*\G����ɍ�J�����b:7���fYJ���1<׋ӂ-X��k�h��`��a]�V��Ƒ�V��X_�U:i���d��w>窔7�<v�Py�Ҙ|/�����3h�'ؙ�VƆ�u �HD�Ut�`e�����)±# ���s�1�� =�* w���,S��X(��s7���6�sD��{�[��9�N	��7��.� ��3�d���#�p�Q�i�x:׊z�!F�*?O�H�N��@5�pb΁a�f��D�Mbp����[%���Mv�y��rB�I/l�	�YWXEf���6��2��w<h��2<��;C-���D�����0i{!��^j�K 1�N2���,46�v��Zn��
�C�E���i�PT����%㝫�?��%�O��
�)Ϣ:Ƭ�z���X�	�����˟9IKp��#��+C��A*E��}��~�hf�8�ϊ�IP���m[?��p*�9��]l'��:�����<�O��uQ���H�~
%�3B�=t�������B�/@���[&�C[@�������4�)�~;]�G�pp-K�0�w��-l
�۵��L&3%Ŧ���!l��m7}�ͦ��<[?���?�Y��m���e����B����>EM����?Dh�8�T<��� �hD��W��B����{(��&�n����pY$[��]T���+o�KK�׿T�dK�b����	 ݽs�Ux.����.��C��������:(�1 G�����DA�,W�t�v��閭���4�'�_�ػ���)!��Z�h)H�nL�7��;$l���PH?������e-�dG�^���)��[�+��-͸�WMu�+��G����2�ӄ��d��I5|J�v95$,�8O�N�2,	���#������C�M�&�v6�s���-ʆo湴o��j����ɦ��6���$��]������b��
T K{������`/����5rM�#�K�zK66�=!������f �]� ��f�K_#)�2ɴ'FN���K�{������6�*���CAٕR���V��?bY��YN��@�98	�{NQ�3&�>|�������T��'�����vE����p�Iw���M���Ш;���(��DYB�nk
���!J5M��Z��m@�5*�֋@XL��"��)u �|�V��9?MAg([��u0:�8���v#h�X*�*?'��l��6kŃB�=Ė��C��@s	A�����Ē�����T�ĮPe�o�� P���h"9�J3�~�i�%).n�b3DS��8x[;f����j���Y��g�R2���`^,q����ө����v����;x���^��9�C�G�uWwN���3���g3���*M��!&�$v'��?���_6�{R���,p�z4�mWC����+V퍽�	ߐR����J���{e<+�����~Ǵh�ab��x��i��VZ�ܪo�1��Ţ����K�G앒ջâџ��|[ �>,Eῷ>�XûpMg�N�������|�t��-ȡxu�̀aH��Y��ꊈUee1�I����e����#ǅo�����8�k�T�i��S��ʤJ�D��k2��Z[q׺��~�9����a��L*Y&���ι��Y?_V���_>rr�3�L�[���?ŕ��ڦ	;O� �O}$"�M�"��bo��X���Ѵ����W�w7�l��:A�#�/v��c�δg����[|�j�x�ADT��F	��C���8+�n�MaP�Tc�AD�T
�W��*K��d�`K�/�'|
w	�U���Aw����}F��#�(a��Ie#ۛ��T'Ϝ���>=�hײ�;ڎ\=<pW-��0HR���rHu\0�<����,��&�ǈK?\�����8�T?�r��kfC�Y�5�6�ȗD�Ƣ_����O�R��Y��H�u>ps�(8^��oT�c�|r��s9��:��h��T��8�D��Mݴ"� �xoӳ 8^��b�v�ַnЃx	�T,����x�F�*^Q�>Á�^#;�s/2�&��	��~���</����w[��}�^
G,�PG��[@��me����u��XB�z��>��e�e�Q��~����^�v��M�Axa_�9��Z4��+?Ċ����ۤ��:*��(�
u��}qM�g�D��ԉ��C(k�sGAP`3	�_>cT��j:�]k�?b�a��(��q�< Fc�H_(��)3�l�iEx��3eT u�?�#HAB��k�M����{�L
���<6�H_��>�Ǯ�ȜK�9�y�)ӎ*�m��|4�^i9v4��.K�6:F���}��K���fk����0r���z9�+[^5H�e+�F�E����?��P�NX��`��\�g���kM�-ѨP]�ؼ���H�5����|ly�^�+y#}'&���&q����*���@�L^ܜND"�2ͥ��i�n����nv]����� �* ��l�e+��1�P�{:�������<�E(����Y��IuU?�v! ikc'���K���4�£>��b�Y�يUq�̻	}��XKἜ�Wc�٧�~��'�0��մ|7
��Ƌr?�"A�MbՏB06�X�9�Z����j	��K�*�ܼ5VQ[T9mP���4R��N� l�����䖹|��⅂K�N��>����m�6'8\�R��4�0��҃���Q�3A���D��]����0\��1xw,���U���[��9�9����>��և�L��q����v}Zv34���K�k��*��7��O�5�?@�d�5���:�;������ж�th΅zƘ�u��d�H����6��w���)�j9Dux�v�'E�@{��Ռ6~U��i���.4EO�Hcy��"�j�,{�zKpG�/M�
���N���o_�a���S�|.%Q;�� 1Ҵ86�o���&/��T!G��d(g�@$���7,iq��|}r�o�zn�ث��� �*��jawӚ��8:.`�S�o��U�٥XS੟w@�����BV�S�E�(�8C��\�y�H>�J��co�ïKB{'�z�(�d
�� ���R�/�n<c�lZ���i~���m�s%���-K} 4 Ѧ@��[f×�~11�/<�;6�Q��>k�[ص��Z��?�'W�9��-S.6ګ�2�@@�$3���2�-Ό���T�q�&�����u�x?��Z��#*$���>��8���Z��Í��hqm�pjCB{$�7��V��!�6�d"?.�7 �E@��ZT:F����c,48����`�����!ס 67�V%�9���/�XWNH�k��.dܦӝ��a�j��D����[�Ɣ�VA:��KĚ�6j�J4�sǣ�h�ҵ�R>����\I�G��N�
�0�����<�m��>.�� u��s�V�_����J �b��
!Elh�d�������H]�d����z�8�!�r�z�ʹ�]X�����fDt+b�S^���@U��-�Sg�/!3�l�W�8���5Y-�1+5�څ|����EƲ���cY��ݹ&��E��,\��"�Z�����&��l���3�JR�`~P�Y�����^�{9��~C���-xÍ<��ډ"|��"Rb?���g��jq:<D�7J��j�A�^��l��;�]˷�l�#\�F�zg�S:69�Y��߻$c���C͜��J��p�}�%]�񳣒�3�;)���D�z� c��J��:>�q���4�g����1�쬓gIX� T��h�!����9sc�K�|�D
w� |��;�v�KA[������ݥ�9�9#Yl�L��֔�����ߙ���x&H��L�/J�O��q���28N�����ww��a�o��U��4u�;q�f���m�E�fH��[@��EJrD�r��!�!�{s�⥰4b!� �Em�a=���k}�?h\4(n�BG1�����#TdHRϑ�S������F۰z�Tq(��%������DU�"(B��u�y"�/��遹{F$�K7-�a	ǭ��ɘ�I��s�X=�["ïAf=��a�cP�����dD�y@K3-b���a��f�!@���V�0ċă.|�η B�B��CT]�jYm.7:�Xص�ʰϯǞ�e �iz��)�V�:��p�i&[ne�tju�"ꂨ�vb0��_�t޶�.�o�V����o�E<+ʒ�@i�}n�:��z��v!�>a��,�j2��}�LR�����X���P�C���V*���*lR��R�����s��*�-����(Am���jC����G�����}�ω�|�-�t	��2W�7���H���p����Z��(�=�1SF���	���bO+.�0x�9lkE�Q����0p�A�~FJL���!�\��k�3<������X�0堈z9=��esr8���@�SX��7��Fg��0x�_{E>��� �yT٘�R	ᜋe�twZT�d��i�ߐ		Ͽ<= ;A{f��C]�����������<B�J�Y�Wf
��?4%��%�.�8���������f�lKb�'1���0(Q����+����9π
��6Y>*��J�+'����>��V�Y�
�!���"Co);������9.Ee���| �4h�S��b��H��t�d�Z+�7į�ˌ?|0b����Z��wJ�';�n�p�/���� /m-���OwwI�Q���%x�5~/ �pcXJ�0����R�F�WVl��~�mIv���S��჉�ē��O��P?2�q��ю�z��n(��my� VKsϞ���<>v�KD����J�PpZʤA?C�������"����0�&���'���!�@�ê4�Ә�m_Sw�΍�y�B�! �������O��;�C�>���FAՐ��6��KOd��6��a�m��xI$^C�`��?b��UA1��V��*��L�<l��6Q3\[ɶ�s!��ǅf���N�^l�	���3sT��AS�u�>-���6�7ό���Q(њ`�K���"�Z��-���6��R�;�9�Pf\V�:]����ϙr�;�L�����z�-n�	T\_�Ek�Y��![�i�(��칇��D�f�$S�hܹ�����^�1l�[�l�P� ��+�.�R���yf$�'E$�\��A=<�U\`]��6g��F�ke���uy��j�'�Ľ�$Y-4C��Qt�B��u=)Aw}ˡ܁Y�b��!��7v!�?�!��okz��(�ލ3�.��ҙ�	`����E:�����9����g`ɭXf���?_8�$"Y�}R(a��sB�@P���������z�W8�@�c���׎��P��L�����mz�3 �%����!g�2�VCv���>0Ĺ�"+9����r������*�'��8�LX�L�Ļ��;L.{�\	��kf�Qe4v���׾�r�.��۱�5ɡ&�̵���|h�G����OW2��{1��7��ԛAb�[-,ᮌF�����cӯ2��-���O�ϛNO��訝����_)b�l��� �7N��i��n*����G�y4&��+b�_qf�t�{}{57Z�zT��g{l�p� TL-K���#�*�4s����l��敃�f�{�����}��U�il`���
��;�G����2��K�:��q�v�� �L��>-�����v�ӣ]��ng��)�%<3�o����(������)�M���C6���㢼�u@&PiE̔��r���Q��]��bI��\�	[�-\��393��Z�i��h�_��>U:y��D/ﳕ��Ɛ"/)�=�������Vj�_'��PE�8{��E2d��~��P�m� m�+��.�佊��i$o��qݡ8�d,z3-�dU\�mb]�����o��q]�ز-����� �J���CD�.����rR��Z�5��cc�N!�rl���h���h��g���e�ઍnx�,��>kd:\�������W��oJ
Ѱ��������'��ɕ(=�*��uy�8���������v!����}��Cx��1ݟ۷ș�LK4����
=9n�z�Ŧ�
�2�Y��/r�������N��$$|�(�0���|>��m�t�[�*�_�y�H�G�"���Ɣ�!��F�YN�3z�쭬�4)L�MQ��BM��7"Q���e��f�!�����~oK�nb��i��#��!��1��?:C��D�����2�B�A������ N��5�s�)l�9�h�F��+��P���Z�Y�S�LE�cd�&~��e�>�O�O5q�B���k"Q��?cQdy�Z���΋o�d�X��=��"�m�Dݚ��?��S�~��e�i�-��]ć�"�B֑:�&��.$�՗�t=qH�'���@�ip ��j���ÿ��������{hѲP�扖����B��']��H�$��E̐�G���:;�ǿ�3iMX����x� \�};�}�w�d�B��������8���-�!�y���}A����qa��2o�[4�f�jZ	q�4�W�4�Yq��	�ƥZ��%�����x%qs�(�,1��7��*Y4���Gz<��Vy��hOWg�h3��H��O���g���k��u��-�>j��Ѝ>�1�76����Éy�$VO�Tm���}�^�!����t_���Lg���"������9~���D�A�7�UMR��T{��lbl���%^�'2L�PZ��������ş��a�"-��'bЏ���P��X�m��MƔ����5���l�&L G��5�b�tbL�R�-���hj
'��P���[�s��!�f�кX�����~���4hCL�go�B���׍���L�"C��˸Y BRhrGce2)���<��9_����2J��lZQ��"ƍ0vշ.V=����fv�n�׵���l��q 1��	�C���V�]��	�QXi�3X)6�d�{+7�0���Ջ�E�%�������ޒ_���zl��ѮC.af�M�:�<L�i+��0�a !�RI�����Nߜ�
����"@�^�-�$G��409<�72_�U��z |5�C�?d�=u�WX�,u��	��xR�]�po��#���sO%�4���x��ɺ�_o�~�s�r::�6sXSs�f^�;�u>ʨ���E`&��f)�#����I7��Z)T�{_�����&4��9>v�H�j&}�����6�[|���;�Q� U�G���ۛ2̈́�6|��<�����5��&m$�E5d��0c�+b��
�.&�2�pS Y#P^�苘Y>�Jɍ �:��%�n@f����P�Q[�R�m����wR{f���o ]���ѯ�X\ٝ�Fֳ�Ҫ���q��x�uf��2J��U8� '����9��&k���M�ڙ#Tb�bw��H
iE��l�Gd����(Q[ޝ�����K�MHFB��ׅ��1㊽��������(a" ;w���E��t���h���P�a�n-7�O3��>�S���{�F�+~�[�~��3�d ���N+���h�Pu���ސ jq��<9)��r�<>daw �+[p}�Bk��S��{�b^J �(�[oM��A5�o��}��=��Z@�e
di3��!x�-!��lޥ��zrKx�'�'j�o*2���s�q]���&)���i=�Q�4& ���Q�˕o����gGV�xn����%r�Y#R�ã�� ��
t0iK>�d|�B��P\��ބO�p>�T�@';Q����9��,�.�d���l��G�����j�*Yu�va1GI( �8���<и.9r7�޸��"�$�Qݼ��4�ڷ��"��4�����gԮ_9V�f��F1Ld
�3Ĝ|7���\�
�F��܎_�He��ch&�f����8*Lm��6
H���������D���E�LIɓJh�t������l���dD
G�،�������1ѿȱ�>�=~p�w�6�K�$�KÓ��B����W�,fB����6��鶇��WJ'��q$�r�(j�͢ ��7&��0��<��7c���<�*���������,���`�V ��	�v򓹢+�mK%(��S�δ�<P�!�s��Lo���Q��9�� �y��$�da p?,��,C����/>��dq�h���J��;�U�{]=q&���E����{���;Mzu�㮈�о<��Pu��b�ޱ?>7�wIN�4c��-�-�H�^^M!G���h#�Z��v��.!��P1��~��!�	e|�b�hp���7�u�?8ƀ��~Ѻ����K��G�U�� �.[L��bqw0�@x�]o
~��i��3�͌_�|��e8S�|o�+�_��Ԙpa�_,p@D�=#(���3��Kv�4\.]���x$z=œw��/�~q�]�w3�#Y�0���f�\S62�]�p+~�n�2�R7@�ț���RU һ�Sc��J���rK��Ȯ7Ɏ
���R>�m��za������<^��-�-��<̴���4;k'��lC[�I��e�^}�W�����K�a��VV��&V�t��N�+�)��7���Qʕ=5��n��7�������c��oi�T?3?���8���i3���Q�W���:�E�&�D��r��r�y����I�La���۫��r�n-'�Qw)����$����;w��ƚ9���l�@��S}���CHC^�?Oc�#<I�F���KO�񈾡!����8���4I�ϿGP��eu�`�u������/S����#������jp��V��(��<7�͓�*�}��:��]�7˭�B�o׾u9�`��Ή���F?>|^p�Է�5����R-��%�~p^ݕ4Z3�֣	S�J�5O��B�Uu��d�F��f0�T]��Fax5�m��R�T�A�:�t�1-xl;+��{t�Z	�C�V�s��������G�$ݺ���
7�s��lV�~Ŕ/]�grjl�����a8��*=��n������%/���SR�y��y�~8�֧�t>p��f7]�]�
+��|�د���G`ÿ�q�Z�iBy�g�:� p�hx�^!Y��3��8����F�I����v����i3c��۹h
؍���ȝ�#�D��͇*6��]�!K=�?p�ᇠi����ʢ�xG�lD:��-~��L�/^�2s�T�l��g��#&��m�|B!i��%y���w��<'���m�?i-�����Z5��]�
w���Sqa�۲w)���-��f�1_:+gl�̌��|����Z�`o?�rE�H��No^ڬ�I�\(�T?�ָ��aQZ��=f�h�/��)� qqZJ�?����n�큁���j�7�}N[��Vܙiq+����6�0
�%�4'g�׳%64Oi�����(��Gow��H�v�Y{��xW�`wd�_�o���F��Y��{��&�k�O�`0	���V���HY-Kr���<ʉ��ޒ4���֗%��0����Ɏ5=q�>�*�̨�P����7�޿y��hK�l L��Z�Ԓ��r	�ͱ4~�������	��P��WQ1P��L�d�Cj%��<�4��W��ZN�m�˴�-�K��6;����V��8E�=O��m��*(ށ�>6��R�sjL��=��_ �|��p��v��*t�9��=oh:K�"� ����a�Ć�/8Ɔ����DE��fn�\��r�$�h���⩗@�| ��_O�@�:��A�%e��{�. ���9��QP�D���J���>Ŭ'c|�>S�@�_��`�Q�/y�i�����2�d[�x�1$n��l#�z�q����$�?b��_cH孎�`B��`]��
w���z�]��<h3Ȕ�T��@#n�LZLD��p���y���59V^9-
sy���1�W�xl� �W`ys����NC�g@1�4A���������u|���veALȡJ>t�HR�ӣ|�%Q�v��d7G�^1lő��f��=��ۂ��{�A*6��q�Τ�\c�$�ٟ�V���V�	���(�"ޟ_�4��|ҫU���	 *]��rM\�1�6^��>�a�8e����I@Al�ew�~���/�&�]
.�<������@/�z���D��0�)O���*��&$K�ٻ���t��A ��4P�A���Avw�W�˗i5o?og���q�f�æ����r���gF��Vg���;����J�>�0��O}�(���Qt���h��g��$�|��I��p��i�Q� �*�z�����DPA" `���Q����m��"9f��ǡ%I|�/�Z��*�"X=p}9RK�$ m�S�4��"�"�Dˀ;is�5��i����$�!�z�U����dY`�����?��3ƁMP�#���*N��D�������~���Jf�^7�=:���Ӝ�\%B�jO,��w��9��e����-���S}�^��aҝ�?��W �3�Fhy�ɚ��>�j�^�n�O�F�^d��z�z"�������u(��8�)D�vlm���$��K����Ij�x��E�8���V8;�3F�G$����t�a�c��9��C��v�z�	�'���l�qbWF,+���z(��<��§u��$��yq'�A����/��Ϻ?i�gCZjc�Jǰ��"T11͑8���c��s�.a��Wf��	�J�e�.�W$�L�1��)'�]Q�?2X���i�Wт�}�u�:���$��M4��G�,Ef<C�S~"%����M�j���Xs$�݄���{���~,����o��[H�a�
D8�ؑ��OVRd�F�4�ٯ�n��:�`{�J0r�m����,�*�p����9��t�g�P( g(��d*H����̂ٙ�ג<VEܣA�!�z���dpXU��vQ`��N8�=4 ��~g/���V� �6��R`���C.&t�Z����HP�6I���w�r�����'�����CL����@�)�����$ߔ%e�<|��Y{ڛ{���~U�ӕ�m��r.� t
p�D��%Յ {<��/p���o�@�?/ �\��Sܵn���1c!�tg��y��)|+�鐸$ ����������l=X�*����(a��J�C�x�S���}�ă�2�YܬV�W�՞o�
��
��5\]�r���X��V�p��N�/�<����~�UX�6a|N����i�MEf!;��A���$%+���(���UH8�PR*���uM�=l@��r��J�L�S:���8���<����R9,e��<���,�(BX^TE��;D�g�x�"�f����ɚ�e�ݽ��\o�p~�@��m��p�>�~㒅G���>X0C��F39����{)l@a+?(���!�C(�k��1e1r��[���TDz��)k@��叔+�ٜ���#1S������ڀJm��H�`h�������a\�+�7��Ib�x��K\��	��z�� V_nέ&c����2��$o&��Ob<M�?k���%�d1�F����E�J���P(��@+F\��5�'r��~�%�%؛�����+$'~)b��Bw :�3�c�&w��tB���� ��!�U��#Lj��F�r���2�(�@l�[L^
s��a_���q��;�ϖO���Q�6wg��N��[���U�N��f�;�ԕh�Qk�n���R˟���D��l�f�>�4�'��!k����^̾�ռ�J?=�q��-�e�]75g%2F9F�lu.�����Y�w򼞺	T������	Xٛ�� E�����dq�q>�R�w�-i���^q�&��~�CCw�1��/X�9�ky� �3��q��)פ�a�m`&T�@�+�/"yȏ�"��Z���Bܨ]1\�����g��ǩ���E�3�	Wt�{�\$�@�]��5K����wG������|��x�$G���U�U|�mG��M�þ2@mD A���1 �=ʕ�i�h͍��o¡gT�U����A�=��3����\b�]����ǓW����[�������*ӧ7�F��[x��$���K�>�_���>h�j�C-��"|v~ǝSs�ߞ��Ďl�N���G>�\��U���Qk�MНrgc!KӀ���sC!CA��1�bB^��[����b��RKc�^i�[Ѕ .��	�zc����MH;b�������l�/�L�ί		W�y�ތ��%^e
���>�$x�{d��`��~U�=�]��x'�z�.c�e��;`���{��H�I$���z��5cL7v+\��,����HL8���g��ڝ���F�ɱ�[���8r2�����s�ׂm�R�v�$��w�&�һ��e��-���h2ڍ��B*u��H�y(<����K/QgW���)4��;��>�3?�$��:�@��a��!������Pz��Lui��Ų��<��A���d����Q�e�Wb��;�M�{����z��J{��{䵲�\���h��
���t]q1��0�=�<�-��?An	~��C̊�L��6����/u��.��~�`8w����U��uӺR2��y�´;��X�S�4&,�ҳ��;�{�xѶ��l�����S�����Ҵ��N������K�l���.����H�+��L�P���8�����:�7Wki����sf#r%�M8X:=3���l2��=�I'uSq��X�:j��5[�s��f�~���?J��씜]ޅG����_�*�Kh�3$:ОSbD ՚蛫���N���k�yI�.
~�̠M�U_?��S���Mlͳk�p��l�g4vXޖx����d���3Z]��꒡QJ���8���8�#�OFL�ӓ,��LLn��)U�����wQ|ة���a/��Re�������f�O���a���$��S��o'�>�'�fGda���2L�v��愕^�m� ����R��=x���0�t8�c�J�)2�Պ�O���(1O����l]ɖ@I�-[�>djĚ�	Dc@J�@��B��C�0���բ,��J�
��w����̃c+�NW�����B_f߉wrꆊH)ړ���t�Z"ץR�ؽ�u��{w�\4��q�,$Lox�0p����m�ec����Q�`�X�0�-l����qP�/��xp�0��ıX�O�=u�|�?[rR0�ߵH(M��މI��<��7wL�+}�o o�T�Ue>�hx��Ї������D�yїщ����kw˓��T�63e���������ry\9Ĩa<�����K�^'zsQH�Aux����&���I��$��y$�j�M�wmZWL'8�|V��!�+;ͦ�������C9dlRU��&SV6�j�ֆ�6�~/�F<�'i�%W�u�P�(�!���,�8wFܭ��?��ĥ�&弌ROW
���SH�盽�w���Ľ�Gs(H��N�GF�=�F��d���f�.~sT��?(l�������/�G�A�%t�\?�7oϷ����3� ���7mq���θ�g,u#��V?Ā�x�'h��˽v[��/M�.f�����{��>�4S��u��,Шb��"� 'c���k��"���Ym#Q��-E�K��d�P�cH%_�q�ح���ذ��8r��;�-����L33���*��@m�r�%��y�C����0�6��O�w��J�_��A��8)�e��Tw�b��ě0*�d(��5}�ƞǸTp��)��Yg�=�PD���v�hO��C�w蹙�����'��c'hY0%/z@���	όm;��G�S	��tځE��X��Ŀo�Vm�h��	�	�K3���oT27(�^X�x���z���/xJg��D(j99�BE�p��W�CYa���ڐQ�z�߱k�be�L���p��EBl�����t���@�)�}�	?�JI�iw���_uY��ZF���0K.@<����(���
�0�?���7��O����w7����Hp�)�8��j����-��N�9||?�N0 ���͝x6�3�F?"P��H��B�J(%�@3���YG��W��DK�.ݱ���0K����^ ���-��m��,�~�f!SI�~(�#���ThҾL����2���4:`p�gڴ�
%�qy�ĝ���?��:��0����Gx8���V�aқOAH��cH?��A<��� Ba=H�k>��}����<zp]+J��� D�s�H�Lxz�Ŀ�U?���:�Đc=uf��L�%��c���C��5�Pr�T���l��ˤ�]U8���������6���;�o�t
j�2)�Ⱦ��%~"�6[�>�Jb�Nw��az]?U6g�Y*ɀo���{���9������Qj��\�g���QU�(�xV�8J�d�����&O�KT��˥�@�d�|9�d%=h�������?��5��*��w�wk�z���k'����?F��t�-�> �cpւY�lv��C��Mw �Ѓ���M!�kS��=55Fb�Gt��#y.��c�,.�Q��y���x%B/#�A���9f��k�Kjh�$��y�����#Z�X��Z$^ 6(��pGup���{�?�����<�
�F��Hm�����~�T#w;-hc���kx�'�������"���km!^;
���_�3Í�]����0 �<�ϰ?N�WDJK�d���d�!W���&�?�6W|�2���a�U5mC ��%��$��lO
x?�i�o��p�h�D��Pc�����/� ��E���і�k�F��$)�H�PC}`�:�6�9C���y�#�|���lZ�@3s�yg"�b���'��FTX��:.f�LH
��ų�� ����y�X��d���Y>�,��Is'�ƹ��/��N���b8�na�j��eJ�z;%�Hs ��	���!aO�!������
���n�����i�U޲�"mҸgk`�ڮjP������F�1gcRdنx�5�eSLu��s���#+�u�5H����\�VB���!J2�}���|�{��|շ����)�H����7�s���[�Gs͓�+{j���Âa��^�B&�j�'mx�'.*M��<M���Q©��K��_)PQޱ"��>��?�*^p���F�ɾ�-٪�5�SU�믔iH(Xk��J�Ёq��o"���&]A]�Z~Yy&�_^s[q�ꌷ��ᶕC�,Zgg����Hͯ���
����&5�l�����O�u�Ϳ��Y�&�5�Xez���x�F�w"�L(��D�Q�k��5oLƅ8݊P��u�Mn����6~�����Sr��57p��S�Rb��_��n?��J��!+�:����k�Ob(��9��C��GWmf��6��p5���F"��)�o��{櫑�0��'vb��
����Y`'i�ȧ�>"%c԰������H_v2�?!+L�ao3�z���Xp��}:X�ao�O�-������6��M�����µJ�?�Cv���a
L�y��ؗ��s.�f����̉:�h��Ǿ|��rO�L'ɽj�5���$0�cQKi�m��憭�޾�<�M9w�-�$%��Rq�=|H�R�����C<�
�*�q֣F���Mͻh�lr�&?L�\�����YК%�����5B�i��[1m��걮��x8�\��!_v����G����fc��6�o52M�2�:E"����>��/e���# ���!gY���vP�t���pi
��B�t��*���fP�Ё�U`E�p�[�RmJ�ֵ�?ãރ��*9ת�2E���`  ���S� �� �$U+�Ԓ�r�G?7�^ᗔ�U��O�!�}�՞o�{�,L�	��!���ev�;�<X���7~!�Ifo�uC������ X�N�2����s7��ˤy�GY�L�y?n��Ȝ+�6���:P�/��#�g <]&��4Q9�E8�V��7E��m%���ac��jEM*/�&��c�J'�[j��N�v��H��dv"��)G)�>�J�4����J~k��E��/�V����V����M���ŏ)���~�γ�
9��Z��ۧ�O��Ǎ
$�i9D���nV���~{}�kG�,��o1k� �	�;�8/����#���7��N~w�	�D%�L$�G�rT���,�4�'�l9��+u���T�*mBE�sD�Fv�LKO~��&�%�x{�׉NKd��$-���#�@�M�ß�E<(���3���_�ձ݅�����,V��	�K#�1lt���$k����>kA�9�N�e`^SV*C���9�d;�c�$�"�'��Pj����{g�X�ѵ �� ���M����)*��m�Y5.��0��a'3F�-1iV�����}��Ói��h�~Zh�u��S��V�ò���M�o��˓I��Z����i�D�]|�(3�1�@���ba��'�כ��J$����+�C�2G�j*�����a�q�VGc�{KuM�[�v�w	�P���Bw�b+�l	��a�-�j��&zrj�0��t-u1Tz'}�l"����?If�u����j,G3u��H!:!e�f��p:���Օ�QNL�XfG� ������	WF�-Ս���6�4���t����,H��z�F;M�u�����-�s�h��|�~�ܴ�X��X�����]��E�=t#�Q�ʡ��+�$r�]-��H��� �}�]8n��?����^�8�+�3���z��+
�+�n�^ݠ�~���n��yr���6�RfY˘,L�g��;��/MoT��d{A�6����\h�L��O��i�+�m��R�U�{e{�3�]�Q@Dx���-�&}��<�[�PF�;���$k�<1�=���Z}k�eh�'.0��a3��i*�X�X�uʹq�Fy�@������QG�-�>��\-�.�'��uV�_�
��Oo�K�=�|d��,8��=M�"̴uG0?2��;-^Κy?'$�G��#��m���H�$�}��$Űn�.���9B���k�Zd��b���qD�?��B?*�&���������B��tT�q+*D'��w�)�?�I�cc@�q�v�Z	L�<D���B�ҩ�;��+ |hӟ�\#���C�R�J*��v{�P��v�5W��޼.��g�f�	� �7J�[މ1I+i2���&63@P-���#����,Ĺ]���	*�� eBIV��4q�3H^(wX��f���2$�e�9v�VԒ	W����PSo�w�ؗ�T�}�P[�5�����GF�/)��9������
��n�]�k@���k�s$���U�-�<e�\���)��0��W�_���uFFD�x�U�g�wY<W^_���C�br��N�f4�Ve��x��b5Д*��M_��+�>D�r�(�I��V|���@P��14��1�^�Q?O��r��Ì:9K���5B�yH��׀=R��)�s?���I�Wiб	#��Ai��ё\�G�=5�A�l�( �>�����i���,ކR�i�e�	S<�V��<"����Q��9���r? �������sͶ(򬝝f<�VEU�K�W����6twHsOQ�iF����}~Я'w͓�(�.����Z�doF��$�T��*�X�ž˒�ݩ�.�0p�D"R]PD���G���/��(%~�Ц�\�p#a-����y(��%�	����F*���s��ou1�"�$�V˄n��'�lFn5y�u`k��k|�SBv84��(C�F��Zӹ���m:�d�P?�_��" S�s!N�U٘�Yh�K�+�]���r<����ك���#���9�=wB���e��.�~��`Uws��80�Ds��cX3�✮�r����*Wz�K� 	�߳������jW��t.�Dbh\Lo�}UO��y<�5�%N̈���w���T��w��c��Y1)����vZ�o�Ô(c�m/���2�'��1�Ğ3��eü��+	NP7#�w�Yϣ�WI��vQ��vZeh�?�"b4���W�Y��\��gX�b�xb��44L@f��PI$%�7�ǟ#fU�� ��Zq���������|�i����bRg^��i�4>��	�:�[�`E�i��ó
%z���ަRk18��4*����xg<��a�����M��{ǾCq)UO�eM�Xptr��z�n;��qQG��-����z�^��G��~�TA�P�VJ`��3xm&e�{�=�"�������-����l���v�g�ږ?������?���! �2/`ŗ`[S-��0×��;#ZG�c2�2!�`td�0W��[A�ǿ���������A�}>��ي����@�����*#��t@8��J���� 0i�M�Z��@J6cP�a��Ǩpf�b��
�����8�,�6��	���pEs�J�1ftj�.�N�~#�{zD�U�w/�Yt+��$~���.��p������R�ͥ� u1��;���#7e6�Q�!�@ma�J�6wo�F�P�E���Ep�tIJB�U�l^O�x�Wq_��w�� X4�����\�q	�Ͼ��#�>g�M[���^A.�$'���}�m[�2����^��[,y&X_Us���i�)2���N�A�+��'�7�"�6##gS�&��������u�vBד�XM��e��l���o� f�V��_���D$�)s~���� ���ئ�7�M:~U9=b�Ó��` f�ū�P	{ͳ�}K��̰�_��;'T�n+(�a9������^NR�����+z-&t�c�}"�P�^++�0�$�������!�::�9�
�a��I۔�[����LPA�kZ����ޒ0��H�k��1t�qP9��%����Z�=$Y�F)�9��hd��j]D}B��cc�Nxm"O�]0No0��ѥQM���^O�#����o�~Hf�c��4�`ʚ���C�s�dv���
8��ؽߪ~�
�?^��W�δ�*���fc��=`W5ϯ��m�	a\%���(k��0YT�)�)�͏-�TSԖ����S,qb3�hN��GQ��i��C�:˳������ʍx���8��Y8إ�>�kcT����lP�o'V��qL���!	�F)$>x����
�u�}pι?tq�ޝZe�I+��]W�;���2G�9�M�'OX�	
�S0��W�_
��!N���+����1lɉT��	{\'�0�%�5S���z�:i(��k��5u�����L���p6ɓ�����Îf�5�T��U����\Y��)�[G~�l��b�{MGl@^"���-k�'QSq�t��	o��C����xs���2�"�ꂑw�/��&��%��Js�d��չ�)b�]_m��پ!}��ify���qh���l��V���*��������x'���pů\z7B���8�1 ���%y��ww^�.��^�n�����+����R�*U�]���_�Y�T����<K0�]��=�&�}�fI'���r_��V��m�kin�!J� Ƈ�چ 0t�<���*�]I��%��=Ep���MCPGM7��1cޙA�gO�Qe��8��bdѸ����a���sYw�ֆ-u���u9����f�zA��	�({qlW�Tȋ(�f��o��=}����y��/-���:t��=[�mN�:�Bs��<죦>y�R��lr5�7K����j���'���݊}qȮ��Bקv;�48f��`t��ˆJ�At�W�C��U_�<a�z�
4U���KRs��@���9���^c�ӭQ���tD��K��*e��<S3�GG�r�U�Щł��/r*@آ�@d��A����pC��E@�wJ��$pJ(�ї�Bv)���q�ʣ|l�Q�zw��o�����72��C��ֲ�G
�i�i7Z ��T�)��g��BZ�r�[���(�B���t�a�Z���te^0/6(e��}dwt��ߑ��/*G2s���I�� ��إ�o~$z�b��;����&fTsi4ЫK�tIy"�Uc�ݭ~�qu��0C����׺���h_Jw�&\KN�`����*�Ʈ_�`�\�m�K5���?むӾ�T3�yG��V�ӦfL���^��.�P$M�#"GlFn�z"\L���������g1��.�ה��ˀG�T�ߒ����4m%ؗ�� p <A�i�c�QОCuQ��e&5e`�PN.P��n1�7�{[$S�)�=�,^����XIC��E�G����1}C��D�?VT����o-�ۥ�t�M��F�W��憈A�{�f�t!����_L�����'�f%ʎFS�²q���׽:A�X�����^p�8�T���T�ӹ��ъc�)��c���%L:�'%�A�o5S�p%s�|��F8`����ΆS{���J�!�ڥf�#f���tAV��h��+���Sߜ�����cMO�k*�h�&�iJX�qy�V��;]�z�EZ�y���A2��L���B����].�}�����`�s�-���9�a.*�ޗ��P!��
�a����Mm��E���Ѕ��O�檩We�ji��z�p�t��!��cb��#�|,����U4(G�΄�����4�����½'"�^���a�! T�%���g�3��7�'� -����$)!:�4ۛ:���%p��_(9 ���s���� s(_Dd���T�9��*�7�*Q�@��n�8��5|I���+%F>dՈR�_�O���ː�f+����kNؔ:�uEHsU
o��T��R�a�]d�4�eP�t(��+	j2��8�`�/~z(:`��s!��sT���df��fj}#�^{K}�0a�x��]�gk��vD{�.�����b
{���w_]�igG�o[ !F�pL��M6ۧ�;��*�C�� �8Np=^�	Ҭ�4��q�EO�� ��b�C�=�2�w��JS�[7B�͋
z� ���x��T��\n��$u���?^�����Z͖�����m�8�S�ޭ��ŕ��a��҅i�]OE6�=�O���xܟ��.x]�qm�+@װQ�la���rCc�vQZ�Ͼ��|�j@���tK�gS�t�+���P���"�^��b����8���Bx�#\����;l��#�\���̀�Nf��ZU硎�i���~h˺�q�n`J��|Y��iѹ��+�.{�G%��ي��O�jo(�Qf\]���!�^ݦj�*���`�VK���!�6�=������"��~؝S�MO�Q�Ԥ���NO�ЗNt�`�Z�slO�&����t*\%(/��y��K:L-���UF�Sr�7���<�(����.��0��FQEG$�*�������E�)���kf��}�?y�����
=��{z�V$=ɁO�D�n�]���O&������-^�z�������Jt<��T�|�d�O�F�`�h�8����t�Y+��ى�8^�H��oO�0�|? 2`�-'����p*��^%m;�_eU��j�ŗ���n��~��"DH���0R�N+��<�=k���v�/k1��<�'p��X���8�&�%�����J���X�z�+	��yo޼�e��3>���+����������͸��zi(�fa��C�'e'�)X�����棧O�V���������Uk�`y�\$ ��i�Z%�M�!��飑ֲ���<���{j�Y1���Fj���<��h�q��Q������E �)=�f��uc��L�Ot���SeJHy�p�����ݍ8�#=���F�jc{̮����J'^3RS�-�;��U���󹢞	��X�n��N���ШN��+�v��\�S�/��zw��ITf�M����r���h��Ӊ	�Ƒ�4`L/��@�
�"pA�c�V���h�*p�{|Q�|P��Z�K��!=��n{�L����΢���@	��n�4Jw�+�f�b?�bE~�O���d��P������Z��
���	dk��/o�0= ����5�O��Z�w�V%{��5��}�1?��f���2K��u`�H�cK�?g��s��%���e��[����["��4nG��S���@�{�,},�$�b1t8L�m5���o`�F�Hu�-&�H�7��K���ذ���bl IQ�~L�'�Pjz���O�Q��������8A���.��V��˗L���t��ݯB�>ԐSp�9�R�e/<c�S�x�O�L�[G��]�K��H�+ϰ� �Ң=f�k�
��!4�Q!��f����H� ��%1��"��B�ۈ8-;/����	�wX�*�$ƌ�䝂���W�`-R�������Yp��)��@_T��CFϚj5��$m1�"��O�_�G<�*�C8�� ��Ro���R;@����2(iu�0���|��pa��#�s���3+o�8�8���@�r�?{������P���cV:��.�L1?������<����2.�r��E���	���!�xͣ5^�Q�c��F�m����(f�m@�o$�CU��t���F��6\b�П���B���҅��1����J��~Z�4)�[��#F�������`�F�N�J��W_m�jK��yS�pZti; !K�� �<|�?�0�������r3�iPZg@���*�� %�^���f>+��s�jM�y���E����d��lZ�p��v��*�K���?"۔�-�q|[b3�Tmr�S�=�q��N>{�Oh�~��Yz:͆S$�2�	jƍ��HO�Ʈ��Ew>1׮8e@��Nr{�'�+ͥ:*���@-��wS�gh.{
Q�}��ڈ�g-�Iߵ��u�"S]���D�+�o�D֣Ý���P(����&�K��kt'�����I��ߏ�����lj
.'�/��/}�S<�R�}e@��)[�L<�Ah���tf�� ].m����m�i�N���@#���Zⳬ�/�"�"��\&V̕y�8�5H`	f�&��q�|,}�!��!M-Ai*�v:?K8�5���M��ʸK��6���4�RyyW�&���Iѳz�;����	:�I- JA�Z��0�S��N�TydEs.�D��%`��K�22b�HUT���ՔӁ��y��W�v�\��t��*��o���|s�BRq57�<xҵB,!���?����a(���:TMA�Y�q�6%bc}���O5_�����;�<��9
�i���#f����b���f��5��ڰ�h�E�=4}9��pgi��̫��!��	�Tk�i`�)����+�éiK[w�Ao�9���%��oNeJ��s�O�b���҄ޢ9zu��??Z?���½��*B��W�՞��9%-ț}u��
fY�+��%(����`v����=�8�`=��ȋ]^����eW"��)<<`��V�z�gtm�����	FVt	Yn��.rӓ�{�b�������q^�|�PXdb��D�Q �-	��O��d�b��{ḣ5���6@B�ީ/��l��yj$aÈ��<~���M#��>C;P���~��Dr�)O�#i�+�f<�T$%���:�0���0n�w�'"�*�AS%�(Y���ۛ�b����С �J�ޥ]��T����'���S�� �1��|���^�����O��y�Մo�|ΰ�,T��G��=�e��-F!�n%[B�2���`��zȉ@��'�G�:�y���8g~u�He��K���r����د�l���^�T�K�?�'@��y��]�A޻�KU7�)��[�Jc oY���I�^G��8����Cr*9�8v�Y-�B,�˝��u$�v������U����q�/�N=��o�?�b���8�<cY�Z�k�2�b8Xq������.n�"c�tm)RC|"t!sܲ�qQ�n��颽�V�����l,tlh�JԒ.�?����h��L������~��=���2�v���k_wLS�t%G<e��]l�$V�w��Gi|-�K��)��4�aD"��fq�g-B����jO?!F���������q���U�㔟k�����I������|�>���P>��faZ7u�qP�g&!�C6�/�Z��LU�X�Bw�d�f5���M�Sl޿%�<)���W���ޚ΀��"�F��~�鐫�x������/�^�����L��W��Ng꺮|�N��^�W-�G��-�"�Ȅ 2�2r�jM���|~-Xꉇn*Q��aV2����vl�� }|k�uz��az�5�O��������Z���4`稸���㙣nE�N5*����4x]3�(h����_t�$���)��C�k�9\T͏��f~)��8cbn-IC�R}�u���<?�4��(��(�os9�1������ʿ6��wb�+'���r��G�&��*S�A�y���oq�/��\*e��n$R���? 	�0����@4>��If��螣�:� X��	���3�sؿ���E�OvXz̡�����X�6�gQ(�ݦ�����;�sX�x8;��}>�E�pS��J�=�à�{	E��QMw(|5d`Gp�����L�
����	�E����x��!<����Sr�fi��QmħZZ홤@{J_.rqY@t\�����h��J��ng0GA``� *�I�p?2�Ϭ����M���zɘ�52}Ylu�f��6�
����}�����ʞ�v%"�Hc8z�GV�ya���[��13!�˜g�<���������7����H��9|�>0���[�0^��jU#�Q��D�pՐykd ��t$i#׉����l����}9��W~;*}Ȋ8�>�/���:�˩�(�r�{�}cy��^5��z�Zmjtۿ��nk�n�I���>."�$p�1��>�m��.���O�8��8zqYX�y�
���i�jÞKɮ��i.��򄽬JM, Y��������/?�~��┬-r'�_!�g���y�r��Q�`'��k^+�<0�2��RCkD�z�d]��E뉑�$n.,ǆG�YXH� #w+/N��Q���I�dQQ_��{��Nf��_R���Y�j�ݒh?	_pg�� ����$�L�a�H��f���쨛���Ʀv�Yϓ�������*��Q����G���.}���㼎¦��3����G�a�S��Pz�;��T��ɍ�J!�f���*j�\^N�<���<��ſ��΍&0��봤�3��f��[���]A��=��{�Ǘ��1�i�k��	Zh�4�4�9����� �ӟEF�R�`����,����'���c��'���L�wWؿ@Llڕ��t�+�	B�3xw*="�xV��aMb���an�!�:f��j����MѨ�:Uo<H�+���ɖ.�g���bZ��(�����^#������V������y��b/�&O���d$�
���MԜ���O�F6�K̛.�@��K��ϸV&5k>�$�y#�Y����R7�������S�d��1I����B����S��/�i�A-t@�d��W����w��$�CҽM:�^��v�!��.��[�{���ږ_ǻ�V���}�}��FZ��>������E���#�-[�E������F%:]_�֠)1���=gd�/*\0��n����͖�)u/��_�7�B@�
l$Eɒ�C�az3�^���?	H��H����Y��g��?��u�6�i
80�O��� �� ���x�,z;RakC2[8y�a����[�L���v]DN�v�W_�c��K��CC| �!H���I�A��_#d" χ<�ȧ�<��6��֯'�����w��"��S���-=����i��0Bn�E�؃:U�F<�W�,���SN��|X���V��E�(�J��܅�%��,��|�ĉ5ﾥ�Dܵ
�gҒ(Mk�������{�F� ����N�����ݤ���
��M$Ml)j� ���VӝV��v~�uh��5���� ��֠��
�{��}�)��~D*Tΰ}�?K�?�u	7�r��?i�`�E���Ix�s�09����R@9��=�1|@3�җ�"�qc���\}�	 ��1��㙭���E"Y�G��6Z�A1�d,�|�̐&��4���y1�!��E� �v[p>K�+��BUC)�ss�|�$kĄ2	�)��'+,ZB��tI-�Ua�M:J�����_c-gňP�$�ݒ~�����YxV�� �z0q���Ƒ �$l��uZSt��x�y����-}�;r���T�i v:V���X�ۑDe���j���'PϤ����Ha��m�=/¬H>u�.��jOz8L��mDj��׫(�9�B��cZS��J�T��J���?�u�jژ#7��z��z����G��w3�Y�6�Z]]~�dG�w�ht-�l�m����݈�2f��k�M=ϷBS`��I��6���9�P�ZH��`��01&�?�D�)����s_냼��L"��?�]���o21�ȡ�!�1�$�i��3up�h��)�J9����e����k�LOG�c;�~�ls�OΕT�)�Z9�
n��V�E;���S�yyk�� �]u�Xf��[�A���`G(�BBj�n����wC5�HX1����������pݶ�����>���}�(9:�N��nsb�h6���dj�9RpU��F<ķ�߈W�r� �
;2� ���>�TR6#{|o)8b٫������~ad�!n-ĺ��;�$�	%�*�}����S�g�c4p>�6s�ю$�B�/��d�/'>!�YE���o����5���%Ș���z���]_vi�1�F�5]��	�b�y|�
�1�c�����+�����{�]O*m��΋�a�=�%	��(/���mllw�V�[�ߤ���	g��b{q�����h��o�c;Ȼ`T��Z-�aiN�g��+|� �4ɗ��ց�塤j��X��o~az-n�AhA��bWp�8a#W�XD�t:r;�]9�y�R@JF��l$4�0r�Z�p�1������0\Z����i��G�G��d�H.g6��~��=�
pXP�*�h��C��<j(�֑�pCpl�`"�B9�sC>�ɩ�j��$Cr�g邭U�uט-����]�&?	��e��?�=��5�cBiߕ'��+)8�DG�:����a!��u��erQ����y�$�ʶ�i.��cٸ��a�P:*uE� R��S���<�D
�ΘyUDN�a��"S���f#�"4�}]�KfO{ ��o�9t #��ɉ��B���*��.m)x��S�X3J�n��3��C���i����ӷ�С֓bT+�Y��8Y���r�2k�)��
����zR҉7�p����C�����/b��DC�&]3?�8��aӣC���W3�̸j�#X�3�ğ=�+��=���jJ���s�h変	����x��O���z.�	�Q!9�B���<8�q�;�	�'�`�`��ȍU�ݫ�9-�9���U/�8��b�%��t���>��aTf�:����U���Ӓ��NN|1RyP}��O�}��VadrΐI�N������?��N�3�3�뱉�!��OI?Yؾ>7X5J�x������Luy�.��Zr��!����q�
��0uKFv�Y!}�貳�Z\&�v��Rk��jݦ��yp�J?������9�/Z"^�؍8AR�l����xn��A: s�[H7;>Dc��Zu)�LJ�Q8��3q�W�)��r����-���}�����J��ۂ[^ ���Y1�������f浡�E#��il�P ���pA�x"(�O
~�=�T�84ڒ��"$b%�т�#V�؍m���{�iw �Z�~6|E"��b.�8瀂�Cݰ?a��b���*�;�9�muV.^Ý�oԡa֚ά�_3q�ql��[�֕�Y8��t!79�4� ��#>x�}���umge�ӣ;�VaT$���x�}O�ѿϳl�Ŵ�d��@��I ��R�o�I�m@�u��!�W��CW�j�\���Ft���?v���'��fy-�gYz@�O���Að�Y�*c��=�ȑcW�rQWƓ
�R�\��%K@��e> 8QKǊ��)��ӓ@+Y�������K���A�_I��U��jd|����A������1����^6��ݬ�:xq��:ܨ/�&>I�]3K�b"������i�o�ȝ�؎�O`�{F�e����zI��������U����Ž�#i�|FD�)p�j!���otD����Sz&�����;;6|Y�X� ��J�F����b�O|� �U���������%�`���Asf�ł��I�E��U����X"D2�p��%�:��	e�S��D	��]w����Fp�0��j>j�Ӏ���&� �GS�z23��ݧYQ�Ǘ�_�����z^'ܸ�������y��p�n\�y?���ͪ�jT��;˽�e�4M+�w�H��p��]�Ɣ���mJ����=Ys��.���NVc��^|����ơJ�p��H��Otc��-��X)��yΪؼ�T+��뇄f�����Ѵb�K����������@ڋ�vv�o|��L�h�tR%���@�/��I ��7��j�S�X#���&��aQ|y��@��L��s�`QED$�<�,XG;@��Y�u�jԷ�9k���!~{��3<��3���Ηv D�rPTF{���.I��Y�jr�W�x*�*��)f2��れC��\_�R�y���9���J���QGe��6�9,m��U�4^�AÛ����1q�,Z�E�xu}.��Y<��%䉁[�%%լ�<�Z}M����57Bru� �)h��6؇�:���S�u*3ːw��8bF�&�CA��,�R�	��.ɍN�;S4=� 5(�	I�����@Iy_3aD����)3��+s�!X�����u4�����cѨӒ����
l	����Jd��N�Hs�᣷:�gl��9�X��`���M{v6F�G~��I
���p����Ҥ�S��GY���&���	�hc�Xs�c�T���&ǎ��L�$��(鮄DC��#I8t-
�ط�q�����Z�FS�4x��(�n-Ғ�է�m���1��7!��z$|N�ȏ�C����/y��Ta�� ��wF�t���e�d�f���'�@
6��L�E�a/�h�V�����K���鑌jz>�6����`�t��,��C��7�Q�ˍQ����|�0���⩓�8Y�q�2I-5�0���Q�Ȑ���Xu�u�D��f�.�zN1'_��;3��	���, m���8K���$W��~ZP��3��q�B��@�ٜChcuR��1�A���.��ܾ��H�Okb�g�=K�;���%r�ܝZ
���ځ�_��vLx�D�������b�VǠV���L�^�Q��t��*��X��x��"(�T����1f�2��%����1*�{�zO�ܐ��/���,'�}=�i�,&u!�_%��1��/Ʌ"j/hz�=�Z\k2���ѽVl]e׋ �j���ay4��H].���3ޖ<�%4m��y��8+�<z̘�,�Yi_7�Ȼ�{n�&�2���|���J�	9ag�/�	�� $���@R���D���n���a���<l�j5h@����1�JO<ފ<P��-r:�yo��2
�N8d��-ǑK&R��?�Ҡ& Z���]�VF�2鶯šVW��[9/�VQ�>d.��2§���+轟�>V���Wh�^]bcb;�$ƴ�\؅[[����k��iS�|�b��RT���|q�6(Q{'U����ݦ��"�HK�UV��:י��7{P=Y�ʄ�Y�Wu8� `-%|��0�:VT��ru��I�cq����xB�d�VY<��������k���w�S,Z�a��vܣp?'}s7~��t6�~�T��&�ˇ_���컝�M9�� ��m����h�F��
�J� Z��/�
�ɇ?���U���H��� ��qM<�/���K/QBv��+w�f���V����G��o /��sE�˥m�P,����:��r��Ն�Rā�~��-��>�?�G�B��ez������r�0�P���ƌvZP�m�pԠ�8�3`���4��]�IP��A�Y6��|�g[��+���^H�}O�qE%���34W�Rk��MR.�i����� e��?�]��s�\1���C��\!�`��vOX�ͩ�_O��?S��v���+M�b8���k9��@��\R����*k�<~��NX���(5� S?L�#���$���ݘ�{������L����Z�)M�=���$�P/��u:����F���d��  ٭eG+-�zD�7��z�X��D	?�i�C8�6m�)��>��\4�߉㧻MP�h������@�#�������7)$�-�bˋQ�;M(l��;e4_G$L���Й/G�Ձ�):B��|�lA��ɥlȂ�!�����������ߩ�1ebQ�����/�J��eq_�4�F$??�h��#�m���b`)bf*��X��xa���q�O���eZf��s�LW�w&o:�n���z?�	���h~YwN~@��}@�"c�� P��+�._.<�3��>�D)l�>;I��(���P�c��sئ���l���&P�E�%�L�̎Ĺ����<��m#{�E�N)|�C��2kY���O��KMx�5����)�ϖ����/#D1��=�4~ǋ,x���8P�n�^�I��ǽ	b`��.Sg�}<@����ٗ�kP�o�����&��d�{�֯��^
>©>�*MW0=���b+b��V��E�az�^j�~~��������-l�ǧز��'t
[�뾽$�7`֛%�G���@Ѓu�J�(ג���H*[C��I��mǓ� �4�``�PC\��EF��	�@����X��dɫ�F�^���u���:3r&�˒� �-ы*�8����B)4!��[�L����j9BK��E�fӺkn*BH�4�&�� �EN��(�eI��3Éc���&#V�_��o}�<?���t��^����`%6�<p6����mß5��|6m�l���軻ϣm0�m[]�R�!��5�?�- cdč"���=�p#�[�T�R�#V*�c��$mi����ʫ�þg1�]�o���|6���4�;�{1��/#����B3-���Y�$e�lDn���>s����Z���֫�>T\�@�s���8�7
>D{���K�H���z�g�M�ow5m�`<�����P~{��ʋ�\�.���DR���#�4�z�%�`�D��./>�+b'��(�g�?����8m`�T���cѱ���S}0�c�	�'�V�,��]�d���2h�|�w�»�J�p�n����z�mf��q�>�����	j����ڿe��{9��)�����tg�^�}��nL$�$W���zUWR��&K�X�c���C�n���!qL��:���Ů,@D��j �`��[9"�����c"#��`��,(m"QU���0@��Whi!0�ˈ��Zh�?�T�������2������߱ʍ�ο���U5�Ӓ�4���a�˯�}C���4����B\�ޔ��1�t��7[��Zp��6�ц�ip��.�nΧ���K�;�����������hl�-7~�!E [*�K���j�|1�M�v�(�в�)��B�fn�����x����� ��0xjM绒(���W��Gu�}[�Co�u��W��S�L�$"��>$���-�YKӼ�/A�<��u'�:W�81���35q�mqB�Ww{��������yF�c��>������	�]r�	j�����|��N����5��f��TU�U�(�kDgI_/�n���>�UU~/����<D4thӠ��K�7$K �a\�����G�/��O(�۵�	F(U�z����`d+c_S>�k�_�	p�����d�N����Onج*�QMԴ�n�����%h�� �;pW���<���E,\~X#}�:���M��?�:��qI��'459�? hJ�B�%�����̵_۟��M��J�.i_�9��4�۴�emH���{�>H���J}����w,aĕcڠ�]��
~5r��N?	������E+$�3Y�����~�)��h4��Z��]�teP���0���H��>������~������FxLy�̈́ȌAQZF�<������,�����)h�@m��\��;)�jD�.&5��Q}�����V�ч�������
!�����'T�kd���L��B5B[���F��C��+%���;��R���)��`2�θ�ϛ��4G4�X�/��%z>���ێ���y�陚����9���F���BW^���LЄ�X�G�i�d�ۮ�K&/�JU"�@��}�1H̳/v\��6��d�*��)T[}m�_򩢱a���s�o����_U" ��l5J8W�7�;�d2�F��ͫ���&<}������,R���vvX�����RcX��`��'1yy�g��$�IP����>y��@�&�wb3���R�d�tޡ�g�p��"������p��e��%�����\���ow(�����or��C�v�`LB�@n������i��Ga"�k�������'��V�Ԉ5l��Л���ͮ�pl
z����w��6PK�pHf�s*���&�ň�wK����>��-����Q]cE�N��׳�S͹�%�]n�a~��{�����b���.txN�x�J0�G�~���@�X/ݡA���V���W2\�G�PGV��$����m����ii�b²��N��H_J�fI,��UQ�cB�q,u��5��������9�\���9(�,�$I&;->�w��3_깅��#����sUߧ�(<k�ޮ�6m[CL7F1��,��*��:� �7�^	3�f�?ś�=���*{���ڤ�4ƌ����gs_�s*��DG�n��7/J�4ep-)����WZc�=�EN���7��kVc�Eƽ9"F�[7�% �{�Z@�U��B�����X�}k	��K��UW�=AV��A��v�[���2�W�9����|�@Х������Ʈ�F�l?������q�WgqReᚋP;�$�G���A�2�>��� k�u	v�^!X*b�Ma�)���V�~d�o8(Cܰ���m!�6S�͟��&���D��d:s�}�Nmu~�e˰�zQ�F���E�ˣv�kDǰ�����
|3�\G��f���I$�D�ݭ�A�|@S`b�����ap�qq+�/�uK	-�u�|ڻ!�b��'	��R�{���vnO� ��*BF�Ǜ>���Φ��/�Ɵ)pR٘�;�[`s'��l���!%��q��Gф��x�e�/ f��7�� �n*:��bV�0�R�����S&�\��Y������nX��9�W嶾����a��U�7� )����	0x�>��s6ls�S�Cr��*l8�YE$G3���n�ѭ��zՖ�`��%/����r�=�cV��M�ؤ����XCJ��h�I㈿A�d�cb7��~{��Iy<�IZ���9q��������*�`�t�h�C�f5Ē�'��}x�v�2<�n�]/0�҄OBM�/#'e�'ۏ$iY�}��'�|�pN�
򤋥���^�����tm�X^���<���<�HV�6�d���^:]��-�[Ԣ�u(I�.���H{�v�]N(�B����u�Vm��k�#7|6��3�V��HU*ɦΌ�-��2s�c��v4��\v�Yq�ë��Y�K{��9и)å]� /���F�<�P�Q�TD�U�b!7��򯹿�� ��8MK��T�vږ:�Ӿ1�d���%(�C���~��nT���6�3�w��k�d&0�<�*^�)��ړ�q�x4��7����()9�E��yE�H��k��? �wK����!x�iHv+�~P��(�CtCױ�4O�Ǖ��*�U�.�:3VX9��Ȑ��nҜ'�Ø_��*3X�Ȥ%�!�|�o+�-h��N��w��t1��A���Gb����uY����7A��95�K�8�g���o�<�АO!F��b�F��U�ĜLW59����[u�%����6�_y�	�(�A82B��#p33�C_���a�
�������X�_>hV�N�I�!*��W�霾 �ʹ|��g��ϒz<�N��@ԣ��v<��oo@�(�����<}�����r�蛠��+(���m�?�w��|N�0�x[�ǚɾjsfS�����:p�*�^�}<H܅��v`�c���T(�<���n4�u�6U�����Y���{�lXF�@�����OQ�7�YDdZ�c�:���\9��4`/	T�����Z�M�"J�r6ũ�<NA�T�F�D_���+쳃�އ�uD�!%2M��NC� ����k)ή��MH�
�l]ls�1P<;KG�/p��j�	M�>G��x0�/�-�[YU[>=���U���^:�̝	�=���	���������^=������;Ma��TS�q>���.,��l��
���Hx�=�Ҫ��*����^�f���g������=ǐ�~:h~j�sG��)i�?coS�4�h.Ѧ��-�-�j��
��H�a�0��:y=6���CB�e��B���NT�<̯��KX*(=�P~$g͓>9-�T����
����<��̋4	k�&vU���[��d��C��E�H�	/]�=��y8(�$8�x_1�D�0���ij�>�\B�rr�[T�uC�u%���[���@@�Z���7Z���"�m$Ͱ`�,� ��jA>�����5)��,�ܦU������w����M����JB�r?dw_����+G��4=l.Q*�����hxP�YU��c��_��QmJ�w�8��e�T��0����K���P3���0/2=F�zņ1�����P���o2~�� �O�~�\�FP�q˫�y|Y�x�����r��C���8	�F���h��Jl�:�?X���In���<J���2p�Ĝ �n��a�P��g(�\�b�"7��G�A�Y��8��e�dSlm�autv='�(�9��H��W�=��x/�����r%l����ſ>m��W��&O��"�E�y���gmq����Z���i@b�.�n���MGd��|?�� ���#�	�7��^3��n��teo�P��F�%
g�I�1��Q
 n�{V���)co�?��U��}�	/�N96���_�Aoi0��!*�����5��{�C��eYw�&t.]wx�|�%e6�Ј��{'=����8�J�5
+����A�� ��6�W�d�0�#\,M�&ͬ�W�k?.?X� 4�`�Nڸ��{g���W�#����ӽ��<��'�J��{3���F7���2����i�y��pmǺ�i&�qc=��/}*�����v���`�O�P�FF�.o�m��{� ߮�'�ݸ�l'y2=Q��������K��	#N4�"�����q���Ko������,�ʥ ������� ��G�4Y�h��!�a:J���9P��z"����K��{�^%�4�?݄-�soyvU�I�r�W|���F��0�4k�n&1xฐ�����N"G�Ȉs�-�F�+�7#�.k+�;_�͹��G��я��y8�+]��F°K�FG~�HHPე��~�0蚇��_3N�C�\ ���Hl���jA�/�_*���(D��P��A���C���>���4̑�Ը���'�x�;C��2��(q�����{�7a���4�����dDb�~�aի��uK�3+7���J6���=�^�U	�"tϟ�8�&��������k�l�ٔѡ�&���5@Dek�Ri���N9X�wL�l0��,r�(>�#��Ɉ��]N��˰Hqˌ0[���¹&��>�:ʜ��\�&�X�'xA�=�l2��|9W�6�[7-Ǚm6��0y�g:��%"Rx����6���醐a�3�
��z|�g?lo�� f��,�	�1
��nPe�;<JK嗒����6Z���@�-�9�__��m���J��� S놉�P/5z�#|EU�O��i��
��ž� �Q��ad�"9�n�]�˷�|�7Pk�w��b�ȭׁc�%X��˦�+oJ�F��1��l��D�@w�	�O^��Vv�Q�/@�R��:�e�Y���&�)P06noV.Q~���1C������t��KSG�W�sX��W�S	W\L% o���Q"s�C��1����"T{��3�q�f��Bqn����!���a�Ζd��*�y��� ��$��7�]���9�T���m]+RP�$�M]e�p_���Nww�&��#}�Eeze
�dI�.���XMk3�}�iN�oI����o���oJ��Eס�sܒ�D�`���}��>�uu-�����L�{�E�L��D���vo-GD�����z�Ac?l����>����XƸ��G�H��@͚�ȅS����?=�����)�ԁ�L�G�����(	�~a��4��n�8/w��p"v��D���8h��1}K_��ʑ��F�cF/��KS�ri���n��,�
�Ն�FBb�w�=
 ]6[�5p������ݛC9a�j����+{L���z��QՌ't�iҴ0�`�+�w�!����&�D667��nB�����2�v��k��1ډ,~�ٹ&܎��_4�s��[-:�)��uu"�6�/��R�rO�6������4�w�R2	�%�Z	�`���1WV8qd�Xmͅ�m$o�>��ھ����RL�4W*�d`�j�%"3ҭxCC�R+:�뢓>�DGCT����':�@��3�-�=}�M���N��ƶj��:���ʧ�8�Rr�X0���;|�-qbJ`�s
���co�>9m*3����άc���1�z�ۛ��¹M)v[ �I���n@�H��,�| ��S�9���B����{FQ�D9*�sZ�5���3��$I����)o>�
���m�8�_3���� ��/<�l��ĝc�72��Sw=kY<��wX�S[����j-U�<���0�֍�i7�Rn�P�)g�LpW9(�����PS�L7�HM�̦��ׇ��%�t&H��Z��鿥{o��9p5�(a�Sw=�p6pUX8z[UY��?���R��y=U�NT��Qm�eyM�J�����z���}��F3z��SH@ۊgUӟQL�Y�@O��р��\fK�Q�W��.�*�p�~���ߨX���P-:���NS��ײ��P]i��OͿ^�#m��(O<kH���X;�_�	+k4�sW�B�D,?wglP�N"}�HN�.]X�����	��,����=!��c��Km�xl,$�X<�(O��2�zW~�����g�M /��������5HT/y��P�y�s���2�.��V#%`/0�ݑ
D�3�y���pӈjFٞ@=�V(���dE�������P�vrI'l��Q��ӅA#