��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1���e}ʲ��cg�t�ϙ�a�:�KR�%���ݧw���ȼ.����[��YR  Z�O�Fk�y
e�T�q}֭��c���ڒ��6�f	�:)`�={㨥�1����fǪB�!�ۖw�*Ƹ�!f�祒[~oJ ���g�-�:�ñ�(p��K�Pߞ�iJE'D�@"�k�W�=)fʎ���YD�$/�\f��ST��@M�R�1i,��%W`�����V�Xq���b�6T���o{��'�"V�*C����)�����n��C�X��Z`��p���Bf�t�8:̬	*]h3`ǌ���x5Nk�C��]� it��
wj�g]��o�Vt@ �6�#E7pz7릙܀��*�!ҬL������������l�6��h�� 7��0�$��N�7:�ϋ�)�A%WE�V�2����k��� �+y5S[��~/!���p7[3���*��x�V.�x���~V
.��R��&����H��&Ml}rČV�i��*-��+x��W���s][Y|I�4BM!.GD%�ީ<1�bn4�<L��&�a\Uj�w��PÊ_��@ p�@Ux�ADD"�~yB7$��ϸѝF�7�'�%J73x���L�W�}�b���6�g�C�x�q|����>i��U��Kȕ�u�Y��>�b�����x�T(��+f��\MJ���<�S���=3I�.E���L���U��zy"e�8���n���e�;�aEtJa�.��M�����Dy��A� �K���U��[�����LtGV퉁�R��%z�� �t��<6�ƈu�$�X�*����܆ɓ��t+`Ӎ*έ3��3,�3JH"������5f�l���ƶ���-Q̺�lh���M!���2az��TuF8��0]D*���L�{\A�!�Z���ބ��e��
���-^Y�?��8�������ٝP�a<u)-),���6���2����\I@k�x L�@p���>lw�`��qes��ݛ]hRRL{���%�l٩U�9�yP�_`y���Xwg~8�����^���}�\�W���V*v-o�ű'�}��0 )����T�� R���$��]����@�>v��,wy��Y}a�ݜ��{4���*����!���!�R^h��9�!P}%�ӻG�n�1?�C5�#�%�Y@~��E��#S6e�:T���"i�7���ܲ�T���k� ~��o�<G�0��F�� ��v6%2	�G����`o���X��*�ɃK
>��&�!���,�W���w�$*h6c��i�T#�_4����壹�dH�ꔢ���Kd�@� ��ke��<+S9��[7���b�?C�"|+�Q8Eڷ�9�rH�w���;`J�����K9����7�����h�C��Н�߆V<����p���1j���_;_�g�v��"���q��(��>�;�!��S���qb���lyN�U�BD�˂��n��r�(�l����[q/���k��m�,_V\��.Ի÷�LG(>B�A+6S�0��s@�1�3�R����N�w⃕_)RۍΚ-��0�e�o���C��(_�E�����ӎ��4���/Up�����K���9���\!(����tc�"W�Y�p���t�AE�9�*�]��U� ܞ��A�!�Z^B�[8ʤ��>��0��uQ�f���\�ֱ5PN��腓?�Z��z���o���tNy�r��)��M�vs[ŔѹU�%R��r��]���Wy G�2ez=�V�G��4�>
ӞtZ�b6�Sۖ���~r�_LN��S%h��Ds��Mv��+[/�^r*d���W���s =v\Pa��$O��A`�+��/�Zgb�	BT��e^�}�'KK-��5;0�c���ED��բ�Ȉ����Ȇ%�D.EFjSO8�e�E�M��AU�G��h�è6�nÖ�M�Z�����V�s��22j�d�?�}�f+xP��4oI��Z�}I3�1�}͟h����Nlս��� �;F1���O�f��	��V���vɏ�_��Q�a�r�3i"��L��M؜�������:�QU�e��\w��ї��ʖ��裱�Odm���q����+���^�O�+��A���h�,t�]� ����Ə��m|]��̻�#s�O[�����ޚ;��A�|�d������ڡ��Q��S6sN�=�B���4E��
ds��`K�D�Nc\9���]��d����+|!�"#�!�>�TK�rhw�]�n&�w�q�{����pTV���k0�MבJ���aȰ�5V��nx�����KNF��?�f���{����&��t0�1 ����*����O{��|���.�.DqONR$���Z��W;�1*u�@sMԳ�p_��F�8����eZ��τ.�6X����Cԍ�4ϲD�$ ���y�ΜC�y4D7�T�����+��MY4aI��g��o���lE=U�B#ׅ���������Y�!t��}@A<z�z�1�o�M�&"��IB�㲕VV�V8f��О�<!�&@���~,�La� �<?��}#m��d��a6�F\B:5*[�p!��M<8��W_R̆LO{���yB� �jEv��D��q�2��#2�r�Tj�2���穆�����fU�a䓽�����"�q0;��E k��>��/[̎$��;��9��	�{>�4@���wڄC5��M��pf򀧌�[�'3�W�J�<�J�m��4��9-O�^�ĥ? +�X��:��?��=�)rv���J�� �ԇ�0?Kf^o��Iޯ��_�]l3'�ସ�=�3�-L̴��������"�Ug?��G��'�R��ǖ��ݤ�Q%���(���܃���yG�FKo5�u�����#/���}�l�PDP�	5�@L,VoZ�n9)�Ȓy:���y �r�?e,(�"n(�3�W�ϔ�L��d��4ϭ�!�Q���%�
�66�5P�M�5�
8K,�x�K��:h���k|�2f�!F\�e�{ױ0E2V#Z5�k&wR��di,�ja�޶\#��|��H���q_�	P��=�1���P�ǲ�ጲpu���eX8y.;X�Q��-m h쾒g�2=���2a�Y�|��P1����.V�yU�y)A��ݡ�"#��G��';�=���R��Ñkm�l�� �iQ���&M���N�ϔEƺ
�g�`��k.uō��xo���*!��Y_���e]#�ι�z����	�&�޿Z����<�8\o]1g�)��/O�Qsㅎۈ}Ls3芓%m'@f���,	-���ؙ��ϴI�[�iYR�Ү����Z��K��	{��(�n��� ���N�x���֒;h���Vc4q&��d���a�%�2}5�mc�jV�Z�����С�:�,\Q��\��&E4��O`���2�'�V�����ѧ$�D�	�u�k�7�8K�VI�8��}$���J` T�L4�,���ٹ��U�m$m��'a؃a���^A�T�I+�aGOrE��E���8��\�Ǯ��Y�T���K�~nD��6�S���d��n�����J���0_gmE$�<b�؃Q7u�O�����1�ٹҜ���F9^KeGtQ��#�>�ף�P��u�O2���h�kS��gc�j}�gs �d)=��ݥt�k������O\ڐ:�7_��ˑ��p�f�P�>��Tj�����9 L�E��M��]L
�����<����$>��#��!\?Y��T�6�)o�~�~he�ΝN>aI�D0Di���;��n�S5�IЕr�L��b�ьF��썭[���r�߿��
�
��I�hzPM�$��Z/s<gwР���(��ƥ��L��*��Y�Z3�=�!cQ4ⷋ�Jz%�K:�P����X��)��rri�}?��K����`�����L�|w3����7N/sJ$��Z�yat�6i�:���bB@���<�'��|K�)�KT������v�n�6��:b��9>�
�u�9m�(c1�):����jp���_���� Ӷ�:�C}X��0x�ש	V[E(������Y	��g-ʮ	f�k�y٠&��!m/�iE�X0�t5�|�L��BEު<��d1�(�v�~��EMjw�AV��}��~˖!��d� ��5�ʴi�~��3�����m�p]dDb��Ξ�3N�.w_5��9� �$��[��񣡑�p�ojh�n��CjHu^���@z�C+�jtmo��&����`r��V��|��ı�{>�����\�R�gD���������"�2��Y���Qn'3 ^Uj�1]Dv嵐"[��U��p�`�{�0��wğ0���\�y}��Eg������ hr�HNhc���CMJ�?�� d�}u�]�Z������i�Ƶ$-�خ���ᄺL�Nb���V���ص�M|��B�;��ܠ�L��~Ć�k6�5�SQ�D����ȫ���
t�CGV���?�c�DA'V	 ӎ)9�;����MG2��KI�S�� 	/m6&w��x&�S޵BL��!��X��Ոխ؎��0^YS9�L�k�0[��#^�]K�xs(�Bam�c���@�\�rv��$��a���ʋV��PM֦:-�2,�-�X�����9�N5i�o9Ǥ:����>�.���#��՟��^�b0��X����XBߚ[����#�!�J�RN�^�
z�r(/g4�dkeV	�tN��i������a{!tG,Н�|DG ���\C��F����3)�}���OJ}��M>�BA�Ҵ��;�abXT(��*c�6��^�<މ��ٻ�D2��WJ��_�I�#��u�7Mȫޞ�q�ӛ��~����L����w)\�M-gr���R�����K/�^1�I>X+;5�E�w�r鈥�dWE�'���s��~����J>*�IL�ĐX�u?��:����r�B�&���-���T��$,��]c�Mϛ2���iG�_g�!B3�A�ӺG�x�3qKX�+��Ͳn;v�=��κg}i&�U���e�J�߲�z4��vܫSnc�@�e5S̚g~�IoY�ޒA�,��s��4�t(u"���;@���%�0_�	
�%����	 B��YJ��ɤ���z-E�]�y{�R)��\w�y*4�_��oi����$��������,�iUq5�9ޛ�������D�J�i�A�ߙUI �2.=�m�[�vs��V�	U���K	A�M  U}��oy����9qF�x'�����N��.E�1�p�.���X�7�7Is�V� X s��˜>]��=q�����U1�ep�)'�B���>�{��u��M��Htɟ���5��W�8��#�>�:c*��O��Y����oQ� |BJ�0���J������+��ա����F/���cI�$���#��j�������[�W��i;2ܬ�Y��L����Cۊ�9'�$D�aM�Z�%��S*J��-ߥ�>��gl��i]�J�%_sYn����^��)��KLgnH�G�*q�=r��gx6]�_ ���N9e���`�34�ё���X3�F2�hÈ�a*��Jۇ�B�n�񯋁ke�t�����ِh�-��Qu�v>6,[/���i�IIXi=������g2�\��# �Uwq�V_F�S��vI@�(�J7��$�� ��/=HK�p�Q�!�B�ePv(�Z�o�\���G�(>�߈��~Ϡ���uO�ў�d�~O�c�����-	�1p�����ݛ�ߩ��r8�I��QW�W�����A��ۇRo�u�hv��k����%� 8e�R�i�n����Ep��Lг�U,��r���8��n/t������^����ݟ����Q�Ѓ�cΊ|�E��c�����'L5�Պ�p&��!���~sr9�T9�|��)LV�A{e Ѹ |ʰ��� ��`1���� �5�=�����c����}��O;ծ����8�S��we@[umM����eA��[��CT\H���<�]��I�š�@ϑ���Wd6@���>���Wi�5���8{�d�ri�.�����H��}��1H�]0
�IrL%B1]�w�Ñ���g�Nok���L>^���C���9�]ǭ��W�>t��L~�0��&P����rϊ>����q������'���ሶ����v ���"<w��̿u���s�|�W�˪�ȆQ�o`=��ϖ����u|��%�"�^aO%�Z�����冝�	&0��T\�
�G��!7�{~ܢ)2\<�ړ��k����Y*xpA���9�A�붒������_�G`t� rv*�M��@M��iHB����܎́%l9^}Q����y��Q��ܖ֋;�nՠ�L���2`S��ٵ�{GS��-�:b �-/O�9�f�f�[��.ݦ�_c���ly�T��^�e�����|�ٵ���z		���34�͙]��2I��s��y5%X�?�ֱi�X�*���$$ۡ�]����S���.�6�U��@���l���`&*ئ�Nŋ����s�����ݴdpv���Sg^O44U� X�~��㭒���u8~!�'Z�V�D]Rqa�B�5������KH�C9:�/�'��[v���$�;�|�t~0���<�`�))qkW�S��|��f��4F����B_�7��}q��Dg�rD?7.j	���gS��w�
�Ơ�82��t�[��݊�%�<����U^=)��4d�ف�6*�ے]������D�<&Je�%��ػo�Ԫ�Ѓ����!TFж �7�6>��y'��6��-R����z���>Fb��Π�¬��3��H�z�]jdt��>Y�L=��d��5*e����Vo��s���2�~��z'�����&_��\���/21 ��� X}�;�Ӑ+�t����Z�ѝ.%�zf���|�b�#���,h�]	"�?������t��t�R�� �,ǒ��Q�Q�?ta��z���� ʫ��Ge�h��ӑP�n�;6�M�OT��Pg��_��5�e�?^Z���&�kE6�(��^��!�uZD��^�x�_��An�,�):q�eT��*\��Qu@����t�K�/"�,	I�B4�7�����>ާ_������Fe�&0����m����t���Z�&�5.�0�O�	z��+���-�Uޗ��Q��H�N�����{�'�g�9�Hn��ĳWmO���ے�e�3"����2<qOev�FG鶎�� ��3��K"��-��/�����}F춒w;�$��Jkc���=��tu,�Zu���.G.�?m	S�j��Z�F�By��E�E+X~�.<"x��j�p��2�{�K�(�>X��mǓD̺P"k盅��m
�x�A�K�1Y-C�gͲL"��8���&�~Dd�γ���s�e,3]�<�t�k9�V��?��5Ҕ��R�Q�5�*GYh]�b�M�����mV��ˬ#� s氯��3��\��)��.2� �+�8��&�"-�#V_��%���)1q~T��c�y��H㘝s���������ٴT}J����^}��������R�&�/J���f%H�B�롄�����l��!��A�`,�i� [����Т��>��C?�}�*$6FTHu�Pm�PIp\&
S��0=�4���n��ϑWt�^[�ܝ�r(.�؀r�U��*=�z6��0Q��w���3<�=JO�]������O�_,��c��%s�����.ӄ��D�3j��8�i���!1]�<rů�����kBps�@��ӏ�2&\��]Z@���Ksg�VwLAT���ie͚�)4n�R
+�)yV���M��u%�����Q��W�Oo���%�s)�v=��hhy\�4�w�e{ӌ+mZ�ƤV�(0�����b�u�6?�X���Z#1�ʓ�m�,���#��VY����s�lI�Q����O�8*�Czu����{�֟���>n|����*x�ⵃ�o'e}2F��Hq9`)��n�n�Lj�&�n��Җ��a�W,|�i��T�Bdt_ɰ;֭����Q
=	�Ae,��f�3��u�Q5�]-������{����Y�e-�G�ۢכ�st����Ó2�D`����&�U�6�����?Ьq�h�-.	m��L笤��0�'r�0d.o�r�J�=��ٕ�T�}�q�줨�(��nɾ Y���Wt�^H��
�Hf,�J��u� OE�[�YK�"�G���QW$�5��>�R�	1͆m�z�E�P(����]P�c�?�Ꙟ��E1Ig�B9��D��un>��l���>���_?���i�z:���`O����&��xqZ\2j&���pi8�^ޙj998O(�b������D!NKd�R ����� �޷�0��I��0%)/U�C�,��׹7)NC��N��Q*Cy���V��}"1PH�&RW��F��u��ERj��"����Y��RvI�v��`�i�e������W��J��������
0_ĝ9>�.�~��I���h��V�-u �5�	S=t��"�t�Z+[�f����q�q����66�c�f+f2Q:&}uoC��K��}ZX&L۱H����&��-�^�O�ޚ����i��e����9P؅ҷ��Gg�"�B#�"m��VԢd@7�!�0������7��wF����d7�H
��r���,y%'xob���1�R� 	�ꪝ�8���iu��u;��K%!��]=$�觟o;�F/��'��
�	h��AvA�aZ[�L�4_�Z(#Hl,8�^���H(�g�?�h���� x�lwM�0���:���X3kZ%�؎I!g+�H߹�)��Sq�u_`�W�*�:���cS֭* 	��֨�idN��.|��ǆE�h{{��M	 ڔ*j -��DEs�������Ɓ��0��@����)�%��rx`kÅHB����\'�ϹV�@��hTD���2�F%�}�a�T������ŵ�2�0�8���%7�����ʣB��P- ��%�@��L���-�S��{�tv�sܪ0?��TO/��}2�Á���XwB��1Јq�����i!��6����ԭ�f�P5�l�L��z�z=ɦ�b���J�A�a��=iZtxs"�ww���L_�����z8�_P�ر���h��r&��S(�K�W�,J�(\�T����Ȩ?�B���p�%����`¹Pp��U��e$�4��#�*��������JЧ�����d9��V��.�A����7��v p3�Jf�R�u��jm�6��UƄ�w���`d�/)۟<��?��ܑۀN�sѶ��궖7��N��9�>jM�:�7��_��wB�<-"%fҵ$d�lN!%���l8�}	,�ƵU_4�u�*E��4���kR6(�"���>1_�@q�����d}���MEи:�).֒��/T��~��Cy�.nL� Ӎ�T�y���WE�}`o�Pr�/I�g������ ��.�ӂ?����(=���[�T3J�h���Iρ[����䪾�o�� �%�O���-:�brY�'��ȱ�œ���4���c�,�������=�͝9?�ɒ�sL��R߅�v�"m�UT�{��͆����^���*]?ۄ������Hm�[��fN6����D?��a�@|C���
�fu�x��=β�(�݂��|�R�^���u��nK���,�CL�7�
�1/��3�e�o��^!�6n6�?'nT[(2D,�wʣ⍄F�j��Ȁx4�wx u�U�0����=S��L��ʞ�=>��~�ӕ��C�X�
S����5��$�<L6�^���J=�>r��0O$5B�FħR���u��+���z,��`�"�����q�ذ��$�oF�Lv[�=��ws	N����8�ՙ8�n�l@�_86����h�h���)q�RЪ@������Pc����g5!�ʘ�� }@q��MTq�G�� ��ћz�`����N;;Y�����lK�n�:�,+�9���;#�5 �|Ʌ���;��6�������F�`�}�c��禈�V2X��P����M�a����0Bf�(�5���|���H"Lt��5¶ٱtB
���/�H�1Lfp�<	3��2t����$��^�#ݘp�����v@�;+Ž����g)�ՖR��L�;좍z��,{x"��S�w���s�B��hG�P]���ٗ�O�AT�]c����!S������M$i����W�$4�-�*z�GD�'𑠯I�?d�L����~��g����O�>V�l�F�%���|$����3����W��ùa���6ࡹRD�G9$3�{�:aNTs!��n�^W{�q���	[�����<ӻ���"As3S$	_�k���Y�.��Z?*�ΑF�v�#�����L�ɍ�W��Y�&6��ޅ�O�U�c�{4b��6�òg����U�`�+4Cn��^.�e�# �vҼ`o��Nbc���9B�Փ`��r<G�2z�f�I���x���Z�ֳ�E9���&�/ ][߉��a��hlo��n*���8V���h�u
{��Y��J\�[M�����D���H65[������C��LNY�N��������F%��䏌�CA
]i�8ݞ��O\��D��e�m��:�JV���Dt�3s��,�$�r�=�s(���l�g��jɸ��B�E%%�A��wd��*;=��t�<�_X�jX�@�脑'<��az�j���X|�9�}�ڐ�7:�Q�Uz��ؾG�5�LUU�^1��Ҳ۩�d{��Qm��~ZuK��0�����B�%wC =)�٥&TyQ2\ӏTCJ�̧��IX�>ѣpΘ/Å��_X�-Z����������pw�7�L�Z�pGva�ag��,���'��V�+/3X���y��b{E��0�?R%��BFv^ ��B7�T��j�{>�K�m��l"<����<�����hJ��)��`5u�E�%�v��M#B�O(�P[3o<��G����b�'��ce����Ũ��4�Ɍa�8�˸��'%�մ�۰�6 ��*x[(��S���Y�=;9��rm�^e;��؟5��_�� �ұ�ZB!;M�R���4�� ��U�|�[�	_���S�~�G�k�ht�{����M�4]�4�q\*޼��Q�7�����J����ҁ�ͼ�n��+ݖ)��$q���S �	o�0�P�%���d@�/��[�q�!�P�:�d�or}OC���V#�~��U#�Ro�1�Ƴ��p$�'Z� �`�� x1��=N�A���[s;\(��+!h��>{5���Q��ik�k ��@�ڕ��NY,��J�q�C9/�M��Jr�nvGPo�)oЬ��+}� NS�����8�6ʚ��\��u�Ak�;��\����i
���+#�^-k��} �"���¼�m3�amP-�Ku��]�i�x��y�Y��%V�F��ɘF�(۲�t�����I�^>��+g�s*L����:�q�v�#�1� �Le�?d�g���h�&�w6�\=p a%M�[ȏ���R��<����)�2|<Km��ata���E79*�\z*��G�[j�x]�AK��)���rL�搉C n�G�_���z�>��jwX�`LΘN�!u���jz~�S J�W��U+r��A�
�A+�i���[�b����[	.�v�<��x:�h�)����Zt��p�y�l�Rʾ���u��}����ey����-�E9�����:!w��9z��D@KE:�A��|�6i�G-Vݖ�ͳ5��AF:6 �>�n��h����7<o���3�&����.K-vO��\����f������q�kF&j���:m����@<��{n�U�lF���{��9�V����=B9:�4�5�CX��iە��le3����t�q��hK�Ua�bIV�O�h�/r]����u�F��i��z�v��Po���BD�|\�1��uG�(����P�P��d;����Ǥ3��m���
��is⿠���w��qȝt/C=��ǗڶIX�a �^W�D1	�G��Y4��;�f�c8;�M�l�ˋC�sz�s�x�;��9��',.ND9��3�T���Od�,���I�n/l��CrO��v�LH.K:O�!,6��x�� I<o���fS8�,e
T4-WxP�Ub㩕����xS�	y�o4�?�K|��J�Q��G�?�������t�$�
�!��Uv������^�6�<��;�!���GjZd�r��V4���JRQ���h80KZ����P��P1sgh�Z+�Z@IRh��$Y+	��([Q�n�*Q���$�Q_d״��}�є����8�O�[M}��L7���A?D�[b��zGV��͹OΨ�u��zX�K� ��sΙ'��ivG�K�5�-��Jj0/���9v] {�	>���X!3@*�u�K�K3檶Q�c��H�ιN���r��.�w���͐4L4L����DZ�;q�Z?AbG��Y�C�k2/�m�R��f�P�$�.�Ά_����1X�6�%}T���f�q���ii��Vb�I(2�'ѳ<d��!�
J�m3�8��0�FL�#��.T�6w�z7R�G��7f���5��??![P�uP��b�{������ut���-����硪��B��~����ugtM'���9dO;�ל�S�m��A��/e&}��Q_���B�Q+II���f�wt^rR�NJA�������b��9� ��x���&-5����C����u���@
8�kِ��f�yv�0	��[�YC.Ć�n��6A�j�.�6ͩ�����&�-4y���'�V�X�R��D7A�h%��Q��8�����>���81"�&�8�ۋ����:���L�Z>1 �p��%FG��g��i/�#����I.�.����%!��~<${�>]}˕���0�y��U�㷚���դ�6?�&1Ou�R_vL
�߳���Iq�9��+d]�.�m�HuA��!�T�����V&L���?�0Z��J��n(_$�j?ȝ��|`ߞ��V`o�5>�(�Ow2�6d�fn���䔅������6EBA&:�׊���It�T��g���}_aк� ��%E�l�MA5�J���I��ꍼy~۸�M�"�SG��&IJrC}Y&�( ^n�E-�uy���
������^��A�����ɣ�.Qg�L� Gw�qy>���@J|�H4rXf��F���9�<��	�i��f�ʆ�YN�\�	ɻ��W�B^�3�G��z� �ns���°����#p�aIJ��yXf����US%U��쓛��% zgXl����rl|�"�Qձ�*_��bSI@I	v�3��\ș3l��߀�2�bI��U@Oە�Ds,c��B�%I['$R�%&��MG�G�g�1��T]��>����(���_����2Ic��׊���^�(��o�%�R��Ж�����������M�-����Ĳ���:�h�ב#Z���<!I�paZ8s��%�5t�e�C� �- 4���U؁t)J�q�R�����}�H�o�C�����)/��)��)Ē4w&褂mY�ƫ�z.Ҭ�R��Lk�����$zf-Xi(�'n�B;o�:�w��.B��|�m���#^2A���?�Aa�g�ѺɅ��z��
V!h����|첫6���om������?
�w9U/��RU��$� }�qM��,������9���5��_���DX�����TV���ě;�RI3�i�nX��e�5I�34pF����^wz�gS����Ի��@ˉ���W��M}ǳt�%R�7�2h~�jhe�ש&�:?��qR���r��tV\��7���h�(��<� <,Y�d!�%/�j�<~Й���ċ���f�\��� [��b�ƙu":�^OD������
�T!|ea�B)�u����Oɏ�y�/ߡ�x��MM�vqҟk�0j��(A�4bq=�z%�e��
�x�)��$M|�:Q�(�n�M����8��a�E����}�o ��Aqd}z:-�(��X�EݠdS7QLa�n�h��%���J�?���!4�U��3�2�(�j�npx��� �C�.3�uj���Y�/�x�R����N������F�o;�aF� �:o�œ�������K�)��woaJ��+�'g���G��#h���j6��[���������Wk� m�Qs�-�~L�z|��V_���C�,�F)����5:�A���E	������j{���t��;���MÄ՜�ʛ���=Q�/#�$�bWuÛ>}B�_5�fY�(f���m?������GB�Bƀ���+B���vFَd��05fN�rC����n���h�[���������!v��2�5ʬ�ھ�Z��Tg�����톽���'Pa�/��#�畑UA5R����W��A���)��h���ڋ)b+�7 �g�L�.p�D��Ч ��>N���*��ziʥc�����]�=�	�9l\y&��5���i�����PX�9q�2NaDa�M�񅢌�(�ԝr�S8]�(�I<�B�K����c���v^��A���Zk���w6���:O�~���Bj�@�#샹��7Cz�}6L��c��~a�Ԗ���%E>�Ʀ�F��Oi��E�Og֬6�0��+�ѯ��}�q���6!��#0ԝ�6e�����S��.ѢR�P�k���_ ''Nf��mD�ϴ��\Bc@������)EB�OԷ�3)9������`��qYvP��8P	'�:Y-�"L��Q����h��	�cnQ�47��X�o�6�%�wHu��
�8�@�����|�ok��˯-�B���X�k���5x�]x�H���':���jP:�c�l]�X���s@�`~[�'t��g�L �zV�+1Fc h���@��3���G钂!���
u�!���p�$`{�� ���>A�Y=C���XC��&�����}uI:c����i��Z�&��/���(���+?(fn�G]��L�6du��F��|P�.���7k���f�/�9���v�Z����u�i��I��C�\|B�N�n��;,�e������r^��%/��g�L��_?��2D�&�O}i#���9�Z�IVch�"}��!�<Q�+���V.Z�!�op�~?Ys�g��/��t��6����[d�TX�`3�����\����V�F���%�o�T�[�������A[쩎�.�:p��됯�Ze��r�	8���a`I�l�"$a�C��<W�҃�� f��O���|jM'z�b٨�Rc�c��G����D����5bQ�#L{�����e�.l&xDr����h3�
0,��8�a���Y�㣠,cx�O�7�N��7V�<��H,�ވWUkn��@k!pI������Zr�e�ҧ)Ǭ��M���"G(��s&����i�Z1�fY��5���u��T� �g�r�м�]g���$d�p�����"0�YV4����K�й�ч@ޡ �=�MBU�h��mn�����-ZlN*��Rg��^6e����0���FP��Y�L�2S�yIz(!j�<վK2�Փ=�����*�����Ota \��9�{o�c=�����zI��[ZQ�q�
�f������O�y��`��1���g�x창Z�O(e�{�@q�K
ם
m���U>I\�R݌ݚ�UKŚ���~J�qL��k��@��g�xZ����yt� ���
L({�{��x�]�Nֵ��7Y��-} ��u]9�O$hp����q��*^IVCZ����[V���c����.�0b�>o����
Us�d"�S���d���>3��qB�z�4�-"����"b���)G�`�� �L\�G��.����O���u���V�W���2+Q� l~0����ސn�=0&@H#��*����O2u��?מGA��Z�*��Z͚�3ǎp�D�/5�G�[A�f�]�� �_R�Ֆ[-$k�r��G>��:Ǌy�i��=u��7+�	Fh�0��������� ���j�*u��$�Ҫ�ņdVA�B�1E�O /
-�ia{@̎9��?�R��z�@R
N��r�֔��ve���`��)@�W.O=�i�Y&���ʔQ�[�k4�n�s�q��N:�}cB��9#��G�A�نd�~t(��n{�I�MN�:�ُ�4![�xY��!��Ү�\Z�Ҥ�<�~4V��?g50�8,�J1z�`�+q��疓���r�:L����3M���_IDtO�V$=	������Ig d���]�.�}:��3{����wr�y�Q�.0r���Ydؕ��PuBHt����Lt�'���|֖�/)�����)���eJ@~ ����A�-7h���{ΟVb����U�]&��r{j�r��~H;W���/\���K3��#���#/}F};Ա��xn)�.�d�c�mŶȶ�J5s<���f��F�m�`� ~,8��{G@�;�R�T[��D۷.���40-0��aP����O:^���<7�ĸO�m���.�1�D��NƖ��C"&��g��o�yз�G|׶��r�fAE�7��s�WŲ�>�Ɋ8�^%@7!m�(!�.ڙ*�u"R3�{&_�;�|����w�7G�r�� �w�Oƕ��|ݽ.�P�5&��	LӠ�����A	5�Ky��6{L[zd�Ú� ��A/�K��u�k�����|It����t+#�^�
Gr	F��]Ĳ{��zd�2>��`F����dw�����f�?Jifr�M���)�u���(ط/%�
����&���+n�����e���T�%jE�����v��`/>O�8(�4`q���*KHֲr2p�2g�]�}�9�т=�1�",nhIs���ɓ��>�S[�&J�PKlB�s5�$�ɛ�ME�Q"=�|��a��=J�˓�Pj-��k4�rO�W���:�y�ɼ�H�+0<Ԋߧ�l�'Ȕ�|Ďn=*sA��8��mg&4��_� ���	��P���s|�TI��XxG�s���Eɉ֙�K	�L���+/��`�������]τ�W�$ٓ�?�,$V���#+:	,u�Xk�Yp���E�>b?E���{Ȍ�� NӁ�
QZ��E��!��e�1�m���FB�S�'�_ը�O�/��(���k��|��+�K,bR��D_�GO(���X''�e|�g��V�Tt�ͭ���4�|y���9��20��G^���P�*��y(�	5��n@�(tC��P�8mRۼ�U-�:�C�3' �RixJ�Q��E88��7T�����{n^8�4}-x��4*�!��i�j� �E�&={Un�(���乢�3���t�a��ag��b�2��ۣ��ظ�?�%�[u�_�p�)��n�<=f!k��Pā����`7Ң�B���Tz���t4���̵�nc����E�H�
 DpH�P~aCy���uˉ������8턹���$�V��\�F�����h7�6�R���YΔ��բ���ɒ�x^vW�G�����A���f���i�)h� yg,�#�F�-�,�S��L�+�=��$��o�u��)���_L*�E�Mٺ���'"Gֶ�S����e�v.�<\��莴��,��;���e;�0�cp8M���؝� Rx�����I?�Y�,��=X0ڣ�bv��ܚ���Q1
��ch�rO��C������sP�TK��.����b�Ya��2y3U�u��=���=ڙM�F�^cU��/��A�	�w�C2�R����q)�?H���V<CT�-�uD��ͭ���pRO?�
�.UA_�||�����Q��?ƌ��+CX�j��.6�4rS�=��Lv`IP���9�Z�@+Y�X�)z�G<���:ىԸf�i�5�[�?��x�Y�����DM̓�(W��SE���9g���Ĺc7bI��S��{	 �pT"$;U�tT��4�
�� ��v���ԡBH}��ﺑHM/F����2��p$m��|#�fF��3�T�A;O!�:O2$����Ht�� O��	�3	�E1)�{Ҙ�~���ng�����Fx\����A�c7%�љ����6�)Eǌ�]�R������^S�9(�j���?~���C�\�#���QD��p8��/9��ґ�Kn�w��^�ۼn��V?xLv0_��Af7Hi��I�7 AL��ܽ��\�}L�݂_��X���N�5��;��ӼR�6I�]��c�F���
�U��&?���и�۸���_xe��v�vP���S\��5��������ϡ[��+Jv�j��z3EXL�;�R�>:�����#�
�}�op��ޣGK���o�����dRFg���<A�O{d���)�-.�#�>�Q�M�� {q
bx��x�`�����ӊ����I󦕪�� ɹ���9����6�]����(�F�#��<òc2)#2��~�ݿF�wTE�̓.��WZyt�s׆S��GI��)L�8	�D����Ӏ��>0��Q���hG�7���
�`G�ּ�φ�\oZ�`4 � �M�pXQ����9~}���S�������Շ��N�.G�k�;H�1��ӆ���Ni=�bH�rs���bXݴQ��;�����_|L�!��&��'<(��ܖ���x
�~�(��g�l���B���y�b�'xv�12�:�ܪ�w�o�	面]�}�B��jX� +w�M"%ۃ�X�2;�x��@|���jm�}�+�ן�
�o}�/�Y�����U�G�r���c�T=a�R�X�H�`Q���qH��ӊ�����<A�=��*�=���X�!�[M�2�|��jQ����+6�)2��#���{nj4�q~zY�+�5ի����!�Y�y(��Tq��/�����LȜƵW�9�7�AM�lPVKɳ�3Q������W�!3=8��K�y�g+����?G���V�΁�2^�D�̃��V�g*4�(��z�� ��	��^A�� �>��Ւω@+�g�t��Iu6�	�?u�s^�gu���e�E�zl�������@4 �!/��d��]���N�����6a���o|��n��'���2Q�zdB�����|��%���?&���HT��*ᬌ���&�,;&�w�>;o�2��J�7���-�đ���c3g��w����@;��\���݋T��(��
�\)�1!��ԥk����U����pGƁ�%`rcn?Q����>��u��6<$��-�nx�┣1��[y����7�P���"HtMыK���=V5�J��qX`��C*@ٵ �r����.�爪q|�y.�rf�,�p�iX���$�,(\dx^��/��ˡH�5��Hg�3kQ�;F� 9�w>�4�nM��o�5�C:����ab 5rf��Q�9�{�R���n�U5*���I�  W�W����/-x�u��c��~�f�P�Z�"��w��XS���5\���)�����{��rN��Q���>��A=���!��,^���0�^�ٞP��^d�t�,��K}��*7�M�d�����2 �zJ�TZ�pm<�z��_�����v���o����,��9u�g5�	H �uԴ�����,��4�5�z�=.09�e�fBۡ����I��7t�9�C�U�.yv���]錆�za-B֔ں�J�CM�kd��n���r��U�)�ɾ�u�fˆ"~M?5�>���ʁk���&bY��o�>ƈ��3 �
��(�GҀ�F+��wP}	��{�SD�S��y�⇃x�����CN@�%�[�S��|��K|�� 8��>wa����.��5�>���oȍ�
�K�>���)��k(��RIC�:s�tu pE�l�ΑP�VL����:B�hkF�G?v�o��N<�Y�7U�|�k�U5��H��>r�\�p��*�1�y ��{�m��oɿGyn��l��r,8�ё��_��!R�h�;k@L-v��-N���*��[n�-���!|��j?�Ϗe��fN%w���.�1�c��ū��R��u��)3��8d�~�^c�K�R�b�,^^}�A#̖�e�d��!w�Ѱ{���� y=�T����0���T�D�Dx\o�}�P�J��=��Mp��7~��"�!����� Fr�;��杮
(?%��_*�� �'ir��@���(�z�i��c�d�����%a��y�}Om�#=��G���yI:F�i� P�;����6n9���b�������%ڠ8��'���uXm$շ���K6�<�dP�]a��c�訤ީ�`ը�C*zOO]�2T�EɆ�޸��+�"G�b���C<��J���q��/2�Sd�(@��AR��	f�x{��+�3��������F�r�2��T���g�2L�m�nLHb�H{���ë��������5J��Q���-9�+AZ�>��p�-�)e�N�2�E�~�:�A4A7��K�@���&��,_g'ؼ nw�v�^�Y
[8O��~x�� {��3�H�Ӑ�3�+N�Y��@T3���]5>R\bX�Y���i��jt��㹩�ݎ���52�2b��%�LʵY����;�
����"����~5P�o&�Z����^�F�\v��������y;G�J�x����16����U+�(�v�"2��{��酘�s��v���K���rT�]��Q�vg�듂�#������Ѻ�j�f��R~��~�}|J�B9 ����jb{˒��9��E�y�-����Q��Y�xf5q�&Bݬ�)��ʺ��^�1ܚ��_�p#/�S���ok"Oᦧ���L���6��w�#�ב�(xf��kY�抍M&L�]X�����Y{pҲ*9%0<fM�{%Li�Su��I(r�����B�(:�2w���8��a�D�N����&29BΝ�<���	�Hː�����6j!C��9|���w�jMv�������u�Q�S;y(3a5�v�]V�2O(n������4���3��t� K��3ٔR�/�*�����P��V�^>��z�b�:�Ĳ�>�QY��.���nc���d��Γm�������ᇚ#,��x�Zj�A^��ڊ��Fg�Q[�P��[�=��2���� �l�(�эY:�[ALI�:����^h։���8Z�HYG���|�f,\YH�j*G������sy}u�9Ǹ9#h��<�������"KK�>�u�7����$=�MﷅPI��ɔ������	o��U�P9����i��4<��poέsX#,��k�P�tcWK�+�,&-ab�3���'��:s7���s�B�� bI��3o�_�Iy�ڞ: kPZ'?�� 2���
�gw�V}so�j!���GH��?l՜��y�ށ�m�\��{�p�PH��A̘W���������߉��q}����S|F���� ���gΏH{�`ĩA��I�Qw�YV|�)��~�v#z_#�
�{6C^�-`d�SƠd^�֐�<�m��7�k�������m�x���IȖ����pB`�l;��q�	��"~�jcߺ�S�
�#i(~s8z�������v�<r"��ٻ��]h�c�ýL)&��7�U~c�Gh�\�h��JR����܁��4��D?(V
���Z�Q��zt��`v�#��_F�>ιO9F�÷߲��4��R�Ne�+���i�GZ�Di��|��|�'�B.䣦G�c��o�]�"�6K�e�跚&�:��Ǳ��6\>�^��^WN@U1�����O~��µ��XJ;�]~���l�Sc��0��X���2�����ݹ������D��4W�^y7��D%a�~���Y��\4_���5ʫ��YM2n��sּŰ_b/�&�¨휹��D)�_�6&WР� ���ơ@q���Lh�vD`����g�ֿ��DU]A촒'�Ӝ�|R}��������oc���{P�"�J�� ���Tp������~�fX(W�L�n0?ᎏKf/w��!���ߎ_�,�&��0�O��h�>,�Z�)�HI r�i�G6��Q��`7��=Q�9���bnhA�����ӑ�d�#�A�a�
��/C�����]���Sw��Hmԕ(�է��1K�1�����{e�|���4r�,.i܇�	��w�t�f�o���npG�3�^��&�ё��pr�,&N!�_��c-⬦� 'O������%�_MC$|�(�s5)�����;�,�|�TT�I��Qh}��w6B��� n�kg[T!ɭv�l�j2E�BMM��}@�`������eO�v �hfo1�j�/8��R}����-�()��r�F���&���D�0&F��W�F�[.U�z̞}������F��+quc�� f$�������`3��5ٲ-�~0����*���<�r�c���=rb|���������ϕY.�Hٔ�}h�f6�$�HBFQ/�)�z��>8�G�u�mX�H1w�Q˔}KI����I6��k7U%�Aew�֭�}�pBi/<"���������� �|3Y�f�2JP*���T���6@��>�;�Fٞˬ��Δ�vۛ�vR�W�ĲS)'�g������Z�OO�h��H��>ş&�Nz~h?$��Z��x2�Q̸��uQ�վْ�i�`�]%��9�X{RQ�8����8�|�(vޔ���$��t���^�P���'���f�l�ޓUX������Lܥbg�SQ,p���nb�����;���������9(4��_C-��+ +`�<�'ҠC6��R������tac�Gv���!�6��ݗ�˾�Q4t�_I%5��!\ ���C3._0Ծ�
xm��CD�$+ڈke�׆��j�v��ݳ���`�{p���#�}�1���f��Q�c��!�z����R6�q����&&�"N�*�0��w 4���I� |��5Q 9�z-A�F�^���@��
S�28aq��e�C]y��r !��yX��b�;��+ےwg�8�&�T��/{Hf%���Y�6Jܺ���Ư�]�sj��S��d���Ň6�6(!�pw�����0�Ŵi`z��iuS�=��*�� g��7| �o�>:�^F�ޏ��{3�#C/�*�H,�����@�p�*��;�q�8R_|����Q[x�](T�j��9�|g��A8&$K�鍸�2�z˥ex�D��g6��K}�nR��*�AK,c��[��L���5�^� $�:!��r	��4~M���y��;�j)��j�iܱ�O�7>a��ȃ~]���c��� �o��N����` ��Y��8�%Zٿ�\�B����d��oƼH톉X�<J*/-�$���Y���#]-��:�c�:��޳H;%}�����O��o�Cd��4cȆ�
��c;����a4�t���Y|�c���S�^�U����Z���#��H�/o�f���[Gך�z��{V@D�.O��b왻��^S���L�U�+B�&E�V�� �3�VP�^[*��M��q^S�f�
��$���*�Xޕ���1�=ڲ�2��p�-Ӕ"����Y���OC����C44� �������R{:���d�8���v�����;X0(B@h�M��Q���d�|��=� ��;�fҩL�����Sp"|�vU�/�FӋ���,#��л��8�V�mw�-�FA
��R�/.�8�k�O/�ԎLl�1�|�G5:_1%�_��b{}n\���?'w��Ga{[ S�8kQkrC�%x�TѾM~r��ffӷ�3Њv�Vz��yުF;O]&��-�P���!ωr��V�T9b<���B�z��K^�f����g�E��<�3:kQb'��:��PE���k������ں�~ӹ�Sݩ�]�JX�6Up�}û��" q��<��j;�V	����.5����KZ�kAl����g�W�t�T^O���Yd��z�<��=FNB��e������Q�= �W���8����	��u���۔��8��B��D�)�`���vڄZ&2 ������dQ��ka�cc7��:]E(�EUD�-�T��;)��;�9��7��y��/l�&�:�0F�	Ƃ���bK�7�޶�.M�4��z��^���a�|�8�AF��v]\s�;����ֿ�\��=��c.N/�[3I;�8��}]����k4/�3n])�J��H.k��;�qT���u�Ӫ��X
fgi/�����2��U*��])�i T���1�Px�Pb�L66W�p����r�{�9RfO��U�|~�R����p\0õ>�F�#<@l~嬢E��o�)h�Ek&p֞�vlm� zr��s%ȝ7�k�B;�����H�I����	�7�2[��u���HM]�w#���9a��wta�q���'�37�	�¨��)wt�O1����7н���!س�^#%�4z��~gi�|�@\��
zIk� ����
?�HM���xx�A�`b�܄x[�4�d4|�aD}$3��FL�sk6�R�k�+��^ڢ0T�.���]X�f�)�bk����9���С
A��ŽI�Tk����4��iK��G�"�}������o���$�i���������x5��
�]�K�r�B <cqQT� K�LIAU@�d�
��Ɇ��=b������*����I�Ѿ�2,6��X*��4�f�7F/ۖ��pi��hQ����cܦSY�qk�{�9��s.)w5(v8��U�����C�S��X���	���=�[VhQ��� 0�*�A '0ʛ�\{�{���k�wپu̗rs
ΠS���(��ɖ�zش�h�!3v�J��kڟ����ͣ������u��LB:W�{r<�|(��͞X��.�^_�X�C̦6��gi.��N�Ԟ�GWf�-���{�Ux�)��	_ά���� U��!o� y-�V�/3������ۘ�#�Zψ(�K��90Jw��eՈP䦟}������g@>뿎�	J�y#����ǻ�2�$��ѾtI8�j����4eX�cSR��B�S=Ͳ(-;�>���0���Ė^:IK������+V�����@T�?-x�@U:��*��'��Bk�ֽ�q�H�t�yr�wFm�������{���	�bnc����ۇ]��X��3�bd��[�C��p8�5�����b,H:�;P��nB�da��P\�<�G���ȇC��٥M��G�[��o�i��� �xܳ��b�W��D�~��s��L�r%�W�j��G|q���4�m���e�Ek=sF`�<$����H�\yi�5��R�XZQr�x���a�[N����N`a�c�S���x^�r�Y��9;B"Y��h��2ϭw^��.����* !�Ňv�����"M�s�{�vt��q��k�ρAJ�s��uua����K 3�{��f^�!���-N��79��m�D>��f�B`��G�S���r��EI�&��'�4�%&��E;�����H]������Ŏ�_��u�!���������W;�4��$IC=�]_E#��AXUUJ����أ���P}@[J�?'fk��z�)��g>b��9��Y��c���S�^�5���؅��-m��Y�!a����^�ȓ��Y�,�SMk�?D-�m�Æf$�9�f�w�ˤ�pl��>F��QAm(������h��������h��{#'˕���⥘im��V����������ZV�1��rjz�?�U�_��z��4�g�Jq�Ǐ�'�k�!w^�������'ní�����GqB$v�؏�h�p�6�B�S�DY΂<?$=��T�
Jn2ҟ}<J6|�+
�otF����D������"��)a�4�r{���{�!���b�v�$��i��ޅ���H�L� ?:�$V�������J����4u�+o�|��.�G#�5�� >B�|�%���g}�e�؝�c��%H������\`ٺ���H�=X�������OΗV���4y��~R��DtS��_��	!�����Jjs�ơ<	i7[8Id
��#�l�i�g�'��o	f��_0D�<�#Q1������(�V��n^	x��̢s�У��a��q�v�5(�&����-^5)�}d޿'S�4<S�-I�+�<���H�#�;��V�ߡ��\,
/���]���(�	G�!*�~l� �:�y^,!/*�K��~NAܿwV��z�D
������v��5��IV,_�v&N��<��"�7�h,c��+v-��U��8�yB�޷#�sJh�C^�����{G�Q�MM��Ǌ�b?�!��,��=��=�ʧ[�������x	�+Ys��]u��=>�h�㇚pYo�;��������H7(�&��0�r��¶�����-��)�Z����$۽<��بK���v{t{N|�5�b[�o) oA�&3���S�o;�l7;tǆVm�(q?��E�'���%��B�WO����q;v
N�](�Ϝ������|�����2��#��A&A>���q~F��	r���x)y6���4WfԊ���������{
Ad�4�]F��W���g�����o.�o}³�)�e�S$N���_�7���%H�� �X������-0m`͝����WD�M��sߔZ\���L���╡-��f�_ĺ~�� H���j_�5�M:̻N6�A�riС���#B�%Yb� C�~s.= ��۞�f ys����m��v����?�ۄR)@���-��i����`�'��F����&.n�5Y�7�����3��~�>��"�A�:Hr�h�+Y9��kg{�|�s�S�È*���蓷Q!�\�W��]�z0��J��F�DZ8v���|���5�=��@n?�5�P��.��j/��j3C;5��"F�t�Q�׎g��x�I]c^�|wM٦��޿��#�r6{�Wդ���C�G,��v¼������z�|�e�X��\�ze�I|��-3�(	:�"�o�`&6ǆ�M��������^�ߗp�]Ժz�̥)��1�z%CG�Ai/��]�_V�cX��ʂ��{�hGv��J�:��M倄�6XyH���� �GK(�e]� ���)�U�l��+<���̎W^�,�O��+ n}Je��e#w�-�{��f��N<���MU[T�(՝oz�a�!�b)s�X?P��z���6�\mr�\�]luoi�Ҧ���v�]�6*_¥�h9y��,;okS�ا�#���RzT4�r!��g��!ÅC��_N���C�	��9�eG����)�U�s��%N
�����U`=B`�����Er|?w��Bx�0"��P�2�FX�a�9�\)^�A������ǿ�{��3BE�%�G�O5�O�sU��'��17l�s�i�8U�ߞ���0R&/�J/s1��h��C�^������m 'b%��N��h,~_�*�ae��D��*N�5�����y�!��ٴ��u�R�C����v��_8�>�谔��\y�Ch?���A�A5������+L��(�3���Qs���@���u;�t�_��J����T���F��(�b�_1B�_7�IЉ��&�'E�D���@{��u�|n��a�BF���MB�Ě�G�:����7�X�8d	�H�1���h��C�a�p*D�Q.J+�9�r����E���**0|,Ow;i]���&���~��ĽǫR��,F3+��M/i��7	}� ���d�cAaM�m�pk�`$��;rج�^�R-������!��v"�c��YMF�e\�Q���7����=�$�	VNcF�2}l��L������3kjV�}�J�1	�Z�������?e��V'�P5RhM�	B�"���u�B���7���LMv�r(PR2:��:<Q����dy*<����*B�$q3p|/d�7V�K
.��.�ӌ���i<����k�꼆��<�Dr�C�I�t���H�f��6�v3Pv�n��U߅����`��e�Ӡ�]���6�a5�p5�r0Ve��`6�ɳ:"��k�����Ȩ���Hh��yok�j��Z��J�̀��ЮQ���M���g�sf~�|a��=�a9:��-�)�򗉙���_�������>r��������!�n�v.�n�f8D�;0��~㜦�zq����^�13]{W�����}T�����ڭc�dU5O��(A| T��P�F\`�.��7�������}	>˓7Y�n�3�D��I�����M��@#E}i����j�0��>�أ��M�i��Q8*���i�y���5���J�FK�0�,�{@U�O��A	s����}c7��;@�yROخ=���Y���ӊ�G5�*VE՞�Ϻ��UJ��]�{�{�������qA�VM1B�Io��lViv�{ԞK����7��c�e	�$�S�u�ΨG+����[#��m�� ��\�߬��7�<�Ma��}�X�T�,��4���ڰ��j�c���<>�pe��ŝc�R��s	}�S�{�`ƺ"�!��f�x�C�?�䯊�KJ+d��gho�Xn8� �%^�1^�@�Z�O���sb5ڑ,�����v��HO5��QP����(�a�QR�n�j2J��0yj�J��(�䊈�;�����)��˦p\!�W���
,���V�zH�p���T�+Z!I�x��[,Tu��Mv�DG���5��5cL�<��Y��n�-e�8o�5�1Ig"�)��R�:��(��4�[��]��5-]i���`�s�)��&Y���6<^���ym��\�fXj�U<�rؔHK�Z!�����|��Rl淶�Yf��2����h�f�|H�o����s��!��GJ�So2���'�4�L���G�[*+=�J�6�j)"�/=�9���z+��d���E�fm�|�{��/�Tj?����0C�D2���W>�Z��l݈��t�xuG�p��Gb �š�
טeX$h��˲?���b��pM��H��)�o~��?��� �zR��/�9���p�X���g���o9�w�v�d�(��x��Av�,�꤁�����3:�j̥��l�*U��zҧc2�A�1kI�W����y"�+�hO��Łi�λqh�;v}�-Y��D�[4���w&!y�OЭ��{{�p�H�������]��D��B�����-]��&g�NY%���M똭�%W)CTE�O8��Ea�E�P��5/w�V�����	�`��j�(
�8��)����j�4[��r� ��2NH��^��)[Dv�b�>���O ?	���r��xt�9�j��	�2֖��;�CI1��lZ�Al������e��ɮ�<��Oa�!~�'�*�wš��Sђ?���>�%��qC�CU�����d�C�׬Z���]����=��D6J�fpii�Z�>"M-�3����O��(��2kC57brɱ��@,D����rD�K�M��n�p�N����W��%�����)�])̼����m��̽����N��Q3�Ҹz	D�j��o�~m�I	�6��Kv�OGDWP��0@k���{�J�׸�fIǌȠe�~����}rwP<�Pٙ� �\E����R���{�.j�lc�Q����\[K�������o����R׌W�ܴ�r�ffh�)�ùѠ���h���'�13�ؤ<���ٿ0�6E�kk��{�.k��X��"��4��ʑ2�ܓ�>�S�ߎ�
��t<5:(��K˃��#��7&t-]e-�Ʒ,�CZ�v|,>%�'�o���;�:��x��굯5
�>�O���L���%0DT�TϷ����1���o]E�Ȏ��CCY��,��~qD��E� ���/𗅰�b%'۞���Jc5Ɠb�?ϩ)�wz�`fE�JKO�Q�%9�O2�c)���pw�8j�<�e�Ga�i���-��uw�6SM��"�Be��	L�Q��U��M47�֊�v����S��#�NqU�5?6}|^�W���U�=�#����)w��>�Hw�w��\G���K��r`Ҝ�F���rkշ��$@�u7l��*�a��7)�]�߶��|KBG � ����>7���}Ѯ;_��(�3�6�[�V�n�����wN�2֠�]���F�2<�[�\s1V��>hc�D�Ʃ�P