��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ��5���5j jQ+���t��-�/����u��̩�Xc��R>G��$b�xA�Fn�z�F�X�Ӊ��q	U�z�qG��f;���,-vl��� 'J:>�V�	��0�7"�%�˝էo%���7J(]�7(MGw�rL�R���<c{��y�y$+{���k��6J?����ye�@��\��q3�!6���J�9�I�ʋ����K�e��t�f(��oǎqz':ݶ32/�.��.N�
s)��9�<�2�B�	>?�����V���c�Kz6]��0;YTHܧp��VS���J�0�L���<�0�q�j��`��Ѕn��-޾�Q7�z��׿�<SP_b�
teuϋ$y}�U��4h!���'N����F*9� z�[�����B�'6$���111��>x/�mD����_�X�5"���B��h�`�I"+F�8 3��R�f����<+:�5����]�-T̖�ߒ"���|�S����'l��]{�`!�к���7��*֨h��3��9v�w�'F��	�;����=6E�EfW"�UB�t ����Å��KKY��Q�&�5�c�Dv��7X��񋕲	+y��h�< a�D��Y?/��Mio��dX��vz��{[�BJ��?qq�:۟�hF���X<�:��/��|�5�9�_�'��0H#��丯����Ҭ���@z��JwHy���F ;��ʻ��ÛV���Q���>��{y5H����z;���Ǳ-�a��!��m�V��Q�J:p% ��[}���*�ֵr�P��ݯD�/�Q���>���ʜąïI�MH��V�"�HMf��$�o��c�AUl��K^�!�p96;�����Y"���p���_�a^!�M-'W�[�r���pU�w�i�)G��mr���l�����Ə�?��X8a�o$�P��L���'���_�H�4�>p���-�ޛ����Xyw'�(�ha���7��j�4��<W\���da���5ib���q]ٱ\i�W<�¢��;1Dv��wC���x���+c^.*�d0iI���DgMS[tz\�	Sڒ�|����ʨٱ��çj��H��9.-D]f��%E$?J�rl�T�LsQ��'b�KT�Y��A�2�`W��W��3g�:�=�aU'�&\�����,�,rT���6~���(�Y�����Dz����e7��.��=��u��1R�N��:���Al�qA��G��N8:ɫЇ��"X�ۑ�#���r~RK�է�9��t�Я��^�R�-ξ
�1�#�+�pTbR�z*'s�*�� �HJ�lJl��8���B���b=�*_�<U�P�vJ���h�@����њ�}�7������{����F��v�-n�K�6�l7ba>t��}�lK�Z���eƒ{�M2�n$�iKV ��4.�Q.�Y3�֑�¨��ݔ����� �z���]_��+iK�2G�4�A������3T�(�Dga�}@zШ�_�og�z�Կ�J���(A�*����b`&�	h�F��/��ȭ�r?z�(G>�@b Z�'H�8!�8�Y�㽀=H�oѤs�7�L�3��7�����Ǳ��t<��s���J	��U5f+�&�����=K�|j���N>�B7�s,�`�u���y�Ȯ0����7U�e �S{1e5�t� ̌��²m	�ng���0z[u�;T����m��W�Y�,Lr�,N�?���F*����ܧX
 ���BJX&�Q�
�O|�%��z�u3\48�;�e
����W�W�@E�SA�6s%"��X�q+�y�d0�U;A_y?�+�e}��	�V�U��E#��C�FB��� �$H9��5U�#8���ƣ���C�t�	#\ar)��\�h�A��YL�����fD����.L��8��OK����P:n�d�lMVb9q���YC��Ⱥ����e{0>u����B!ɭl��/�Ŵj�)A/�Y�_(T�_��U~��b�$߱����l�"�������1$X	-��n%9���"�u4����g��}��!� �Db`S<�����8D�m�"�R�����[fVڍ�+"
^&[�ޖ=���o��-�g�c���(M�O\eB#�xcf�J�Ƴ8�	pm����/坠�k�u��!B�W�Q������͊� И���w�?6/�a�Yi�3����~���0�\/��cXw���pV�j@mdY�3�Kt"v�����z4B彈]r"���2��=!�\�rPãZm|JzS�8��b���I�ȡy�"��JP��3�8��(A��/��j�J����?-�y<�B#�a�'ۡ��n���%�y�����:�3�(�����E�E�`�����x�4�Dg63�*H�lր�3A�β�3*E��v�A�
��)��A�{��d�����72�oظ��|�:�Y*74��nq��.�}�Q���Pڈu^lzi#&�<���;�a��p��ͮT:������2LWS���5 ����Бn1�=�΃�鱳�iB��D�`��q���s�u�����x=�Ä�3�(�Vu�Bآ2W�b	X`t��șpP	ٻ��	�qUǰ\. E
� �<�V����ȸ���p=4�� H���g.���7����QB^G�~z����0�kg؎ފ@����1��1�zId{s�J+��A��l6o��YL9�
��>�3����G9����o�Q�Fc愾�����W�ҝ� �1n�k���U�Ө<e�b����68�I���9_�6�w+�D������)�S �R�L��i-r�8s�O�Za���g3T����MM=�/��Q���g]����
S�o/�Z~���	.*L_��+�S�W�Q�fӺuYR Ѱa��y��ߪ�P� }:6��OtS�����{)x��k.s�
�){���֊]�(�#�z���1o�G!��o^��
]����h�x(��Qڂ����sF�(��ۖ>�X��+S��|�s���0	]�����N%�*���m]�[��ӄZ�:��c�������A�W�Xg�k��(4�M'o��v�7�DS�G9h�zI��;8�;������ce���Ca�nٌ�Kt UnW�ݝ�u�w��������[�~���y� �_�\p^뙾KQ�h���
�沵��1v��s��Q�l`������'�̆w5�*��*h�	����5[��[a�oa_�M5h�9�~SIB�/V��
5L���,�Hx���6�9�X!��M�w��B_s�0�Ǣ�TUFf?b�Wnc�*���~Ő�D���ܜҬ����H�m�s��R"�+o��6���	���#
U�ڤ	'9�i�q�pJ����|E�ps�hRMD�#Jm����>ۯ,h�pz�lIx���d.�3�+1����>u���5����! o�s*ȓ�f�Ȗ
�1CqH���ImW)4�	Ѡ����]��Tx��pB3��|=b�?m{{�D�@��:�-n��ZX�q����/TE��!g�v�,$�&�y!� �@������a̱:Hɳ��7jb���h�R]ƚ.L:%�Y04č�>�8�U*��r��+��ջӲ=G±B��K�)�_�����b���&c�V����M�G[A=��k�d9l'Y��r�V	�&Fn�& 3�T�=sQ���4�QI�����%ǡ~x�D�Q�?S*���I�oD���U�O�|�`�m�6��p�ɣ��z$�C�(mbGм�����>�ldY�d�b��&�U��M�eL�:���C)�|����1v��ϑ`x�|Th@�M�	�o��ʥQ���b2�d͒������s�d V���lo���4w^��b��-�؀�*��rG�������wߙ�)���$yo��0G	�1��	Z� �'�c�����4����oN�!�;>�f��u	�Wփ_������L��	��T��	�K�wVtfoc/ �7�Y<(�<5.P&y�P�
E(`.4��T ��Su7�W��L�eu�Bq�G��o+fª ��q�R5��|u9����Skq���
�ԏ4Q#-�0� �zdZ��G���R4V�?���Q����ޒ�b�_A|`��@�ӵ�ٰU����2p���N}G!(!t��~���"a5��%HD,(�d�!�+����*����\����ܓ�h��2	�7��ڝ��,���7��;� �HGS�P.(Yׯ���\��7Ɂ��]�