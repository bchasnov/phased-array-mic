��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\����q�?��e�I8�b�Ǽ$��"����ׯ1�V0���ጌ0�4a4�#��d-c��zi��t��{�b~?bbÔ^��~�"rF�W��$��dp}�t�a�Ds/l��}�$glܹٖ�GB���sU�t^+s��[�����/uҵWЊ�]<�4���r{>��!������D�Z!~[TH��9h�)�"[a%S-"��T��>�&{r	�ަ:�G�Ɉ kR��̍ h�Jf�<BBl������vr��QO5WH�]�6W��\^���ޤ2{�ͪm�̺C���;���o�R w�'�2:d10���M��G$1�;v�cq�<��a�j�gjT��N؉O���}�Fy^�W��$ۧ�K�0]7�L|E�D}e����RĻ�Sݛ�u�\��&k������|$v'�"2h���|i1��V���&��M�PH0P���#uJG�ٞ&9
iI��iн�����#'����_a�ނ�(�i�i�b�C�^q	>.�&�z�����ްs#/@�UQr�'p�Y�pA�x҉��J�V	�/��${u_�PM�� ����Z��Hɮ0�lk_�"Qn!��c���Dt�U����ׇ�D{��AɊ��DyM�rUm���X�,�A k����[�[�bǨa�g��YD�
d)��������	a8_����; 1��������"t���ڴFy5`��8)�n�h����x�����̞���y�:�-��|^¨*�)�s	v�^pw��DV�R�d�>{�lG����&��oZ�B�,2�]U�J�3�Y
��'�{C�d���iZ3�m�rڿ�w.��Z_�������f�1F��B����/�A��^�9��� ���[.zoY!�(��W�\�-��x$J^Q��a-�Y�X�L��;I��^����mH�1�駶��,}r���F�MJw1e�V�/�T?�jV����@}|��o2�b�KU?��X��t9oRT���xzK�<6Y)6���Gtރ�d�0m2���sk貔��LZ�B_���sGQL���;<�πe����|Y.���Hݤ*��.�4�����|H �V�<���<�㴬�|,d��W딞kEc�ܭ�62u��a�D��sŁ	i5����� ��7t*z�$��F/�Gil� ���)��y�M�~P��Cs���3]Z��wrb�<�߂O9�C����퍷�,X� ;D�c������H۳|ϱ,e`�-�\�7�7Ih���4�!�ERT�E`�8H�����5�׋dej\�4�&G�]3>'�����Q9�~� 1\�b#Y���=�R*Pdx����zf-�~z���~ g��8�r�q�yS�� �*8&�.�y=B&��|���D�Z4a���4���H�(��6�}T���D��Y��f������Iq������(�� ��
g[�6�ƨ{��WkDB4����
@yu ����:�! Ĩh9��,�������	��GHbgƸO���r���ӆ�����m.�/�`�z�p���=�${�P+]��ZQ,�UOѨ��/�u]xM�벱s@���HhZKZ8 �ޔu�w ܿx.4A1c��x� 툽�e;cCE�K��pV)�	h���6��(!|�s���hZ����!A�m�µk7/^��ބ=`Sڿ�S�X��Ep%�St=ˇ�,7t3�ҜXY"��z{�)���e(�tQx��ˑ�c��l�ύ�[�R�Y�T�4��-C����+��<7��sH��]�J���G�������V��}�Y��3t�=�5Ac6B�l�G���w�1u����C|��e�����g��!���"�0�R�WV���p6�핝��hI���eQm��,�U���J�������Q�t�j9�#����&�IZ�'o_Ť�������H�~���c9�?��<V�3Q�o����+�n�"x曂k��T�76��˟4"�����_�����>��k�����:lp�+�4��R1d4����7 V��p�=$���]��:M���iيF+M�VI��X[�$�i��Y���iF[��x��&|B7|�
6DFr%}�V��_v�/<��x���1�t�k�&�,���0�6�UX�+)5�,,�?�O��h�2,��Px=L�����^T��B˰� ��H�E�k����k��#y��M7I�^�I~�_a�c�
�D	?.w^�mhX�c�|R�����1��
rʲ�p��U@�q�K�l�~��6�VM#0B�@���k����?c�\��H��{u��L���&϶#p7����I�Tgb1���$p!E�`-��Pn�P$)6�� ��O6[E����?K(�ԗDU�@�8��M!w�ڧ���P�b��PE����W- L�������ٍDŐ��[a�H������@���ڼ�@x���x4��SJkEАK��HXH6�^���Q��Q5�*�e-<�@�b��dǳ��?��uD���M�$��	neq�  TQ;頒����h�x�F��99�_�6X�l���pP���Z!�ϳH�<k;�����%52��3��lS
7�jIo�ްLI�N�ՇN��w����G��`�����c�� ���n��?�xAw:�N��z���_o�A��Y��J5&�C9�?X\O���ׅ9���n<�W���Z�R~�4�Z��e7Na�����;C�~X��:W�f!|��z�_���~o�F���R
F�V|U���Z����|y�w�챝�7����ɠh9}_��V��3�.��$��D�&���U����Q�29�z�(�}��yE�`��̢:�>T�;"!����ԯ�wY+s'ah_�gv�� ����$k{�C4�� �6��T��J���X�HxҨ#@�*��k�YKs*w]��R�u2�Č�;I�J��rh8]ϖ�x��L��{<��<gx���]2WVZy�ʲf��"���q��sB�D��>���;��k�(�E�o���$kToP{AO}���Lఋw�܉�E���o'=�x1D���l<BI��(�՜�����e�~������FI�vvd�l?���\4��������&WU�c7�p$�2���Fҳ5J'�Θb���K8̭ƉzA/Gbn�+�K�k��07&k�`Z�!�8s�X���f�f�	��M@m��6�C�$ܑ��'�j�����^���c�uN��˳g� ~x$��X��B�}ݓ��lgB���,�0�`@lN��\s׏+7 ���J�f��7���; ���Wo���ųNr�`O�%V
�
]x ��\}��m�P���4kX���t�*��E�>�/
s�����
=e۸��	����۠g���'o��jb�H[
�"��C\�#�[�/=$�fK��1��x�i���-�,n,_s��	gߘ�l9��\�	�V:��aD"���̋ �����E����*ӿ�����K9"�#�Q��< ���ع���ڣW))�З�����j���P�\�$l;�r-��g��5ƱҤ!��A���F�O�<r}O��69B>I^r)ze���^�y2�|�;�-VtCӲb;�x�0��~p���l�U~i1�Rv+(��:Cz���`ϙi4�1\�R���ĩ�ݦ����� Y%��	�8m��*���,�/���  ����=��;����;�Pм�Dg{ٮ��X+�6�21Z#�7��Os����!�I�+�:G�^��a�	�J�VEu�)��v�O{a�w������#����ͩ��zg�kS�-9B��(�/���QѹUj��ְ��mHm�a3����/Jw�实��L�:�FO�`҆�<�\��Q��s������`X)�7�tu7 �i_���Nha'c{�E�?�v���Ģ���[�jM�Pmi��{R�/������~���S�:L���K#7k���w�q_�5�G��"��e��A��.�#��^�DYY/\F��X�e�m>����L؉?���zRt���hJJ:!nz_ت���qkw\.���
�hSq-v&��I��"��ŏIF��i�bN:5Ä>�?��nH�%�/��f�������C�$ �pR���B��W$y���F��Cv�
�����5	f���n8�W���6�j�[@o���q̝	�y�B�H=�E7�ᅆ���z3�Wt�g(Ǜ`���Z������7�v(g��|�%�C�(a�4�-^��Q`��h��7����tB�D,"d�F���"�A��b��;�&�l�V[��i��l���3�o�3쐿;����V;9���g)F}^n;�(0��������Z�OR|x+��cȁ]���y����ꗥ�ʜ_�A=L�Z5��=��/�d�;����зc?�_�l.�KV��i"�~-X[�S�e�P�0xv�0LB�X�
���E������_�\̂�Nu���	�����m��`�Sѽ̃9�|݀�( Egu���߉��B5e x�J���@��w���~2��Z3���p���s��D�PZ�uV�8D܄GB���Y��z�'V��D�E~��Ő�e�GϢF���9JJ�4"BC��3�Q����Z���A%w#t�O�DQok��T������h9���
Gl_"޺J)���ǂy �`iH��gj�������O��(��\��{��VZ��F�0;r@��?T�^�/��.�i0�m.3��0]���#֔]�k3(jk\p߮(�6��e{�(�7�.5�L;����6�4H�"S�.
�M�Sy�o���2)�{E#�{~*�W_Fm~���E��c�TL_=�{Z���w��a�,�R��f��[?u(�~���\���u~6�s�H�;����T��G7G̩^�V�����v�ƭ���8e�2���q�����4��z%�~G�	ˢs?F���,�xl��(d}?��Q��WK;)/E��Ʌ��d�8�-^c�J�����x/�e^Ո���e9n(�f����>�ǧ����$v�B����pC�U�Y�]�L���TKu��v�V��Tm�W=|��G(=�y�N#������&��&ٰ��܇!:�w��+�+�|��4�V�>�+ld�����ob��h�	�P)OI�\j��l�+�@�{�P�(gJ(D��5Q�->Xd(���m.&������C7f��}�ީ�Y҆xY��l"���:�+����T2�9��xFM/���Yg���<9A��X��.��X;�n8i� r�j�7UBBEǐ�'�@钞�����Q��|y����O�pm�ڹh^�Q�"��UtE~=AƵ��I�c��>���٬Q�Y�����ei�L����w㼞�1��~>I ?>�~Z܈�l~��PA��:w�të��Gw3"�?�Ë>xɴdp+��V��4^8E���-���	w6m����&��J,��7��J��~%qhQqJuu���-R��#����Imv�d�Y�����N�����ךR��;Ȓ�i�'p�u�R(��'B��6<����w�X��p%���6X�"��fVh'Bx�ƃ�O�Zl}�`��i��C�{jK��*�-SG�(H
�rꕭ�O�9�I<���A���
�YR!P��3V�#&���\�D$^�j�p5P⑵3��K���.�2&��75���ƪ��B�	�PW􁳣pc.����Q۬�s�/�K�]�mV��� �7*Q�Vk�&��H�f��S�Hҏ[��ٵM��߰4�O�Ϝr�	r@�������&�N���`8�I��;\$�`�"{��r�������i��3��0�����1y��Cl�������ߎx�n��A��Ъ��v��CV�q��EyE����n,L��@h���&�7�~e����S���we}���d�%���u��%x��D/T�30M���4�=�xQP�`N�̣A;1Z�"s"�OC:��[��1���,r*�HwrL�Jm���K�5�v�g�H��`�ĔҪ�]$j�B4w�X��ﭰ?nP;��0�~��r�<�6��{���,���b�A�HF�����̓���1[���������<���Qp�@+��]�|c�/�V��r�LS+~����>��aG�u	G�U��r�`6����WX
�����i��}2uJΝL�F&�4~;&�;Yc$�7"IHS~g��Q�|���[]����a�Q����0W�C���GO����<.��� y�x�zs�,����!Ml��2;4VpT�X�Z���*k�E�]0Q�M:�MB:[���?�����Ơ�]���H`��]W;��Z�@VB�:�l�cq�],rwi��l�Q:̱���E�bʀ7��Y�g���?"��o�!�%���$���^�3y/�~�o���V� �����x6f� �.(	�l���@0���,VW(��*�ɹz�
���pw�Xm�!�lvs�E�0��m?�m�z�b�s��lC���^��G���p\�ΐG�l_�%���f,_���&�G���
��߀�u����m?�'�����;�kBn��r����K���-!����aY�@��� �{��6���0,�� 8ǣ�[p�H҄=�04~��聄*1�
����7����N%$aѫ4c�߬�m�9_6��y��jo%���\o �o��.��*��:�$[�f �T?Z��Yǒ�������k�t�-?:̇ߧ�ǿ��͍����@�S#:e|������]ͫJx��0�.t|˝�g�t�A&t�8��Ӹ�y9_�TΜؐ{<>�\�n�kF�.�������:�U)������jH_F�[�ص6�������`iF�9�fD����<P�wڒᏕ�=l&���~G�rI�8��Z�����W��#�/cqD1��KMj�(��� �y]����;<}^��/�������-[���G�����[��'����^�=%�.과4�����})�/���#jY,>�PEi�sg����C`��s<?��L7��r�\^d+�$"&�80+�Y��B�Wr�w��S��n�`{�Ѳ���3�4�k�5]w���נ��7נ�%�VZn���rF�s��tC���	f���,#k�_�y(����s�܈.��}�um2�5wf~�Ҭ1{
�	���O�Lv@Q��	~��l �����L���9��=[T,_{@�HIH�\e�ő�����Ux_�ۦ�#��rb�!��0g��,���M��#,76X\��j��l��h7����4O��}P�u(���$�<f���3��u�Oұ�Ĵ~�M����pD���ӻ�C{9�(JVo����]�@]|��u��۱i�$x�����Z��=�͗#N{w'����D������ ��^�W&�T9�z#�&��-�$ p5z]	Z��!��_D���@�+nAW���̔��5)_�q\��w(��;	��|�8K��lݠ�M��z�7[zs�1��_gR��˕㏮#�8���{t�ExR�w��'5+�.^��A�97�{r�<1�ד����B���c�3B
z���VDq�.�^�iՎ�ָ�,�C+n���
	2ߒo��PJY��y����
����]�#5u���3A�"� �r���΍'�H9P������@5�]:���/6��z��EL�8����8�:|�G.�R���Sfٍ���D���W�����͛�K�'qT���d����R�`���Cʈk�y?c�D�"zȰe�l��L����C�� ȶ�A,��M��6'U����F)��!�c��#���D�W�̾��l���ž{���x�s*�2�q኏+��$�Rgd�����S��m[�"�`j��T�� AѺ�A�P&9��5��(��vR8S;={�A�M.ǝGnA���?�+L$�3K����:��Yqt0��l �����p��Aɶ7H��]��Yah�teVMGW7��r������1�{= ]A1�6�^����sQ�O]@V�;'e,���4���*̈́��[���wx�Ab����¨�>�9?���y�+Z9*���8�2���a�&���ۆ��E���*��]aF��i��}Ȋ�s@a���7�4�� �׃ڰ�+�p1��O1���{�#�� �����V ���͆�w���VG��Q?L~��ۻ��È����,c�h(�)��j�[8d��w�$@[LD�B�����2����3��#J	.,�@'�Vy�2i�G��V�.�3@�\�~�*w9����f��b�"Q��[!h���E�jT��8�՟���T�:Z����������T�A{T��$����e����h��/�%.�f"�/�G��~����Җ�����7��r?����)�6oޜ�=�u�"X��О/�щc��ˡ��tnQv�������ov��*��Y�ģ��M��`���;1e��m�*L���XO�t�橝y�J�F`$U��4Y>�m�K�K	�Á"������e����|z'��/K�:'��1�+y6�-Y4�+R/(��G1�_�>18X)A�rQ�����d6�˴7�[��8	"m�����_����r/�E��D��pRV.m퍰�v>�G�[�;3Fݵ�e$���w���� Gg�}(O��`%hs^(�;�M�a�EM�zh#%��R�@�+b���$n[O�p�M���c��L�pf\O͸����$5MC�OHÑ������	���^��`���� q����OG"ƴ�%3��?��R''���y��Բ�M��
�C�M.��\�8����ԅ����#� {��h������?�z¡Y�]$��l%1sĭh �l8�-�u&B/^�w����B
i��0��H;�F,ݣ�$r#�������[>�*�Ȃ��l� ճf�kY��'�-���K �����0��&��]t��i���\�-����Vu�K��R���=�o.]A�1�}��y"������T'��ɜ�;�?S;�b���V�S⒎`�C�:�c�ߝꣂ��O{��Y#�عs`=��������j	���?��d�N�< ��n}�I����c��#�V-�"�F�RB��k�A���6<,�-��X1��ɭ`��^.�Sq��tHe���B!
z��K!���;�<n윥U�3�(VaǚJjk�8�o^k.d��E3������,;�j�qE�Hq�����U^�1A�_�툚�^��?}����� T8����l��r)W$��e|�LW��3Q��k��r�[�ɩ���SMw�rьP7m��Ю�>�����=1@7}&g(�H����Q�?�E�h�ܚ�����ax��q��!x\���L� @���w[Bo��C�B���/�e�Jku�� �A�l���`�j�)�fV��Q6.Ɂ�`��Y؅RT�P��%���C$lI@bm��.�'�aA�6L/�`kG��`�l�<.���Uz׭>��uf_V#x�M��,��c���r��S#A��"�3بj�y����Lނ}@�pK1��L���� ��!�e�NpzKH����:�����ʘ�m�UE׊�%����'��ٺ�G�-�?��G�9�	]�U���)pO�J�!�4�`,o��3���x���7��Z��͸3�&�����QS��lc�/��Lb�iD�9̇�vj/Dr������L�\JT�JrH��.��Ta�'�%����viK]3��	@��#���~�q
s�f��7����|�J��5�x�5+�=�����mZqX���~V�hA�蠹(��(����Onc�)f�\���	�v�;��d�>��/�6I��[ޮ��v����b�^`!�� ��9p �?`i��9��5�y"9vz�%]���I�`9Y ���f�c��W�m-W�̂\⨲����,�����Z���Q����HL�w���W��2vE����r*�O��<Ĩ}�x�{U���:��&�-�ߣBl=2��n�FĻ� ���v�Ӛ�\�@@0��z�).)�*�Ѫ'�n�ȸaozr�����Ҭò�=�Q��nX��AW@�[������CR� ��졸�ҠRI�0�3�_�u��}[j�-���ƭh{�[��d��1M�6�*�,�_������ڞ�}+4F��S�jz%�{+��ě���^CH�R�@�p~����ў��P�L;�l6��ix!H�VP�y9M�3�.LxJ�ކ�3�;ϫ�
A��*/�pjQ
]�9c���1$Ǭ�s�6�&�b�'Y�J�` }	*�������D�꬈��f��!��IYԣXok���Y���Ҝ�H=a��$�o�{�J�H���~��5@�[-$�����q3'?�~@�N��/d��X�Z��3E�-��E7�O���M�(�	�Y)N!��i�W.@L��K�cI�rㅱ���ЧaL*bG;�*/����,���|��+�X�,���#x��s���?J���oI��� ��������ef��S��^5;��m߫�m�d����|H���:�PxQI�YP�ٟD�,�	EP��4�9L��(wO�sΡOo�O�FҊ]F;�{
A^G���pp��Y��iF���)-)�g&���*���NNw�t�p�A��?��v�ُ���!�J �F�|C�S�e<x�"��pNV3f�|�oD�H��Hqu��s���,�Gdij������3�ٶ I��.���
�)��x���l��ԟ��F/ƪűf���������D:��E9���k�v&H�Z��*�����e��X1��͉��H�w֍V8�Vv%S��8�+!pǩ���#��!�+xѯO݃��o�1�����-��E��m舔�PI�b��x�I�\L��	�-��<Y�c�|�\^�W6�~��V-01���1-�|��ۘ!1���Y�]<��V"�^���Eq&���%��Y^��6�xϯ�W��o�y�c��g�d�#��-~�����}�D]��<��p�:ӣW�Ab�`��g�\O�󕈢��Z�5&���+`�{2�s���
5�j����[W��p/�g���+���+�G���+�I��*�Yͦ>��*��I>�����Ǵ=��
4���(hq|��;�ot?l΍���@��@|g�G�K���qe�gPJ�,�rv��Z��
�D�/�ՙ���.�5L�;���B��Z��T걸��o�p%��2l6(7D���彜�m]h'��P��	�4����?�c��j|�2&�F���C��&�|������譹Jcf��W�FR��(��]����=��Ou�A�̦���Y,�?�Ygߙ2��FߣG�y~�aF���8�<��!� +�W��M-19�|�zů�D:�]>���I����i�S��h�Y2&�PG;�&������c)�$�A�۟�d+����2Z�Ru�(�?p�D���z�G��hJř?����W&�Q� 0�Ӧ��v2�!ftm}/�����ޖ��p^S9 Q���q�B����t���!l�a�|<C�8��R* W*���rã⢮�Sr��N��Z���8x���kt����Z[٬���8���.w�@6e����I�8C�C��M���s읶��U'>��L�	��*}�9��4o) �jb��o(���?�?��ki*X[�7~%�)�@v�� Ds�t���Az`)���P��"�ͯ{���gb)��O>八�k|�GW|��f��A�`�b���
�P������U^G��*�����+�1�����	�i�"�}'e?��| �Nʐ��c;�Q�+%/d�F/
���ϛ�r ��:L*�&�#B�����}D<m�ɦ2���E*�]���S�.+S��?P�\g�)���U�]���k+�c�N�|܅��͆�1�B2W��j&�zVļa~gf�^e=�l�����K��W��+�����r�K@W�ˊ�'���ʭ ���{��H9�	��L�b�f�2%�䬙NC#��jhl��I�N36K��R۪�^�{"�@����u�f#	�Eλ������$����:qE��P�1�y��zݡ�)Xڬ��p_�e%E�Pg�q�>�㌮l[���
�Q0�B��v�
�
Dm�*��h������=��s�^��H��|��z�c��	D���TmI����g�^滑��> <�Kyz,�4Yo�_Mq�G`O�A[�8��ܝ]F����W�Ц�{�MT�a�0�`�ɠ��J?dO�u��h*'����bf�f$�Y;!�݌ӓ������ˡ�F|�p(@ᒕ�g����Y���ś�^��s0h�`8%1���<�=��cǵ�\�>��媂�H�H�|��%q�686bl�V�:z�����HP�о�P�a���/�-A�y�$>?�o�[4s�95{%�:Ԫ��6ӌz?���t�cl%O�k/��i8\o9��b�%�;bvЯ�$\dV�BB�"�{N�Os�V:խ�\�]IҜ�cJ��ANcZ��&(/�+}o�IBx���3&�~܀v��w��c�~M�5�j {���s����|�W�b����{v�����a�n�TD��8r#��e9�@侽�[�=g��Fw��|�9���ؠ��k#xE�F~�0f�����D:�[%��G6����h~'R|=�U\�Y�X�03�3�xq>��Pӏ84�$0cl����e���*m	�fo6ф�_��D���t�>Z��l:�CRۉㄋ��;Q�6}�U��'Xg}�.�y�+h���8j���Q�~�;4D�������
_��rٯa��x|��������]}�	ÿ���$�޶��;��A�D�g�@#�p��6�vO�K�2� ��=1�� 8�:��YƧZn��¦�l;����}��W��b�͘�m�b�-h�%��o\�M��,�EP��Z,��f���p�+�{�L���-�é|��M��-ϩ��o�_]�K�� 2���7�.�U0 �;`�enq._����Ug�@?�=%K>"��L���u�`���2X5e�"�s"ۃ$�:���
��eB�vvމ��R��ͧh��n�����|�H��߅�X���.iw�˼���"`��޸.�����x�Υ��Hcо7��r_9���/�2Q[`[Y����qr�J�y+o#7���؋�������k1S4�����
GF�lk,ݱ2��� ׯ���l	5v?�,�+��ӟ���7�d�ܕ��a
�D�3��l���Y����T�W����8e?�`�D�n��v�������Z1�gI������K&i�,��<E٤��b-슩[(�>����LI�#���L�}��G��z