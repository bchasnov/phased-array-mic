��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|e����M`p�M����N��-o��i�*s�"O��@*&1��ys��5�Il����<��q��	+8jUT�c��&�%pc����C�������6ĺ�E��;s���c�Ă.��5�&7�]/�n�Au(�v�Z"��g��԰f�ϡ���K�o�ꯍ1%K'�;	V�qB�@2*Tx�&�;K��q�<g^��_D����0"����!%�.B���[��z�n�[����#���P� |�|�Ҭ���*N~�%Uf�D�<��='5�w;�u:^�g7лP�̣�R�X�l9� �!!
�V|^5�:Gy0UExE��G��w�B)Z�����/���^T]�)M�{��edL��|��)�'�d~v��9r��P.�b��BE��� �ǈ���j�@@�fq%� �n �牺%�^e�_��S��8e�@]"��b���+?��ƻ����ڣ���cd�)�^��>�h�|5׽�.��)��q� �`��]�7*��5�q�V׺�7�a����3]?W�3�AH:�CTb�k�:G��g9Ϫ<���+ϓ��5]b�q���&,��NP��S��������3�.7F�����Z��/4�3�>���n��N����Q�AUw��Nu���^�C]�Vt��j�欌q�d
JQX~{O�_��×��6�c*����b����j�*3��bU��>i�W�/?Kȇ��!s��1g�yU��Y{�ٞMc�6�Ss�A]������@�_m�0��bq�}7�py�:S�����O	��[����?���r���=���s���K���o��O&�L�׽c:��Y��� 'А	υ<��x���R���c���s�9g�|lQ�q�g
x�R9�x���A�<S�'V���߻�va6�V��h�81�m��ق[���GZE�̎�h��������`�c�����A:�Rʏ��L�*:�b�
��+��Ь���g���O�scr"�$G��M��N��;@�J�Q�������«fN"�����/T����U��e�qc�!a�»�,�~	���K���I���!�Ӗ�PWXQ�UK�v/R�y��) #_*�$1ܹR$עW3�S��6��k�c,\���L�ڣI8N�]��6z�
ӯ��.\�o���Oj�*ĵ	R��I����W3�Q�}$�|�[M�H/7tk�W�%�`�/(P������L�OLڹ���c��I9���������0�,�o��"B��c��P�����!�W�0^g�L�&r�]�
"�hy��0�؟���yS��
UV�9��c�S�R�^X��!
�AC��N(��Q~]#M�;{D��JQ���O�\�.mR�:e�1$zpo"Jz��[oQ-��P���� �a`����Q�J���{�v�� �S/�-��C;��qUF���|�*�����:�XD���G���Sd���:�-��,n�9��t$��}9ũ�*E��iԾ	��VJ�,� E���3xF�����#�K]��4�P�V������c_�wo*�jGskT�:��N�6s��8��Q��yk�� Y�������,��h2R���b�}�dxP��n-�|��h��z3�1��d�������W�O�!�P�#����]��ϿJ��k-)O�5���r�Rvc��������W��{�so|D`�.��o�����{��?�P	����Ea�Ś2�g²��	V��� k0�e�F.�s7C�p�-(;t��AfМ���|����A)��PwC�Xz1�t6m��8�҇��<^�:�y��2��qj��&�֫s���#sI39m:���_Tv�ù����8J+�:p�����,�rվ{	����P(�`M��)�%<9�LR+q�����?I�A��G`���rǔx��v�]l��@�EiH�%��M�p�O�G8i�k7�K=Ő���4����B5ھ�P'K���:�w��w��^�p��k�P��:��ݎB�Z���0��Y3"��BU{��$���qg��B@�� �K��u	|�d*�մ��YE)<W�T��~"�XxY�VI�����,ا��;�N���'��Y�~7���|-;2N<��([�4ȩ<06IP�I1Z����ٞ�Z3�X왪N��uZ7ﰂw#�ܙ�:Is�����F���1��V���0y�v�O�AO.�cx�C%A��t��yu�9oE���a+�k�X����>M d�[��y�Vs��չ�]�3�Mo�y5����VP��r�zlUG%��}��ÿё2-�A]�N^����}�?�K}�����S��\Y���C6�l���8]��7Q��K#K�ohY��F�<����(4�	�	���0?�6���-�B�����`�s.�ha���ۋD9Q��y>�����֍�dِ'����Ҋ?1L�u/��b��tv�PS��`��Wꄩ��c���&Ǐ�S�{ ?f?�p��۞�����-�w%�ڋܙD�A��7�[�j$�UӶ#ݓ�Q��H�O˲�vK�Tr��X��y�m��g<�9_|�>�0�ő�6o�S@B4]K���l�S�d����g����J���s�#�AЇT���Ze�����a�� �Ҿ�!!P�ނIj\79?�T ��W�פ~�F.�!��+y	�D^�,	cXH$j����� g?��j���:�M��!�̨@��y�ܨ����I���8l�	��F�#˔|��.GC+U�̲'%����}��%2B�M;���]��!����Q�.���U�\3@ug$�K޺��f456��w�Q(����c��!Z��i�@R-O�],���#���D�� �=GO�,)+��Ы|-3�L�/r���բ����`��&�j�p��6� e̿�[�8�Uc����Ѵ,y��M��� D����n��?\�T�*��^R�b���#��&{�����Z�M�N�&:%�!U��U8�&C�W
������CYS�Rk{��SϘ�(������n}�w5�4��ܥj,��c�{}su���D�T��q]��v�V��3M竒�c�&�/e ӵ{4�6Ô��{^��[��!�J�H�W�1�Ո��`F��iG:ʌ�����y�F�O.������[�`�(��z3PJөT�yC.~�#sҭ�F�_��h���l�#ʚ��o0�!��Sq-ኣ��) E8�jޜ|>��gw�
F�G�J}���j�Q�6ԤTf��G9	���wr��`�#+t"�*�D["��k���<����J��*'��d�0��X=R��-\s�r�;M�TC��Z�;��h��b8�[�X]5h��8�?��}5p;��f#R��,���D�w5���~�@S� ��Ң�i�S$�iȲT�U�O�F�"KFP.�͸�����C � DԊ�܅�1<ZLٶ�� �[Z��8L����9r�ՉJK�l�h�|e����{n��R���ebC��v��I�u���
+c6��;��W�������X @n��M�=���<��+�@�����D_���s`�ҷ���5��{D �Fx�n��ǝt'��VC�w�0���M���.&���Nwc������3��DXj�2�����N)I��z����3���n�y�_��X7-?<x�5�Č�y��UV)(��d�N@�"��ז��hN��a��p��{"�I$��U�4]�����l c��O:�V�۳��t�\}Z�I�����u @�;wA��d_�v-`ٔ� ���ה)X[bx����9,������5�r�c4S�Pj�j�����=J3bd��rԄĀ�d$#fxt<�V4�kf�Vg��/�?�l����%kJh2|�<f��$S��{��Q�I���Bt���`�77̟��Z���\I����J]���,P��r6��q�I��q&��o�P&����Q3�0�࿸D� ����B� �3	�6"U�M�dĽ�LH��Amp�ڬ��u��R@1��8	zrG�y�! ���ݵ}ķ,�0�Uk�1۬-��`���/�q�-f(�\��$*�;����ն6<u\����k�����~��0�$��~�G/BJ�g��1���`�\�%�c��xN��� @=��V>O0�2��m�Ӆ6�\~ݯ_��NUq���`cc����d��}�n��5d7��*,�����j�ӟ�H�YV%�9�X��ҫ}82�s�ūޮ6�J���ƍ�͡iSclظ�J�jv���i�8�c5����:�r��`[���k�k�����1��г2��;���g)1�����廇�NHX���a꿝[�$��� э�?��A���U���N;a��d���b��ȯ��	�}ZVI�{y5��>�x�i�Go����D`�\.C���ڊ�9��r�,}�Դ'uw�J��R��]R��Y�
�(���h�V���[WeY�)AWCB�v�3��>U� #����EvxiWY25xp ��${G����}�/L��}�������ۂ|s�p�ݳ���wlT�����뿧f<6�ir%�{w�[�dn��A~rC�n�� ��l�����Ud�
�F��_�$s�^|�<�e�/ۜ���/R����fW�+b�r0����Z�o6���%�f�޼��qB1� $�:����D%�rn�<�Q�7��/�2�}ѧ�G�/ ����uv��r�\�:���p����LN�]� X7�O}��J>k^�q��vD���#���6*x�բ�)�Q�=d�<u"u�G�Uw�ԉ`"g�GN������uBC��� Zwj�AH��`�R����0Z=6>c�2��������Et��z�f�z�4:��6F��C�ق�%=gb����E�jԜ�xI�b�%��%v������/���D�c��E; �^}EE+������3�b�xE����+n~�S� \?��3̿)��=��B@zi��c6�M����-���fW�1CJ�Qѷ{�8�6C�e�c^���_���)r�"�bf��C�$A�̪�.GM-�!�՛@-�-:����ju%#�Ǧ����s�x�A�݀A��{[���3��_G��~��Z�؜��&�Ί��0�E�s-�d(>���Zv\���R7����Y�|{����-�h�4�D� ϴoL���
�K:<�Tu�t�#�/��ʷ���z����X����!L����v��(3u ���
����]w5'��E:> ���	[_�d�2���z_��C�r|� T�'����EC���r2e���G�����+F��=�k�����$��J�3�/f��«I�,���e��m�{CՊ�82�ӗ��0\��Awj�(-EXa�̻��L��K}���H�1x0�P=��ѹT{�"�h-���O4$�y�9c��a�������)���,�:ʣ�^*������������Ŏ�?�)7p*O��j���q�m��e�K�8�Ba�g�{�1͐���3��(�1��O�ձBKi�{GO2LP_�n�1��F2�;k�ʩ��X��i�a:��f g?�~�8�~�͠B������&�6*�!��.������7a�U:��E�_}v4�Hͩ����HU�X�+Y��S��v)rT�S��ZB��_�O'�V#{505�^h�GV���	�e���:���<��esG~���Q�Uz0�R=���X�:&���ӣP*��E�, `տ�P���:�o�u�v&R��$NrYg�������mo$���b�+&���E]���G^���-�ʙ��Բ2���G��=� C�\Ĕp�����ѽ��5s��o��'�}��[a�-���;MBV�O��0HD��{ϽPj伭�TrP沕$���穸����7���KF����{Z��o|�RE$,���3��1��5���K=��������9�6C���y��*��o
�o\+ �k�s�����X��>n�;��|ɺ�h��l4�R�� Kۢ�' ���i���i�<�7q��ΰ�У��&%�n��6R��r)L��h��,�J=$����.���y����CJ@�N�5ǲ�pR��o\$f�0���OKO�+)�Ɲ����E�c�C�«���;Aa��v��h)Y*�Ҥ�w�d�wI�
�Q���6�W��u�SnN[�����nE4ӂu9�i�-�]S�~��WJ�������D#�w����60ldU��5N�����H�a@ ����yw��jX��-4�r�*\n�[T���g����?���gv$���F�ær��6Fq	g�JFLJ����r\��Q$�B���$�{������Pxq>q3J���q`�m�'��TR���@^����#��bn��;�P�*��,�e��
	��$�q#�식�<�ڵ�fg'�6xn�"���9U������9�L
Æإi�7\��v0�>�|en���PU�����/�l������8���B���w�7��L��72�����в���<$�A���H��cg��9������.(����s-��P��k�iy'�ob��݋Y+Z>7��:} �t�M��C���m��r]G*WQ ������cWDI�һ�����0"����һ��r�1u�v���/m��<3�~��|�y�t��9�(5[�<s$hۻ#�#Dp�F�"rW:�r=�స�����b*F<�Os�L�ОR �U�I�**�Qz �ݳh|�s���`E ���+�ݞ�Sw�Aڿ�-�.)i�T]=��v�k�F�K�f*E}����¢�u
���R��Q��@�)%���q�ty�Ϊ��t��sKA`o�����ō��g�A����,ӛ��a)O�hg���V[d�n����x^g-JC�׮�Tǅ��k�-�'�xMϏ2:Qàp��OA���*t�Lͽ����6��紉��m��?	ōy�52.S9Z��q���9c$c�q���SU6t�7Z�LtՔE�N�X=Ry�� �z�~��e���2ܿ8�A �
�" eⓢ�L�ц�|���^�5�W�>�(�c	h"x�[:�n�}���᧫*Ġؤ��O*wq�r��'c,v
ܗ�mzy���������K��k��+٣? H�h�ui��H��)k��3y��U��ރ�`@��(����-6�k���^w�ᘏ�]�:�j��W�a}g!`n	�mYIx'�m��P(�q��+������k �������?���6&D�{}��2���*�ibOA9&�v�Y�@�B�y,���]��5<b����)�*Z(Gd��@�����I��{��Bi��a4e����9��'�>
p�w����ⓟ5>gi�7�+���_v\;�X��]�Y�� �Ҵ�����4��ru�/�p#�1�ש��ȏ�yE�Y�c�ۭ	^���V����Oel�G'�\�B��&$�/���{a�\i��L��#T���ko��N��f�Af��{�߈q4���!�0[��6##ܭU|T���y���T�ipc�Չ���Á0҉ҏ߿��_ܐYr���rZo��6,������A���-�OyR��n����,�l��l񲑖k*���̒��2MTgDoX����"��Y��6��%<�B;D�+nO���dK�+�_��x������Z�\�����uTV�y�ԭTH�j���֒���f�r7�#Uhct@/`;�ûojX�P�
�?2EJ����SW5'���ouDM v;�kD �^|���D���>-�c�� K1�����e�s;)��;]��X�l��y�yza9p��ubq��s!�o."��W�bS�f6�z����$'#�BfƪV%��c6!��nl?�UT�%3�UݙA���F|��I�MF5�ťT;��h��}���wJ���$�귌}����f�kR"�0������1��4C-�׵��n'C�yUyI��� h[!ZΓ~�.�� � �|+�؞k��c:��`\��'����e��?g�����q@hr�^����Y�}�N��to`��E<�"ȍ��VЂw�+�Cj }���&砩�1$�k�e~s8�0
��Ǚs��Ŵ��3�T<�m����	����a%K�3�ʄ ���󅛺���дo=�u%`P�o�v�jw��"��R���FU���9	��.��iW�0uh��{��7 RV�vS�>��`�޷^�\ˇ�Rz��!*���jm��O�����rc�soQNw�/f�s�O���4>d���GnM}�ʸ�j��2�M0���������d=��O=�ne<����Q�����{�˷�,��+��ִ:�7��.吾-r��[�je�MC`w��G>�OM� E�5a����V����2�����?'�X-=���~���������'֖H+�q �~%Ǐ��3N���4S،z��D@��B�Z�f@F)a:�N�ʆ������c�!����w��ѣ�"�O�<��?��T��3��u��c����e�L�d��W[nĞcMj������3�-�a�.�[xr�?�����I�钯̀6o�����j�E.oyy�.�lo�1�H}B�������+��p�5y+��৛�����=� ^��� ���S;s��,������	2-C"�,���W����&Մ5gѶ{ dOri�$U��#t=���ʤؑ�u��-<�B���av(���*��dJ�� {L�UP�[ ~��s�6�8�Q�@�ͥ.k03��Ƕ��Vn�/���Q��O��@�ܛ�ٯ=8;�T����$�4�2-@1�D�Dǫ���R�����2��?^O�2�� $��a�Y�6_vCk�����C�ďυ���C�O7�g]��{��E":���@��}_;�uEx��#),���Z"��A�?�*Al/�����$�)L�H��S�bHvg޸kB�ŝ���c����TR�h�j�����Y�E;�;d��24�f���W�FOB^��?�AXdҜ�q���a���q��ȴ�����/�/�3}ὨB&R����J'C`�-�Ǿ�%��/������:�o2�cC��ir���EZ�l��Ed�T�+�k����r�&|;8m�{��������C�ÍgWJ�'�������( |d�ݚ${.���x��a�������=f7T�����M��`P��B�c�V��'�I�m�b��=�p�(�-jTsh%���q����VnnP��>����l>C(�eW7-d'���V`�D��DRwIp��0�};CСpl�ΈZ�7�o�z^5�����f
�+�5�ETWb�A����)ۜB�Wgm��dav5�%ƶM`�g
�cm��X���Ci�W^,�t�+9akٷ�g�c���P��3�ikk"���L	pי�I}%���Re	�E@5�L�8�_�ɃS5ł�r�:�������E��d�q�|�J.���<�\�W�.�%:=�cAP�Ѓ�B^��[�y�FԖ�z�Nذ�r��ἴ���#*����t\(g�	���}������O��41�B�*M8<0�$v�.�?zE��kT��+�'ai��٣�"X�S��ث���:�f�w��˸�wC
5��_O����޴��yِ�k�~���#�Ь���G1we��`"`Uqc@�̆�
�GK��R>�7Č"�r�6�1�ުF1ԉ��L?�j�4na�˭=L�ݕj�HAMW�|?Xf���y��_G���b{|�8��g=�kTE}b����nM~�)�A)�B}��|�ip}�ܙ���{W�ܛ��!P+t=�B�
��ۖ����/���G3l���fG* �khf�u�OhRAiHF���e<��L��Y+�x<H���h&?Lv��
����h&�j���?l4@y#������qFٵ����Qk9��i1�k�n6�Q�����Ct܆��F��.!����Q�*��\8�ly��_�=��^����S�	�T[���cpaՉR��%�Q{#���qSF�ϒ��k��yǬ9~�j��nzU���)ZM,��7cs��f���u��Mg���c��By�Կ��P��u0ƨ	��h�]��x��Y�#���}R��=�����ߦ
ËM ��Wp�pT}nE]y��˷-����y���h� �B���羂�{�ߣ�Be�o��G.�vS;�R���0�>�4#I��v�S�k��P����>h��ܨ񺤡�y�l�A����lag�����#Q>��:$l�F��}0ǻ�]��nƅ;#���|����[Žy�������'�� ����m6K&FHBR�:�0���~Y���nx�`UJL��&��Ne���	�@o��5P �ps9vL�Sk-md#���6��\��ў��~~*yx,������Ov8BG*аg�`�B�?Y��'>No0?��3�2��8\��24�a��.��un��?��cKGa�:�}ǝ��9�o)�1�m���~j+�	��#�^T%�yrا(�9��KXS��e�`,�<�QfB��{q���T=�c��������J����<��5���`�f���^��f��Vr�#z�Y/@')��PV�|}�p�P[�NC>��-/�i,��.ὓ�ql��#/����;��I}��L�=wy���_��Z���#b�T������Q7���Ɇ�m��@�����l_,�1�E�~!�����BF�\`]iseM�6�i�� ���~���qa5�x��|�1��JS'�V�r](���7�,��~��,�[	���֫����ز��U�a01�U����\d|�?�o�P"ӪffW� � �/lZd�y1]iD(�E=ͻ���Sؤ����K|�~e�»���5�f�WZ�j��+�;1���Yx����jA(¸�b��L�B�J�-�׈ù������4A~?�wW՞*8�V�-&����j��g�H�;�MԤ��z�>���@�E$Ndկ��k,[��x꓄$17U,��`ͺ�p��J��ÿdN��`.�8�3����WXʇ磦��Hr�I�<�����m'�F�*����{!XRг�_����Ҷ�x�Sz�,S�6�k���#�r�� �"�v6u]�����s����)_��kߏ9^<	��������6��\����g�H3 ڄL�{*MV�s���/uE.��ಀ��K��	1W��L �O:&a��8���Ar&���W�y&q\�WC����LO����F���U(L ����6*���Sן2wx�]�RZ�	Ӭ_�큠Rɚ�Nk���]Y��c��,�" n�x�ڜD$��,�S轳�(�^�@֞��xm���F�ȥ3��ɺ����e0D���� ��)5� 6.u�4;\�C�"�l쉱�X]O�0������e��&�3���^봎��^�8���R���9c����h���#p�ʚ΍M��@;�YL��#_7�n�^�(�`X��5 We�(Q�T��|���`|k�. �"�g5ǖ��T�p7��=~�Sr�o�����B`�������~uP���adWS��&bY��a�h�5���Z�Hv�C�H�3����Q�Qz��:ʤ��U�����'^bD�"� �(�*p�0��
 ��'T�����3����]t�\������"�|*��Ly�$v��,�!r.<^ ��NwH��;D�����HO<�Y�x���M��wKh[?�����7̙�����%+�|Y@�������Ū7L$������4\h�"��;�8b��2d��݃Y�#Iؖ�N�q˃�05�ɨT�p�]ߍ��KN��� ���]�w�c���5]�)š;�B��T�_���_�@�P'�����#p[�_�F�M�[�:���H���1��m��9�M����G��ݕ��I��r���u���X���S����>{�h���5�˴�6Ph7fQ��g_7f9�����``yS��N��JץX�W�H�NPj���ȣ2��iw�(�=�����Kg���6����}���j���4�A����jl�-�S ���������-�|�.�!�Xyi"[4-ºd���n�Yc�Z-�︢�����" ':wOH�-ȬŁf�.��y��"��y+��ܳu5�Iù�Y���atj��x�se�&�u2R#}� E�Е�0T��#/^�����vw��I�CAfB��b������_	���V�h�L�X����:���D��%��<�����m��s-�eJMϷ?���<`g������<-�-(�>�#�]�탞�4�����Bο����&~�(��2�sR��EDY��T��*$z�� ����lon c���6����W�7��߾�y����k�Uk���X���x�
*´/$��'׺!P5ݬ[�R�/D�a���[K|����wD�[�4n|;�f4��/��6p��-�Θbȍ@G�)d�+I"4����ne�,��B���ލ���:���4�|�M����Hz������P���+�΅�8�n٬A�R����*��r�w�H�F�W�Qŀ�PE=u
.�S3�"�8h��V�|�)gm�5�O���>.=�U�>\�����-THw��jQ�J轒1&�17�o�n��^B�ć�k4�H�0':��l���7���J8^Z�&�ڡn~�Ac�ccӧ��l��+W,?�kE6}շ@~��ΟG(2�Qm�2
���d�t������zP��Z�^���n�S���RQ�P�����]���~��V�F�~��P�������==���A�'��6�~[(�ibD ֖���)�oE�s=��-RH�G$
�v��H�h�_/�R����3])B_؂��%�90N�#�$L�����?����J��Fk�6��Q�d&ﮫ�}�9ċ���s<�7G��h�����Ǆ�֥6�k��I3-7�s #���KD��R��y��-Q���lC���'7�.<��-l�: q�ı� �bd
�j�ڞS����Q�]p셒����&_#Gw?�����1�]׽�X�\[��1�́���F����~�d�Za���Ku0%URCG����HI�X�%��e&�	����Fޡ�;G�����w�!y7�^�
��>HT����*VEÐ��ZZ� B֗C�����dz҃?LT�EC�ޚ}g�bz�yeLN�mDO-Cڽs�ki�^˧0���`�3<�(��8K���r�4���x�ۼ;���N�m�	��_V��=�emZ�a]VFM�l��e�$��<`�zv-Q�C�)�덥�d��pv��	����eD0���Љ�J\��	����`O���饧ekW�oL����)�����J�&�G�2ap��Ң�7���&'u<I�	�tK�,KR�F�I�B>�~CZHH�b�݊hP?���(���츸y֭msc������.Jm�:19��ТDW@	�7eʓ�!�+p-ˉv޳r �~=�> �Y�Y��%䏪�I�8P��&ńX��*�''J������Zf�?_4�������J�N��'��m+��=B��`��*"�Z��^0��@�|�B�+Y9 �W�&	X��a�*R&pg�S����Y���_�/R�S1ߢ3L&�E�D�2AsmY����H��gOc���1fy�C}ww�s�8�M��˅l�T��5[f��c���{����<]ߦȣ��#��Jw��jc�&��kMu�j�43�����vc`bf-��9����6��|FM�􄋱��7(�"�������������_�!�S�;4�Ygq�C%	@3��?��k�Hd����
�۹R�~5�=�\5�ŝ�(�����"͏sBI�S�_Izw���&v�.[��<F:���z���/�d�Vy��SS�ט`d<���I ;�)��:$Z�w�k�C:�5�J����T�p���oY\�����kv=�����i�޲���Z��ZN����_ILDe�H[(��a��GO�9i��v�w�����w Ռ>.`���Z:���?�}dO�lذK�Yz��?F��t���P�)�RN*�ǋ�Cy�����_��.����A'|�����do�	��f�o��"��d����Uc���?8�%Aė/�[���3�>��0�:˾�Ӡ}
�����e�!pCv�u0��>�+�qs��mv5�5h���* RJ
Pm�D�d��l`(kP���q�ȧ��5`:jh_��-#�:��X#>�X;�-�%���n�,x��xB6`�����E����4���Y6����R�#��ǙY-rx�{+���fy�lDI�Zބ�5�	�M��Z�W���mE��t�댚��g����I��Ow{.�&�0�O��2�mG��Q;y��2@�4�L�O�tR��_ �x3d��@�MVM��Pen��3�*�͡��i\��&�zk�M@�#�W&N,F{�չ��F5OQ#��q�2	�>*�
��~����-�j��0 x�&�k�T������k+T�Ꞩg�=�X�����0r����~Ć�8��h�߮�����z>�p7�[Q鷮�f^�]�t�g�#q=1&r�h����X�^�mUi�-����"}�`#���F�U%��~�m�z�a�Գu
�:f���5���#�:B*F������o��OR}�P�T�5u�p��
9�X���G@�K&���a��~T�A��4�5ǌ��d$�.�)$�Eӳ�T��t���[����!��+<k/�2]]#�+��Fc�h�?�����O~I�֭|L�n��)�bтK�"N�]~�  o�S����#3gٰ^�im��﵌�O���Ee��@X��Dc�?�	40w�����cal��%t��xfE�_0M	�/������!k���uz�M Tk�:R��QB����꨷� H�9�L��a�F�(��&*:�T6��[�=�3ܱ�S�|m�j��2|bZ6���S�Ԃ�R�TZ��c�>����_�!Q���*�z����2m�Z��g�^�L�p{��p���xT�Vp���e�!l��[	mn5Ɔ���b�e~}��յ�J}���ź�GQ;a�2b�Y��F(�2�s��*��x����q3�S�|\�䌝�G�+i�$иTz4ߊ�s�z�	�a��'rv@�[FD��������ﮭ���\j)�-*7gL��K
o�l����KV [f��� ��mf���s�� C�-T;���[�P�1U�|�vҿ�ƥz�E,�6� �%N�����7D�}qΠO�K?�V_��E�+h�]+�@
����*v�������?
��H˟`x�r�,����y�1�c������V
Ϩ�r�j���1۬��ww�[N�9E�Z�J1X��4�LyȬ{璕֭
��� ��wҿ�Uί3o}�߉�K�j9~��
r?���
3*?��Wu"��9�xW��p������S�a���LUtߓlb��L�tb���Q���O�3�`3oM0�gyh�֟w�K�ȼ<l8����}���A]r�����}�T���-�ZB��j�jך��h�p8�3  �њC����,kf:���SLlSq��]�y�`~%6��%�g_�a���;�P���B��V�03�`�
ԁ�	�D�Rh��4)ƫ�P�o��UKpſcX< B��˻�i�:ە�.>5�@�ZՄB���[� ��UG���'H�ܺ�C�N��g�?}�jTɵ��L��Sy#c�h��D/۫�ӥ����Ab��u��'z��r��ͦ ���{��h�P�o��p��,%�j4W���;�	���G��z9>">p�����y�8C��c\�~z^C��݅�9�z��I�ݝ��"��?�� �Z����_���QnzOb�.v��.�u��l��z���N�Y �@pQ�zz��t�c����dOޝ�/��`����YO-&or�%�t�@?c_���B� �rq�y��^b��Eq
����$�b�y)�V]XS.Zɭw��EƷw����p�,Ol�͈ɥ������*����b�,}ԙw(��N2�-�Q{�*���$�R�[Ϝ�NTp)�(� ��>r�>�S�6ti&s ��A���EY�-����1�ٸ��ϑ����M��fx`u���H.�s�������}ºښۋ��:��S�Է��U�ᱷ�+z�P+�Dp}e�<��U�hν��M�5��#5���l�gH��xU�%�@��^i��?�W���L�w49�6�)9��@�c�3&���VT��?��}�r@E�����U�u�Ik�#a&al�w\Xb���[�O޴�?�A�rv�w��f��[���Z "��8�>�K��g6O��w�H��bIE����Yf(� ��|��O���wA9߾�
2��+�'�졏����)ۄBd��dR9l2'�}	��ܺF��`� ���<��I�s3�7rT_�k������k�US���Uv:%G�%��6^��7ү�߾J"u{������F^��*�����L �P�S��@DE���&g��Q�ػ���
����@�Eb?�����oæJ�'��Z��j�.�%偦U�*[g
���Ⱥ�\��q�i��23t���P����F3K��x1
֌�QSK1J�z]NKw,Q�=A�� O0-�
s�����$l�T���1� �q����� y��ۣy?g�#�g;c�`or�?N��Z��M����(�����S6KBk�b��`��8p{]3cM /�mk��h>ؐ�2$�f��A�$ 7)�\�pm���'֏&�}VY���.��j�4f��KQjo��ڹ,�?�7�P���D�^q�'��7!��ۙ�)�/ƺv+p���5`L�>S��0 ��L��N��H�y|�6����/zv��E�6�Gd��r��sΤG�'�(m�~���2m��@�@X�8B@��l�w�9O��ed��FC�/٦`*�����/v�y��~�#̅X�]�"d� �l��W=(��G'+�|��v��5�t܏C�%�f�3�����
$k7��\L�G��P��[���
��MU|JBF���6�-:Sg6��ө��0�e/���
�kY���o}��[?���7pe�o5O����~���W:��HKD,!8�va��U���Tm����-�u���!�&�F@��'�TAq�ޢ~pW�׀�O;RȤ��8�:��
K�r+��'Ts������N܋U�/
���ȥ:ہey} ��c��r��ˮпQ�kt��HO�m&�j'��
��PH�X5 �_J�x��R;�8��Ys5+�󡮩,�����,p��Е�ߵb�+�	Cz�7�eZ	s;�'��)w�����~i�!�<�]ҹ<�5ޢIvL���b����(0�h]U�޸(��QOk�jc>��K\�-H�ϐ�"Ud�Q��i؅�HQ�g��D��D�'�5�+�^SHh>N���e��1T#�ŢaC&2��}���VK���	������ύ�I!���!�뢁���Zt�e�X�I�^�"�~�-⴨�s��q�X�n�%	�������-�\O+���H�m�xE��Mx��� 8��Ғĥ	%�ҧ�v�n�I�*2+C�v�,5SjW�G�`Rb��n~X	×t�\P��^X�3�;�*�K��9��PG%U�X.�5R�_�s*Y �P��r���Z�`��
�P�`�Ч^�m�.�*��Jf��n��jE��V)�m%�$Y�o}�����B8f�z�IF���[؅�qL�`�tcDKN�76�z�S��ʛ�Wլ޳��X�"��d�3���4N�}�1PJEvf�����T����Q�AP*X��b��L�&\ә���6���n�0�<M��<�O9=v>�ϰ���J�x�λ�li->ǟak��?gf~}A@��W��k�}dZ��U�އ$]w���E�P�w#�3/mf1l��͎�*�ej����!{{rޘE��^�C7����D�f��<<�=/smHi�������$H׋�u�e�'�c�m��x7�=�8�m���XX4Ͷ�F���u����vS���I��+�Ho.��*�OQ�ka1��b柂Ԛ�����Z�Z^���YZ�{�	I9VvX�0�dU�td%�S6�
O�����Ǹ��
�NJ�����\�������ݒ�Ǎ���+�����7r>|�rOkZ%�	K����;����l��Ɠ�G����	���˵�0�"�Kӆ�#"C8��4��!Gs��!�eN�_�2�创��/K&tei�.�f����IB�fո�h��10�z}2�n=�b�>��3l� Q�����C|Tc����jK=�ޕ~�{c�z<2�La��[�eR9�s����L5�S0C�ۑdrE�,����)�"���X���X�h{%��_:!�U�f�r{nY	��A�݂'JQ���rP���_��0��$銱�s���RTt=�iQ��?�;��=����4�,��Q��sN�LD��8Y�;L>[�,�"B3�9O��~�N�L˞޴�}�3K[fDe��3zL�� ��Hj�� ��v�$�;���T��"�yrmTuX3�4a�������;`��Nn�@��nk��v{0/���V9�R��P�I��;��fl.Fe
�V���>߮�������k���<�w��S,v�*�=�[^8s�$���ɳ�Ʌp���(���,I_8���r5�v�A4�����(/5	�HG)��7<FOc�L�f�"B/�����S���7������Bvxf�ƣ�2�[.��]\P�a�O�fd� 3{Y�7`U~�JG������	�Ry�匠7�b��c����R�6�{�8���<���
Y]����}�+y�����a�U o���B���晆 n^��އ�N(6]�Ɣ#��*�#|KIPV� ��"��î�[�G���(sD*?�ʇ��"h�8����/�K�ԩ���j���)u�c����r�p�,/�����ά�:y���i��[l��cˏ�w�܂GM<�K�w�OLjD����&M����l�r5��' �~u�謂n�T�}D3�B5�~-�D�V �J�/�p.�py&�qC'��`��L.EUZ5CӰ�"��{��"��k9�T������J��r�۟
�+{�I2��2���6�8�"������ z'�K��퍾�	5�o9�pt筵f�'�bŕ<�(E��j����UVl)���_l^^��� 㑌���]�Wڔ%���)Iu 	���x��~����=��_&�!�&��lI�v:n�B�%���a�)^��!�GS�x��(K~.M&]l�+�q�D��q�rպ�Pٻ�P�o�����(���=>���!?���]�:܄����Ր���
��Br�S���}�a��4���&��_B���~�(ԶX��4�oOGKɪm�%+$j�T������_}�-i6�]N"'��^C���Ex	X�a6�r�9(����8��\	��כ��ig��Q�ы��=tSذ��[L���ixj˰$���T�'a�n�o�u�iB���6�#ݶ�r��ޙ�
$�\eNg��c�3<�ek�E��L-v�����4�X��^B.ֽ�J�R��f��ٲ%�)��k̕���8�
;�z��v��ʯ	HB����+O��N&�W��&�<w�,�D��)�uҦ��VH��e���ԣ_��;�
��;���Ⱥ/�*�ֵ`�����e�y�=-���WP6���L]#�����S���B�uI�[S+���s�ɄT��1� �m�{B K�9�c1��=�ٟԴcc*�'܈�s��
_�<ޘ��Ot<7,��E�X�X�(��<��V��'8���с�+Y��*�)�-;H�t�k��L?2h[�?���K���yj3��S7
޺'LI9��S���$H�6��̂����9K �8��?����1�v?{p��)��ۈ"����I�nr}@J�d�,WD%����L7��s��+�&c����-�c��5���3�_�s<:I0ϟ^��������Tp	��㙗���!�[���>��8�b�r�S����`E���n��,��`�d%#!Q��+B�I=0ݟe�S��Y�$o��d��4͌萖?�ѬS�!�	�ʵ89?��*M���)�6GT��9����RuL��
gS��_u�C�sv�<(0��\��ď?��2N;d��:8�c9�T��94�pJ�z���v���o��s��00��b�o�TGX祹 soe�P��,�Z�lU��?؃�=X���!{Zt�Epd=m�r�`����m��\Ӱ�? �_�8����IA1���UF�2KQ�*�0;�n�+r�y�����d�(.��q#��n���}�SYhE�BxL��A�o-TVÜ����	n�g�Q�ן���n��"0<��Pw�͂��yHP~TTl	�>9- #y�f��TVSѿq"�`�oU�,\�6�*���+���s�?��[�e	"�-ٯ�)�|1���'c�l�#�q�RU5��"�vbs�sL]�z"�4`q^y�@.�)�.[�h:���0yOv�(bx*�vj/S����[�?ֲ�؅�T�~`�(�e~��V����v��ϓ|(�S:2�p��bK^�8f$��tx�A��Ǔ�7��}���״E�������Qf��� M�F�KHB�[�,~�qf=r�(D[4.�f��9h@>)w�&��=��%@m=�%�O���s;. �kE����Ϣ�j2�㒶q]��s�5����{0���5=B��k�}�T�ۼ��U׭D�J�KZX8�$HN�%�e0�����{�:�j�J��z;�zO*~Kv�W� d
�p�z��{@F3��E�O�C��v����七K/����<3�]�����/��_��l��r$S����Fy��M�}�_��.Ԝ�-�7�3� J�:�	z�'�80��gq�
&���M-�� ù>&�Qzǌs��I_Z�O�H�<6qqPϊ�c<.҃GU]�m���r$�⧉�	�n\�����[��l��e
r���k���m��D���
{��z\�I���2w��p���J���ܷ)���]�fF�Nd8tF���7�
x��6K�Т���q�	]P��<1	�L�!�I%AAcLm�|	�'��٥�G�����y��k���3Zj�&���	(W�|X��J�(���ްF�U�E@<���[ڥ��s�s|�"@
�n8�ru˯$j����P��L�IEK�O���ɿG�S�������{3Y0� #5� �����B�ntL��S��k_3�#e�u�U7,����ljN�������#�D^��|���J�o��s4��g�6�x%QQ�b��w
22��~}�<!�����e}���H8�(�-"j?ed?����g�b�`|����͢��#?r���D�ݶ'>�m!�*�aj���ȂK!�5��7w&՟���!��R�,PW��H8.5dSh�r>���vc����K^�'a�9��)��<\���l���T�x<�xR"�S4���BI�H��(}C��� ���X���w�,�����O��+��I�Q��G�:f����Ey�������l�/k�J���~)݃��eև��],7� �>=�ܷe����wh�)M4�c�#�ǰL��F�'���1��/vH�t�/J�P�''�Z�q4Q��z4�u��_���ѷ44��@��R����p�K��p�Z����	[�h����vǀ?�Q`��Iem����ݚ�׀Ccl܀�2l�
��v��d��x�{�؂?�)�+Ko"9 �AUѮ�Cb�#_,���8����Y�ڹ�JK��3~����F�.bq���9+7�I�fݲ�����+�����h���d�}��=R��O�d���1G��[�`�\��0�6�bd�p��M��mO�NHPê�j��|Qaz��a���t6E��C�����q%�%Q��U�Ժ�B�+�<b��N�z_"�h������ᙠ��}V́x��G��0�z�7^,�2?#P��]mF���Δ{��k�4�s9*X�YQ	+8Yx��r@̀N��2AE_�ɚ�la6.Z����u��C��S<W�*�RX��nP�oW*;̎��4z�w���Tl��9��`�X�q)؅F��LΜlԉև��X$X�+m/?|�-bsL������v�M������D�g^�:���4�n�	��\�{w�[��E���jB�m���Juq�n�p\T������a���u�{�Z��stD���84`r�MJM����yW��yu�����ȼ��_������3�}AT\�b��������?��|�'[��|�
 ��G�@�rqv����^�ͽbs�Āx�h_,$�;��G]�jڼY�?�N�$�����H+Ԯ�A�ICa��Z������j��Ո��5��;l��|�X���jeGb�.�{����8Y�t�s����6��0���< �Z���	9������T���`��?֑��~�y7�"���]S#�w�d��YvP�E���<����l�u>=�J�we�'����f�/�}�s�O}v��H<(f�(4t|���C��c�ߞzC����Z5�-�^�v�/�%�b���s^���?y�7K�"iv�}+)�E-'Ȗ���5i���	��$�<�`r*�L�З�_C�c��+! �u�7γ ی�_ө^&p�0d�
G���&j��qkp�����l���+�[w;�9 !iOK���j!�?�wx�w�(�,�v�J�O��
/b�:�_�����vA&W���s���-�kk��l��%����O��<\����4g�c��]�(7H$R�m���h���#,�&��C� �vʼY'�ğ��\��ͺ /�-
D��Q
�q�ѳ�A-X�w`��|w{�v����f �a�U!v�?5�S�3�(ZH��_-���k_�WY�b,^"^������[z�b�@TGLG]�{9�~�-�0]�J�w�s�E�]����a���/�(��|��8�4蛐�У�"�8�SQA��,�,G�'���߱��v
<�bC��?�W����r�.D<򵾣���6S*4%dY�F��:[���&�[�14{h�Q�>'M!�Yme�I��ርXb��"(��E���k*��^(���jں0�<o���pg�I/�&[��cs�����?N���R}y� r��Nqa/�sE5�Y�R��Ʒ�(x���j�׻��&�K� *Y�Fϡ���P0�<5rf1>��I�ĥ��i`�qL���'��F���"x(}�����%� F�}����O���1��"���J��(`���n[7�y�[�U:��L�	7.��Rۖ�O"��Ñ��\�$��4J�_��m[�K|�ћ䏅�O����l����4͇l���q+qDSu,�q�i�SBZC'��!)M]��y�:����ݣ/}��L�׹�lQT�#\��_kQ`��>O�(ؕB3�R	�IKu��m�mr��vo�����p����0bbC���G'�E��&�I��QN���� B��nB=�Ւ[��w���x���xV�1� �!�U��/��&�;��Wc�P�o��S���E
B
�BKB����v�K��;�������0_eq'R���!H���K�0B�MW���s�!p�Jʚ�(g"}�A�Ĝ�7�������ݽCNvZ�Kl���{���~,���sa �;��6Q���n��]�?[��L�MQN4m<�O���}+��ByjQ���0�6XJ(([W�y��6C���2�>]�V>;ZC./e��b��+��SҎ�J]�F$9�?�F�A�E�f�s�7�!�뛆���ea%��LY�,:%�k��\n^���<G�C����Rj4��Y�`��`��=]c��P:��1njƋSpLۆ��T��UϹA)�QYfg>�[Q�B�Vݱ���2��e�z�ǆ���x��n��ŠR�	�22�I:f�F�T`����56A��X�bG��}�.�^�%��/e���0�EZ��ֵ��|ߙt4�Axx���
�NS?3�G'D�!H���ju��P�H!��Mo��g(�~�\Ι�{0�
�[->�Ĳ��Or�mq��U��zc�$��/QS/�7���a�4.Vc�Y���K"rm<5�4=f��k��L�]�<R��4��͠a^f�݅'�l��(��&�U��=�F� ��EZO��;�I!�jh�E����&�7����0rQ8�Hє0��=ځ,ǒ�/�#�eBU�G��-Y ����硠�x���Y�ˤ��5��U{�<9��(�q�f�(���-�����̀�4n�J�l��Y�ϣ�c>Si� |1�1 �����gH7�Qg�U�AcVά�o��
��n�?j�]��NcՕo/[R�p��ZV�$}��iC�at���u��4Z�tk>9�^7�\��7�Gs���q#�&#Ϡ��:p�
��x�/���ew8���3)�B�jCIܓ m�'R�Ɓ���L�T0��ޯ>�������{HT��d���6�<̴O�^4����>�)R1��YGH��E�V���Ц��8L��lZ�9�$�������e���� 똎��ޠ��r��"�Vuߒ�tS.0�3 	�5&�fk�D8�&b�6�9ҙY��[ı��ޤ�q�[���`�r�/�=��!ZX`U�Z]_�惮3�}7P�7���|�3M�D�=���)G�A�y�����k�\bW��S:�{�`ߗrCrͶ�� ��o?�&s6�������{�� ���� ⤆x�bM�F�L1�^|a��gv_�i��3;"�ra�K�a�����6�(��W��o�Ǫ�-�-'�D�f���,���!xX����@Bh�R��
�{7�"x�9�y��W��y�EW���,�fE�.��j"vP����U~y?h����j��C��6���q�	��a�;SO�q��� �����<�J��j���a��*�jR�t�n��57�t甾�Q�
|�K"R�������t�K�%!��h�!a���"��)7�c�	��k����tǿ�j66��-b7���q�՛�H�
��w��7���n� �Ä��:����Wh+�aX�3E�s"\���X�� ����m���<T��/�T��h|�(�V<�j���U�YM-�l�@��A� p�&/�b{6į�;�yG/��o}�������)?QK�[��1����(6��N�m����#���!�dO�;P �5;��]��"blT�5����\LB�psX�-�F��$o;c�(I=�����w���3�=��b XRb&c��z����y���0�E:��\mf�;�+�� ҁ䟟�c�a�,�рA�*�nF�'¹�!i�-T���Q��f%��[لhN��'�_SZD���u���ŻW��.#j�N U�`Q|�>��j��0S�����#�\C��x�f�3�h8!����G�����c Ғ����Nrx�8��r�	�ˠ�\l��g^(�ff�ITX+]�ԁ�.��$�e�TF	 F���3wS�6q��Sc@��9iq��4Q�� �!�s��\��#���.V�-5{#�u���l�_G�nA�˩�=6�D�~x��~U\E�q+˯�,񶶃Q�,?���tn����aD�<�*i����vQ3|�L��;: �E�w���+ѴSN�����k��l� "B��8�v�D�i@>w�H�j�(R�� z.3ք�bLkC�Ӟ�p�c�r�!�����8�� �����+*�$,��Ki��K̋��mj�ڃ����xd������� YŤeE��]���_�\���?b+�UY��Pr����8\�Y������p'�0�f��Sjp"�,�@U>�X�[ 5���ڼ%�x�)�ݓ��O��Yo�û
R��y�$�9�=օ�4-L�6S2؀�o V� �R&�� ����k�#�w�	,Vz?t�O�D����qh�m�����B��*�/ |�H_i�: