��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\����q�?��e�I8�b�Ǽ$��"����ׯ1�V0������ ������n�R�~�S���"�[:nθGs���o" ��w�8�>��:�g&�V����k�${#�u"7)��hq�9=��6�X���oG���{Y�<G�͕ʋ�����m��m�sI��L˸Kj�{K�u�!�/�����ؙh���Po��lC(D�<��C���W~�yg7괤N�ٻ|5W���k�|�l%�������lR�>J���܌��������&�`�֩K���I�b�Y͆X������?��,>���$ ���a�⇏�,YC���(K9x�Tb�	��yp.K֕��p�,Y�>2ʍ�(Q�TN;oS�^-�W�F�`o�Qs6,���N�i�(����ʪ�Y��K`��b�xP��i�PxX�L��j���H��m��K.I���G�$��{�ʏm��Ȁ-��r{E��bm�W�+����ޜ��*�k�������
���궒�y��"�q�r�,�*��-]Y�\M���1��&j�y���7�`�ӡ�.��a�ad�Z
��An�������gGg�Uꕒ	VO��G��W\��}�[�[i/.�}b6��������#W}��*��+l
K_���H�1���~d�9h7�� �b�[���m�/�p�1e%��C8t���{^��Te=K�@2b%�S��Թ�ݳ���;���A���[}'��зH hs��iJsy&a�ǃY�77{���&��/%�8e�jOt�w��V�����}�D��gl熑���o�����=�%Z���B7�B���)2CJ��Z�4�s�����A׀NV:�Xu�����O �k�~�3>�-_a�mm�i��)7 5%& ���@�6�}��k��_�#�͉)�����>HK��[�H�x��L������C�K~o�=���ݗAo���!�S`�O���L���M�u��BĊ���oER�O�>E)?���Amiԯ� �|6y��y���j�5�J	��������K$V�')�0n8��7p�烄��k��Կ�����/�$hd*}z��Klw�c��'�a�7X�SO���]:O^%6���rX)�,�X�8T�:�r�����L�چ�����}�b���|Bhx!osI"����q>zE�Yd�Hxp)����M���OT�����j�߮Oh�Y \o���(���g
���2���1x�I��� k5D��s��5q|���~�t �%�3�4�ߊ��A���� *�i��f�U��!Ƒkɞ��w�s�y*�X�|�^:h!S���|�o{�y�9��Cc-;�X�U�Ǳr�IQl�@���M�X���co�K-��Hm�f��9��*��j�F���4H�%U��&�����U�i�ȏ3�����������K�2���t�g(�tF�:���W�Iઽ��R���g�Oh��
œ�r��t�Rs�,^5ត	�(��zj?QЌ�M���ѻ`@=���߽=d�W��^���cI%n[
����%0�Z����D��m�lc΁(�ߪ�2t.��;��L+|1�-��O��Zc�>l��-�u��|.ٔ�A5�3-f4��ŏ�
�pl�!<:@n�U�j��p�Z�i��O���k3	LM{ㆩ�Tt�0$5��z�½�v�P\���}q*��ﾞ!g\�YG)����X�&yk�l]ޏq��� �5�� x�Ŧ�~�΃���F�mL۶�K�L����������oS7z��͞�6}��b�V����D���Ԑ��CsRV5jE[���+�%(��.�Hd���#�ör^���ru������������?�(C}�C(���fI>�Dnq�1 �?�)߾��u�cdy�?	�eH�
�~a7/��*7�<l�Y��V��a��F��]k�"]M)iM�-��'�M��z�Ra߹m΂�^Ð���O��n���6�y�L���26���|��4�yEDQ.Wm�k�&~�S^�(5��u�m�:��@L.�F9)Ƣ���Au�����}a�5I��6OM�5�f8/r^I{r�|�n<���v����ж,a!lY̺�x��n����vځ%��9�;]�u�3"D��Ws[�w����6�?l ���F�8��VTV��^+ �[Q���Fo�Gi�m\�.F��TT��))�����3�����E���k�w�����sOO���֣P�O��MpX�%�j�Z�Gd������{��ǐ1�x���3<r~k`2�L��@��v��w���JS�J�4:���&�qd�U���6��`Sn#[��YŅ���3��$�e���tS ����҂����A���D�kU#$u���׼kE�I����%-7�<�7�'��L�T���a�.ӣ힞k�v�x���U�`�9��Ҕ
�"�K�#;�gB38�+��N�jh^G�w�ބ|��U�f^,��^���)zg:v�jT7a��ћeeu���o���W9��=���>�V
�ʧj+���R�?����pV�V�3���*;�K���������[I3�d`�}��{G;�U���6�b��m���@�j/�GA9i{x]o{�p�03z��뢯(m��q&�y���of7.�kqHn&3O���܏�.}	��n��*s���ɞ�+��I�$<�-X�i�)����n�m�%J&�wB]}��N_�u�v�}b���U���ꈏ_�tϨ�Ⴏu�H[ �����;p�1RP��HI?�l5��;9��="�Ak��?íf��ׂ��y�0���� �? �$4ȼ
:x��eVz��uރ1���?a���H�� �r�s��n� ���
q}��t��y��){��ۗ_f9=�^��U��������SR�a�����c~� y�!��L$���!������`��:�8@W�;hju��k�h'�I��6zl���\�2J�_��ɑ.ć�)+���]��\X�;��:F'=6ĠO����"��x6�PnZ��>�t�uzh����ߪT��J-8�,����R ���xt�_lzj��'-��0N�Qh�A�����ЀjyG�=	�ʨ�+J��폏��$,��&c����`����؏:ٹP0�zMnM�6=|1}��Z�Ł 6^�1�r7��}�1��k��HH��F�!l��7��l$�(��t:Q�����W�ۀ��Gq�<��5��AHĈ�g�􆻡፹G����[s�Hhά��)(IFc* ����k��헾ҍT�wI7GqQ�z9Y#��tlU�K��8"	t�D�x#f��`���;�gL���s�B:��f�,�-VĨ��3�7:UV����)�$�u^Ìl���L���?k0�x�q�*�o�7z���U�#b҂����=�(�R
����<�N�P+���_]r~YIGɱ��,I7���`�L��BX��D����,F 
�����t������@,��0���8��vu�o$�MN�(;�V�{���:�Ww��I��-jp��q] i�8Yz��AA��z>�n�Y=8h�t`�0�]��Y։ha�Y?��L�ƘE�R��Ύ;r|�PJ����MVz�.m�-�M6��_FC�������U��ݗI�`�E����=�3  �n�[��� �Ɨ\�PE ����0р�<gK�˙(υ��te�n�W~�+�蠟
��q^�*�t}I�ɪę[�}�RZ�DGT��:������^~��P��f��qW��[5J�Z�H�F��8���8��7Q*ڻ�VU����h�����,�r�_gʌY��ŕe�"�'H�߾-l&03��4�g�ondv�6�l�9���qc,�i���4��������e���+e��Y�뛼M��Wl���s�N�^T"v�3�L�C�A;���������T���d+��Q^+yf�p�Z����ax��IJ)�	F����#�M	[G�J?l�Z�:�!�j7���n���I1!	,�������[�@j�D�I6�}pv��'2P�JU�[�)s��;�ҁ)���y]~������n��@���QC/լ_A 0�)���;>3�An��q����;5���X6҇��cn���8t��~�D�������ȥoo�"��3������3~/	�, ^���=���D��v7�\�@�s5��> ^4�,g�u�vä�&(Z@�s�P�	�9��oA$f��0Yǿmp#�C��p��ٗ,��P'�զ��BM$D�淆��R �7D,�u)T��Ȗ?$'�j`���yA)������TY˧�&��N-�À���^���y����>��ڤ��,��X�L%�b+�;q���U�D������3�Ƕ{h�ۿW�	��E���.2W�<0 �$�,%�<��xپxx��-���Z�S��9c�kkl �,U�RR�
قP��ʈ����ՙv��{����Ѻ$����.ã+:kж���q���W��2 ��n�H��Ē0�_6ĭ�v�p�sg1������O��5��\L��4����p�Jh\)������}*;��9���������%e���
|��nP'���J��H�']�c9��Q�G�{�'9����i?@��C��Ou�h]VU]U7���U	�3W ��� ��zȼ���M���O^��^�x�w�2R"FT�����%JG,�q��
��)��@l��� ���q���oTtt�����J�ֻS���驽ؒ;pӉL�k�H��[����7��!;�M��)�� �ݳMf5�I�DL�hV��.���Y��wAj��i!�`I\�`F�������³r��d�xǀw��2����v��T^w�;ftr�����LT1�K�����[��
.\�X�u���d��	��C��0��$�E�G~�k�Ҋ�N������0����CĮr3�˜�4�N���"ի����o�^)H�1��`�h��0�9�1�E�+�����S����0�~I�H�A��z�|�*oTi_܋4�"��W�D= �`Z�*rxS�;r�}�;N,d���s��
o߁(�Ա��6wd�Y�p�
	����1�'C7P޿�z��f/ƽ9�4�	�2{���X�vي�߅o��L �L���dm��������"o��C���`���f�s[����z����W���Jr�gx2oB�Uq�r"�<��Hs_����>��%�lzu	h{T3
M�U�J��K!6A��'[(�B� �< ��u!�8v0;R��� &�g�l~�\��8�u~�ؘ����Ǚخ����^��u ���Ae�#�D����[.po�9?��W;��a]7�1���}[����جzw�����q�jݙo߄[�	O �]dX
|��z�3�+���כ����_J�؂5u�ViJ�3Y(�����BIX8B�՟CYr�m�������c[�gQ�b�y|� O�ж�Y���ۊ��� P&�$��[Ks4v�qȓC\����j�m'Ve)|Vg	�|���(�,8��'�|�";X~�O�\g�rY����*�d�c���� �GJw�x�=p�9�|f&)|bǕ'�����6�z����v�Qd\D!m����M�#�k��Q�$��F �aP+�*S`�1����ɳ�c��6��T�% ɻ|���1GP9)p�z�=�qL'='V�{��̘��\�OMt��E�(�����Lvz5�s���Uخ�YOh��y�����h�A����;�Q(t�3����e��_=!#^Ѫ�jֈ��_;h]E����~����`�݋����z�]!MRR!s�c:�ŧ��4�73���N��P��ix'3�"�B�%�sm\~��s���>�%�=Ix�O�EW�E�oR���V�t�:T���+����F���qp+��䲲)�\W��A?#}Sn0&8v{�g]yjƲDs�)^1�'IUMO��ʈ��A��yݡ��)f�|��>�i���]�3	5�/�! �2�8:��P����c�nQ
��a��ƩE�k$Ԯ�3L�M�^̂�?�Ji/��CΙ��r�aX��g�
���}��=5�M}�����Z��Fbcҁ�[)�m�Ï����O��{�D�0]����$��wb��&�v�
����LO��Ff��;0FE��1HY��~���&ZX�En�z2oʣL �k����j~{�p9fI�YS�V�����_�f��&�b��y_�/^� 0�<g���	"5�N��
. 'YF*�d�������'���J�ݺ<m2������� #�}EaՇ��6��Y.z�o'�d�"�oNL���:p�'���o����o.b���3dGkY�`9��Y�:��C*���4r �����݃#�u%ˑ����K�Z�������H�\Jo����B���L�k�>�9���{70A�z�����P=)Ҧp;����e'�]��qNF|��m@9��,�&��ۜ�U����ot	�Uӯ֡�8��>*��ƚR�[w2���������aP����t�?U�����s`��ł�V�ٗF$9�J�q7T��-o�]�����o.oUom<�dhc6pgh�{9�v�F.�ouQH϶�{j�B�졛�vӏPlY��:Ľ��`���.q�o&(9�*�L�Azb�(�G�������M2���cA��H��V��qabv��J�9i��CK�՗�[��|\�d-<�Ċ��P�t_� X��v�2v�)V�D0�o	�`���w��&���S���m�A��!lJ꟮�i���,��T���'%l�Fג`�m��dH�$�Bգ����C��R�}롻+zs�j�����ck{ ��V+`�,�"��]:��G�10�ѝL�qD8o1��A�l�;��i���Am���9�{��#mP?�B��N��s�Lo�v�y$�3_ì�kJ&��l�Kl��1�0d��]f�
�C��P��c���d��un	
�L2<�JC�~r�p�w��ǥ�@�L;���BRP����M�2�o��W�|Ȓ��лB-����iu���D���QI'L�&��u��'�n9�����0(e:mt5P��!6��2u�(�.hb��r��t/%0U�	r�y��}��%$�_�//b��>e<�Q��)�\��-��F��_3�:@J�/c����H�-�v��r�4���E�	�ͮO���Q,j����oy���
��0w8X�x)v��2�i�ⱙ���Ôi)Zٻ�kX��Y��4dS���˔����NI��}?��H�)�Ʈ�Eg�e~��m	^Z�Z�G ������:�����Zjg�aY*#�7=�
>W�/O�C����Є� #<�?#�)�?��{~�w�%�xi�U�i���Ψ�� ѷ�����I�D�RcF�ߛ����ԱH.4!�!X�p𰞌@�-Q�JO1���E(F,U������QAe5<�z�e4�fC< ��X1���y��$8Ty;���˶��#{{�D䧎�}��U:��J%1�em��u۠�o��[f�'�~���ُ�u��0� )�(�K�0��LU9��3 �A �����O�zj[FNm�Ȕ�@I��{&��9p��M��V�4�dH�k�}�;4
�(U�.��� ��?kO���Q�!�������s����z�Q���8	bvn�U����j�4���M�R��Q��pq���*`Eր��}�j�I���͉n ?^�4�Z-�5���� :�z^f �:�)��~�����,i�E�/XCR����a�M�d�R��Ƞsy�����r5�u��\.�K6X�|'#�)#FZ-����3(�A�$����'G�U��C��i��gʙ@ k�����=�ɬ�^F[Z��#�<��MVq�CSO5J�"~K*{`<��uc�ֳ��/Ə�M��"&�n�z,3ų#x�c|��vz�@;����IwL��H8rj Ԭ(�Y8�!��Lf��z#����"ڜJ�����3�P�r3M���ޘ#�-���zՏ�&��Dyw�5�v���:���t�q�?a'Q��������sy\!��s�ㄘ�mC<�u��rbd�l���E�  IC+���~n�(P!m�p�	lToJ��||	���	9��i6���
�#�9�+9�[͏�?�N�8�k����o������.���8[�zv�x������J���!���A�����k	����uTw�D	:l������Xq��x�X�+k![XUN�^��Eǖ#��]@^��m�u�X�֣��g�u�\�3�62O7Uee�_�PT�b#��R�W����W��bg�J�����	�	|�６L�HG��~�
^4'�ވ�H�֦���k��]����1�v����NM���0��H�\b��v'^@�A�b��:�S��p�p�묽�	GX�<����D�`ú���)3:����vVC�+��Ru+%�Y1�����݀{��y�?�|�zO��#�F��;�j#*�(Ti�Lf��(rL-���U�Z[>��Z�^i���+�i��‸�\�?W��yY	��D�}�	xI�jh�1/�Y�r@���6(+J}�G�A�z4Bm�nXFO1��ȹ��3�<߂$���
�#u�T�F՝�~��^���O��а�d582���Xx�7_ϛ�ZqE|bd��^-��6w�P&Z��пK��W�����;�;aB	���DG"���>��os�A������=7ճ�Z��x.W9���K�{ܨ/Z��0Ƃ����Ǝ�����E��G@����]���U�ǽH�џ�'pF~ܐϮ�{y1|��D^˸l�n�z�1s�T�F	S0��gwp^�+��GU�3���
��\W?-�y~G[N���dŏKW���S�φ� kv�_�ɐ�Vh���ql��6�pCK��V=Q~Y�M�.�d��l�3���c��Pۻ$g�A�o�7�"��;������ִm"�g`��"��FK�9�n13���m�����C"�b�頥G=��/:�g�VLu������}p(��v�n5`�M�~�ǭ
��ɉ��s�W�&��⭂Yy�s�B��B��I[���n,���t*��A�MP���h])�E5��ԣ�#!o=#�_m�Psk⤄<3g�#T����sv�T�_0+	��4�2�B �0���{g���d�,(U{��[�i��G�������h �Ei��AU���&֬����e�	(q-'5�+�z�c.2������E����Lji]{V��w[v����n�R��n��W�q+?�<P�LI:�`i/��t��l���⼷����*T��eIE����E��#JP�����t��׻�&Վ�M���*��i���pZ�fԪ�߰h|!�ĳ�(Q���G��Ċ��A�d��r�˅R� Uحd`��J?�� ����S}�����IƐ�D�wA)k�=�|���CwI��#��I`����R�~�S[��5%��� �T�O����g�|�M�귙�ƺs$�����d[6��#��9n��V��6�������q�v���Y�h�! ���0���֋�FkQ��ϰ��߂V����x�%�99�����Af|��ݘ( ��q��rk��q�e�M��}5N���No&]&���ǿ�B�.�J��j���(d�(e�W�G�o��P��:��M��]hj����nj��`�9��c<}�N�p���˟�ѱ��o���
�%x���]�sŴ�d .�Q� �m~gI"�6T�KA�֑{�&_��	P�)��&H��<�&ʝ�Pq��?m�Ԑ��DXP��������x�P�Zh{&�L��RU`�81��%P5u8'!*��:u��%��q��Ը��t���l�9����B��?����� ����5���as�X�n�����DGm����w:��c�a�(.3`�~�̴/���)�S�X6#Q��ϲ�೻25��l��O��O�H۞����nu�MJ�qb�_LJ0���e�+h��bA"�	�ک͒�50}TSQz�� ��'C��np3RD,�� fz�����&��諊�;M�g�Aw�O��7Ox���>���BjuPK��`���h��w/�"��;�+i{#���M
��߈����k��L{k��' �,�R竲d��R?)�BT�gي�\���R'	NRpt_m �������`N�W�pW�ώ+�v��d��J�Cyt�`��y���._2l���Un,��e�!��$��	�9s�Y�����3�w ^��o�hZ{c�9G(q����G���sV��|�	"����`}��j��uG�J�߫�o(.��<���J^VB���E��p^� ]�����$�t��ѐ���0����Äː��A����m�^��4z���<��I�V���OYCP�k�a��T��R��]���A����!6�E\B���`�4���ZW�n�g�S%ߕ��c���}Ȟ�m~Yr?鹾��:�'.YeS?q�,.�n��Q�&Tڙ�Y��7`.�'��G3��LC`��b�����@!���	`�g�5��z	K��-��� ��#���R���8��BS`I##��n��A<6�����=��Ugr���`r.�X�����w@��Go>,�E������Ԥ���O�%*AgZlu��Ͱ��uF�`bw���VJ�|KN���cy��z���K��Ǚ ��P�=��,>�����Ƽ.�9���9H». �[RMэG�e��4��C���~�%#m3��X�(M���[u��-��)W5Q���h4q��E���D �9>� ���r� Q ���]4��B|�<zԱ#�	}T�.7�LW�p�"�e�ߛ���fۮ�9A�_�c�rb���Q*4&��ɚ^x�����Wk|��sׅ�F����T�#r��>�88�G>	��f���sx�m:@=���������*@�C#�3��?�\�P�e~�I���o٢�0!5\}]-��L�R���WXK���cGOIp+�`�˾C��9�����.��g[ Ш6OW
$k�Cc�N��z��gQ6�T�q�V-@hv���EM���X���,ڦa>�q�����eC��5(�bmO=��:���~�_��Ֆ�EN���:�#)O,G������F�g��^��ƓI�8:%����_o�Àe�������,����2�V�'�^LK�͚ҳ���U��k݅u�����T�ۢ���#p�'��<��ycF2o�Q�bo]}3*�2�����S�[>�{я��RBQ#ٖ�w�]ŗ���a�_`[5Ƅ�իe�n+}�T0�4���O^��"�.M���jS� �+
�=LwXw�<��<�_��C�RCa��	m�8s{g�NHY�iH:l悧K���C��U*�>_`�eH��5"�݈��d����n��U�|c��۴$�'�{���F�Sߖ�8�=�v��.����;�Х���V^ʜ/C�|��3dG������ǁl�7"H9�Ө��`Ѥ�5L��J�cE��IV���1���$��[)��ė�yz�_�;E_Y�Z:4��T�	�y=	�G����__d�/0mxz��s�
	,^�l�]^��6�"�_�lǵ
5M�qOޅ{��Y��i���(���'�V�}��� #n�s ����6Ez�M�|��`�M2��9J�Q'#�k�?G�T�P.y]��zN${?�%Q�����D"[gB���a0�LK�'��sy΃��4s��8	H�.�{��4-�Ѵ�)��v�}�V�/����O�����a'(h��G���~�pq�(*���b	IL�C�0����2h̫�(�w��ZW�޻&��Y������s�z'����ٗ�>���\������$I%�V�2UA��\�Pq���f�ov��k-�������-?f��ǥ��A)��N����Hֽ��1kh��mM��Q�§/l���4��O�Re|U�+�Z�,h���+�|��4t��;���݈���������]%�v�d�4�s�������� ��C;���[��qs�]�m/�6?:"���:�ѽ�#=W(q�z�T�����RO)��ǻw+�Z����c�ͧtT�¬^B��{}b�C��#9��02&��e2AK��׮�*�FV,S�^p�[�����J��	Wzx��9��� i#0f�~8�*	b��$�7pʢkRb����/)����*J�'g����<��i�e;M%������Ë���Cɀ��	+tt<FT?߂Y�H�HcX�*mD��0������G(��a���cO�_�%��|�O�f��W�{X��_w+�*���[�vXgR �<��U`/\�.��X�����Л�QϾt���%�w����b�9�����"9�_��+���1�Ԑ�6o�Y?c<F%�G��n7��E�ɡ�� ������g*�ѝ����L���D��K�P��T'c�5T{�rU�b��h=e�X��p:'^<�K�Ev[�t.Wd��r��Q�֌�N�{��&&�/���,y{fKOe�Ax:BUT�쮀㧜����Ak��oJΔy�;���0���� 4M�ݍ��7���&d�% ��8i�>����9�2��C�����E����N�V3:$v���V�&/�t���$��tN��y#�r��� �hH���t*��]��j7լwL_���+WU�����=�]��0. �!�yx%�Xi+����A6h�����=����	? `��+�C�+�-��ǒ=Z&Z2b��*$��n�z��p�&�z�̅'i��5��
$��ض͊���@&-~��S�H�a�m��#A��^���c/���d�F|'mi�P��b
gP�IE4�x�/�kA��D�e0����;���&_S�B܆nI�u����{TUe@���˿���-���#�G���}�b�k�m��_��cB��0�[����bU��S��S�"m�]O�J��Z�%/��PEь�����PgKԴ����
����#Y�*���^�Yȫ���%�[s�	~\I�m1=�`j�4eK�pau�2����k{�j'ߘe�������{y1�b�(�$7fwcm��C��\�]]r��q�0����#&�rZ��T�W����]sv��ֱ��c`��kB�ˋfb��1S&�����F����-�vgӖ�U����� ��b�	��@0�^�ûǛITK�k{�3�������.�$�+�BƁn'��]\Ol�ʰet�2�#ذu�
ש��{��%��[E��?���+	�w�12���I�Z�^�Y~�Ǌ�O�?u���ʆ}gW��T`?�Ľ��gbf�t��4(�S�QDRP\�2�����Q�'�c<��$/�1v���ғ��53��XG��t4��I�
g��\�,��om
�퍯l<���Q{�WM��2�Į��k56��&����z9�*c���u�sEj�����Q�N��V=$p��Ns�n;�w})�&��_1�`E�(����1*�*��&�XF�@�}B��܅h����ab�2�n*�.�A��:�2�������{:�PK�g�Y����y�w)m^�O.lEAt�\��@dT�-҄`�Y�c)�Lh
����8U(��GN� �����6Z���7��l��s�9*��B|1����q+}���nO�h�٦g�C�� kw�U��d���2�
ŵ����gw���;����Q�q�$<p�TA���*
���ւ$c�.��|G��]�P����WU��;	��dc�g�`�a~�,�o�m�gc��c��q.3�˞�(�W���i�k�Q>}@G�T���Զ�(�֦VPc���/1� �&[p�Sa��?\��G�!�i�p���-��N�'K��3�d�0����p}+a��7���I��'�ؤ��U�����1�^��j�nÖ�0=��zo���M��x��ٿ����I������^�kf��j��dl;��j=J���C�ZB�}W2��Xn4��G�o4��X,j�QX����ݓ��ЙG��J@8���ڢT�d���۵I���x�_�M����Zsn8%/ZA��h���OR��aaZD�>�Z���Dyֵ��8a�����N�,4�IQ
XQ�D�vƷ�����ūi�Rg؝'��A��D7)?o����OE4���1���s�9.�ew;Ħ�h`OC�N{�aX?�Iwz��b��Y%��y�F�Cbtls$��sX�)iF}�=�B���*;a��SVƊx7u�M���U�Bs�jc�c�q�D �>*F0{є�T	h+��B��j#��g�̌��;���'%$�>�*!���[hPQ
���ێ����+Q�ӭ� j�ް���!�P"a�C�Ttσ�g���5���~�ڼ�r�#���ii|��4�H�}h�N}���"��3�N���O�}��ڐ�f�SR��|P
ޔ�*�QmeK3uD��'XsK'��>�M+w���]�W��jy����tí���d�7T�@E����
��
��{�x#�M�KՈ��3�G�g>��Rљ��u��v����E��D�N1�(i��QUM��>����Xq��v��t9-%@�24ö���}:[�ڈ�@���X��l2Z�χ���{a�n�	G�ס<��nl/��Sf���x+��@�.�s�/fH�ē�no_�kR��y�:��y(ص_xwu�����uI�&N~���
(}-�$��{C�?4���8p��˩�	W��h�=�,a(�(H�*�w���WQ��f8�_q�������٤�f��C���ԷٴDM�,<7)�{�y�z=����Vz<�l'3�;���� �2{���0;�CY��z�����Z�c�@R� �X
�T2��������T�jYG��C˥E���甜�:t=p��Xi� ���	Д��.9ߠ�|`h�s���rC
-�c���%�|������҉������xNm]�X�o���*p�2�olo�ɩv+P���q\HUL�.����£`y�:@��)�R�M�s���>,C��J����MT �稡>�2k��]s��y���m8�}:�r۝��\�/.���!�7G���#����נ�Z�Q�+p�t빊4K�z�EB�e��9� ����$��zSZ)��<�8�C)l��t�S��.������QcPl.}M"/�;dG��Z���p��P�6��
q"�S
��0zi#!���6�h�i�u�0mc�*�G8�1	�)�|�l�/��_4���@B���
	N�|N��k�vc xD?=�1U����E��~2U�gM�N&3_�{�� ط<Z�#�a9?\h�����%��4D�6x9}B�BNϕ[��h.�N�M&|첨��6��qQ˨�y�X��x�^�q��ҩ�)��e�ON�	�x�y��џ�2�NOD{��B?8t��˴:�0�9��m�!��>^+0I^Ԑ����i7��r"���Y�S�1{�F�� ^w��R�?)D-���:j5Ckm�,�	p99	����:��\h�!�u�X&3	�Md�5��b�0���h����QU��9Oa��mcE$ݥA(1���](�,ψ !|y@K�=Yk|&�������K�7�86���&,��Ut�xDG�w�Zڵ|-��K�zԽ |��80�a	�&��S��̊���k���f q�ԩj�+B�qi�8}{%�Fo"X�:���;5dɮ��*�����y�=6��2��:֣b�^\ʘ�-�u��0B_�oO��'jU��3�q��1睙�@��05eA��!�3������n���B���/	3M��iТ�#e�4n�'-�\�ۡ�?QO�&�Q\xbÙ��~������Y�z��o�i�*�����P&��:_��:qhC9;\Ԉ���oֽ�@?
>Ղ�F	�`��܉'j��VX^�9�|����n2�'~A�p�p�*���&�ֱ�Ӕ�-�^6���5P� �IR�ꢌ����� Xg!����*w�)�%h��C�1O��95&����Ǆ)�����mp�M� 
�Ȑ�_�x�yr����ua�DS���C��9-�Hg��JN��ڤ�͚��n]�^��c��Hy��3��:P,�~�C�4� /8)ء�$V�ި��_#���i�jd	T*���aC���V�K�ds*z�j�F��IR���s]�(�<d2�׆`��tӨ�F�9��S&�5Y]�=�Z��?_ѯc!I��g�g�2+�ذ�ӿ�?�27�����<�Y���I���㭨Z<���}�1����m�	��D���q3�t�G)��:s��x�ۀ�5N�-t%��Yr�\I�X�HrpF��D�Yݨ/���6��^��N+#������s�Ǭ6��-~����K�-+�����d�+񸊮��p����`AͼY��\��ab��~�/��$G����,��'��������ф
���f��,����v֙���c|,ך8�I���U���!j�D��O������i�����r���`����tb�e	�p/�&,��Xg5Ta�R
2i�_�T@n^Կ��!}�@@��]ے���N:��*ƕK��_� M<Ơu �s�@7��UP=���P�Ę����33���� üp����6�`Z�'�5�}DD�������&�/Z�x'��X�Ǎd=���9��M�AO�"U�B>\��'Z������|~��'SQ֠���J�Χ�А�^���ϱ�KБeY�\E�����(�>�ьvd������H|���#�
�W#n?s�~��U\�);?��E`�S%�{<Y�W�*
�Sf�b�ڊ98�|����97�ΆI��'��9V[�đE=`wA��Υj,7�k#��Qq�E��C��c��\ԯEo?�O��s$�����#De��s�ʪkł|s���V�����V�%o�U��R�Yŗ%ͬO-w@�ۻ��7�&y���v�2y;�>BKn�}�r8ݾq\���L��lP���SB�b��: �
}�bͿړz�	ⵀ�XA��MpԳ*�)_q��|�h��0�9W�>�F�4/=��e&����
�30��'<*P=ɡ2��=�6\J��T��F�����K��U]�D+'�����L���~���-�����@eE��a�7 ���=���k!/-��p���	C�(�g��1�UgF�i`d��6����LG	�j3`C:�.�!�A�B�*�I��4����M���i�ϯx�S�A���J���޹�
 ӫ.���>�M�E��x�d��ѳz�d��YC�2�:���y�`�VKW�'��р��]SܺafQ����k	2G�ُ�۵�E���:�#��.�O%������.��c��.�d�?z���1:���f��ݦ�<$8آX�:��܉�L��qT�j���TA�Ά�]ۢ�q�Vy�m���Gʜ�v���!�$`���=�	�,+�r��?�!{nsh»�{Ƚ�hJ�0H^O}���#%��0���ۜF�ǣ�Ue��^A�F��hW�д���R�������������6@��L6��#�n���}~H���O%��'qPOdӑ�0t��r|9�SpՓ�Μ(���9��
�>�9�,��gHY�C��Q��mD l����n>Y{م�����@�T�`'N}9��3n�v�/Ǖ>(���4r��}U�q�I�4Dm�P%IZgq�Ƭ/(���%& H���K+�jrЍ��-X ���-�eyIΞ��;�eOF]:Wk��rE/��x��ntY@k���T>��o.��1���if�M5�	N�*Ú
'o�Q�%����lmr"������9����s�R2�5h��+���#�s��������%-�b1����6zΫ��؛$C_qx����]4��u��2��!&���@M^w#�]����dˍ��[F��_��!�"�*��lR�|��󖂃�I����%Ϸ&��E3A�b),:0^������������A�y稭Pp��]У�i�	�;{�����W�=�q��hNg`}�1f"u���zM� �q�hTZE�Ba�߾�T����kB\��s������e�}����"������HG&] Y�iȼC�r]�����Ғ�~@�7��}u�4�Z\�L�tѥ
�R�+�,0����1��; y�宔�n�f��O���d���^~�BGi
f�9�5{�=E�����X�\S���x�Cڏ2Z�����͢�$��Ž
š���Dype\vύ*ج�M逕��<Q@��Q�\�����3a�}5��Ck��V u8�� :;qkG�&� s�����u���߈�q�G��n[�(�D?�;���}H�~�7���6�z#<�N�����LƷ�>0ӗ����r�*X����+�Z�� ZG���R�xc�A��)}?>;�9�Jg3�5}��01���I��$���|7L��M��j�`����+�γM���,�%)(曣Ӭ�e���h�y��uT�·w�	������7�`yͤ��<�Z���WBxH�kY�~��"e�L��M<�`�Y�is��km�B:��V휼��.~ې	��]�41����Ȅhr ����B0���_����r.a�I�i4��F��z��$���K�X��o�]d�ʖ<��h��|h;.?�rza���zzƅWG�b83HD�B��2�}�L&l}0�n/]G��=	��oǐZ�����4��<"�n���.TS��'�[@|o��XǀtlG���h��H��S��� ����oV�=;�9��j5w�w�]����DtdH��{�i>�G�j��$����Co38��rV��Ɓʹ�fj�f|�~��wĎ"���b0r���@6y��*c3�>-('�,w���_[�c���eյ���y�˫ʻ��v��<{�C�^�u���� ��D'���CUh���';tjg��k�����F��8��ף8dcI~��w:����i�Ln" F�RA��w
��ֺ>L�_c�r2�2R-i�Αr��u��P�W޼�_[��ʪ�Fx���y�{���������B�����b��d��|�߿lq���A�K#>l�V�/��%i�*@��Z�i/\5��OJ��_��ڙK���+�a�K_Q�؆--q��~c�-��F.Ǻ�OR����xCQO'.�}h^&T?��V|�}47߭󡙂
�~�I!olG�xz� 0E�����^o��V!p�]��?�޻���?y���7��Vr颉s:n[<J庪2Z>;�I/.d����*�k8 ́�za;O��BR�L�m)^*̈́cHD2e��yu�-pD*��d�{!?����
�{Ϋ)����$�i�vS�3ު�$���>qr��|�?����hf�Fhn�p�O�ǅ3�5yb���Xj�&"��0�y+,G���\�`�����J�C:�s�l�M$��9��K��8���@-m3��p�F;�ˉ�WKm���<��-���&틐�����6�_B��f��t���'�����$<��H��&�n⪶
t�|o�toH�K8 6l�Wv�%g��7�����Q�����	��U�j.	 ˔�.
�6�_�p<č�����mG�iqb-����W��v.&V���W��m�ѿ:�kF�)p|��eC]!�%qOo4 ��ӱ=0��
UͦTZm!��Y�FU�J���ԍ�@T�`W�& ���E�i�np._.|��eC��>o.AJϮ�މ>k�oG����7wr���\���-s�ǳ��yQ1�
��6�B�Q���$O�$�-1���p
��Z�־���#��P������.�s+��ۙR�qhb/��@�f��'��xR�nVL�4�R����D�F��c���x�:��9{�|����A�Q�hU�o��T�B����s�7 хB�-�SO/|�j@�� ��=�j]��=Kҿ�˔�3b��u�Z���-���Y��O�f ��HZT[��/'���r�n��zI~2!pg����iB=���_+G�Wp�����n���_�0sJ���[S<�	�@���MIU��mMc�d��!T��T�'�S+:�$�c��U��s��؅����k��V�(�:�<1����}"n���▯��rWM�6sK�Ǖj��.�l�9@Q�X���Z��D���L���n�R���ܠ��#k�_��"�$=����a�J~pg��s��V��y�����0GQ���̖�~F�u���a!Yt�@CU���Vhe��o�����;�&�U��ꙭ�c��&���9z����t-�]{G<&߬�N�c\zpF���#��]����l}�.�;g\��\�4�f��H9��-���;X�i��8�&\�i���Z�L�h��䨹�z���H?k�-ߔF����KY��;)�ձ���Vb��W����c�W2�@��Jj�$�ƀ~��<������b���ntO���|a��[��������c/���!���:������ᢝا���u�=o)�����m�Z<2�{Mp��í��4|�J�ٴ[���SI\
{q����Cg!;?L�T�LHd3F��"��1߲�������~�K<�Щ�	�ƥ�Uy �s�<%�Q���M�P���̢����M��夠8�x���P	�+�g�������K�nՅ���)�pLp:j�(�]w�ͦ(�<��T�,��L0�	@B�q�i^|�߉�M"�*�g�9�Iu���7 ��vd+��a:�LW?+����b(�r�� �R~k��W��5�s�>I!)��N���X�q��F�Z��E�g?eb���Q�{������ѕz�U5��31�זC��5
����R�4�=�;��ȥͽ� @H�.:i�ʿ�!C�V[�H�(N�6G�>�����z�I]�jH�|��ѱ��\ys�0+�VBH����i1p��.Z�w�mm_3��QŇ'�s�+������1�FRC{v�,�8���m��mv�<�\q���{��<��Qx[�=�*���|�4b�LH�J��(o9&C��U��fE�����{��eԏ��+�k�c�y޳Ef�̄y���c�v���,�5�Q��=A;}%-\94;���aԼ���'��7J��w������+�R�ɶ� �a> ӟZK|W� ��9MU���~i�]à챉:�����;�I����P�x���~���z2�k�޺k_��0A/����k(��*^����V�̾�5����e��K�#�%�p�s�s�~V�"��<���|�gL�"²`O8�T�z9΋C�h��B����vz�
{��{�=�xQ��%��r:�s��>t~5	�E��v�𐳡���:2�y嗵����'x���ĭ�>�牰��(������ ���δ���g��iw�����ÿ��me�"��4Я���S��
�Ҷ�����(�$�u��|.�����#�ʩ��[��.9��b7{B�3T�6���������2��S}h�7 ~4=#P�5�Hi�w�ѷjB�;�y�|F¡�FT|B����F��-���2�+~��E�ց��W��-/�����XaCSfo��C6۠p[���p�	ޤĖd�@�E򃔱��	�}ʕ'\+�̓�����q�,�dO"��6� �^�q��4��#zz�����%T!���7LTt�;�I1�۱�޺��3�7�`NFw��N��1��3�M���}�O�T��U{����ʽʒ���Q�����Kt2��>�7��"M��:"��I;�QU0��d=W��̠�hG��h}��x�Rb�	��n��`jz��{@�C=b����
�s��E��7��D��ͺy+�8p��4���)��圊;U��w2<��FӲ@
N�zeum��󢳦֕~|Ѧ�0��=��+�5.�^�>��ow(;M,�*�e� �tt����炷�Sz�H��e-�N��H�ڗ�f�lY�j)_9���P�幃��7������`���u����L�a4�!�3.�ޚ*&G�LpӸw+# ��̎�u���M�o���gG���a>0�ѕ� ����!����콈� Oxwᣱ�ɂ�[5�鐯�g7
Q��SA�� ���Ų����H���R?���@:�ļyQ�!�3�^|Pｐ���C߆���\�py��S��f7.N�]��#NO�|�u�oL���ޮwHs�~�١劵�a+�t��Y�|�TF����C�zl��y��ūa�<Pg'W�q�[���߭d��~P�#�I�}��1��p���>vz�IW���(�[��G}s�{C�,i]����ey���D&��N��7RF2��K�K��ы�]�p^�(|J90���D������ȟoʍZ���Z��<��Ď/�%Ss�؀c�R�
�����J����H��'�b�?�o)��0;]�Wr��U����c����o�|�׸�?T���熱c]��Uw������:*�:�,��Rr���� �Q ��g;ӎ��\|��6�O�g�����)/_��
?e$C�$������ʕl��_��A�U��7�{��(w7/�O>��c���q�Tr&ᬁ��g���UlR(�2��c�S1�*�m`�SŁL��m��("����PiR����%��U���CO�g�hk���e�1#I�om���7�=3�R:�~�[�*�yjs�X�;k��.����g���X=����a#�#6L���4Δ���Y��U�m{���)�B<si�_�Ȟ�b��gn�[����������U���' 3諊��T,�6wC̠١Ώ9�u��e��uN�fΉ�s���B��G��fg �O5޽~���g#��59-4�w�J��!��=����U3��l��)�i�G��Mp�Pk�T_#z�՝�{ ���x;r�I4�X��,w:GJ�x<|�Ҫ�#���2������܋�7	���
tf塧Z��_�r[2r�*T�G3��k2U �Y~��%��'{�IVnƎ
S��F����ngxH��w'�x���8�,ݭg�it�g~�TW�^����8�;�ɹ���t�5\8�Brv�Z�d?�U�@�ȸ�����|��x}�Gڵ!���t�?%��v�P�"��&:,ќ�b�s�/=
�h�n���e��o-��ψ"���[i���q�e�	l5&!���ۅHd+6��[�='�OEJ���z_��Z�bH���8`���E9��5���Ʉ�HD*V�U$|	3p���C/����q����U���m�\��|z<��W�i��]7����Ҏ.$��W����^���=��C��Jh�>�t��S���΋���(���NZ��:��ӑ���2� �-���ߥ���[�i
HE�ď-�����-�)��H_H��R6K�YM�1�.�U�(	t��DJ�~׏?"m�|��m���L�TƑ
V/"������UDI�w}|�T�7����?Q������y�
��������o�P��Tz_Q[��8:C\��ms9���p틴Y����3���s�Ո�>ӝ�v�wnU_�i[�/qE��N�9!�3p*���>�ϰN ̰�?��EY��3}^���]��k���P�N'�}���#��J��4�Fa�&M�~�wD�4�,�H�O�=�-�S�C��\,-JE�4m��)I�`��IH��7��0�i9�#�F�+���1�D�\&�����A���tA'����4�q>]X�aT?�
���t����ɐ���UG���&�A�m�mp��i�}t�bdl���I�e�QM�K�/ɐ\(ۜ'�>�ɺ��_���J��{��	[�y�J3�����.�<A
����(w-�e*�)�T�'�ʕɍpGj�Ͻ�%%J��̙�S�)��Bv�O�%	Nx~�S�r��IyJ�00~�=��Z���[<����#et�?ln����"i�j@��&�p�����{�צ���߷�(�x^e�\���AǸ��Vl�NX����ۚra��糣X�Q��3=�s�Y��X����s$�'�a���bI���:��b����v�_�W�ƚnU�.�pzZ�&�YڧsV�T0�%��<�B`�gڜ�b/�F�6������P�%��<`�����o]b��X�c�;��~%����8ʶ�DtP_�Ln�p�GL���m�hZU	8���ֵp�_���<C>p�sW%ˀU���Z"�[6 P�!Q�ܤm�]�K�B�w;1?��/qv�h[�(��Η�W�Cy���8�:���6c�z'����d�h��0�\�s�
�k�3�vk�R�̰�K�`[�a���2���(�۳z�2�1>���rG�⊟�%l.8P��#�H���d敘9[`=K�����iT�b�����0��pp��������04�d��9��>`	Ik%  q�ݟ�y�]�ھe퐠�q��l��$��U!T�)�z����J�ԿQ�[��]�*�}H���>��ަ���T��l����q
�
چ�b��	�e?{�$������ⱔ�DxL�#�P�é��n��qA�0�D96��]Be��Ӣ�4��]�B�SI-����)H��H+t){Oq��1�sU���JY&�U�팣(d�[Y`3
>�TL@���T��	�T�T'�s����w����VRwA1RהY,�`Ca���Lj�{u����f��*�c�tfL&c�%r#K}�c�>{4��#}^3�\�X���-/t�4t+Rc�qf�آ��zVZ�p�	C\9o��{�Ƒ�
�� ^����*5�J
�C���&�8���U1{���ϸ�taT��zN:V1�NC��k�.�y�mηN1E�Rf��b�� ���n��P�h�f��0��j�t�a�����w1�6�L���'1.v��DMCt�Z���[��q����\I?�t���B�?��i۳�}���2?�@�:�E�[߼)����-���'��[&S{�xk[�Wx���7�|��_V巿S��Efp�ːl��'��w�iéR�χ��k��vf`��o�x����LWv-�i�i�<���r-�u��� ��	�����V��K G�M�z��g<������"����a����?�ޑ���Ʃ-��L��
�pe�W�5F��6f,���|$����:�M+DZ.41l��ȞFO�c����M���S=y��@�nP���5��RY���o�"!�N��H&�'�O7o���,
�{
^<������׏K�{y�]MR�4��4٩\�M����C��~�wiI�@���HQ�n�;8ЎY�����rfEߒje� k��yͱ��$l�1ײ����U��f;�(�5���A&�!��h���t�K�B*s��ݚLR��"x������:������h@�%���ｬWO����ה�ˮ�!�#�w�U�^�P�h�ߝ�K�)�͐M�8�YJ���Nm4��O������f-S�(���X��Ӡ)9�s��V:�{�g���"��D]���<�K��Զ{@6��e>;���)#���v�*C)p�O����l�M�������,���H�� 1h΀t���дK�~[�
�r�]eU���ڜ��2%�P$6���g�Z%�29!�8������q���Z5+��2��v��ƴ�xݖ�7ڤ��f�݌8����0�����'4�����3?�K�J��ʒ�	�76�();�����������
HTt���'�L��mp���-���y��x1)f��HZ�6����k��Ң�C�D���u�1�,�ȴ�7��[rn]\�48=���Y���l��(���q�3�S;�[�&k����lh�n����hq#�"cB�n�`&h�Db)�0�d�NP��Y;�^���>ʡ�>{J{������I/9Q�"ȏh��g6#�h�be�}?	P]5}��aT1��닄˸��+ޯ~b�.J��`�B��ɀ���%��L�g�\yY(�sdar/�#6Xc�����0v��s�MxPS�R�r�,�8���c �Z��>	߿�)����4�����T���^c�;||���8���	�x��I���`2hi���X�)�1p�Z9�a�R����L�7(7���Z$5"���g��/MF"��K���7��5�2.Y��]�}��J�A%C�����e�H��q��`vT�P���/��>%�4ا#����/?n���,>��5��a]�*^ҵ�
H�6�f�'p��߃��PYΚ�	���E��Qj�ŕ�Б����ߛ�����ԭިhuȡ�yk]��[ P۸�eoyȝ����dO� �}[o��������Y�I��P����'S���	�o�H�HѲϘ:]i	B2`r6�]���u�ӥ�4~�+Ƥ�������څY-��F~`*�ؙܽ�^�3j�,�����ac~�Bft��r�~ˌ�Q-������E���+�}H���tc��S��9�ޢ�>{�>\���)W��u��}�,��S�t�&�h.�� � �4��VaUc������Oyqj�ȃ�9%>� N�aM��am�R^tZ�1c�qK�΍'����#Ѻ��&�w����ݙ������+D�0�y��r4QfGKx�u����gn�iB�L�TqH|anꔯǱ�P���vj[�TQ+S�$=����0��[�^bg9�����L�>�ѭ�ZL)��߮�M��~n����#ϯ����Ci���\Y�}��t e�J�����Ǉ�2�������5ہ��h6�k�[bօ�c��*~P��,�Xb+{�ҧKҹ��a5O�T�� -4�ff�X���sh���S�	��b&֤gE|m*uzQX�`���Ԯ%/�����f�Wg;ܴ�5��j�T��J�p'��v,����z���aS��5x����)1��8Ҽ���M��H�ω@�I��W�i��/�ߔ�Q_0Dz�\V{��V�*5�}�d����S�(�����%�@56l�VY�S�I�Ek���J�i!ɍ�LxT�� ��u�
��uZ+I4��w�%T�@R��#�@ۛn�՗B� ��;-顆�:���✆��1����H��r�?\�ɾ	�Y����JZ�@��&��Ա�iuT�s����lo!�U�<N�Ϯ��<1�4���t��BE)�߅Q�u=�`RD��;�24���z`O����克H���w�]�Truǟi2-��J��Z��;�	h�.�qk�h�,I�o&ev�5W���
�����={��� Kim��,>�1�8��
�j��[ͼ�)�\�>,�`PP����ڥ(
��zѝ\�B��֟��+� ���~�S���!J��[�Ăl�uPؑ=$>���mݨ�~�)π��b��DI%�]�ppM��5��7�/�kH�X���_���Y��>A�V��c��
�}9����5}%�4ID�f$6�S��7��3�Bƭ����7o-G�
Ɯ�4o�$h�@�7$ua8�n�x�Pa�?
Hd����f�{�"+�g��z�"g��\��L-���]�Й&�-����\I��xzp�_o*�j����T���C�s�<���mh��sO�eLC�����?W��ـ�#����ú�̰x�7|��UK�Yb�3�С��G�e��曙�ǡ�b�P7sX�/��-�n�fQo���
������ x�i�*#��Zߡy�i�M�
-%j���:<0�0�4R\a��&L�i_�F7���+������wQu����v6��� ��Q&�n��\�I�L2�b�N��V�9�t�c���7�,j;J�����掩vc]����gH��L�q1#тW��#�k$�]X�����%�Ÿ�l�1�ߕ���-iW���YY@P��kJNP��e����ؿ}K��4l��X0̷f�zn��l�p��֍��
J,nВ�T�Ħ�Xϰ�]�Hm;ء���%�'�[.2�r��� �޾	%��O^l*�R���ߡjU1�5��Jf�i�;{[�b^E������:@�f7��4+�^x�8W�a{����~�h�@������RO���ҁ-b�wL�b���2�Ӵ3�;���#��
�T@�&��^���|�2z��U�8���,�(�͕�_n���G�s7)���0���vF�6��p�L�"Dy�¨7�(���2젘�	9� R�)êe��7���i�{[�f�n��7X�c�RP$� c�Ijce����W!B�CŰ"��8���V�Co�"�49��.-��W�/v;�غ��Ҝ%g$�я\E�ä��2� ��D�A�6Cg�"���E	BDg��P���Jq�{�b�$�yn)���Z`��x#�,�����>�M^ /�2^_>[mf�G;Ot�|j3�]Rn#�@,�a��4�������zH�~m�����^�n����qN;{�{?����X�g�ؒ�WX���[]��<�O��D��\)�,2��"�>��t�8��[�n�+�=I٬϶#����aM�aW~������sW� �m3������yŴ�܉ai&8b2��[d�R��LE���A(�>��8~kW��VB��R-�0�|�����Qq�����&$�G�Pʳ�)OLVA��E���̝�`�֢�⬙e?:?r��X���@��R������W�_V�����l̍+R��;�lɢXA����Z�#�G}�E8����A5'�^�2;��o�^F���d�x,�b���B�H�G�5>�I�˔��g��l)cT)q'O��*^�Wl�q!҂����)T
�4`�?*��(msg �ֵ�&�s�W�L����Y<P��K�$��љX-T���󙐸�Y��>h���ԝ�0�]�����H���r>П�ν67t#�*<z�b���ͮIV%-���
����A�,���5+;���R��)�U.�I?��ɖY͎h�'8 ���CLNo?]7*���:�}E����ciϋ���Ȉ���x���Z� |ds��)���9���6�]
(	0���a�GS �9���%%�7[��;��}�=~e����t��9��e�r���,n^�Nȿ�*ˢ_?�c�~��Bg�Hۛ�F���ћ7`�`�B�/d7�bk>�˵�2z-��g �O[��ǉ����#^�i���f�V-$�dH�]��E6Y�5f�>���>��|���Z��l��V�pw�,qI+��N��K�(L^{�9hi��2�i�ɑR"�a��P�����m��)kc6(D}jvƵ9�n6��'!vM��G=�k��b����dX����J��A:w!l�~��WiM�������1�G��"H��4W��u�v�p3B���8;!'�l��w41��nE`�i�Ct4��^��Ey�å��=7�q��"ԛ�׶�C9����u�zz�b%�L�c�R��~#��ǌ^.��;�Z�B�w�'F��a�*ޫŪΰ&�m={GK~��� ��(?E�,�EZ��6����5?��P�a�%A�-+�ykW\Pw)���Y��p��6�N[�Bp\�H{��)��B���d|�XF#�I��v|K�9W��y�*��⸀��bNq9Zs+���9�� �Z ��s�Dd��?�&�������극"��^rݾo �ᚡ�Z�h|,��zkA�t��T���6Npje�3��t��XOp�|�(IW�2o�p��*�$��8kq����Z;m �|>�CA�
8}º��]��b�C�lg�~ks�m�a~�L��篦�%<6�������
Ѱ4�_:&l�ј[M��=��4Q�m��k�_^��{�	�,�踜��E�m����u�2Y�e��䗧t�xMR�7�҅{H�M`tG��kΧ�yJ�SU5୐Aa}��"4����G�Y����E"d��y�Իf~+%�9���O�Z�$���S��S���y�J�v���H�҄^K0Yai��^�ĭ|��|{塣b���#׼ڴ;)��l<�Z>�1�rZ����ۼ)L��/����~\�xlָ��C �Ճ��)zY��%�A[L�阵N���DP��
w�#��8��Kv�&[
DTl��Q5Z��m��Bb[�O�-�V٫`%v��Dz�^ "`?]��g�"�U.�<h���4�[^(��b���&0U��I�yU��5�� y���5 G��P�s6�j�"��1H��S/Ve1ޘ�òXo��&7�Ar�$�>�꼬������̊�F%��̍�/k�N�cc�H���j�f�r��m9���t�	�!^T���R��uל�Է�N�����3�h�+4�[�)�"6K9(t���ug�2��Ol�m=+�=�9�����8ڥn'~B���'Fd�VdV��#��^������%�2�Ή'�O#مb�*�rm��p�]�g*���$&Y �����S�)ԋ��ݤ F_�+���:�Y3�X��~ώ+��"iI�@�c�9u�r@K�,'���wmFèFͅ��e��Z �=��		k*ó���?�N��8^^찜`���NL�}���o�UN�0����4c�����4*^�D�B.��u}W$	�2� :�۱�u�m���+ٳ&�slI�n*�B�4�^���t�<3�>�]�q"�i�-х?�C�y����.��@@�O�ۅI������&���|ܚ9A�_��|_�%���=�g���ɪ�Z}�N�yxg����N�_�K�X�i��>,$��X�1�Y�1՚f"�*���S<�	5Ec�νE˨/ �������W�ͧ�G=�0�;�4>X�B���75�8Ry��X:^�1���j��Oe��_��B}a9��A2������w22�A1�"5`'���<�&��M 0?�`v ���q[�.\RF8D��2��bGU�P-������d���>_�:!�=��n��Z��ĥ�.@٭a_�$GJb��ݺ0�`#lՏD����M7���~v�ֶ1�O)���::��T����<�q<;�m���������=	�l�(P!֛%E]�Q,q�8[��/2/�����L�A���/׀�b� X!#0������-+s�&M�a^
�e禬�v*XG�a:13e���^�}:���22��"p �-�V�^���iF`<�QHվ���}6��z^ݐ�z*Ɍ%������G��i97�r����"��ow� �0K^u*k�k���~Mth殇&K3���jУ�� ��a=)��R��48t{q��XD�!;ɬ}B!��nwѤy�Ũ�V��C����U���el-*��q����ӑ/�-#�ݠUEGv^;�w-�����Tw�F��T��;,�"�)���b�Z~�&O���jMI��iA���F��*M2�S�9��!��Uw�n�-#=�����G��uw�Z��N'
`�v�l�^L�<v�"�� ��7W^���.A�8��"�� ?���ک^ =|)s��N~ʿ��$̿A��a��jy����'�)����軗���.��ѐ��(2��V�i�;��&'ڌH>g���Ɓ�%�qғM�{�� |�+�.����(�z�EZ�����>��Nuq���#��,�|\w���������~���uEe䝿�#�P*�pV�������Py~j�etD�|�N�ѽ�_���[���<��$���2�z�SZٰ�K�]��=eE!r ��URа�R���I�s���)�fi��ؕH���:�Q~��aq�
���`2��� ��Q<L��w箬�M�6����T8lc3i�R�!U{!Ք)�˅�x`�ɴ�c��� IutWl��G��%Z.9����*��#������>�0��ʽ��|�O�o����V���;5�X[��9 �hW0L��8��ϝ����x^�O��������b�uXT��h�_O-VFK�GZe���sݑ���p�1��Y@�k�X��L�E��,�y��=�f�!�_ɬ/1�WGm��o�����m�G|ݓS
�"� ;�LOPDW����$�H�rt����D��W��K��(�P@����E��"w��ic���l�:&�+i�^5[��g����l�O��v���`l\P���似1���|}+ב6��S�$7�n=pY�?�ʥ�+GO*�kj��HVx���;���hJ΀	w��w��.lF��`d���*��P[R���L�<e�R�B�
~K����dր�e%���Ð��v�y$m���~A�'XUf{�Ri��>�k���P�3�[���]�|��M6o�����+�x<�1DA�p�������lTK���o<�9�\t���/Q�$��ky�!�wG�0U�t΁��A��>v�UDh,!�,)�-X`)��d�ǺU����A��d9�}T*+H�A����kk��z�!��*�AG�P�|ԝ����ܒ�D����!���
���[T˳wx ǚ�u�Y�u�A#�=t`ң|KM�F�[x}����V�3���t�����«ez�|N�E������v�7��y܉�C�#N�J��b��vN����-�i��Йx�x��#@0�t�)�ꦞL&��>�Z�Q6��oh��M����$M���=,Y�%}�d�n �Y���zI����r=��h��������|\�~�2���-�HJk����6����P)�T��^@#�8�̺����e�	c�&���2�b�Ko���i��.���Gn�z��?�� 9��[N��U��X��ط�g�6�.#6������<zf����v�2�"���;�y^��<M���v�2����΋���HݙB�\� r�Ӂ��l}�>Um W���n�{y�ʖO�/\�f���]�0��LG�����d N�0?|��3�_O�z-�\!&+���+�%l8@��� ��/+[LP�#��O��/����Wei0|i��0 ��o0%�x��Q(��dy��`5���w�޸���S�şė��ָ/���\|�b�-��C2��p�}̌�H&tJ/���\��0$�C�Y~����v�T�(E�ʼ�����-�Z���r󶚱�)�^�������Զ�`I�P��Li�
���<�`\`�҉���DpՌY�[�p�䠸[�����c�˛����zB``�L#��EkG��%��C�h��T����B���of2[΁��n��'���\]xw�7o�'��&�/��7z�aM��������Rl��<0��)���z��6������z�r ]H�7#)��	�$�H�ޝ�B8�FgЁ�U�8��}c�r ��WDa'b"��4�~�J.�k��w�L��+�!�Y��²"-c�3�Qy!��UJp��M�Pfy�9��W�?+T<����:�E\�m��e��Y�r�ݕ�z&� ���a��[�jRf������9�J���(_2�d�ʒ�~\m����=^h����G.z���S����ɛ����S��?�Ҙ�C�����ᐗ����!�N����S_�����T[�R��t�D=�^��U+���L��\m4�J^/�ݫt���@���ʰ�a��G�D.�4�Q��ut��Zs�En�G)]�k�Q���LBI�(c��Y�-�x4���1�ͨ��2(��/$V�z�ڦ���Գ�mi�K"L;XH�s�6<ƫps��j8N�.*P�	�:������:��Tցk�yE��v��a�{'�5sk�����4�"@���t8�*yM_P*~W�Kk��Smw�����Exx�{2�S�>-�c'߫�1��	A+�d�zјC�к�?�D�� �Ӏ0�����ۈ�<9 �GP�8�'Q}ܓ?+u�v0M�fo�-�|5|׸U4ݣ[�=��}�/.BI����D|��&�fwq'b=�h��O(k׉�����F�0а����Ð�G��+�C��1S�A��AӢ$s|DJ�	fQָ�n+�o�e����&��6+)ވ̝��d!���CW�gBɬ��(6/��_5�x2�0h�.�4�KJ���t�ױ-����TD�-��] eu���u��M~�OE��t�+�P^*w����.>3e�[���٤�K��������|������gڛ������W\�a��|[�L,���{4�]�4��
�r�98A�S��Bpn���,��}���F��P�
�&�W��5W���G�|u�}�UO�HB��;�2&�u�~UѤ3�Ů^y9�}��0��M�_����!$�|�Z4�e��x��d�a(:�R�p��GǍ��֢�����v�|�O`(�Ƃz'*�q�l@��%��e�'��&y'(�c�X��݂�ݐP��z�x(��i�-��@�(դH��] �����F�'L�eV�j���ꥄs[�P/w�Y�|~�"� ��'H ���h��!��D�bB�K�1�F�韩6���
�0OB�)?h�_��MUR_1=Ơ�*s���_��OLR��nd����[���Nš)�loGy Y��2��[J7�0%�I�������F��ӄ6]�!�jr����t���CG9j��BN����f��I��Z�d"�T�
�z8��8�2��Vg0����A�?^��0����%����%Cs����4�<�aj4Ғ�Hv�MNrFK���oM�`�g@
yI�*�&�o�;E�e����%/Iy_���;�}���\ٗ�d'嫝�JЇ�n�� �o�C�~�s*�C��)�pv�����%����ko�N��V��G�Q.���v_$���~�G�ъrg��rZ*z減��|�у
��ف�6zWh�����捍H+beWüQMG��E�
��IT�히G�n����0}E�-k6�kk�ܳ�%/���GF4���_�B�;��@�%�f�J���^�����rO�����%�����-r��R�ܳ<�M��l�������YQ��y�]-��5&zh$,Sآ�F�N��c�<�A0�{�u��Z�HX�F�h�����6�#R�蔾ww-=�j&踿K��<R��:k*k_����/�wي��s��r���b��FA��V�;$�^]���⠗'�=+2��'��6D@$u�:Gu�2��p�C���51��wp�)�$ر��ڒ�SahT���Ϯ���%~`��X�~_�{�Ɇy��s��$�D�H$�u��t�q���%��xNS��9���V5e��m��dFs<c}p���÷�\�ޫ�l�d�yD�ėb�7EM�
ި��G�K^�%���*~y�ĉ9��^8���G���LV���of�}�6�:U,�p�e0���; ���XV��K�XM0�W�O���8Oo����h���R���19\,�G�n���_�kӉצ>Á�^ӂ<|i�l��90���ć��+ P�=��9T|��++�m�v����Mc��H��NԼ�S�@�����
�c(�\���$��1<Ԣ�h�Kh��tydL;���%'��BK��Pu=��>���ئ'�2\��Z����"��a ����ү��r��o��T�kj�@}3<��`yč���dRG���}٣@Dy���d�_�R�O���o7L�u86�v�x4}��6%��4t����^�
{by� �O���>�QZ��[��=�K��
�f��,��; A�B�3�����VI�԰�Zfy���^�/w�4Р%FIu-���e�ȉآMJ���Xr���D�LPˣ��F��E4��$�[d�����kb?l�t����uNm9����)I������ ����KP�sMZ�B�E�����4_<�t9��<�+���%�a1L&�Sm�F�͗n���	���y����3q��E+��RJb8X��\{&>H�7ݘ��@��y���9����zȻZ��>�������F���1v֞�?d���iC��C����0�I�hc`�M��$��";��i��霶�[�<U��!����+V��*�Űϧ����y�,����G�g�UpA;5�f����{��hM����Z����bಒuBV����{����
����Rׁ�U�ƶ���Q��h*����Np��d��¡��a.u�AE�i�ި�����ޏ�9U�?��"ŵSK�;�̿��UF
��.M�C6z�# ��񪇟��Sgw�=8�[y�Z��QU��i����:_�∙�;�7@NJ����J��M�5�N�b�V��߷�ҏÒ��E�YeA�%�I�G����#�τ%~@��8b���KQ'��_2����>�� qK�(���B�A�A$��rާ�c�VD{��8B15�"e.����3�z��&���c����Sj�o/��{��Ϳ�'[�c�]~Ɗ�A�]e..�2��b��e�s�Ո`�cP\�8p��Y�YJ)��cӲ��5ѐq`�γ�
����9��%��wD�z4�rcY��uQR�͆w��׹Æ�(ns�Ju�7��R�3�. �u\v�;�Q��z� �`}�����]�wg�"_�$H�����묨��V�q��n�{���
�U���^R`�&t�(�(��2_��f`�
`l���*|K��[�ɛט��!�+�����N�8Wtf��G=�s�	��`�z���oP?h\�qV9�%�@c��Q(/ЯU�.����5w)�)�Wp.#;�[�Bu���XUhR��C�(�g�1����
�6���]����*/��WFk�lz
���
B��z]�/���u@��Tq�\��x���M`���H�INؾ�l��i��\<��a�i�g��u^������g5�e��1?��w�J��V�H�@�2�0�t��o�����W}����8�}I!�0S��%��⡹�o>]M�cV���XDs_����?2s��Y�����=�Ǩ}#�~R���:q��Ɩ��w��"��5{6{�.O/v'?nd�r�lV��������uS?�$y��1Ąz���oz/ҿ�QB�1L��8�.7	ݩ̇Af��J��u(������ ����9V�i߮8�kt�H���Y�T���ݙP"��D8�ZQ�ђG�~0�F���ٕ̅�_��AT4�F`�1;=3�!(����2�-n�H�Ɲ��"����L���zDsDV=��,�+����G�	��q����.�}�W�)�,�q� Z�����v���v���sB&�b��pu�@�ㅍ��¹��S���,S�w�� :l�����\��u�-?�5��?#�j��KVJ�~7%q2��W����4
�s	��Cb��o9�[:�G��
��=��m��{���0�!|Y�ݏry��鵖bHév������=ԗ��`�t����K��B*HC��VFVg����i�j�l��l�2�*-��1~ߪݘ$(�d3�U�������7:�}�]"M�w����}�H���6�z�G�w�I :랴k���f�L�Md�U�{�b���vl1�D��JT/hJ��ο-� �Q��6n�:�g1!����Û���)���������=ôU:����΢A=Pe6��
a�K� �g�����@��?�����||�L���Z7��<EKnU��+7���o	�٣OY%+�K__��s�4l�KL�6.��z;�����d����۳�4��c��gv��@NȲ���>�&e�j@f<��gML3���ΰ,��#�Ű�A�1�d������}�Q���4�_�ʟDU�|o���yc��J��]x���U��h���TQ��E���\M�W@�tt�7g�ɒ}���R��$��8�;���	��H4kn@���QM+�,~D5�vQ��	����b~7g7��@�2��1���d��<�-3{���V�(�i�Q��t�Lț����l��>��&�H�\���V��m�u)b�kو�|F�C�����-0��[v˼�y����gT��a\����-�0�y�p�]i�e�� {:L��u['�;�n�8q�V����Z����\�]Ҥb~"� ���^m��m�.�~~�� �ʬp;��1Q���ѯ�^=/ ��/��֯����A�����ƝY�[�=&h��9�|3 .m�.�0���YZ�t��g���:�.e[��9�����"YK�rf�q����d$�;4�q���ڈ�?��q������Nm�t^s��~)Y����@9�A�!�𣾎�qT���Y��w�ghWf
-,��$]n��t�� �[��ʩu�@�;�s�"�� 	t�,U�if7����L��x$G��R�Q��ݎ�?��8Y�T񩱭��_䑌#���aq�Y�ko���MtT���{>{UOx��/��.��垧z:>���k�:���N�8�UETV��vӷ�D�Gua+�>�%�!Z^oդL4�)y͕F C�_Z+�������J3��|�A�ԯt�<��{[^��H�;C�X�<|��b�R�i#l�6ha(��s@�kl���_�&���x����z}RRG8��H
�r�"�����c�5ʠ_��\��n� oJ�#���_�f�_�u�q1�ɳ�C��M�
�0�:9��(��68�����9>tz�FR4s�`��VV�NS�?\�5��S9mf�y1	�y�V��p
��b���a��E�3��$\U�]6P� ��J�Qe����Mf�,���A^�x2���F�O��o�]���UL?@p'���y/�@n{8P�<��I�!٩f�Pu	�?Q�-f��Ր��+�v �����[Hɉ����G~�ߪĄ�X���myL���������L>�M�:�*j����� :��:��K)>�$J�\>�Z��g@y���,�e���-!"�e@8U� �GR[[!�I��{�<� a�ۇ��8�(�Sа㕷*b�Sa��� �4������ߜ�b�� 1���i�t08���Dx�S	8�(fo��S\�9���W+�|y����wʅ#"B�)PYa�T@�;R��7��K��C�Z'_k^c���}A����E����^�.�R�lDdj�7��ʾz�|3�[E�~��"�����S���s�'���&��G
TV���kj䰀�AX�"(3�`)�f5=�,�G�x������y~A$����QP�@U�4c9���M��L�*�{z��Va�s�����z��3�+�H��������2�v��#-�S7�t��|�P�({�I������k@є�\����S�vgA�ըx�zP�����Z�S�j�bm�N�Z7�fN\�i���!H̱Gx��to�:օ��%�Q��:��$��s�v�Ed �Tn$�,�ڠ�3�2"�N�~4��>p��kS��a��G�*�5'���)wG}�JD1�"O�C3-��*6��k����[�M�E�Յ��M=���@���T��������(��ǳ�	��m�􇀞|`�o��ɲ=G������/��f�<�I8�<*�dh���d���<(y��mG�@�#o8K1�"a�H=�̱�*��
z�?g)�?L��K'�sŹ ȪI�ş6�tX�@��rą�6y��+kO��ѵ_��z\D�>��'Z{Ԭ8�!~�3��8��K`��P�M�Nc8������[�@+Ƹ��Rϝ�<�~F�c�(B�҉r�s]��Huv��0���{�J�(L+�0�o$��:<p���K������ �#t��:�Ѕ
c��>{��M�ׁ׆&��|JG��>�va�x�����}F���L)�`Fp�����a���;g�����@������..`��r+5�L�wܒ�x���1DZ�|�'\Z��\�؇��v��޸�Ib8k>ij�f(	��F�T�GN�)��p��/
:�>���b��D�M�eP�I����'���vë�6]NkP4{��Hg�ٰY�f��p&�I�M1���}-'��R8�εM5gb��af������P9�l��<�/F&b,7��2m)!��t���F,]�@�9��^>��dg�C��D_�������^�vi�)��7��Y��'��8���3��`Vo����Fʂ�ꄻ���Ÿ�1e����𔭒��v��S�2�*h-e�ؐ�U��H)�k��R��=oؽst�R�/I���~6�-��� �s���/�%�yhx��g��v�0uLIt���[����{5n�޻t��t��Il���2�]sI?���ܼt�u#6M L~�����<_���w��I�c��P��4^���-��m5���`�1���� �t\O��A")�chܬ�g�F���	;
rY] Oeف�dL�+�@'��0����F�a�&j��+��|&/�u�*��@a"�f�� R��X��d[L���E4�����I�}�Gk>���ckvA��wӞΔ}�S��w`�}�x�l��{���fn9"r�,��*�CM��u����E\�{g����*��7)�.9��,���a�.����,?. ��& �/[�F���1�˜�r��vG��6&'�B�e[D�`����.Q`����-��V��e�H�%d恑b�4c�aFP���x\�F���=+� V�~���,�8�ش7�޸Z�,`����v�E{�f��.-p8�D�Ð���34��KHތ�ѳ�-8s�oz��KJ(`��E��"��fUi��E���i�� ��	 G��U�.�Lkk}"����LO��j�y��m�)�M�򴿋ƴ��=���×�gz_pCl��\�w�%Y�g�G��,��0�(�½�%��W�~�bJ�φZC&�́a��&�\��sw�5�<�.[�v�ʮ�`�^��t���{'n�j����_�
�ƥ@�h`$�Qԉ�1إK������hq���9PN�]j���˒��2T)`B8����tJN-�]���)�+���_�;f�<Cpq��l����ڲ���.��Cp����|��.b�+�Ff)�J�`�`�9p`DIS�-֦��d�|���}S�B��֕�[�=��Mzl�Z]s��ԯ���rZ����$���I�S�� ����+�o[
zՓu&|�C���R5e���"*DG�zm�8�_hJ�0F����3�|ٽ��o���+sl���A��]?���aoẈR3�/�H
��+q������\n��P��Y�/.��̚x"���A�h:E/	�F|�|���sa�J'�~N���@R��)�A\�y?�	��.7��!yUG�{x$NQ7��.�Q\<.W��i�-�ax�ݮ�k��~$�X���Kp���c�b�Y�����{��|����"�'���4�>q�w�L ���j"��
�@�\����ם�KW�h�����/��,��ǫ�1> t������yAy�`���������϶KN�R-g�9��%+�c�Ú�
�:umn�I�"�MUrzJr�c�ݵ�n�O�:9kA���- �*;�$A����"��M��ȧϝ`(���H�zTg�
�
�3𐺞ƲW��y�}`�xu�#ƣ(��@1��xg�z2�	6�/��
8,���_2��1o� *-SQk������gT�hb�!S���$չ�{tG��.y���g�YuM��Ij&]b���
W�{!Ȱ��N�p���aDU`.�H�,	�H�ky���h�u^�b�������in���|7�c~�I�z��CK�U����%	AO3b�O3_��K$⇬�ӭ�{8�L;GJx
G�磞�"��H9�ϲ4��n.�rU\1�� n|�: ^��|uú��0PJ�Dj����̺Xd�~��G��!5��1��nj�p��\�[����B�^���}���6���y 	���_��ſ��OX�ԇ��<D�Fe��g:�j���&�O�����]8}}Ιg_��0�/z�/�&iRmJ�Аӵ��x�> �����bÇXn&6%����d�s�Un�P_Y��EÌaɭDzk�K���h�I,����7\�H73�O�ڶ%�R���vԻ"e��MR9�� �[�W���8my��2v��R���&ܪ��r�r���|�a.�J�D���"f���n,�4WZV9s-�Z�ҏ�>{��ƃԗ����Ҙ����sMK��8�"�0�=��>���0*F~p1t/Щ����$7�<���4E`LW��x
}���o5�#yW��`LPƈm�|��@|�"IWXrم6��v�A��v3�Y_��cR�	>ҹ���L��F_��+���/9,���W�-+�a�ɦJ���'�Q7
���r��{�[�R�;l:�'DhFoHQ"Ng���#;�,��X­'�llƙ:�z���Ja��j��c����8�#����6C�U�vQ6�Gn{U�i@Ǡ�>�	�XtD\��w�� ��3խG�9n͉
׌���M*���Qݣ\g�/�:y=k���װ)�� ��0��-=�XtuJ	�Ze#�s��|�``�}�5�I���t�k*Qoq��N�]�`3Ux��v�AZ't�G �B��T�K
!����Pz���|�}M ���B�+ �N��ݱ��0_�W�1S�`~g}�}��?��i��!���OJ3�6�K���#O.���C��i*%b�?Ɲ]��MJ�6��+0��JW6c�塞������Du��h�3zs>hDj��϶c���a��]�H�&c5c	dj�
��g�Hv�Lf(Y"z��~rl�Q���pv��
O0��+��f�~av���/��.;91I�;�S��r����gV��(��{d���ؒ,��{��2I�O�{�"�G1ŏ�������z;���Y򙃰��a+�+)�2s�DƁ��u���D(�)���t0��� �����3��t�n��e֒q��3��*��tW�0�D-�u"!��5h�i��OG��<����L��Y�fb8�.v`�2,�jʎr����JF-�w$�u;�K���'"�i�
B�|���=��@ 0�����yq��@�d��۫o|�&��(�� t�]� Ŕ��{p߃ �#fKĤ���v�DI�sQ�����3!*�/�m�V$�6���|M���(La^������(\B�m�� B�,o�uI�����3�>��{�~�P>���M[_֪�wS)����w�T�~Vt~�x�����U��sH����)��?Uj�*&�l�E��x����|/f�c}ܦ�5Fl���<���[�^��F�o�x����B���E<Њ�<k��Ra�$�}��hq(��fQ1N&���[��DGn�z�np-�"֐�R�ɘnz?�is�u�Ö�����ܝH_C��2V��e��+
V�н�L^�K�f��4#k�cP)0���3��tL���f*
��vHF�����/���	e�����H��?d]+�	��U����X�V�ڬ%;�Gn��un`��_�3�n cP����aQӎ�|�YoT�g�G��J��ٕ��c-��
X�v��il�c%��{�$��ػ��u��I3hSU?dY�K���O
��(�:7�+h�p���㳾!øT�7����Q�ቡ��[��hc�':�yoܥ*�p����L��I]���PB���F�1��\ ���{2�tDAɺ���=���$�n�
��\2/�����	�Α�Х�f�o(,�{��=1$�|h�c҆cG��I-"���~6_�bBF� ��]�X�;=@�Rݣ�Z� h׋Γ��Ֆ	�μ@h��F�If{�D�������}��/v�/�v/,��H���b��R�@>B~��1����/YH�p�]C��P�CzY�b��������� /Z���Z��@O�{���,����F����$z�}zE
��<B���7Q �מ�����v04��'�&B�+���o��Jr�7eF>�ʷ�����:���ٳ�4ݎ��۵�:���f����6�4�#\�76A�<�ݱa�8�_m��2uB��e���/�Q�;<�IJVV�K4\$�}�<����ru�ؠGl�Wf�n�Z��� �?�Y��8N�Wh�F<DGX� �M�2$��IƏy��2��s�FRlP��r&KY
�Ck�@܅
�h�AC�SM�����s���K�Ȓw�p'/x���o*��Ԩ���N��0�Y���v��e"��`�_xi��в�0i 3|.�b~�.%Q���/�a&�Ns	�tJ�*��������<a�];&�
W�H���2c$0$�y��^�0�ئ�E3��`��5���#}ջ���U_�T1*���R7jZ�����m�&5.�	����R^�^�pZ	-� A"�#l�g06��񦚵�6��Grʎ��p���=ǘP���Wl��k����et�]�y��<}4�0�U*"� �M7g|f�}<ZSт=7��m!p�ƭԟe*�Α٩����&�|k
���"�΂�������K�З��fW���������SX:��J�%��!q"=���u�v�S7��J��+�rZ~N]B��F"^8�J�d���c�C���	����"1�~,��X�c`ӚN(nX"�M�'�FE��X�����	]*�.����^P-7S}��`O���U����oɠ�Y��^6k���t�&)E��G�WY�tO��Ɛ�,15i�I ��.3A��+��4}�w��<M�#�7�
6� 0{��74x�9I��ɉ/��3W�����X�զFS���H� ߓQ�A���l��Q=2����>/��A0��ڀCe��̬����w���\�C��h]��fOi�w�����j�hxфyS���.��@�E剧H^��IqN�����f�d��}`��P �� /��v`}�;'���=}�wg�}͊��l)�o��ʄ���M���������G��s����R/*��6�!��;���7{��Sݓ�����}A�?�be��f��L�½L�v��˹�p��*��g`v��E|@�H�0D��~%�WN�Ln\ݽ!ˮ���>���ͥ�*�^����0�I�a[��FXh�p�ōh�O�tm%�C��c������"Q9����ϗ�u�d������v�/�7}a�jKO"';����9aE񅜥1;&	�`n�C���EC��T���L��|�1�8���6-lS���	��/D�G7�7w�%���tpp�0�ʟn��PY���?�p�e�ϥ�b"2��ߚ��Dj����lYNnPq�w����]�����N���[��P����'ԋg��Qk#�^�r;�z�P��z��[�Y�C�f��B686�M��Ѻ X����FPi|%?�XL┅�ր�@�����F��b,��@KdY�<��x��X�����+��B����f%�I�Y��YD����WA7��^�$Z���?I4n������-��#�"�q�q67/��SO��g�6��&y�4j@{e���Ɵn��;p/��;�lYh�~��eȢmz�Q�%W�GeXt���Jݵ�-.�F�6�S��}c��a���r#Q4�/��$XR���uxe���&U-7�o+R�QqUBۡD�F2m�Y@`�`�0a�9F�$[[�y��G?�6���p�ؠ�ޙFL#�S�M���i�E9G/7�Q���x��౟��S�!)Sb����!�|t�(�����<Gqr�&=%6���pN�a���� l=m�,�Ã=d���L("Q<6�г-N������9�q�����E�޵A� �-V�А&�_�:�%�v����F����kE���=i$>bz�Qb�Ch��V��jB���ߊ�'�բ���3�����t��Q��s�Nw:��G�s	�5�s�4��u;M�����)3��97!�8��ʯs��!r�k�7�$v�L��n7��X'?K�L�ve��@��/oޜ�H���0{�0ӓ�f��*�:t2!�Em�C��qF����@�|{~|���*�����dr���S<ŏ�8�3.�#O)+��4F�ZG�����vK��]qţ�����usR��v�-½�,�j�b'�|���������?BPFg�(l(��m��p��k����,�)A�
oạ�gb��K��w�u���+:��N��>����;#6���r�Vǆ`jZ�	Ŗ��;;�b��P��Ԡ�0ejta75Am�i��}�
7*��a����3%����d�ڧ8��c���5=k[���܊����0a�@��1F��������,%�@�F0GR�~��Z�hTI����,�)��b��W�D<�,��3��O� N�J��<�Z'ֆgF^��ƃL����51)�&0���$;n���QuQiߴ�C���Tqݜ-AJ��`�]�T�c]�B�4��	sk�U0H��ڪ�P��b�L�L8��ͽ���o"���!��c+����
	MM�ϾA�����
�(�Kr
���ef�T:0��B�'}5Y� ��[E�xn�C?ew�"�L`9n�)ޖ��Բ��3$��	]��yڜֽ{ACՕ6!��ɟfr��u5\Ma�f2iuA���삙5�����7��E��M��>�Pym�ed�0w��B|һ��ڡ��΍����AX�1�:�T��X�M�"q�5��s��|_�L��4��7�:U�k�jn�.����O�mB�S�1�錚��gs�1�B�nlO��X�2�n|�,z���-x�E�`���.�m��:�|�l�#����`����һ �	��[I��Lh�P^"H.�ϼ�4CL��OMq���Q6�4�ЯR����5��'�= ���ES
4r���Ũ�/0�:�
��d|j�����JO���a�i�	饵�{/&p��t^�*O�oJ&y�������#9�O��o���Pm�ϕ��Ϲ���L<���K���K�̗xl��g���*�Н�m�J�����;��p��^�uc�z'����%y-_�I���O(��I_���Q�

K�(An�[�׎F�#���)������4��O�$��}e�Ct�QXo�,C������E��R��vk��Fn����}e����?ZB��| B뚜��er��w��vqߡ����@�	qAM!��>&�v5^�Y)�8����~[uK����?����C��P=�ׅR��'~��e�@��Q�\�o؞sTX��!xߠ8�{r�!��sr���?$	<b��N�%�I�Y�K�S���L�?����o�Q{S���s��yƆl4y��eH���Dɚ��vy����b���������:3b{�i���q����J�޹�@�=|S���k4��D��زڍJ[�. ,�S���� ���ЊtMpن���I_ P�(M�'�݋9� Ҋ�����j�M"0�X����l��թo�u1�
���i0���BZ��H��|ԓ��鏊��z�<�H)7���e�BJ�7t!!|��A�B7�vX�!�*40�ό�2�n�v���N�ɔ`�����Y�&����v���CN�9޻0�i�i���d���,�K<����L�!JVa�!�(��7�g�A ݈U֌d_��Yy8�`Er@!��5���_W-`����.����ӪH����&R�;=�+!�@��	3�^�^G�;Y�]���2W� 7=��������0�� �� �:L���r�p�I��������gX$\��(t�@3��5�L~�_$�!�-���D�kC��jִ�|��Ԟ�"}?�3
~^�V� /�p�}�3"���]�B'�?fu�D��䒒��f�\���p����`dܧDaf����@'�®�BP;A�h�wzW���:�ƻ�ό&��H/T���9t\��M��m�E��?�:���ޑ<� �E�!&�Q?�DLǫ���>>y�7��(5r]�U.�4�%Z�t�N5�R!~����fn�7�똲�`�3ѪjG6���G��|��O�UN��u�񁊲U�z5�O�����L�x�?*���&,N�
~����>x8VM.��O�W��u�ԓ�1O�O[H��Tf|�:odib���Ac�[͓�U7�֘�j����^�'�#�����j  ���{�C��(�*�R�ݪ:�vHS[�u��B=�u��2�xB�ѫ�]�y���,�jKX�i�z�V��%}��9��]Dg2����Dn�1�Y�,�{ <{���E�h����,v�60�Na���=�5�F �I�Nܥ���[�	�R�P�i�p%hc��N!� ���g��<�R`ɳ�(�7 �p�eb�j�6nށ)��OZ���S���p��Y�: H�c�q*vm�a��[��14�X(�l���9ǽ��V�67ϟ�b�}�]s�j��k��ETk�x�BPrrş������s�"��G����slvB��p���S����2�M���J�'4d� �u>�gznM����j�0��=8$�������į�b�~U�������UR��c;&��$��BNM_[y3 �kRy��Ѻp[�2[�B\����MĦ�fz]� gV_��Λ|z_�$R�1X�n�Uȸ�	��B�%�Z��e���g�s�9��(�O���8\��HV��(���^Vc��n]�F"�3�*�zE���4��4G���>*�£�J�A���zmm����f�\v|zG�M0��)ur�'����M}�$@���yEnF��D�#L3U��%��ߣĘ�@@Bu֣�i �ᅎ<����H�����m�y�X�Xӧݮ��y�0��g�{�SlW��w��֢dMb��b����&^�����i��QO��d}qADd��®���+��?���r�{�[n�s*q;�~�t{a>)�laO˒�C��<dPlC�!O5Tג���4������Z�_���G���������D�/Щ&�9I�LOo��X���d��j&N�F����FK�:�e�ډ����������뱿�ly��
�lt[��t�xM� �A��DЗ��~��va� �	۞tF1�-�8m�&��-�u8G̡R	�uw3,������%�)�s�����~�o߇�p-��.�q�
>��e���]!G��M�]d�_YrL�;_6p1Q�rw+���]�w]�嶢Wcy��+����D
�" �D�0�B��s�O!�ECń,I��f�:�W�JA�PN�c��Lc���j��0�qH�yl{)V��������>\�H�a�wԾ)������^x& 7cC�^�ƭ�W���t{�]�}-�� �B;w�(1�(ȭ[�Y6��x��tK��U���I.�y�V ����xT��1�/c�%u�=��'g-���[r�q2%F���S(Dx%5��R*3���]�|3���g�o4]�����F����/�|�Q��tЌ\HL,d���=g�|ݠ�`��F2_ԞB���"�4���&����+Q�fV(�/ݮ&��;J��-���~3l���z`\9bN�5�^�S�ԕMUp�)�ȧ|Bl�?��V ol� 
�=��Do�6Bm5&<Io>�x,W![��=2<���i�����-�I�ڷӉB���(x�>4��C?1��?9�����������s��ݮ�}���|�C1�Mú�W1w
�jP�O�'��i;M�qx{m`��{�Td��f�q9`	��9�J���p���n&v0�22&�:8�!Z��_��l�H�3I��w�"FT��������`Ob�u�:��r=p����&�nӗ�z�#m�Sp��S+���'�)bȄ�T=6؀�-�F��o���R�Z��Ix�5����i���1CN/im�!��)��8������$���lr-��rD6/H8��)��E���N6���n���c�Om*��@&�,��%�?%����B���\��b6<ó�a6<��<��0٘P�&蝥�˰'�n���I5�唐/%��	d�el_?ݹ�z6�zp�D.ދus� )m�kO O�3�ޞ�p�疑c5��9\�����ܙ%�� =ҡJl%	DF�暩߬G���BI�0�a}Zф�݈�^��?�S̼�T,䐊�r����G���O���j$�������T}͊�J�azdS���og�C �M}�ʏ�ӝ�'���
(�7�?葃O�"u��G�g��������C���w@��2z��Jk�)>[�] >]l�%�7�>�����td/��~Oge\�S�_�{��hH�J.�0Zq��^��Y1�ae�1 �Y�]�I{,��T��~o������1�3zP�k4�y'��Ѕ��k3B?*6z�y���i37���G��|�w�QV�8�_�ӕR���6(��0v�C��x���t�Z|ժ� ui�'�l����uX�B 9)J�b�����-��L�y	�5�]�h��p�Sg1��x����Y􍧥��I*zS�~%oI�JU�7��v(��*d_�e}�S:0i	:z��X}��^���-�X�g���QL���i�_��נ��~�_��q]酼V��O)���(:ɱ��壘#9��;/��SE�N!u"�/|͊S�{�a�ʔ��[�X�/�x>֘]�V�I�n� ۞I�?���}�{e���(������|lb�<z�)���z[.C�@�Y�Xh��)���R�j7���rd���̾�%r�l��Jq��Yt�Ag��Yc��G�͍{�&��LY�˗;��|���!U��RX�4�Q7�z�����1>�c!�)�q\ܫLɧ�K��8���A�`>=�Xk�o�M0�i,�8�o:fՉl�\�����U�d|�(��4��d�����١���U�d/��[c|�r��\�T��yK����%�k�P��Br�t�����ɒ�T4�C�W����E�qE�#��Tņ�5�7%�����"{Qa�����E���<�` ZT4��))NIp�����c��0)�\���w�J��:q&s����L�M7O;t� ��
y	�~$�u1��_�˘�ɵ�N�+,=�%fh�\�� X�o�}ocq�	٪�1aw�5�p����B�~�V/�]3r�0�5Rz�hy�ZDp�������=S�C�/��X�`�w�� 3�C
�ǘI����Ƕ��\�l�����QKI��w3᥅7� ���=���v�ldV�l���݌FEN�$]�$�о�dϪ�y�M���� �5�	�F^�x�YPO4ke�{������-w����L�N�zQ�
1�'��^�Haf���U��/���H�ǉI�&���S�-K����)��8�R�r��Bv����p��;�d���@���fr[7��7�	���`9λY絫w~#��3!��4�L�hsf�<�(�9�/3��Lzb��4�;���I�l��`D|�
{!i��v�!��i���$�0d��9���Y��}��"*d�KB9d�r�CM}=����@�O(�z�C�[�)��k�����m�}<�9�����k��Cg��-�|b1A�6�u�3�+�),��h���ZAI���CAn��(�/7�E��q�Ju!����s�.��хWQ">cl�lۣ]����I$�©a���G�q^B��-V�B�ZB�GrB���3���:��"�2�M{�"T��F��(3���f0��na�R���R�R`|^�e
ޱ-,�j�Z���]�L�ו�t/�	��m���e��]5�E�OM�1(�T��q�P���;��H�*��M����1_��2�>�W1.���� wxXx��b6�`=)�Pv�}8��w�NS�[C\�k���Նr�W�'���� �7�fl�l� d����lz�2P�1�K�u�~�� (�'X�����x��N���T���L5�O+������o�n�%���e��T]���eN�`��ͬl:B�����z����0mj�S�����.�K��k�[��	�t�Ln���|
��Dr��PX¹��}Q��Ƞ�#,�G�p�^ ���m\ܣ(Ϡal�W�0{�(���;JmU��}�T�T�LXr�M�T�!�~�1+��9�%���xmgn.�c,��@�m�?�i09ᣕ�� ��ӌq����78���+F�Q��!_�a����8��;�J��.�3W-7�	C�����`[� �Ҹٞ���O�[З�7�D����h�b�@g!���VH�1J�� ��.�A�O�:ٕHc����#����ME�+n�P�1��ai�Kl�6M���-ð9���K'�9%DyxY�zO&�#)��k$�B�*O�)������W{�D7ݕ���T��K_�W���7_��z8N�_3�$�C�j[��6g:J��;SW�&	\U7iT��V�R�^t|�����!>�{�>����_A?�_Y�;{�d}B>�9���69�MH0pL�)���^ �9��h�d+�;�������bu�a27Ҩ�N!���d%FS�V��T����<_d/U�[s�es�/�Ȓ�(	��:C��!9_`[
�̅
�,>�a�����_w�v���>ǹS�AJۑ��#���r�L�����e�[�H���ߧ�mՈ k�(�'�@7LO�����]j����n��f���~��n�ü��G� ۴�$ձp0�A�$��!LT�S=�D4��eoV�z"g����O ��Ғ��1À(3�}�F*�D]��v�pZ�Vׁ�4�j��}��ZA*A!��������>mZc��U�4墣�n�ob*�"Ry��Dh�U���,�m�gܣ4���.��[�WdB���Wd0-ݫN�[��n�?�9�Ò-�;M�3��?�����/_s�����ѯ�/��đs.�UPL�W{f$C��C�*p�C=�L�'�����[ԜyJPa7�,��OQi�����>O����?Z>7��ѽ��u�2��"�S��[�4��G*�7� �C!�|�?gՙ��r��<�̚�@"*l�!�:��i�S�@a׸K�=�lK^�X0�A�I��� �x�oGÆ>���!�RLm�h�q�E/CV8Tڋս?A2���s4�2���x�������Dd�Le��a���t?��"���җ��c�xV	��>yl�F��Vőu��/�~�c����q�jW$a٪3ljL7�VYX56\��A�Z\g�������'���c��m��>���V}��51�?K]��Ql<��&�sj����e�/)�ye�ϷPP�aÑ�F�Iy�bplC���x�e��jm��iGLVEi`��>j������4|�f�n���Br�+`D��
�$2���k�n��*\7m��ʛ���΁��t��>���&��e����u������r���ƴj*�"F�h��Ȭ��x�%ޤߥ�:������:	�_v���5���4դ��Ī���fx���*��=4��oeA�ܳ��bN�MU��u�1skT�6�bNS���򥓁���~o|�%�X;�fʝn�lt�~99�tk�#��×��0�i�(�Ӏa�6�×L�+����Ɵ��K�P��7_ʹ(�`��O�*��S�^J�������|����@c ���o����5�v1>�6�W%&���rFYW�!ݺC���4�I��M
�S%1��^������aK���G� �8��w��Q8!1�HV�ޡ�	N�ڙVӡ[�;�T�B�f%Y_5^���Mb��39�ʠ�9a��k%��{<��v���#����+PEo���c?Kb�������=�M`�F��|h�#�O}�[��y+������sZ	�8��f�	��;
٬�����{6��[���B�N����]7��ْ}k�9;<7�y�������uQ�f�qlS���1����Z���6�n�v$}���� H�JOI:�Sߦ���Ϣț��1TD<\B7��@�b˕�l�(aOBn�^b���hTE߆նH��'�
�P����xK��qsu:�d��jXOz�Q%}��{����IZ�fOZ=�HA\��2��"6��K}!���W>�ڞ&�L+�p��?�} .�����	?L�ũ�����+�UE��+(HR�(�Mw��qؠ>1����y�{�"}�%�7DY�!F��5�-E5��[����������ؿ�b}Z����O#�E�n&�c�]�%��t�,�$v_�/��W���n`�������/籜ȴ*�	Ď����йh��P�=Ef5đ��M��\�?=��ǧM/H�azg�M���}~��EĩB,V�7�����	���D�r2�8�Yz�z�S���M��E׸�Y�\�5]R?9�����	@%1T�� ��Ip3�7��r�����7�/M�eS/��djH
�-懔���o�&��5�����o���/6k�h��D2)���y����<��2'K�#'��z��E��{`W�NH�w����7�Y]{RB�xj㌽�+O�S��_�\Jp�fh�� a��D���|��e�IB���J���A/��9�x�E�b�.,��m��.ab
�Ā���M����׿>l�7�3�&����;PsJ�'����Ry�bt|yvZ���\(
���[�Uf�T�"��*B����B�c?ujg�`�_��,r'�>b5f�V����P��6O�;�,C�2w����
i)�H	YֶgKo��������r���3���В�#��,�u���u��&���~F�����LXN�������Ήۘ#$�����r�0&�kiAa6��,n}�A�mI��P��~���l��'*�_(�P��<�v�V����=�����R��j�C�qu���z:��;��m�{��w�A.i��|}�nI���1m�X��z��~����	T��ms�u�x�9���,Xۊ\��X����Z�)��v�` ����"�����,�H�V����s���t|�l���7�V��HEڿ23���~E^���5������Vݬ�姎~��bG)�3GiQ7H������G�aoېx��^�59��WN*w��A����[�P�C����fx%HQl�UA������o�������I�b
l���C|�כ���ܤ�����^�{���Л���h^�����Hw,q4�2�M_V����!hN-C��e�N�C�˞�?����\ 1�e�et�q��<�fb?�BF�Ek&u Ƀ3�S������I('�������,�.@�z�R�������w�7_�`aeܧ:
	�3�v��b)m�������k.`�0Z�nA�[K;eZ#�<_���L~XmC��$�c����ґ?E�ɥ���0Q \&�Í��5�Z���A_4;�I�<X]F�-����e������І�����VE��߮��� ��J3hP���@ۅ�>��X�R�D�;�T�[�cC���Q5�C���x���]�P7vZ�Q�����&���������3�a�8�AȤ�e�)��{I��r�I�\ ę��9�1pj 뮫?/�6�&��8�T���G:$��Ғ��Lֿպߝl��:��a��[� �6I��RH����S$��-a�g��mzw�L�_H}�Wa�'������3��=vyz�Xbh�2|2V%�i�1*Y�:��c��]Gs�e}C��j�g# ��T�3lE`7n{;�3.o�G'%�-?Y!j�"���P���9��j߫i�Y�I�4B�� I������F�g�X	bl�XzWZ[�"n�*�#���vt,\�������H<�7w��P�97m�c�d�I���WE��?�X��ۼlր��x�]�k���Lu���VD�y���ʳ3q�g�t�z"�k�-�Ok�lAH�%.bl,�$����f '�ik%u	'k�S���V�`C�����[y7���Xon���	�HKM�V�`��˺�!Is�Mb ��R����a�Cʂ��x�/Y�Ŵ�`0��k����Q���S4.�bn|�������%��OZBd�r��]���6�@0�Y�O9T�p�9|<b�`�c�k�����8P�J��h��l1x��{e�H���~I��N�ن���pB�r���>R�pv��v�A�D8��.�:uY�!�{jJ��ꌊ�l����Qw�BL-���x�aq�lr���'檾��뚆:_�9��$�]��hC9\ؐ�yU����'��%ޔ:�;����ڤ� �(}�e�=$樑_�x��T�;T��뿊x7������sz�ea!r9�{[c-���|
6�M���QC՗ю�&���pZ��m~�|H�92Q���`<3��,۫=EK��5�R�ġu!��r�=��׌lU�<��g`g��蕫�U�(;�'�P.���1	��i�%c��F�eM�j1(G���y.�b���
�ڹ�C!aA>y�&��
Y -�M3i	���jw7d�D�׻yDO�ߠ91���N�@@'�ˡ�Jő�G�E��[��l�������>�c�b�t\��a����ͼ�'{T�~c�' mh�a[���DY���M߿�f�T��G/C=���q �#���8����"��^�s|�v�kUP0 �f�D����N�,��4x=�s	l�1Ib�-<H���1x$D���RAs0�)?�CШ���Z�ܶ�c�V�Y*�M�84gt$?c�,G������R�\$�q��1>y<U�W"��b�8Qv#<�ǝ����X�_IU��\Z@նÛ!���a�Yޒ�I7I0 #��l�k�0y�R��}��rL�P��I�&��d.n��e��+����Ea=~����G��e��N�S]�-}H����r�R��J��~!��=L�ȝk@�`��Xgq��s�ª��7�
�񳎓 �(�?�|�I~��bN��G��U�h���tot��,�V��K!{��]��ƹ1��w�D�z�pw��&�5G�r��~�4Z�[���¨o��$��~E��H)_��IhW�C�͚�"yB��f�N�O�,��?�Tyo�b�ne��$\�kh�����4>���/aĲ �q�
��5�&y��̯�<[ޮ]��r�U���@��|z��hn�F�uH�=��~K{AZ����_WQ��jz�<`�an-�|1�ʬ��O�m�c�sb�9�!��
j�h${!�1$�F�K;L>1�L;�<��ƛ����/��vQ� �E�y4���ᐭ��jO� �G�l����E�Lu����o��E��~&�QG_���J��'p�-����Qd
�u�俢SV&YO�f���OI�+,��3'ؒ�?�fԹ=~��R��'lA�y��ξO��ةi�xr7���I�}���j:��%�"�z�A�͟2�'c�ӫ��ʋ����b	���ErsP�i��e)�g]����H���K>^[��I�����941X4n}�F��T.����>KJ��t'���9΂�x��?~U?$I+d��h��<��l�9��g������_�|ܭFfj�=7.���CȔ�Ht���IV�(��2��'���:l�f�t�����i��H�������q\�ԧ.��"��]�R����@���\n}�}���9t
o�7&�3�JB�/��X�JM%t~��}��~6����z��ư�����U b�>�Y* 	ͨkZ*>;�']�EC�u^RY�e�m��:<�%�t��)9� D�@\ ��2v�R|_'�b
����C����\Z��}�a��-��/��jm%p������;彙G��o]�K��#[徵��I�S�}�u�u���g�}�3���8�����J�o�1&ô�����{��e���$rp�׻�����>.�+}�\yy�T1�B��8�����Zu
2g�+�B�Ɯ�W�!<���B_`�\��%�8^�ٛ����/�-Y��z���L>��9ruR]��"�u�i�c�}�!J�E)=��,4�-ȀI�2j�X��)�v��7�����R-�U���y#��c�D��S;�nG�����|�Vi�G(�d����ZŜ��mms�/3[���&�P��a��G��N_�֊��p���H��5I�Kы{ ����V��:!J���A��>#���=J���(�v�Ҳ�<*��b�����h��Ԥv�ߕ=�&���N�U����[�ȁ�aqy��D�HyRE��Q�G����)>s��ef�?*-�?��"I��BF���l�=G�P��)�ݢ�9�b'#dY��&���)8�4#�A?�?&:�	��Hs���gز�#r.+�*󀁢�&� ��H��I�W��2z x��gɾ1�~�� k��_��_�����-nc�t���U�S"��%Cp+L~.�C��H�g�C�<�+��}�'c�A=,��0�K���
��HH�zt�.P�0���¹Tm�A[�h%��J+k���8M���Z?c]�Xr��#����@� �����j��@J1�4��aRdƝ3|����V=��ͯۋ�C�� ^@I � q��;D�whhZ�h���2���W�B���l]�;4{�թ��)���y�k��G��1����h���c���(v3�p�J1TIw��ZM�w�tT�A �NNpQ.mF+�n������i�c	j��ԃ���cVX=��.R���'[W��+5L_�ٹ˭���$���.�~��l�r��O�cj�L�x\I���;/��uO�q\pG?�X����͈7�W�l�n�q{�rt5]T�ď�]ʻ/�f�B?�v�00�F�p�eJ�9c�[�cr�D�9���E��Ѷ�E�>{]�U�Y��?7]����T�<[��ѣ����Ч2�MMh��"��f�5*"Zw�B|S7oTio���t �[������!2.,���?m��)cUOj k;����@�J��:���4z���cNb̚�D:1����V,�p�9Tjc�_��&*��^}7�%���A6�msW��<�wI'h�'�J�6�e+��[�U�0嚈� (y�%/o�_������&����G�WrQ�YB�����N���gX*�����G��cՀ��F��öo��]����Ea2a�m&�ơh���:fJ[v������@	�,qLP �Շ�wZ�k�]!+K�>@����w̝o,"%W�5�i��B���EE�0���Q�����e8���?,��y���q�J�ң����=U�#�1B�����b�o��]�M��[�c&�4(�젅^?�(��g�Vn4�3Dh�@&ܡq�z ��ĵ�+�� )r��9�xZ�~RK�=/��
���DzM��I~Дg�]dZ�D .,Յ���P�)>H"�t?��u�C5na�)�Hm�cj���E���i�yo�`�_�{e��퇘� ��Bl��VW�<Mc]�A�V�>#e��$���^J�<y
D�Xr��-T���&�2&M�2��JGһ~����$:�!Gn��\�2�	������D/о	��;��]iZq|1+0rbڸj+ob�,�ݴ��jmn��#ꪚY���KX��}�۸ϮcT�$>8�f�/�`b�f}�sG�#��kV.����f;ެ�W�J�Tt�lՑ�q����	}ķ��3f�M�张���� �_!������	 �i��x�B��(O<$����d�X��q�Z��X��P[@;Ȋh���Z�g7=�s=�����;vtf���_�!�0��5HN����d��J
aavt�Sv��H��Ӛ�lKց��uW�����7;��0��	�S��с~�O��&_x�{BQf�
ē�c�>�����3��F;�$�nK�ܗj !8~�@��sK
��dC��!f&l:��R�����<�0��w���[���������c�}�04D�eCK�����͉'�}�8:�e�C"�0�;R��b�mӿ`G�j�6UTDr�LAm���u���x�0jo������h���6U׼�꘸��%�K;Sr����x�l�+�� [���KY���`r�k�Ѵ��y����^k�B�:�Ğ��|%�MoQ>sh��.��ch�|�/B�Ҷ�W!���K����p�̶=TP��o�����#3ny�U�崯�g�o�X��?�Uf��K�J�ޫ8b�:L�v�7��[�By�7�~8�CsE�"��qN�<���pd6�Tk^��1Ͷ��&/�d�@��Gn��BqH�;3H�xc"%w+'�-M{y��d��V��y������^�d�����2���H$�W�VI廀����]�����.	��=ߴ��¹KoU0�
Z�=>7�
Sk��-k�r4=�mY�+,�s_d��y�F�/y9j*w��v�Z�dO�v�;>AP/��e#hh��0*�=���7�r�%�V�[<�B��R��Dծ�	7f�+�ea�tٍ�լ�+�Q`ZC�����z�KElBl��F�1�$ �Ii$-QKGG�i�pG�5�_�.�1�$����Q��V��6K3�R`i���c����A�ђ~.�9�����"Ar����X<V2�����4�	�qq^��R|�̓2U���^(n>�\���@�^pp�T �np��3_
]���ڙN�1�ԃ8ت<��'gl#�*4�x�K1 kH�MB�����e���ј�Cp�[��È�D�b���$����2������{�{s�LvtU�Bx=!96�X�T>�Ӓ	K/Iv�i��  uu�H񞨐��|w�����87���_�^�`�;��.���[� TƩ�092��a5;�x�j����r�����-v��n(M��<��� Dk��4&�ůkd$�,cg�1�o�����_m5�zlZx#�8��sF'��.[��J6lf� 5F6i6��F�3(���)�	�r<�q G��o��_S�.N��,�H.#�|�}J0H�՞	u�)�`�a�X�mh�\,�6��Z�"&�B.1�OD�%B*�Sv����P�?L"jZ�K�V˔� nE]���үTD�94=���,� �G�1HOY{�ѡ��X�"�`�R�~9v�߱�|��� ��yZ�W3��M�f���G	�9�$	f�|��ji2rCL��H<؋��>��|��f��I}�g?Oh�N\���W,P���q �2�E�0P
�����P5��Xc�<�geR�Ʒ�+���^1���i k�aAD�s�*c�@]�D���L��>��gY�K9�!�?tR��B}�PW����&"�$�	�BИ��]svZ�M�所�prq���&)k���`	m��n�LSl�.z�%�J���=�-���*���~�E+C�Ts��6��D�~A�.�t�����Lz_U�S�nW����ׂ��Bǋ7U|�(��`���`���-����pN�6Q/V��l@e�1J��c̋���1&$}���A�v$���9�[=�ߍ�y 2�&YX3ǥ��p�j-�������ꪸ��'��d�S������I���6n�MNU���@�z|����x�N_]
�ѱ���7&L']�:��)��P���3�?�����m��4�48B�'�γ�ν�F�Ɋ��׍�[��:���_y�c'{��3�{'��*�N'����I���&��<:�gT��?Sv0�0x=$���?T�7�/$i�͆ږ����?0�C�d�=JPJ���;��
RȘ���k��U��񒤼M�CB���ME*����܋�E;f����̽�zY�o$��5Ws�� ��#�9x)0g� ����܄���E.�&\�P��T,@=Q~U-���}���%jF��@b�~ӱ�U���-,��+5&3�h�z�3��1Tk{������~��?���V��"��e_>xd�Dz$����*�����g��5�q��d���r�Å��jRf�ުWiY�Sa�Y�/�����Լ56��}}��~%mY��-Hy��c�;S�w FG%���|c���Z8`|�9��E�#xsJ~��|���¦k'9�R�̌.�g|�)���j��a�P�<��f��L_%����?�wk���ٰ�4����+P�L��c���aV�G��o�F��`�9GK���YY�9d�`Ӳ�����`v�������t`�������7t6aԷ,���}l��r�r4�~v��~+(qF"������OO(�'A��NuHF��nT>��~/�HS�:qo�0I2�C����
&��B�<Zu��l3�`���M4A�&>C�8>�|˙G��ˇ!C>]��Ƕ{�e�x�vO7��V�xLz:�B���$�mA1g&k ���z�fT����A���M��- f��-���'� rǜ���~3"��a$
�H�R�.�0�M� {$��I*��Y�@�zFZ���F�������(7��{�3�{7fH�����2������a^�1�Qk��w���D�s�y���t|_�{���]�4�d�C���%���;�K34Hm����r�2a8���Ws}��J����A�L �E�-x6a`lv�N�lu�
^�К�=<	p�W�8GR���ˍY�0v��� �(�M�3�wC*�\�E��b~���6D��X�e�Rk؟��?4~��V��0�?-SDIpQ��$������ʦ��nW#J)��<CxZɅ�A�1��0��f��ɦt�!Ȗ��U�F'�vT ���T���.M4_��X���7��P�c�Br�ʃ���kZ���r�hV��x�Ӊel����}�Q�ȚD��Xo���xN�A�ܲk��y䈰mV>�)�2��%�n���)�����y&j�p<$E�vpmd�)[D�00�%�~R@z��B`c+������Q$>�ݥB+��w��jXO4�G�t��19�%9�d�1G@HX�C��|𫨅�jre�Ҭ	�KA��צ�9z�.�п�v�RW����z4}ܖϹ��=V]R�ꖋH�l�W��ti��:n���kW�_(A�ZYy�􄇍:���9��h����$�Wݖ�G����o����,�_N4��-�����E�i`�5���e���4���Q#��� ˌ*�<>��]9�r� C'��� ����'V��f9.,��L7y��3���a�}Ĩ�7ՠ_�ʯw_������,��"i���*��Y��h�o������'GI��r[8H�Y v�����ٓ|�+.{ªt����#Pb�Pz��P>�Zx���uC7�mu���� 7I~ݬŋ�*Y�bRy�k�@��s����yx詝�.Tk�ʒ@¦�f#�TCj��,t�k&��{�vq8��ϧ޺db�g��������T�����5�`EZ���և��5�S��1����J���y@�f�*�>Pa���)�����N�B;�QTi�X����e�M@�G6`ᝌ����,?E	��6>04��A��ks|�䘀�e��U;a��k,QڶyU��ԻK`�EJ�>�5.N�_W�|@"I`+$��'|Y�� ̞��ҝ�N�&����^k��.�`X�
��L� % B�t��yg�z�*��s��t�vhh�W��b2��[��7,�}��ts��؟��S�EY B�A�E٣���8O�G �����"ȼ�
�*R@G�O��"�ͣe&�N��j�d��:��(h��Q�� Z���DǺV��8�_4����7W�`��� �I�vjTl^sh�O�!�u����mὈT�9}��O+g���Y�-&�l0=2�����G��=����4�b�sԀ���������{ۑ���#'�H��]g�c;�g��I���?�4�촮��)�'I��'1������͓�8ӳ���$u轙���h0��K6QI`���a�D'D�y�,!c��(v��k�>�N'�I�\�/iQ'sW����� � �kI�ϏS�����P����%�2-�yq�-uM�st��`W&W=�8��[��%���OO���&q�{������R9#����Hg~j�������?�$7���4=���Ƭ��\� �2��|���M�� M���	2��>G�{A��7�mbD����C���]y�;�z���d\k�-t7߆�~�(i�r����8�&Ok���ˮ�(����'��_��X)�l�^��LV�U%�J�s?`�U�2U� �F��\i����;ݘ�N�rz}6��6������ �e��,�|��ږ�0���Y[��I�t�>
����&I̓낃��'��Y� 	$*��� ��M$0��e�Q�"*g�C���� �Ќ�����D��qp!p��mx�@i-��!�#i�z�64�V�-�3����幚u -�2��Ү9����\o��F�؞5�t�1Ӯ�[���!���eǀ�Q�1�:\���sd��b� 񕬑��ӆ+P&R�Tp��琽A���*d��^Eu)+zJ�|���_�k�Н,C�5�@\��{�g�@��L�"����[�2����2��!9�̰�z��?���AL(����j`ҿ��mD���n��@�J_�1Q1���$vY}�R]�~�1ʗ���7��3�!|s���I)|J�|H�O��C֐����;�l��M�/Ml��"+���
Jg�ʮ�т��-Zb}9��w�:Bj"*jZ`5��&MVChx�ǯY���!:2[��D�	�{s2���7|��=$�y)� /�f5���L���π�s'�'�Ӹ��orQONJe����n��Lm$�Ć��^n���D��;�2 �eHjN�>\�5�~�H��w�H�C ���� �ŉR�"D��2k�4MF��y��z"eٜ2a��)z��نqSϙ���� �I)�W��^�`�.,��M�Mۅ���y8kAˡ�z`���6�,��)���H]q����kh�Bh�p�̠I�������]�9p�L6sв�w���_P���]�B�I$�ʻ���y馛3IQ&`�$�1o�j��@�DlyVV�c����<&�-���K�m��V�5�H@���{�j��=�&����[�"Q��u�Ԧ��r9�;g=���c`XƏ�o^���M�=@��lvF�|�A��Zt���?��C��{��dw����}�"��=?�]ea�5]�Y�������DF���m+B�Ӯ�{D��J��K>.a��}��]��N���̹��ZwfG�G���~���<ς���xE������ԡE_����4�Xaf���g��.����+���}�:R=�3u!-b�F��q����%=�Z�o��jS�
�i�b`�F�m
�tk1+zr"H�>�KK��z%���z>�����`�:��q �km s�ݪg��D�+Ilk����r�1,Rk�	I]$�~�OiEf׽6��. 
�[K��)VR��/'�vQ=��~��QGU�P0�oy][M)nB������
���.C:��SQ^�DvU������f����H>��0��q�7���dK�x�NM.���'�B@�e���5����,�V�K��P��Ӣ�٤�f<٘kzP�K�#�?�OѰ*��!E�\��D��L.�=�K*��C�j@#5����3�d*B3m	w���q܋)wBE� �I}�v ��9� ��8ژ�y��q��	z�0I`.����S4h��Ev5R,�e{�6��U�Q�	�d��O����DU~�hT�������5�L3�R ��t ���4
��w]7:�Y�����Gw���n՛�$��p�Rܜ':=�
(M�\D=.�}cp���$�:@���K7w��q�(�U���>�a%����ycr�g4� BB�c:��P�3t��@�����!�y�tn軎�5�������v�m�>�K�Gt�/���u�Q27�ҁ43<��9{���u��μ���9�2��pң��j)���ZR#�<� !�SA(������D���* �ʤ���1�9�	k� ���l�|�|�R/�[�~b��IM w���{m�Z�tا*Z�j�:m���G�+s�L�#n���eh>��wl�����=cI��z"c����)���u�����bmy��Ƙ+��UcM�A H���i9��%�;DE9��Vݪ��}�]4j�7\|2��ϓ�B��}�y�N FQs_���i����& {��o�S(F�l72���x�.��>e{��;
���{De�ɨ�8�F�i#K�٦����J�$��<{���	��yLgW&4�Aj4�ob$N��Xd��!�{���IPٸ���p}�=bJ�G�L�dS�.�&��wED$�o��,��-��\�{���SI��xW��s5��o�j���#�l��M'��߸��Gw`_��R�"�jC�}WN3�$�֩��2���!I���Ck���!&��� ��N�����g�D�E�_G�vi�-:M|$6�2�_tR��0���}�f�{�`@���|t�s|�so�V��[m��ߔ�#��`W�Z��9�t�3��͜��r�I6��h%���@լ�6�,���e�F<��f��:�4����g�\+��d[3|���ɜ]S�ֆ��EIC�/H? ����7����m��X�)=�d_^Cn�c���5�8��BkS+��01r/���m�f�����9�:"�z
��3@ǲ�����w���ŗ�ߐr~Dk6H(�Ꝕ��[>�Jjʱ��%�c�]ν���Ml�G�-:[/��]<̦��N-��=�Sc%�4�R?;��'�-ºE�B��n�L b�_Y�7��� 'd5�Z�o>5Ő�e��=�gm""�u.�ك��K3���fِL{�m��Z_A��CT%&"�)���M�5��#ϊ}%{��*�W���H'1 ��������F�z����9��u�'����|�_��4ã 발�n��`}�蛞m��{��U��m���A"�=�W\4���D<7�iy,.���r �H*�j-ǩn�sg�36Cp'��ۧ�\�Jj�L��iO�^����@�(�ɼ�RP喡�8c�T�%��1(��T��3u��HΚ�؊-h��-Qćv�7�.Z�^�y9H�(ꭱ��^_���h٭�w�Ws�F�[xE/Xq����5����M�[���)�v�"�ߛڌ�AQ���ʔW�<٩t[�3�Gy�إ�/��υ�6�
{Q�2��d$�v��HD��l�ؿ_�mL�������>�A�u^����Y�b���Y�������T��d'�9�I�c�����^�=Cˇ�4Q�T�x���װJ���=Ũ�^�Zd0�\�N$�͠��:�}��f�_�@��S����]q�K@o��ĳ��I8�<�\�s��a,���;���/�pO�k���d�܁��v���уQǛ��>҃ю�`ͮ�LR�vːG���ta3e=����	D�E�hj�,c�o��R1����oL���ƜLl!u�U1#x�Ş'�'�T�G2�5	�B���Ӫ�YX��Y�B��;:m�5� ���m�h��Oim�Ԏ�+�������_]�15�+,*�9��K0���È
�1%��|�W��	���^�~������])xvS}��<v^7��l��;�nk$�BԣL���>󉎔�����QQ�;�ჲ�Y�@�M"m�Y�ʅ���iS�E�Մ���xyU�S �^���c~���v�30gJPFZ��޾��	�XZ^:$�	��Ġd Q��c�T���S�>��4ϓ��We�N��(�ڱ%M_L�_�KuKD}|�����*r������++>�?`�1�N��vh�#}^�)g}������l=H�z@��~E�މN�1���&_��$�.��#�^�p/DWD��ߌ2NQ���Ҡ��rP
]��J�Kp�a��|˾�~�;����ǒt��z)kU��#���^	��2�"ܨe���_����(_�h�/P�8�O3�s,l���k����_��	!�%���5 �����3�ֽ�j���>k���@���<y�V�&`�E��{2D��
�m���f���Э��Z�"s�C0	�j	�{~JP�3�6�'`Rګ��mLЅ,WUQ�O�����Z`6��Ap&�*e��HnT2�A �!��C�2�j�"�X��_��8g�<5���w@<	)cJ���A�[!��M<O�4����0R�׈�ڳ�:���R๔_AO����+�%䔵%t���fҒ���P vg~�6I���Z��p���B�v:�9�h���m�
R�9�@����Si�g��=>��q�J�7�p8.�j�L�zp�},^T�ፇ��N��d'	"�p	�ߙ�+�M���č;���Ϫ��ٟ�W0�����c=�7�^Is������by�춃g���&voi@� ��f��C�u'�k�;\"�o��,�@:����F����tr�cR�˝i7E`�Bg���u�����]��1��y����"Z#�q��@"�ū��n�P���)&�w�x�۔y8�V�!|$���u��6S+�.�����pj��0z

s������ϗ���m��;s+���j����}o�����>��ȑ��DK�A�Y�SQ���j@�`�Y ��|&.:A|�@m���� )�]�i8C���yI��x)T�ve;�g�zX��^����X}̤�
��z�p�D|�x��U����վ��Qo�n�^Y3q�����hvI�Vb���B�X��i!�W��	[�v�b>�3,nS��;��5/Z*
���5��H9rӫ��4���.�.n�0��~^�Ű���wǬ���v��Ρ?<�����]���+b��rd'W��
 ����?d��	�z�]4Rp�Y6Q+�w���� ��:����𧦙c�M�֟J$�Q�{t�{��B��b�^�̞<�����t�o����fM{�bt(�i�;<4y���;�+�%�bX�-$�EӠhI�R�
�T_�Ԣ���d�q&���`2�,#[�����3���n��~$�5�
S� %��)�*�7Z)�K���v&�4H�����Rdz�!�N�:Pa��)�/�TUc��TL}x�����A�Ǧ��R�.�����P�&L�{�e~тbm�D�r�XӧÌ�j-����$���VZ���e����l��Cy��SJ�,����4�u�%p5��q�G���O�6H�`�fpس�[��P�k�KN��7G �ɥ�� ������e|7��a-�-/�ԩN�t���/��9=L��n\*���+$Z �	*���+��P��0:{̈́�Q@�j���Z�^��S��u j�]m��}�S �M��]�Z���f-4����w��mUr2�˔>W����&h�1O$cW;e RF�8�%NN��iY�Z����c��$Odd�z*���e�a�۸xO����]�{ �A�6��Yf�i8~�CĐ֙�~�^(d�h76���UDVe��Mǚ�}��x�u��b�w�I*O����J[�0[6���/2��x1���E���Ƞ�3�#�y(��N��'LTd+g�m�<mC7E�l�����Ru&���4��*݃gr���f�hޕ�B��X
����j��fs�� (�Ӗ���J��ƚ���!�5(1�?��DS4[�?%�v-�C����ul
�B��ngu�-����ad9��V�=�4X��2jԸj�w�w�ۆ/���t�5V��|���9��r�[�O:´��;>Z~��	���E���D#�NH�m��L��<��)9QG���f��00��\�]�3�/�h�n�u4�Y��ԅ�:����7؟ڿǼ������g ��c�[6�F�uT����hK��!�8)���6���a��0�kvlSC�`F#O�b�:{_j�� ��s�_Ji�}K���Y�^^���'e^A�x�M�q�F����ιc��&�Ɋ����'�iD������>��b�]����"��=[[����p��R��>�w����C9�9��>�����#�a�ܳ����ɀN����(�H��jaM_62Bn@�ܯ�Z2����.��6H����H�i��u�J��^(*f\@����������p����G�Z`�l,q7o��L(nG�L-�%B�4tX�jjP�j��{k��=�p�W��ܵD��Ũ )_��f�d0Z ,0{�y������au	}~��h���*A2a>�^�Q�.	ƽ5wR�8�	!�}���Jŏ��<�$�O��Yv�1��"��Iq�>��c��E��QR����v��
H�\��w�:F���	E�'�����/��w��vuΛ�w�u0�+���:��`J0��^��+ǲ��)c�@�`>��P�_���"-�p��Ed�-w8C!��\TJ�,��5맭���V���r,Wς&�H�vȂk��fa9W�ĕeF��f�=6�9��Z���@���I���ߞ��+����I#1�Y�j-��#��Y��ѵS�SB�>�2Qn|�S�����n�x}�H��=�����rx��7>6����<�Tvh%ʫn؜H�M�=���;����l7��f��O���������~Ģ{@�:/�΁����Ŧ�FW �0\h����;@�����ӭ���f^ŏ���.\���ލjOF��i�D����Z����à��ju���"�&�3� b��'��A��K�7�F�#@j�kҼ@�B�����;}B��l��_�%�}��v�T^�����B�e�d+��/�|t�b��ĆWe�B���o��OO��5��WU1 ��P��.9K��	շ%8������$�M�[�~�8�U�Wo���W�i�HOC�X��`�R���
��$�Mi� 9�n�?�>��B���K��:!��k�&�Je:ŭXf��A��u��(���nO{"�?��74��8��z$2�R�M��V,�؃(�A�SEߪv�u�8��0
6�����أy��(EW=�7�i5l:SyF� �.ێ�� ���Dxx��	4��!���K(V<��}~��ӓU�3˂~�)�e©���{]HJb��x��9 ��c��-&��5j�п�۪N%��p5�;g�y�ӱ�����s��*V�ڜM1dW,���F�*�-Mx�k���!4�92�'-�[�;WqŶ7�۔�e��5��y4��Z�����љ�wc��A
�z�I!���?����������h-�d�a+���K`>3S�Ʈ���]e_��/�m�N�ά,�!�;<<'Y� 5��C��7g:(�����MQ�b0ʋ��x(v�;Q�g�'�#u^���Ie���ΰ����m*��n��!�:C���2��B�8ڲ|0�&f^zU>�ֿ��~���Hl{�Ոy�M�4oEj�f�I�����\��5����>�P�O�s�`���fjh��.����YY5?/Un;N�Q;�\zgLy�j��\;�S�ӽ�-�R���^��zk����I)p P$^S���t|<vEv,�}�X�6~���n7$2�\����('	�Fѐ�A��9Mfʢ(~�!��6{��h�M ÁP5#����ㅦZ�4�����4���I�Z��՛$�ˣ���ɽf��ެ�e�9�>����V������1��YJk���B	����y�whv����OEl�^��H�	���br���#�����4�6���s=�E�?MQ5�@ 6��<B_�9���<}�m�Y�^�D",Bυc�pʔ��8��,��,CedX�lV��ȴ�GZjt	�j���fA�I�5QTTX����`z2�,?)y��@��v;��+CE����㑪��{��G��zǦ/\�����D���eH�W}�X�K?,�H�:����C�};f�{n�'�E���E��}�9�O5���o�]G�S@���e���̔yî�1�o��9G�s�N5�Dt�>ښP��xtȭ���l�sŴ���A0��!V��ޣ��������!;�>?V���Ǻ��Sb�72�T�e�uW�:���g,i�ˮ_� �,̒�v�+��$\��P��0�Ҝ�(#�]���'|<��YݐO��_7��P?rH �z�}���@=��'�&��i �9H��� Q��'2���>�A�+0��u�&l�f�M:��H��vX��6����L�6n�����݌QO[�
�����x�JgV�p��Q�&�����G��)J�Y"���"��-���o��w
8(�����x��{S�2�\��BF��)K�b?p��Nq���k��@s�~�*�&ˣ���Şg��?P�V�����)��6aq����,-wp-p�Z��:��(�`�%-韴%l�PN����p�c>
qͰBֆj6� ���;��H� �s�q���ᡤ7va�q�Z<4 �8��1@��#�=OY�#!��Dc�+}�w�k�n4�L](E�Ins��7�"B�%����]��Kpq"�v$^]���qt-���ֽ�A�R��Qq���ǎ�`��C�,8y�U�[����9�9��PWu���/�7��4oР0fR�5��������,{�ͨ���yJ��*$pFn���i��75VT����M�^(>�}�J�.Z.q]���Zݹ:��/�\8!�FUB�Ӵ�EM���;��"����1y訜�L5��U�V�I4��`7�A)�Gú���kfŇ�RcR𗝌�<xиa�,|��	����|��5�8;�}��R�`v||v�#�ɴԧ�4�����Eb|����OeU�є�Q�O���o��Kf�rл+�ߚ3�
ĝ�@�\<�����l�y�_�W��	@�hH*�/j����e������ذ����X�����]
�!攛T*����%���b�4���C{�2��-W��] g�C?q�ߺ":e�PR9�[$f��f@2P/�N����A�M3Z�bx_
��xX�<��@�k�O6�dg��������o�rC�#0�RX0���e��z�g�]Z���[q�?��WF.*mo��J[����Y���:D����4��#^�9:�C����5�x9���=$�(��e$Ɋ����d�щ��m�e	�,ל�|���`�13_��aX���丐ǮW:��ؽz����p���[ܯH�UK��V�٫@�0��X�j��Yg���l-�?qG�����9��a<�O���1ϧq<���YK��r7�Ѓ䮟�%�R[���E\�1{�x&�:�n��V��{���	o����i~7����kܙ�3d"E0VF4��z7zHQ���2u��Kdi����_Ec܈�����Y��E����<r]I��u�@��y�f��(����}��b$z�Z�߀spxʏD2)c�UgN����v�vQ�n�<E�A*�?6%���@�Sf�)�� aT�Te���H
�К�<xwC�M���6?�2���&��6��o�朌ڦgէ<Q?�U禖�2��ڠ6a?e.ԝ]!���D�L���wlD^�L25¦Ol�ڹ�:�rfH0E��9gGo��[T,��z���C�%�Le����|��+����$N�Hb|�c�*W���E�_���5'&�1R\Bg6���天<��kb2~��r:	}�E?uH�����iMm�gqHs����{Z>�O�e�TI��\�����/m	�
;�5��Z���Uz0M.�Q	M����%إi�2���Ao�lS�_m�^e��g#�{N W�i[��K!k�1���i�j'���U�-D�z�Tn�m�茗O�˩̋��{Qr����P�<���"lt�z\�:���ڷ�H�(�5���A���*�)h[P������H�p��J%1�d�E�x�gVٟ���#�+\H��y��9Bgl�Y�nciRs��h�Zh�-L�q��`���ɂ�	l���+�L���G�y�w`O�Ǚ�&�� ����10��C��2��7�,��R�^C�I�%�^�6N���5��axj��bݐOL�a���˧�|��(��#e��UV��q�Lk�1
���WQm����ԃ��j�]��~�_yj4��#.��qo��\)%���k�*9�qdء<` ͺPKnv���i������. ��taP�"�\Ϙ)�֩j�����dSo���uSMʬ��������=����(E��������V~��.����G��`m��+��Y�(��>�ܫ���.�V�y?��
�X��_�C��?t5vF��b\D���ꁡ����ն�ӻ6�Sl#y8g�J�d]䣠��k���A��ߡ����iĖl�IM6R�����O�i��g˂�� ,����ܞ%��d `ݛ�f�~�m�Ó+����X��Wa�M��r������i��?�5��A㱇�p{�K�>��w�0��4�Ih��i}��[�YXh7"6u������1��m-V�D摞gs��[J'�!~�C�%e������������'Bss�%�o���l�;s��*M�%��OE��!4�s�6@=a��e�/��0�dTF����/�ƻ[$���c��e=w�5��_P��d��c�Ȫo��k\*=��({����M`HZ�7�l��@Tk�Ⱦ�k6���#�ދBW���j�?�C�u�� 7m��_�1ް��t~gDO�y�G�����6���	�QI��L/Lb����@ q�z��Z?A��E���W�S�`���t^�9���Q�a`���,��z���E��.�~�EHIҺ����2Rc�we@���e��I�g�:�jo%SoY3Y��(%�$��OV����R��XZ�V��*$����tv1�t��Vl��5p�(I�7��*�u-�1���R�,�y�ɪ�9&��T��<.@�=p^�>	m$Ҝ([4���q�\t{C���R��(�X�'�gE�_��,&·�U9�,���L��g`ą"�X���un|��%� Xf�
�7��<b$�)�Il �^�/ұY��~:Y��:�f��!�7 �v��#���"����%���sD�fKH�ӿ�ʂ�e}=<ӳI�����f@P�!�s����z�;҃�x�z�� �-^C�� Y±�F(�U[ҋy��^��X��[I�<��4g�`m���T���	��W�)T��c�6����X���<�L�UxP��<\��|�Zw0Z�I�uϮ��N�y�5վ�O�R����� ~�_�Jb�fuk�0D�0�vǡ�v�¤��Sf����^�>0TG޳F���F�,c�뛔�����b}1S���$hR;���1S^r���lu݋%.j8��"�p���-M<I�m��	:������܄�b����rI�`�	)���>M��eŮk$arن��U�h�����_���Ϋ�A���k2՟�:BjZ�H��TOp��0Kˎ�C��<3lˀ��2_�����y;Tm��|��_'6aZ�QΠelx��k�(��^��2���b`�B|�*D�Z���ԒR����8����L˷��<�?Eu~�T��FvjD����N�U����E�y���Q�T���I� ������!��Qn�ș5)��+�8H��Woih^Ţ�&�7:Lǵ`C\�)3M�[���jj�( ¸��U������u�?�,������=����
�u�gaC^�H����G�=|]��޳�L-]�먜���J��I�:�������ymAT��q��4t�%2z8WTMZ?��Y�}�t`�ן���qc�Te�o��N��m*�0)]�D)�W����J�� �w<bҺ��<�'.�`���4��Vg��m9���F�1_�f�|�&5T��DbGTvb�@6u���w�����7w�=#��Ï�{&g~	߶�7�_vU.���H �va'�~ͪo�?e/����Q-<���S��tj`al��U����z����w��V�pN(ҽt69O�����N;%��\�*��?��V�vMh,x������P���1�F�W-a:v���WR~�a}xy�機&M�v%ܺh%��wi�ȅ�Y����xV���
�4l+����N"hf:�P�}e���U�Wl�E��7���q���M$NYV�,�C�q�a>E\	�	蜂m{�Zs�Jm�}��,K���n���&�~R�q���:ܑ̊�S���Z}�~�"#��"�7#����w &>�O��B���.M��m?f�v"G���cip�yS��(E�گ�Q*Wy?�DS�"Ɏw�2Ґe�fgᾠbȽ�(��xq����./���	��Z�6`��.-�-�wn�2&�{�b��Ū���^������z^0�sR�Ȼ�P��s�R��f���v/�����K��TA>��2o��1��2Q��������=���D	76J�z�N	w��n���sI�g�|y�r���eQ����X�9Q,���_H<�^"�}���nm���c �CV1������zp������g/=���#����P�\x3N���W��<��5V���;L�E0�k���͟���F\4gC��ڷ������.v�r����_���oc]1���M�񪞵�����-Nqk  ����$8�j�	��4�[��j���q��j��ְ/:���\v	�
�5_��U����%-y=��[�{���Ȗ\U����-���m���'܎��P;����O�T�s29�[�5B0���C�@�H��E�pҙ-��D��o�e�������P0X����`y�<$5��k�o}�,K��-D)�:�+�&1���5��b�ŹF 3)�1}.���S�BXi��p�we#�V��.Ψo羷��bh}�o�|[��(p�6z��w�m�)g��[Ůy3%s����|}�F��	_%J�# �L���x��9���Tm�_��r�k�0�������+����2s�)UP{ܔa����_-�QI	wKe'�����~֛�sc��H!�8ǐ�Ke�����|ߤ�Ϭ%�Ƕ 4��xGO�u4Z����_ǈ�%�@�ڵ�1�����F��|�ٜ�v�Z%��jw�Ah³��"�J�]dk� �.�WI�W�Kɒ��=��U//I�I�K���1�2���s�x�2U��e'3f��_h�y<bz.����Ef=�&�.y�R�{WaL�sLi�{\Ab�'U�y�bZ�S?*k��J��IJ����z'�E܄D���x�x���F@�"�����^q|�c�R��i� �z�'V�>�<_����fa̾�����>�Bv]�~E��iҰY�D[ߋ�0g�)5�s�ݷ�<c�%{J�6�7��8����ݾ:��3������c���{����ﺊM⣞�0"�!y��&^���~3�r2�/�)�m��Mi
�S�x
�n?-�J?��y��n�9�艝�(�p�8:n�����s��_C��`�u������Q��g$�b[��'�I�\����~�K���E��|�Ѵ�DLI��U}�Z����(���D/fG�3���n�K�5���t3O
cպi` ���X��Ыջ(�[��ڍ�\����h�Q����Q)�>DLX27��p��>�a�;*`��a#��_m,ëKCD�mJ_M�����FtS����V\R�0���1&�/�F;t#є؀��&`�m[�������@CZ�������:=qYN�*���9���&�*���v��X{c{?�V9�Sʛ^�����p����)�jЛZ!����Fl̞��Bt���4�}wԉ��U��_�v��d[z�`K�].�z9���o��ڒ5���$a�
�Y�!=J{�����yA��yC��T�x]P�N�h6zk(k����d�v%7���?�3:en��`%#�Lb5~�����b��܅�>p��R� Gidm��3�"�.~A�i��D9�%м���ڔ�)�ϸ�āSρB1x_4j��g�y}s���*�^Ԏ�4D�l�=$R΅]U�D�m&ϓ5is�	j��-G~�����N�
=��6"a,<ri@	��uf&�*�/�f.��Kg%��*��dDT�8��#G����Cࡶ�=z�،^��K }�8�h���_b4�^��I~0���#z�L6�Y��(Ji0V���G5@�`l�#з��J֔a;��������8\%��W��0'���5���ܪ��E�Ł n��qF��O�jɓ�iZ���b�E�ޚ8��yD%h.9GӌU��a�o�*�s�
wBl�0:����@g'⻙�Ļ<!�E#N�]��yg�HYg'.��#P�"1����/�X����1�25���q?����tX_uu��5�`�
�A�.�*������<XpU��
�i�򓘱��gI<iC+���c����Z#Z�P�TL����z�\h�c���:;�YY%��v��f��U
h�;��SF�1�M��e'"�����+�2g�o+��A����/�
�OIA:�Gα�?>7��2�u
��vAgc��9���_�n�O�Z�K~1�,����'��&1���9߽�O
�4�!���Eë������[3G�(O�*(	��g0��Ue�qHte������}�
�"���w�e�֛��r�%�ט/��j=�v�kݪ��K�f_@��>��QP�Gj�4����<��q]�� �s�c*Oq�`P�
��zK�	�G�E���y0�;Y�]���ٕ�.S�6z�]t}�o:/���V�)���cY�a/�n�*���"{kB7�g����k�:�9��|����#���=H���uIV8�4w���d�R�,��g���9�a��K��s$���:<L�;<fX�f�+�#�UK�K��v��8�ݭ�\s�'TJ����t�̱��*�(�u�LK����i϶x����j ^s{���ʤ��o�=�D丯}�k`��������+35�wj/��J[��ݰ�!�;(+԰����V��ңF���<˘��3R�I�]��v_��xPun���Pͥg�{���\�+�\I��W����]D�p���I	M�cݦ�ڂQ<6�?m��U����*6�r]0�fn���j�9B]�L'l���/�}8��1H��p��K�f�-�hz��[۪�d����u��觬�b�0�:<��	ʎ)4�,^������-�ő{rly ��m�L�TʍY+`Rͧ_�M�ti!��Qz�� &�}�̆�7�8�Ь�+��C0N���o:�� ���);��T��������\G��vih��d+��_[���0#NIj��4�h�����Aa�H5'$mk��62Y��r���iIG,��,;�$����J$\l�o1����ɩ.�'�],De�)�r�|�-�Ȁϻ���zH݉��n�__�M��d�~䣃�T��,H;;�(�3����������q�yBZ�7�8��g�YQ��~�m��_�I�\��$��	v.\}"�D}��I\�5k(��ѹ�1sQ:�_*������U��}a=���|QJ����{t��:�0��t���{�CX=\Ž��	Ε��0��h�X#����:��Ѹ�]� m�&ǼQ֠pW��֌���E�d4d�&������E*]�P �[F��!�+��ʸ�K�
�f�b{i�ԈϏհ����Ķ~W� ���,��!032�z���Qn�(�:pw�B����Q#K���&�'k����,='zAU㉅�h7 yn�裧�;����G���2Yf�lE׿*�� �\殉��<���.��*���k,�*n��S�"?�/F���^N�澫5#:��=Ŗ���Vټ!�Q��:�v+Lf4�7��]gQ��@as�5�0u�H9\4�i��(���EJ`�c<Š2�ı�=�>U����5�����ޚ���ҵ�FUxn��ڋ��2��/�w��Eh:e��b���[TK���:���&�ܦ��_�y�T>��7�
,Lᖹ���Ŷ��ˍq�N@(N����q��(1���R��+c9ʋƠ;"u��]c^��p\��X ��ń[���#E)�~BN�ԝ/R��c���gxvp���e���䟢�����㴎�P:�X����h���o:�&tHH6�K�h;��9�-��:W4����/LFv)�����ܛ���26��,/�C��g���Ӛ�9�x�9��s�3k揾[������h[��r��š� laV�˗'�!w�;����&O]R��<����Sp�^�W���dw Nxˁ�����h��,�`�LAi8��0�8���uU�����u��4�Pd��!�_glW�cڴ���ԶK �{lQÖ��p�s��m�Se0��ׁI��0I�/O�X��4~(���%2ƥ�p�x�E��T�6���_-�eq�]�0��]���e�.��krt��v���,#��sݶ�y��{�Q��b�Fg-ە�W�b:��Op�(���h�_Md��غ7����#�O�̙�P!V����SH�����5����ל�:X�X2$�Ĥ��:��qfČ��<�T��LvO��=W�\�;�O{[q��`A�������٤z�>t���a�����?J��}�2{T�g�}������3��)1h�.c.��ݯ�7$��#H��Kjq��7��
��5խm��G�@U7����Os�3���/�(}1xPkޭvBP�TMXf�F!�s����_���n��\��T��m�����%T�0`-A��%����n�,�89�5�>�%壆�X?F�=f��f.�IN�D�A�W�l��b���׊�͉z�O��՘��/�+���RZr���p�Ͻ1ޔ�Ɖ�@]��P�M�OܛB���		�J/��B�Kb�{�	��I�����Z�^����{i��;nUTI�F�4D�/}��(q�_��D5C��s@�[�d�]S�|(߰(�=�X��'�G;��^jԘ�RD�ⁱv�y]C����m28�}B�`ϊ�j���������!��?i��_������7-6�<:M��Q�_��]Z�ϼ�~��)Qb��J��4�����
�xp�i�~�z0����������z�l�KY=a�؎_��EMSwc�,�g�{��N�&
��v�.�Qӷ,D�6z�5��غnZ�R�	���k:��[�f���Rc�.&�4�>�G�uEg��#��,�����y������r�G�
��`�׎Zb��^\q�<X�vi�f����a�M�����:+.�gĳ���/�v�(��*Z���H�T ��|j�_0��Xd�έ���t� �?.��yCe�^[��V`��r���>3r�{�ɶ�3�߻}؂�=�0m�/vR��2Y��?xa�P�:-ZH�$�����n;-���&�����E~?���i��Բ,=E�.�&����\1ɋF7֬H((��%����ݳn�]��-�'R?6������w��39O�-��N8:�$J��,�( �Q^���Bק�K�'h��&o�a̉��}�������%l4�R�|�s�7��;����:�v��{�g����o����>��eB�,$D���p��.Y��c7�n�~�)���*�3��$���g�����v�B�^�;���Yw�AU=Q}7���j������|�׳>����N���g�vl��q��l�'���ܧ�k�^�}!mԺ�F�������ۄ7��{
�3w�jwXq�~l��Q��P#ǯ[���u��x KSԱ��3^xw����\��J��?!FŪy�MIm��&���DY���&�F]�=@>�oX���-�� ��fd���Ox`���#�X*W���˷�T,��O Zc�����<"�EvcR�y�K��8�YG���A�{��:��\�44Fu��G�,�٧!�b�N��L��z�gn/������9�r��
��,f�_���Z��&z%8(v�h*h��7�QE%�JJLU��&"�ӯ1�����#1e0��Kp����RDv���h�r��+h=��,36�R���9�W7
�
�Fo+�q���`��H�"�?!I�p�N�o`��7�]ߒ/�U��:�e9y<��o<
i����*����$�c��m�[���nE�4��$Yv��T�>x�k���ҡo���	w��o�S������I���({��}(����2
�*������V���Ou4#� ޮ���wps������_&��!��0��SQ�3z�`��?���}�V�E�-��) u!���Rl����ٿK:�+�+�e��MF��p��N�Jws��'H:|��G�_�v��|�6Y5��KB��F�O�p��&S�`!�)K�B��H߄�Z&>� �8p!��5�B|�cA��F���;y��k�7D>R&y��Zܮ���k_��о"X9Y����GH.�..D�b٣��g����D��t�<�����������QR�z{$Ѷ��g�
t�Xv���O��d	�L_����43�^��9Sg?s9�݃��[�?|�!��H��L>�9>��J�����u2�#q$^�~=0]L��]��Eu@��UL��5$��h ��o�"�t֊��I#�QM������M"�a��Æ��>S�~��������n:Q���u��ғ�H��5>AH�v�R�.����gY|�$����j �e�0��T�o8c�4�;�c0n�V8K��_Ɵce�.��q��j�q�U2������]��6���U>$}t}�
�d$��P�S��m���.�R�\_��c�,m#�e.�Y�<����\/Z��0eэ�����s"^KP��������>ɠU�w��0 ������!�9�̰��Ǉ�R�n�ZVa�9EIЂ��)�����B�+���F���$�mr�a(�w�3��<�PR ��[����h�G��̞P�w��P�?YL��.��h������a!��۾FLE���	�����h6�DM!���Ūͻ��6;+rґ~<[:PqTĦlu�?3c8�Jpy��rl$o�cG
�MLɳ%��7�JEfS4���(���n�@�Q�x޷��g���8�C>e�����;�I�`L�O�0�^�+!������p]p:��(�Me{��vԤP�{R?��`�+��8�$��*��`�/~�};�S�D���ceUi��[Q-�����18d�@�P��E�bM�{���@��n=�XG���_.$��UbxO����\�oE��3�=���}r$��V��"��r�"P(�]�X^��9�_Tr��B�{�ju�K�rV��<�Ѱ�o�(^@
^�Q�FUKq��xf��ck�,О�!w�ˤ
񱁟��yڛ B�mHm�S��hꕣ��M����*�>29`P@��;�!��d��]�L�C8x3��+�l�����oc��ў.�}�X���<�,@�67&M� ��ڂw�k7o� z'�3$�b�k��U�.+c%
'�x�O��a��Y�!W�$�Xa �����EY���[��|N����ÕE\wo� bt�'� ���>���&���ֶ �pC|Ͳ=A�[EvwH��7�-$S����y�|b�Ӱ]�YI�D����e_C�y���f��>[�J��_=����3_���y]��Y�_�� k1L���Z4b�߬=*r����B�+de�.�y���s��}c��@`��w���R���)7&���6y�%��z��8��f��(�lR���Ïm]%�ߜ����S`���T���8��rg4�{l�}�	/{��خ��Jy�fz֎8Һ���ʓ�n��l'R�S:J�̕�^���8;�ٰc�<S[��������:$ķZ�1i�z)�|)��钻�|��Vc�k0���%�y�����~� �w$�V��xWF,\�Hb5�eD*�r�+N���m<�-e�/9���\B29l��E�P���煞g��m��3/�Y�m���ά@�H���!�.�4���Q;^LfDf��l^�p^6�B��k��@q��1_sy���2�~{�:K�"y�q��hb���g��Θ���T Vh�@Y��^� I�#ešqTN�c�PPR�lʰ���}@��nJV%ش��@��x��{Q�5z�ΞnB@8�bY��;\&��M>-?;
�{q�fg}���+q�@�d�E��E��H�5�Y�Q w�Q�5�$��y�,x�-�pL/Δ�n"}�C�o�_�Z�V/��4<���~X�i���X[dHH��AN�Y~hVs��Q4�k(-�,�	vdн�ӄB��f͛�-�WWL�����6
)xʼ�Hω0�Lw����b����9���}Y����`"�Db6+�2����i���/��.��n>�7����c����Ӹ��غ~��خG��H������q%+Z���Ɔ����4�vy(��$������Pm`���N�z��/�rz;nC�0m�;��pS��?���Nx�S-��J��KR8���o��F��W��6���k:�RH���[&x`I �0�ժB	�<������N�/��!�-�S�J���D��B:_���?5�(Q��p�C<`C�S���X������E돍A���o}�ٝa�?N�h^'��0K�h=� �Q�Em�g�S�ˆ�I��A��r����gwɣ��Vi�Z&����wrU|<]פ��25	���I��&�I��[�<�c2�M׺�Ή%���c�ԌY����cpG�Z{zу:�9���f�)1-!L��E�ߏ��	?���l��3
~,�Ҁo������Uh@��[��0Ѳ�M���3���z@&��B�kc b>~g��F�A�I��F�3fϸ<�+����Ԣ�ƶ$b�[̏�R聾ȺSj�h,Â�z�:lO�N;�Qm�A�l�S�\	h?������>�C�,�*;9#���.��qn����;v��3�]ͽ�|��1+�D�@Ғ��M����Z�����M\G?��N�By�Ϡ1�x�x�1-��0g9�fXG�`�^�Z,���t�#h����Ϧ�s
�%9�E��t�������~�e�;s�h���[
�A��s�*���^��GX��{�Q�s���*vh��x>��D��-@��1�� y��g�JlK�Ug�i�H�H1JH���Y��cq��[��m�'"��ܨ�4�p��b�+�5��l�IH*��mQU���l��P��'?�m0�0_�HE��\�x�{�.�Ӏ��xJ�O�����d	��k��t)�YaCU�����$x��^�eotO���]���1�pM[��1Ht-s�i؀Q�����c� 1x�}T3>�+�Ҥ<mS$�Z�Rb~P���[C�b҇n1�q�<}�Қ����s}ݯ>5���i0�%�1�D����a���|s�օ�ρ�c;ZB��E��P�LY����d�P���~!��-��7�#�&&�NKCp4Ѯ�Xj6�-i`,�8ݧ��/��}`���M^�ј�^����T���.��i�ٍ̢O��k!��3{���:��Z�
=_͵as��(�W�W��Me2����D��
�7�~���Q��Ap_��!U�|���ǯ�����WI
�� �#�ʿ5��R?|�޻A�}_��y�����:&��w�}� �A8��p��a("tڊI��a��ߐS��7V���1A�~M�f��\Ձ�"`��3MM�nҌ�!J1W��%����Y��r}N�%̴�QRv�A�9]-�1Ħ��R�c�)]�)Q�Ě6�\̄B��79:"�z��T��
�pQ��NL�b���W��ya�T�i��%���:
>! ���GL�G@<��
��J��|�軚��P�����x�Rw�N�[
L����^���P�d���i�YhP�:�ZSf4tXE��D�>�27j��莵a o�R�ؔ|������kCQ�9��g՜LZEb�(�da=�{m����a�I��U9����1������!֝��c�M��[���hK� %�JD7���)_)�U���(�dV�X�{�#� �\L���K��͏�<�� ����1������i�D�+�ĉ�5AE�M;x����ѫ���@�D�G��k�dAVyB&E��'vR%��^��9�[�-!6-�Z��~ۊ?Nt�Ȏ���$ؔd���8w���]�v��
w�-�:�X���Ѕfap�;~Hj�H65B �f��nP�l�WT�Z%+�m���B�w����bH5�ݭ5��7���u/��p dz����9ΌYpA&<S/�&ݣ1\f9#-����w�c�@��2����|�#;�̮��-q8�2����/@�X��2s;Ը�<}J,�����	=e�^t�̩`\<k��C���*�U��=26��j��h }���y3ږ��sb���e�~b~A�}YTk�'|��xdɅ�%-��+s�c<�hC�%URl���55���ᘮ�x|��1�9�ij�e	�>ް�L���+HK�y�qՃ%��[+��>�����HU�yq=�w��/���9�]��l�=Vy� ���
U2S�L\��g�3C�a��U�Ι�<����g�xhis�Hd۩ ML�D�l[TA�1���G��Dd�p:j��#���/#9	M鑯.>���{�P^sM�RP�M����rJ^����G]h����­E�U��q#��s�u�:AR���ƪ�Wqְ�V�Q��i[�j1�;�^$4��LK��E�����.���z@W7�mL4Vm�+]Ռu(ۨɴ�0�����P����_r��*2�Bx�ڂ�]Qݰ+�j��6\��ތ|���C*�F��4N����\��A1�����T[dK�k��I�6�3�e��Sgߟ��/nERL��w�S�h�#�x�4��N.vV��JQ|k�����W�X���$����d���ubS��:��OjI��5e�{�1��7�tO�[��
���V�l?�_O���W=�v�Ed_.}��A����!�8�JWB��N>���D�-)=�8��63*�1�2��]1QG4v���{#��B���\�t��b}�Ɉ��ֲ�f#�T��o�n�ҍ�.Ƭ���
.������牴�yuz����E>�%���۶�γ���95�>�ex��?q�z�c�^(���$"�4�l;���w"� =���DNuy�-�̆��X� �u��PY]z�c?�c��:ě���|.tC@WG�%S��:�dc6 E#Idn�}�)�.`Mu�s]�P�@��Jd����c�QB:r�ugxl�=�m��8�?f�&�t��v�>}��o������=r�B����$ٱ�;K�Ej1�+;�H�����\vg�e"�^�Y���I��+R C{M�J΋y���ȴ�߱��1�|*�eͰ����bO�}�N��>.z;;u�RP��M��>������6r�yGI%T���2͊6����s�.¢V��w�j�A/��oX���y�G츝'_F����A�f/GJ��B(�,�1��3�5�L��cI���@�c~�PW{�Z�5��x���יh�T�ԬW�-������pa���J�lP ���lx'�/8$|�$���N`M_BQ2��u*��j�E7���s �u#)]��?vǼ�i��qE�ɡb�%�N|��kT�)Q!9���P�J���@r�W�d���M�zw�o�J��O���c���"�:0)I�	A8X �se�*m<���)
��xҤg�V2�J!����VU Q	{��<��
�$��ɤ�\T�(��c�Oz�P@4r��79>v�4Z�|�r���K��O�!���B҂�/��f�w���^yW�^�.�n��*N���<�g?]D��&�;`�j�Ųs#�κᓡSEIN��Zr���!R��0��Z��,׍�m}��}���=�vs��"�|�G=0��F�/S������;?��@�ߑ6&�����߆�օPS�H��oP�����w�ͳjf��S�r�l�&=�ʿ�`���Hy���`#���D�k�~ ֐7Ȅ���=11�g��w���I���a�����W�T���}:\7[åߌA�~����/X�~&%�@k3�nH��s<��gI���^G
%�H�Ƶt;���.�H��&�$�خ�m��4n"�^Y>�sr�.4�s��8J�u�$�n��CR�8:ݩ97B9�w�$8\
ᒂ�>>L4w�b�+��ĭ��@Ypj���_yA�@���&��/���@H]�dV����F������<�d�%4�έ�!|r��" F9I���-28��q#ȆPC�u��R�_q��н�s��%N����L�߿���F��T���d�R�'j/�k�!�u���^'lC�\�%0=Ch�2&�=�[�Р�w����Ka�*A�k�5%?�u��2Aq���H�
e�e���o�`ݨ����P�������X���<J^�g�!�js��!�jg���I��C(Y�J�R���+
��{^A|���kG�:�;�O�EÂbD��L፡�="��Q$8���VL��%�B /�A�ޥǿ?�W�IfCHA�̜�/U�%��R9L��w_��C��g�̝�D.�24/�ٰ�RH�J��sOagY+��Io���cs�Q	g�
�
띕�����}�Ul��BUe,�����7{]O�N�S�0vq$'�����F|m����t ��K�rgA;E(�T;���nǸ�7�&��C�{f0�Η�������Mv��?����;+���[��0�4�C�4��ӥ������nJ��A�yC����$@��s��8q0���9��ԛ4�uB @��~C	F��|��/qZ�駭ldY��2�2��u���7>��������z�#�c}VT�(@=rE�K:ԧ��͜�f'h-�\_dT�,M꽜�ߒl��},�gz�T��I��`���3zX:/ݹ��%�\�>nsDF���X(�i�r�πW��_ձS�yC�	4�?VAB������k��z���:mߕ��i8���=w�%ؖ ���3fD�p\�l�a(X���d���VZ��q+O)����[��)&1>�h�f�\Õ1�+�Kd���7����5AF��V������� �����ֱ3r����F/����ox�
��U�'E�?i0vݡ|x�����|�~�:_�z����;���_"+�2�n���Ҫ-�<ğ����wI�z�:�H����Y*���I]x�יVZ���S�-
P�&��D� Jo�<1Uו\/�wDjA/p��8���8�o[� ��F� \�}m���W?�W|ؒ��/�*�F�+��[$�����q��?�B�6ing��~SLQD���}$��p�d�-� E3�7�P�K��wF4B�Vނ��Cȇ9<�K��$mI��Xwb�C�u�/����~}����Z����H��U��?<��=V8�P\<q�FҏC�=_,G�X��ʏzJ��]ʧ��R0�.���n0%�F�ж͗^ɀ����J�*2�
Z~��Y�?i4s�8��t�������"��]�K�ro?�w�SR���6���.��n�^]����CjU]e��O�/�b��F�cxrS��<G���$�W٭���D`�J(23�R�m�_k>�2FzZ@�`*�Y��)@�X��X���4 �ue�Gͳ��+��2������d]J�D��?DK����\+��Z����h{���b=�x!�>�&ä�:��n8-P�Ik��#����
3���р35<�m$�sCf8�xJ9������::9�be�s!ﰇ�k�x��͒��bIȿ��dx�^ךti�����U"u�dU�(�`�K�����j4�Ue�M1�8����M�
�2�8_�T��N�ӳ�^La4D�P8w��iQ{�`��I���ED{���mH�>nMdx8`]bu9�.��+H�q�X�]f<v+D �1����ƕ1�;?O�O�ހ���� �=��Ԛ ��;i�`/��*-K��<�	��*�[������Z�Tc����1���7u�����-�u��{$�L��ڀ��cH50�w2����ܾ�Y)-i~�m�;���7r�0!�`�$ޔ�ԏ�^E��P�ez~C',��hM�ʺ�>� �=�S�Ȕ�gc�1,�u��n�f�hLb����4鄩�	�p'f�t��̋����8Z[C.F��vKh���YF��:J �����NAaOw�
�Ig����7�N�x��X&��-+;�Q�ȁ�� �E���25���@����EU�r��׳��B�,f!��+���yɄ���[|2௫�=�Xg�c0���M̄�����s�˥i���/��z}��[3\*�䀸��k}�;댉�ը�W��~���S�hA�&����m[Z-aJ��,�� s,YR��@���ӟ\#h�/|'�J�}�W��U���n! ��C�����G���4F=-��T�;��#�Fz��+{����i�grĳ_=	�K��ch� ����ˉ�I���v\odI�,��P( �U�������`�W�{��k�{Ec��):U����za�kMɇ4�6ZH@�����0����E0e�P��V�D��Q�	tD�h�Ӣ-Nm���ʖ�R@�tJ: �[��iK��e�e �,�{%���  �z�:d�����h���c
#�����ۑg��� ������F9]\��Qu�P��R*��z;8���%l�I�� ���ހ6��VJ����Ϸ��nB��45$������Dp���b��*�tm	��*e�hKP�~���1�:�����4xi1��?��(N�s���8�R�nK�&f�����C�1���4��bY�Jތձ�oȀ��r�+E�s\�8IPnk�,��n>�O�)�?�(*A_L��7k���HJL��.-W7���}��s�3��'���0��� ��}_�ꚹ;C$�� ���h���/õ�����M�$$�h2C�f��.K��O㎇C����|+�T�p����L��N�kMWk�����W�}{"�1~Z���+�Ts�&��L���;��q���s�f ��Ms_H�)���Ӛ����<�)N޼&���t��ӄ&;V���K#������c�Rw�,)�ۈ^��˛1 ���Ȣ��#�S�'a>__�'�$��Q+*��z�\�d�S�l�8@�Uҁ�os{۩��lm&�B�bal�HV�����ķ�t�y������������tI>럮5�����!�y����C�2gޒ�Α�OS���]�K�P�=�QQ3�q���������J�KԮ%�����<�}��W*�����WVY]�|G���H_��/.KB�e�ݗ�ザ��ˋ"t&���qQH�t·f�H�RF�
��a2yu�B��;���f+�G'��Cj���r�ўs'#��֬�I��ؗl��,�a��O�^�%?���1/��L��+6�B����I�K�F��$��%{��X ��Ԝ�C\�L�?�����V�=il��T7�ど��8Q%�?ؤ��V!Jq�/d�*��1��H���~�v��f�zcm<%y2�I���!H {&�[g�7�s��0'�R���uS�[]J�U�kf�
�VR:Ǌ��J�2Y�M	.nX0��c����9��Մ�-4*�V���}v��p������N�#,0VA�a�`��v$�#�H���/��v0�
�G���9G��%2�h�!�mA(��u)~�o�3\��H���Q�z��r�،N�xo�{p��Iv�����O��?W����N�.�Ww�f��b�����a�*|�����>���ÿ��ڜ�F0�a�WxZ=�
\��:��R����ɳ�{l���Sd�J���C����f�_��I8N!<g���3K,�3NV�̌�֘I;˒�A�2Z�ܨ�1a�9��Y�A�G]�Nl�F���trHU��f�n��m
yh�;]Զ��
�X ����s���7�(C��4��"�=��캩qCÜ5Ti��
U��\�����W�Y~��������n�a`:�Н@ǰ�[I����/^
q�M�^���P���Ml�(��ZP9]b=�d��԰GR�|%7��jI�qZ��H��٧��bh��	{b�K�F�9��S4�P*0��S6V*Z�q��,��2d5�8�3UYC`������2�]�gk{LC�t�\��	<mC>p"yd]O�',T@�o*ǯ���=�O��������?��Nj�-<!�B�=Ž�?Zh�+n�Ak��4W��:�3$��$�ՠ�ᖠQ�B5�:(�0ӧ���i*:�ٺ/_� Ĺ����o]r�=�M�g'YH��ͩP|��)����8��*93[ͼQ��#�2�MwK���X%p�v�h�^�4�D�;�+��ܩr���S�ّ�Tc��dߪ=�b���	��`H�h޻�N�%p��J�\$�E�����Pz&1DtJ�c���2V�n�[B�Ā,���-����^��g&�%[�;c� �x�F-��L}�{�')�?{l1���I���)�
Tm��@x��/�S=�UAkJ�� ���*����ǻ#v���S�x.��W�lEo-0
%b=�5%uOl��8���/���������?�'�'��U�.�L��Cޖ�`o�.ۛ��{RG��K֤��S���3	<�J .��[P>T��}�����$�$��[$�x�Mu:�m\'�����BiD�2Aq��"�+��p)*gj�z��eM��~�t�K��(����V�"�]�/�pI���\�q�P��؃;�3�-Ь�-#�&
*�_�5��[��ӎ���)����e��Y���ͷ�-~��za}����2ވ��v���Dk��2����U~�*���p��'�,���΍�	��.�����?6����6��QT]2����Xwl��É�v~�88g��5.�Sf<c}Z�s��?T�a���*>�.�he30ʠ�A��S+o	#��Z^�V`��p�� �/JF��6��BT6U�r�b����u^�'�?#���e���3/�M3���=�}��?��_�1�:�]�ߣ�I^&�k��h	;��7�9�=�C�De$9��ؿ�M!&��s�]B�m�gT��w�a�aGr�������>�����TkYTrϽ�z{8%ms���w��z�B����^�B��
�-WG��+#��d���Vj���r��,��r�)�V��ٖ�YC��h�������LU�@[���[���o���.���DN�����k���p��.��lw=ǟ��u�-�z����\dFeǙ��L���;�S���Ⱄ�_H ���1���Rw<���P��b��6�>�[�5�0>�"O�H��v&[>����!�]k���M\ZM|�ę1������	��}<�4�h]��Mawִ����o^V����[ŻD钑ۈ�cQ��٨�pH@�ͣ��LS���s�^�����ŝH�W�1R?����&Xj*��dR� `����GN8���e��ˇ8pv�_5?��8�&q�s�Q�{� ,���C���Ng�^ ��0�IOK� �R�|���,�!�}+RI��lЈ�_w�����ܲ`z)(�4�BaF彣��n�M'��ޟ��'S\�;$�4��*�j2p�u��4s�6���{��2�9]�!*Q�)�B��vpfZ���t�z���;T��߼���P�D
�g�⭠��1^� }3@�)V,�������k������нI�E�
�kJ&��s��v��K^��5�O��j�]8���{���L��8���	��Z�������Qv�x�i7%)u���N)4B-[SB�9L@��n0f�ok_��v�OZ9�&��yqo8�iO:�)� ���߉�k(�efx����*�3�ʰ�M7����d��F?58j���qc[�oW%�ł�d8�XŇ�v�4���T�w-F�v�DS��F��� �|�@.��OҀ�RD�r����\ݔx�P�^�"�+���˗'+Pab��b�'y5����"���w�^��pQ�,���eх��L��J�Tw3��f|܃�P�'!��v�L�U��$������`]��m�Wͽ�K;����+]@|���W���Ѽ����[V@��W⹋ [�W���\/��!���sy�����X�T�:)�c�! ]�XQR�
��Uv��1��h�(kY
K�Y"����߽��i}���v�f`(DGV��	�}S���4��>!��.�l�֘}�$gi��-$<!�c�����K3���&�F�'9l����)]A����z���l����!zj�:x�FCwݎ"�Mg�e3%�����W������j>�3p��t*,3��S�����V����%���M��-}�����,�Ɉ�6o[]���쥾��ɸMi�_��������N��O��Pf�qJ��+�}=��m���vF�ڭ��>k�l��OaMf#�ұ��|+ ���\�d��H',����0�C-ޯe�Vw!-8G�a;c�+�K6+u/ү��ʥMDH^��Q@S;�����	1�}:B�b�a	dO��kd�g�1�6���J#l��B�U�P�Fuܹ/QI%#����[LS[���yNq�� Z�)ԁ���7�5|�Q����/�[���գ��^~�����Yx�^B	vXا#�M��B��Z�,<�?R�Sq�9���c�Dk7����||�ߡF'\��j�)7������$���_�y��z�������h� 	�ށeٙ�KW΀��.�����oYe��������x�h�6e~-�G��1��(�<��#���|�q��q::F58A=OL�X.���Nx8��2
0hFw��s�<�ډe��.���C�P���2٬Щ'������2�w*f���YȖD/��U��s.��WmK�i)Ѹ�`Wj��G�"�ૌ +TE}Q�����Ɵ����i�R�<♇�SEYJi0O��?�kt^�d�	�D"=��N/R�у�ųA�#�l�m��ENT��LV�+��ԄE�y`cG^�m�,7=�_E��p���1����!u1��y��f���%�G�>b^<T���l"Wq��3���X���|�IԶ �J��qa3�º��g�%�,D@NVjE�L��LYr��;hO����;����д�CT�CR[ⱅ>#�����x����N2CO]�ឦ*3�^��9�b�Ά��$�J�&"�pM�5�]�?�pZ;��� ����&.���aj�j�|��c�螽��S� ���;��@+���i ����5�R��0C����6c�d�"���+\�V(E #�v�I#aw/��>�ý�P�������7p�Jw�,�t�wr�