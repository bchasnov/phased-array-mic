��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1���e}ʲ��cg�t�ϙ�a�:�KR�%���ݧw���ȼ��W��d#�w��<����A����Z!eҤC�5s�"x�{S� ��x�v�U�b2U�fr_�`,�p7�.ۋn�8ZQc�ڳ���;���`���i���GW�;��Ԅ�wo�/C�v4]�?�S7�4VX^{��'n�u��ͽ
o�+c��T�������"��ɴ�Vx��n���1��1F��f��Z���%��`j��ʨ�2ټ���!n��f	�e����Q�|ypZ��n822e��,�&� �1B��#%���-#�0��o=w[}(�g�U��y{�}�:V�`����sivy�p�S*Ρ��.�j/���b�y���<U��"~o�wp�^���Hhn2Ss�/�����V׎��Pl��8�&���fB������%<�כ C���r-���|x��c��#3�2f�8r���|�ݰ�m�#4X��?��qٴ����ěS�m �6�p��
���k؏�M%�5ES��� �}��F�v�Z�ق��J>+�<=b4�� Ҥ�l��8�M���Y|��4���r6��"gw�'y����"�� ���-n�#���;�$�A���w�/��z�qp�߮�S�mସm>���gz?�L�Y/�����Q� �Z���	L�
��Ug��tC�y�q:�_`��=kz0�)Aۥ��l�7��P:�Y��D����q�z�,:D^��+�H���r}-~2ZJ����<�N�V�`C3�2m�FRʜ@����]m�#�R��y���Xf���@o� ���%l�y��MzhFx�����t��J ad/'p�D�x�����.ˇ�z�\bO�
����!m��k��=7 ���zߨf5��g��4Ē���*\\&p��^sZ�Br�U��8�rD|�e(ZQm�t��W�,����UTOځ{�+�fa�����?�&��BF+�������m���Kq����%Ǆ��ދg�]�:y/k�ؗ"b��_r2�N;zO���\`��0c���~JI� ~����\�i��
�y���03y&+Q�a	q�c"2L����*��D�_��\��Po���v[o��CDP�^����]�:.Ͽ�&�x���`��(�qǬ���_;�$F��?��q��|��&�`좢��7���B:c�b�of��}��
�Cu�0��մ��|��J�Č���-. [�;;���7�Y��
T�*��]F�-4�:5��{���d끌.�# �%� ���ѢZ�A@~jW�<�@���X���N����1]�S�[�f�~�)��Q��7�Hv�E��U�>��M�g�נ�I*�{v���r���F=՞�i�I��� Y���^�����J7���̲bc�mb�\w2E���y��=~�]�c��W1�~2����n���yo*���?� O�G�Վ�JŌI=�Y���O�<�0��'d���cł�~U��2Y3e�9�Qd$[,
:�8�>�b�os�u!�Z���/���G٣�*r_�m�x��|BiM܅s&���?���]���v���^9���`�9���ڵm6����˹G�Ɓ���y�	���C��Hw
fF�ݾ�C�|��T7�.T1�9,ц�q���^!�c���a{��MajqڈXH�Q�}�	��E\�,7��+����sS���H�D������gkam�s6�� I�|L�w��L#���)�i�H�{:�=�1���P{�-]^-�$D��V����	���j>���q�k���֩����;O/j̑h��<�}�$�M�C���0���)
:Em%�pG�+d�x^p�_P�5@��˾S�r��Q�V�Ƶ�"�4��c�<rxV�R1/�E�Ro���MO�H���~��=�J`����U��� )�v��~z�M�y��j���F��dÔ�e8`���֠i���n�T�??�|U;����]A�w�C��������z] oUFm��S���w��BM*�w.��ȹC�(sy��մ���Y1w�k���e.ᴱ!�"Rư��#���\�g9�}4��EbV�1��1u*3Ŋ�6�{���ke�z��c�T�ʹ��Y�a��5K��)�!ة��Lk)��Z���oн�c��\���PQ�p��^/�Q�T�i�Gl��W},�1�,l�7�=��[�=U�¸�44H#��'o柱 �x�>q�/:�� �.���m4q��@�k� r������t��)pe��5�˔Cg�*��D���S�*r�C@-��4o�=�Te. �� |*hM`����g�e�*��̈́���mUH�s4�{��i��R�\0	�}"L�T.�A�N�u�q^�i���俴ga9��s]��)	Y��!��� ��J���o����ڋ&��Q��l��}�x�|�f	�C���"�,!��	�ӕ��E�R��-�K��kp�Ѣ�&��h��a��+�:􈴑.{��p3!�1�U��~���O�FD��q�еf\��'g�O�o�����B�QF���')�S��(w��n��Ś�8�>�?<Ɵ��I�U�%{��`T�f��|p���Ằ�ع�~C{�u������]�ϖ(9�4I�:�?���^.`��W��<�(��d&;ء5˄�����6a���NJLd�	Iί�*�;88�r�,z�r> u�v��!䦷��4A�Mw�ϰ F����^�|��~��?R��a�P9�����W2#�v�Q�����6���%���~��/�[�-����.��s%�2��r�i<]L����oDB�����:���j���Q'sZ��K̀FX�F����GKm昮LW���b_���,�&���Ҫ�J��s6�Ņ�	�#���hnK|�L����[P�m�� �|y67����8/�d�e�t|��.�v�FgJC�Gb�h6��O�;��L4ٴ�_����C~�P-��cț~�^�}X �XGĩn)��H�G��C�)���2��j��͘�u�?n=Y�I�<�e��-5[�L�����J�J���������ʛ��0?c!a+BO��C�{���f#	\ch��Q��]L�@L8^� ��#΀@Y�lP՘s�a���Kz�ª��{L##k�N+A
����;�y�~ć���j�,��@O~�b��z���*��|ёmM#�����n�S���pȨ_�R�Cy��"�+�
�7�K�[���7��1��O��ƨ?�Հ*�ڷ_	�����z b@���_`����-;�{�1�;�A��
�0�l�>�!cB��E`C;�!�?X��2xay�:�����`� K�Rv���St�6u�(`��Ue`�'�Q��A[��itՖ��7�
�[�k�ep}�JNs�14&g�1�Z�Q�~��:1Ɓ���T�B��I�����TǙd��9��ov�W̡�F<}t(߷.�S�(ٗ���L�A�p	��/�9�ޮ�d,QW�$�'}���kPL�H���Bd.H�-|/���y��H�yqN}A4u�G����M䑳GY�Ϧi�Ć
f p�O�&�t� �7B<�Ս
1S��3�G� jT�VC��g�M~&�*C�a"$D�Mڦoo��]��������u{��6�O���B���rV7�|60�aN>�$!�]P#��t?ENß�S_���U¶�iK�5�P��$�j�!��U����_���0Fy	���-P�Oɞ���e�ґI|k�b]�B%ɭ��٤&���ya�C#�ē[��QPƌ��fd�E��-v��&}X���^!��tS�
Y����U����,��F��m%*���ЙIm���V$�f������H�#�{��
(�wcN��w&���I�,o�H�b��L��C$�
v�Ԁz���sS���3&���h��!�n�
uV鄀��3�jfߨ��*ks9�T�[&�w��f+�����>e> &�ي��o~Pⶵ�Ue�\{�d1(�����K�OSrDWV�(�Ⱦ	Q�d��^<���a��	8R�	��z���)�~VLox<�
:��e
\��,A�Uw�ot�W�c�A#�)��Z6��x���ӑ��t�{�}6h���(�\b}�U��5P�_��]x��f���ؓ��_���az҇��֨45"�Ŏވ��֑�tzv�l֧��LTw����4L���K��o�	�����\6�N/UC���&�g�Y��:��#�p�!�m1�_c4��i��K��@U51^Dۍ�d~����K�5|Z��&�&n�$�LED�zz�i�$�Ǳ'�ӡ���ݨe�+8�Y���F���f�kI;��H�&�H���`.�nK��&��c"�څ���3��<��k��T�k\�W�1!�&8���g�r�B�%�ڿ i`�Q+5p$�-���v|B���"b�F�l�z��=��$�`��o�ɖ���"UչE� �˧�8<"է�(�)����e�`��S=�!$(/���~R�{���F�n��Ө�R�����	F��9�Q�(��oq��mP8�d����D�i��s�w���$��k�C�;@K���=ް�B�v��`@��ꭧ<�=���#}��-'�n�`8K+u�o$U�ރ�05��TFF�Žz���TM�N�����2�̫D�\�Tt����8�k:J-�#�d���b,Z���v�_� �ߒ޵��^u�� n
6Ĉ>�����k�D98��Q��f�Rm���Bw�`���.D���i�1�j��#|�k���u�D�588�0��8|�E�h�7��0Q�S����<X�ʤ���Ѓd�6���*�9t�MȈ�H���;�#��~�Ag��� h{!u�u�c;}�xv�T����@��[����M��Ԅ��k�a&[9�N�����i��}a�:�-�_e�*wp����1���ٵ��"��31�_��"%4>�P$�q6�EjY�@�Jބz�R��K.4�{L�M�J��#z�n��r���2%:��Sn���}
��(Q�ڲ<pnP��e��c��|�����ɘ���(�D]�A�"v�7O�v�k��L�l�҅7+
�c����8D���rv�Cr�e�_�;$2�f%|x6RP���h���t"�VA1�{Xx\=��k����1�K�uB�)<^��?0���t�Ue?@mu(�|�v ��1F�⮨��[��K�XG�b-¶E�oa�i��	01oȱm�Ι^^d��}��x4|����aH�Z V�,^�������/VO�(�Y5��$�3�ws�y��i|'����N_K����4O�:�_��w�)r���|�Wt1f|
ֳ�$n�����]�ҧc�"9��QggA~��q��X���;M/�/�}��,[^�%S(�����3wi�o���j�n���_��C0�ؙ���~��x�rGQ)��-gEk_�)����Q���!cu�2df@a���K���Ǆ}�'I���V�ㆲ�mf�v�"����V�|i���v۶�r�>j�ojaN�r8�N�Ih�]u�$�xf�j<bZ�ewz �iJ��,7u�Us�Tq]�[�m�,�5�����N�����!WOL�|}3(�֣tZ�׃7��2{I��|˵�"Z:���R����!�a.@E�����gy������C`��!y��������������_�"C��U,9D%��p�ڍݬ��h] �^�Qv�i�����^�8�M��]�e�x�������E6��;� �pt���D�	U�C��&���6s�	��v�n?���7|ڽN�ȆF�p��K%o��P��F9��vSg���f��$�S�%���|v���sx$Z�D:��z�4|�^(�W��%�.��}����` ��������e���lJQZ��f1�׸$�����".�a�EQ#<��U��������de`j=�Zs�K/�㋑SSK�頖���S�-A�\1��d�8ML�C)�$ۣ���~��� 8�����,�O�AgeߵWۻ#l�sp�M���]
� =~�&�8y���b���|{��	�Pq�3�(�^[d�����@��$��*AHR\X"eس���u^"��ۗj���jV]Y�e���n���p��?�~�F�K=��B��[Q�B��AZ�jm&$6�m�ɧ3�0K%�:Ӹ��. X�Pϗ��$���X39�C�A��<S�P�eQ��h/�j�^��/TcY:�����Ǎ+%ѡ: $�u�-Đ��{���f����e���S+e���u2������VW���c�j�ݒp@�Є#4�ڜ�>��x��[�xѾ��=�2��A�},���m"K`�#�)7q��N�2�+�-��]A�<q}d���7�{���I�@{���3����{�9t�4�9Uyb8fr�t�j��b�̢��-�ɽ|o�i7KS(Y�&���=5��.��:�@��LD��d��]:����َH��:*e/O��� ��Ë&-[� ��	֘x�S(�9����U����|��j��)��y��V^�Rn�oJ��'�M��nN4���Ǆ��I>�Cj��B���L�-�5�9oc��e�]/������&�	�a�𦖈>@���u�as_Npݥ%�t�$�.�n�"M:g�6����;�"܄	����K��4%���/�llrieM�"ߧ��	<��YYb��P�i�k�w̆��������t/�	-���6�9p��G𞧝���G8=��Z;R������a�M;i�\,�?$�xW�a�hS�*�V�U�s_�������������W����N]����#���t!�]�=.�B�\.޳�5��������܀���9�h�N��1��.��>�5����a�U�2{���:S�reC�Y���� ��4W$-�VY6��ߠ�Z@��U�A�7��lD�ӑ뒘i�+�J퀤�B�]��|iԗ����2���IAkVg��Ŋ	s��!��6��V7^mJ'��H�ͩw �,�?Bseu������U�"ɈǨ�4��`�^gƙ.�J�3��a�_a��l%|���G�^�6��h"���s΄�I��D6�^'�{��%��E����Z�@�Wt�2���Jl\fLh��]�֛w+o=&-���!�º7wJ!Q��6����0�Y$�ˏF��t�=ڄ�t�l�:��eϐ��Gz�s���w������*�Y�t�no��n�H�) k�uo�\�Њ�(䰌�o&La��
�E�Ԇ��%�1��Z����d�����IH�xG����\��n�<��cᱤ]�rQg�|K&nv_��,1��k���W�ژ�y��c7�Aj[����IE�Maw�~n0Ā��м����y��Z�Q~͒�*u��aZr\�/1d=yU�Q���!�Zإ�\a��������a�g��]gl�h�Є^��U�q��~�ҍ���zD�	��o4����p�#��%V�B�͓��z�0Eb�2��9�rlC}:��K%\�F�q��*�]6��f��Oj� =��Y��Y'�/vT����vQ�-#�4irU77�����l�*�}�e��7A@�z�X�GE(Wj�?V��"B�#n�Z�`:cP��7�Wӌ�=��u1D�"D��P����iF&�.7���A�:v��@2�x���	';���@����֔�H:K��teW�.@(Dh��#�:ˁ�7N1�FHP�%q�b��4�/�����k%���OO��3��t��$A�)4#��*�x�Y�[����g��G�܁���>wV���(����.�ohO�t��]�S��_Ȫ�c���!�9y�J�]��^����X�z��rq�/���Y���B��	3i�o�Ѷ��� f�\}K���O�������X�
�{�!{M��Ɖ��~ŵ��K�k/��:�5�!N{�~;b�0���:r�K�"���$�B
�K���
v��^��գ�W�3������� ����آ�\��y�}*�Q1*�I[<`h'3!#�E0S� <1�X���3��j|[�4e:��������B��,��Wܗ�� q��x�)�k7����#n��vP��B�g���u#1:�����?�2��[�:�:/3ƴ{)�x�
�'��
�/��
��p�֒�Y���D<F�p(<ni��P���%Bl�:�9F�/RA�%�I
=�1>�_\���Ņ�����A"�[Ƃ`>`�)�U*Q����b������$�'/���QVvƐ۹��I �H���'
�!H�l����[X]��с�;�Ī"��w��O~qKͺ��CD�p-�5S��7x1���,����Y�{S�ֵA��f7V�Չ�3/�m�S��c�De�Y�BWi�+��Dvm�V��^mM�Oz�k���}]|�3�0�r,���0��w��=���fKǩ���J[�}"}����dd���j'٩M@�@S��P9��X'Y��}]ov�ToO�wyya���E2�u�\�<��rE&Gy#'�TA�l����?x,m���+܁檌�h�ru� �aV����7��y�A�Q�!+Uy�p�����`���[�/h�"J��ب�Wز���"�g�*��bo9}�����TӇ�w(ֽ�����Fh��[ ���Q�䝇7��?��ݸ��\�gG������� �<���L��L����i�xo��M2M��.$e�}�6�^ܴj1H�z
�Y��φ(=ޝq��D+��ZY�����1���=o2&��3X�,� '�\a��գpu#�2ec�/�J���et�5
Q@}i`����[p�W��W8x�0?�5I�h߀��a�Pز�#`P�K�X��#\gB\C�;��d5��|��z�P��!��1(��ٿ�{�*��	�}��O��hc���dc&^Y�j��zG���q{SN��=�Y���b����C������oD�tXz��<}��z�&w�yx��>\Ox��	��_��e�Y�T+�,��R���x���������͙e��u��5�w���G�i�s�����V�}k��ŝI������9�8|���㱪�p&dΰ�Qى��-���"�lR �k),j�EcLF`��!���>iy �bH�� "�+��f�����h&,��Y�.�n�Fb9Y�>�](�{��4������O��O@�H�d�����n�		�H �5�m�M�ֿL������8��?��/R�r�٫����m@#���S�X��I�Ĥ�����қ���٠U��0��փ|Ν��cZ�r뀳�Z��zg�����y/Z���$�`K��<�����x�Hb�l> 
S0|��<P���zU����%ρ4�n"T0��h�1���[*}�o����l9|�7��}���mJ�q��3��n\c���X��H�Tw�")=�8��j�"	+�m�.@�k������W������^��=�d{2�swC���e7;4��zw 2J�����H���@�J�f��$�Ш��G��N�|��I�e$�����'�CQ��ї
O��1�_���}�C�G�Lx��"��%����i=���D�|8��%��@+�-��� l�4���6ߖE���SG�A�Q/��?�<�����!�VĘ<���7f���6݆���Tb��]�7&Kؼ����令�f�����-x��.(rMMܯy\���uQ�B<��%	@��G�I$m��n E�����W������J�)�B����2(
B\zjzpT�*~X,T��r�U��xdq�#�d��E#�2{7�X�F�,?\�Q�U�s-��q���45N���h=�����m��$Ҙ�H����B��.�"ܮm��2��O��xVs�,T�[tdA�N�7!���`���-0�򇖿}�C�U��S��H�SH��_��?c���c�����Hn©��2�=��Ɵ����ghS'9#_�x����c��47��[���(���i�*�e����"?�sժ�8/ÃD�CY(sBfy�T)�D�����L��P�������:�r2�1pZK�~�qv��G"Lɰc�Ӎ'��̌W��{TJ5@�N��{3Ś��^%^u�\���m�OP$Qu��r~�j=�.ﻦ�K�B.�F�����+C�YB��������@���"=��rE�ɬO�]���kY��	��l����W�\=�h ����'v<h n��@�l-�F6ul5d�\ ���t��Us�	c��c����fU�jH.�$2�V+��p��L_�{A���c�4�׭y(����a����޿������z�1l;��չ�e�������D¢��Ԙ|���XB[�<Po�\!=�����a�]���2���� GP$;����iXԔ]@��=u�o�\�Q���>T���Y)Db�����ܽ�. X]6��s<vj�jYt}��.Hofr������\��F��)UȽn!7:2�5�_��sۮ�t@k�х��Z��qr+`@��̃���<"���5A{�'�*m ������k[);���uL!�Nd�P��H���"ߵEuA����O�S�'E9�#C≂�9S&�@1$�iq�?uk�374�A-��:
�k���ҸWDS�����/�|Z���w��(���M��3FE=������!Ĕbfd�>�YL��C����>A(�^O
3��3�**�֙�^}�9F]��:o=��6���c#Yj �Ҹh)k}��&*��Cp庼�� yu:������{g+|��?���W4�}�T�-̦�QrNNo���W�����U�=K�w���R+��t�
>������S���1�g�8t��QQ���Hb'LY��-��)zx/ћJ�b�cRV.8�����񅵱��y����|j�v�1Fu�P�>:ݣ�Xf�����]:��	)�Ge)�MG�<�y�t�j!ŵ}X�g&|I]Su������3c���Z���!���\]��y��'Ўj��B���u2_Ŕ^��پ0|��I�h���01#�5��/�\����4�!��I@~�N�e�c�q�3�~�pX]���S�{��'��^:��"�ԖFl;:��T�ג�қ~|�\^>}�(�4qI+�����[ɞƵ�=�[V t#��V����j�݃\�񪟮KMl͵��\��q�����n��z��%�I�FMA��D��/�s��Ց+�g�5�����>u{gPT�ȹq�*M��5��$��SIN+^-�+��m��-���oi��Q�B��e�]�G�IQ��ݏ�����d�?��M���8��uj�����h�!x��t�!�xYx�x�z��C_̤2Oߖ��e~i�W-S�塌�?��Dߝ���B�? ���,-hw�֓m�<��ƧI������7@ɦs�#�����у�����m�ˉ;^8��xO��w���P|%��������ݎ���ȯ�!�{�V�3Lm�܏�%�"N~���mZ;V/e7�RO��}ӥ*#i����E�V`�	S�h��U�G}�E^3x;�Ή䋆�"kik�L�Ϥ��K:hۄ%�d�%���J�cX�Q��1L.[`�:�V���Ӆ�jk��>�gR�8O�D�S_�Di��=[�R(Z[<�Ht�����ƈwf,E���٬ch�2��kQ��DJ�w�5��U��Nq7G�s�ɜ�6�t!�3�|�������M����My�/��Y��Cv^:%��$u�~��9E@��y�`����t(Y�G��ykʏć�����|s�AZ��z��yct�J�� �*�S� ��k�4�H���M�F��w��%��a��U��Da	���h�χ+$��r)��u��/�}\�[�����Y"+��WAL��?:H�Q7,f�{����C!��.[��bA��V0 ��i����J�G��$�ݴ�TDo%U�!�J`	7lH��%��6!��p�f�22hX�~��Ϙ��b��w�Q�/dY�*t\�m�n���6H��:U�Q�Ӻgb.���:�u���땂 �?yEɣ�SAv�yh@íC�e~��e����L�қn�N{�]�h*��Nһ��m��E����X���a_��E>���-vR���P����]#g�q��.���
ƭ�ğ���|I)��d�Q����'�©9F3��V8�W濏t�&ۅ��4ɷ_�]ս��eK��Z�*�\%U��A���Y{��\#c��l;�E����;>�2Ϧ���*��:��4�S����I^4��RSr~��+:^���Ba��wR%k��JJjA�{���#p���D�w�&�:O:��[��ĺ��^�
̕Xm�B޹�]*|��⌢��;�3>��w��vݦ�Cu7��կ=~��)�ؘ#v�,�7����B~��o1l� T_�0<�p�b�vn.�p��bV%Z@��>������Ƌf�W�,]/�1�3^�d���	�\�|�4��O�E�חd~�߼eAg�Z$5�g^�nx�� b��|���D:��-5�|��^��w�T���lhYjY�#;��b���3���/���O�/[ë��u(\ &o�*S�GZ[�%����v:��b��R�e���C6���s�����2W����zۿJ4.J��T�,Z$c�0����̣�yEC�gg�w����?*XQ
y7��$p�ڌ��rFA9�rH����>%�\�r�>� @�����dʭ�1�GvF�ܶ�9��*9�y�C�\Ǩ��]����}��u�śJ����!�";B��bO�M�#JV��/���7սd.�ÒLTu��_�i���.��� F[��l�'ʏ�`���[����-�����|}�D]s�Lz>t�