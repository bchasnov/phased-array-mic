��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|��V�^�Z�RRQ�����ܕ~5����iվQf�q��wG�5㺊-&y�(ӕ�'�oA�!4bå=y�v"-�G��p��/��+�rs�P=�މd.�`��~R�)	B�n>�|�8:3#��v�&��O	qs&*�I���h�+��n\�?�,w��!�_./��$c`���j��4ᤠ����	S�+x�7۰X+Q��\��\���5�7�2+�4C�.Vl�.�4`�A��ݒ�rY��ݖ#�z\�2�:�dV��~]�DE↘85(��� ��@]���̮�8'��!�Y���c�S��$n�����Qx���x�܋��#2�u[AU}��Y��&�!X\a�50�ix�h&x�~�3�[iO��7�(�S�;�������T�{rc��5�� �9`m:����KA�i�����2=��)pX���D�ld�B���g�9������̢<8E�l�$�|���æ�O���H�b� �
��j�tOe�!W�h�o���~_+`upd�ԷZg�M����5�w���PS��������,�~��ܽ��>c����mƮ�f1}�^W"ԓo���#С�@�E�tn����@1:Ì���)wn��g.[�~^K�+�xz;���`6y�zI�l�8g���+4�D��ցȒ�l�Qc����z8�'�7}��
n^N�u�s���-��n�-�n�>�^�𪘳Jra�kyT�,�fef�2�v�}lT�S���˃u���xT���Bϛ<����Zƫ���b�C$�IXsT0z�5z`�ӯ�����!���c��T��J��]���mQ&ߊ;ɅݵRܷ������X:6{��N�}��fKDu~ĭ�"7�S��R<�7���rΐ�C��U%8Wوb�u���,أ��;�^A�B�<��=�NLWm�Z^��}����ж�3�\\����$a\~�z���S�6�㴣��E^{49 �I�phH��u0U�qB�&�G�k:�Q0$o&�5�ʸ��ۉ�O�gp��3#S�2yG����Ќ4TO{3w��ڬ?���N��ꂒT�AȌ3E�Ri�0�����m�[�}�E���<��'qy�*q�̷M-`zR�O���/nAR��n�ʱc���֮���͛�J���K�FQ}�u��6���Ǭ!��a�����K���R��^���⹟x����TUt��Qk���CV5�^���՗0C�6�6?��Orܴ��#C�9.�ݾh��w�
��%�����F�f�*"3�q�J2(���~�k�TeR�R��e�{I���[�($5Q�ͻQ�fɕ���l���:��0��n���P����ۡ�k[!l�-�^���Ά���r�	��5%D����;oo��$%�4��^��`�m�����[�з��[&�L���e�{�Eg�E/�S��a�J!!�?Ze!��,�������v���4�&�@I���=�h�� X2,�Ψ�l�vE�Ӏ9�y�'�!I��KpC#�Ŝ�[�Z��" ���'�yU՜*���@T��R���{
L�=���i($^���|n���ޯ ����� ���y�1��ݗ�#�e�u3-�all��B�f~}<f���I=,�����:η�\΄��j��UX���&5Զ�xV0[��z�},�唫݋� J�X��1��䪜F�Q΃>:��E�ow����eI;#2���Y�/\��Ҹ oԇ�S˿��>tҭߏp-�탸3�E<��>Z��z�۩���\��B�V8�OǕls�5�8q�yBC<dW{Q"B�z��%k�^Ph��9C��WՇSOد/��^ʝ�P{WlM���f��7�U̪0��I�wP�"��<�ZB�
����92N�c#��;�jp~{w ��3�#Ir�J�<�m]F�_s����d�[1���.+0U�g����8#J�E� ��/�l6��tDlق5�_j��$���^g�M��:h�Rh=�g+}��fA�e4�֐�h&���&��2?_�Y���A�n=j�M�&'v�@}\j����E�ýU��#�|���<p����*�����*��4�R���lA<�Ll5Ez�b͋��B.wp��~2(E���1�T�Vn��0����D�ޢ�'T�J(��	V]*5�[sF[����
�3=Er1�|`Ȃ\��i�����f`�G�fc%�����>�k���Z���o����*uy˓I�ȓw��n�D
��`���'!�8�q���u� ���X��&��5�����c �3�q��Bה\L�_C�UW�K�M�����(8 H>���/��0X���GFO&6ڂ*�!$#�QrĠ�N��V�?��vY��-�(�@�u�+��`U�bF.Pr����&h�ӏ���%�w�&UD�0��I��[y���S������I焽r�=��5���D%"���zw�8Eo̓Qz:/N�-���gx�6*�/�3g�u��~J�I0�-��T��uV�k���s�4Hb�_'<�`!TV������E���_�#D���k�s���T��.����@k�k;z���<����K|����אt0_{�$����ܛ5��+�>x9��������)�i��W����1w��_��	��"�BC��j0J��������;�@�l�ۡ�ݘ�|4��誑-�ß�X�vY����[���9���z�R�Я�BQ��d�(lV��p�
hN�*\A�O�{���{��m��[�y]K,��+��jte���T�����|�o�FtB�D@nԄR�\#��3"z�i�%>-�Z.��u�#��P�����n�[���]�k�A���MCu��v�c��:,n&y�Ջ��q9.�������!B,��Iv�2i��0�����ߪ�'���PE�Ex���/�_\m(I�"+󗢬���4�ҭ�^>�,K�i�wI�/�
 �R���l0k+A���	�?2+XT��y4�����U�`�t�5�V99Z�*�2�g�0�<�� E����iG��ܳM9 kbm����~N-�o!c�r�QGNx�a��	��1��Dh�Z��#�FI_7�p��	�~}T^��	8��R����F��r9��i��?O�+~�;_�[�܉HM�`Lb8�[�e�Kr�え+�m$9*�6�i)IІ����f�5�EՒ^�$��e/���l�E� yRыy�E�c�3(F
�SE4��z�Ԛ}4�ˠf���\?5-�h�N<L���v��DaHJ.wɿ��`�`����I�Q�E�!��~0��LE�5/,�H�"r�;����_��K���KS������-��.ixL���`S¶��D����u�錐�~��o`Ϯ�.2b! �xzJ܇�M�*1:�]m�LVt���S�Y
�n2%��٫���@�\��;9�W��8�:��h�m<4}��8���-���^{1a[p5a	x3�,��&��b�h�k	\M����O6X` ~Yr�j��A����Be/Pzr� ��S/���:��d[r>�n�_RK�-�!�ydV����f�o ��e���%���k<�2{r�*��E�.����ӂ�W 	}ԗ��LB��/���hֿ�ӊ�F:i�WWO�r����%�W��'�g����bZ���r��_�m`q/����Q�'���A�/Ҁ�y��3���YbA���;��0�0{̥;��Q{9)�0��@��Dqb旮�;�ۻU��*�k�a0��(���{`�ؽ�Pt�#���b��G4ر]�"��g�FHc'�G!+�M�f$&�K�u�vDw}17q	*`�j�OMW���Yxw���~ޢC�_+�p�ŕ>�����$���M��k��ib�|8_�C&���0k��K���.G԰��0�p���و�N�,��+h@D>�ͼ=Gv��i�@���e��8�q�3+.ַ��}�LBQ9�B0��| � ���3�]L�li�x���q�63|c�Eq�cg#��M���ܫa�9Ab��8mk3�Cr�/���߈���J�fÇj�b����ءuG�^5$��w{e����i��ҹ��'W���ul��w<���A�X�i�7I��1�G�"�8d������3V��bΆD=R���̝�9'���Jf�g�ő�7��R��9���K�#t0b�=(+��?f�Z�����)lbp�aZ�/�-��);*��2v�M��|8CK������`����>w�wOɵi2���F�
�ϭ�8l��7�~�c�s2�� �����r�����
��6�3ȶg��VY0+m ��w�MJP�>��Nŝ�n�o�?-��Tf����1CH7UԉL)�u��YP�`�
ܬ��\r����"s���9d��jDiZ6��[��V�!Y�Ā���:�,7XCP�]#�R�?�d�%
�L�r���v��Q�7>͖��&�M,����~�m�I{J>̜'��`8�#�M�I5`�;~51Ҫ�")Oe�uz
����4��a�\�S��Q;�yo��R_t�ǁ@�-�)@�U:㟆^�i�V>DX�u@�l�rmY6ɼAW��'�٘j��o,T�j�J�)7�?HXh�9��^�F݆���Cs�]鱘".������X��a8cR>��	���F��Nj��F嫙�OY�Z��2n_�q���Pt���$L�D7������q����fpAu�������CД]���3@��-#��`^y}���-�4ػ����'ĭ&���qk���W�U�XM>�V�B���tٝ��Y��j�����Cv�H_�
���n�"Da���A��Q0qh��}�[�j�s���$�3nN�6F�^��| ~N���%��8���t��[3�e��}��ź���*���|��)��*��&�K�!�B����7�(N_v�A��=(E0��w��%���-V�[���H%���H6�� �"Yv��{���8�m:б��9s��P��7KA�ԡ?�svQ��Z���f�Z�@DhW'U��WF}U*�3��d^/�_��Z�L˒�Eݝ���� Ԅ�����ueS��l!q��>��fWq��ź[�u�/����Sx�r� �o|mأ#�'Y�����p���ԘI0�54*+Ń�����PJ�1v:��1ԉ!�S�퐉=?�(Ň�*�d����;�?�/�Uű!Y�A/��G\���ǉ����\�)_g:�:wI������g�#����pqhZc��9�������+�bmR���k�������`��i{���lJZ��SV����l�I3!�w?3��y���1}� �=m34�w9	=Mb�~�tȚ Ύՠ^0G�[S!>@�L�1��k�=%vh8��/��7�����ֿ�Z�ſG�QG���6v_zϻ2���	�iR��Aw�8����Ԙq��e�!������_�r�x���}�}�1h��OĪ����_&
b��0�TYn�����M��.%\m��6�l��L�4�k�����	��w�xy�X0į�������$<�Q7�φIe����3=�1Im�]Y
�Y�_��]���H������l핹�o��!����L����>���J��R?��t���5���}�;�>���BElR�DO>�>���C��z;Ԕ�	M���
z��_�~H�*�[��2(랲ל�]���&�`,����u�r���J`�v��	���>�Ͽ	=��$H��G�X�J��� (���n*<K�9��KǺ�����MGb�/�M�
� ��`��60r~�8/T�	��x��C�5$�W������F" ���H-\]��r�XVH��w��EQ{jg	{��������x�7Sl�N5�p�0t��eejڥ�PG� �L��(�<��f�b��j�7�Ow`jۉSD6b����"��0A��A��(��V�*����X%栫�@و!�J���:��c*�}Y�q�÷��9ޭWX$4w��0h�}G��2���wN^((1�`2���LЎL��q��wsg������b�ͣy�������Q�2K{l��>�<��z!�F��J�;�=b�.�d5]��`#��B�RP ǈ��>�~�G����C��д�2/:{�yI�I��VE_��|W�~���$s�.k4�B{�pYA�z��'�Ҁ�@��X�֤��?�Nޗ�'��l��p�}oI�_p*�?W����!��=P�~�]�4�����1����3�t��װ�����A_�n�X�ċb&�>�n7ˏ[J��jA遨c,ݖ��>��G�d;
��>��	ꌎ�4V.���$`4�ႵL��"s�"�i��N���C��t�T���P�,i �Bb��g���������2��[�M�.��N�
0��+��Ľ ������]�Y�e�A��w��̼��$��)�����?(���i߱R�zG����� �
���?�]���<.V�#�SƠ��6���kи!o3(��W��x�뭡���n?��kMl�u�x�I���p�~�n�+〄�	����'��f����)f�{af���U����8p��0��ն�O����c }�њ��*�� ��?�y�D�=�����&�Ӡ����é�A�F9���+"����=�89���>���~��#��v��4��)���e݈xB��'��YpD*c��-�:˂���:.\O'a����'.-\��P�;�Bw�����T���C&Pv<�	�M�	�S�\�˚g��2'��{��xٔ�z�y�l�ˇş��� �3�g�#`��q�|�&�ə$�=eqG�ki�0}|h:!���#l�\骟�[�t$M�tpqd�<)y��?Gu7� d0O*ǪM�i.#�������ҵס�Hm�Y��#_�:	����	Y�d�]�i������ՕnQ}N�(��)&5�\��������m w���Ȥ���/R��4u5B�FY@W�X놠n�i�h�n�|��!)ш��M�:c� ��H�2f�
�<!)�dxq��� R�G���8�G0H�\x�}G5�f����Y�Z
2��}�$S�t�(�J�,Uܴ�z܊����}����9�l�M�=�qn\���=�``:�!P�ݾ�A�	VNBF�E*�YZZ5��؇���I��^>8#��i���!.��1��@LyN+%�I7�b���,8*eg��'(0���j�=,��U�6G&.&��ф�������3��� �g1���#٘a�jr�9����7y�t�	��1��Ij�kW�r�y���mÜqS��
��G��:����$���/�Y����hl5�[�ܧ�޹�p���`T�x��1��zH�~�M�O�~mr'5ڴ���6�/fz��ۿ�7	� �Y��I�V�~�7�G�	���+J�[����L��S�Q9�w|�Y}`τ���Y�RY�[�:q���&�]|�i^j�9�)g�Zh�Kҫ���(��G���:�-h����cn�|���C��j�C�Z��ſ�T�;�$0��9_N�ESDܓ�O�ȯA�/����~�˾	 �������S���vwaׅx����7o�z|@�=Hδr+Ր��p�qu��� =L�mV�8\]�M��L�S����VK�i�@ɞ8����q�d!�0hN�U�6�1S0���j4�҂�u����f/@#��	`�M0�`�5�rNݚ,
֒�(sJ���Wj