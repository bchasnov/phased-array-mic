��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\����q�?��e�I8�b�Ǽ$��"����ׯ1�V0���9��";/sE��ƛj�4y7
y���e���}���y��!��q>ы��x�F��\����S�۷�`��{{\�vt�6k� �זň6�WӉ8��o�Ϣ}�ᗑ�),�w����H���S��g�F/"1��+��ܶ��"�Wǚ����"�$j7�8Q��*��M��>	PW�l:}	�B-?ޜ����_���
���z���)�eq���ݧ�ja��e��ǞaV-5��ꙔU���$�=k�m��{V]�$�RL���ݷa�˰6�H�.(��h���~g:��J<n����_y�l~���9�>��]W��Ap��A�VŒ��)Ӧ�B�ܛ��Q[�v��҅�p[DHl�J���N�XZ�����&���u��'��=?"��J���&�l�UEa�T3ѥe�H��=���P�����8�s��irD�u�<K�2�Ş=f����Bh�4�b�ƅ�	P�0�f
G#�>*�T���5�?�z�����}��po(�������.��5@����o�g����$���CkP�� kb�#�
�7��͞�R�d-O8�r`o�˟r�BD,os� �>�Z�Q�������2�v.�HZdbi��q¹9Wdm���iCk��`Ig~����7�5�sF�{�2a��H�T�1����5eŮ���/E�����B��2�� }�h�B]��|��ٱ�ڶ���.��i)�}B�G�]�G#�[#,��O)ף��������*�<��A���K�1��Qy�p��6ԝI�Sv�E�Ʋ�̪�t�=��o�'����X��������G�]U�8�A\�a��b�ҷ}� �<~��R7�
l����$�X��|+���*�1�g��)�_B���N�����s\�Bu>�p�N��t���'�����=,�f��Vt�W.*U�+Q
N��.29-�7i�Sj����<�������)���x���-C9�'�MtU��l��{�
M�/ަK?�ʞ�w%]�3E^�t��)(F��k�D���g�S�i!�n���S�~�N�x�]��q���pG~��H;nL"����{�sX�/��Ute�1���j׫�f����!��posz�!b���1x��ݬ�i�^�ؗ*#�_񳽜���˛O�Pzan6��p�/�2�����	���	 �Rű�P-��*A~�y��������5�Lce �yq�s�nu
��m2FWu6��"26�
8������w|�h��1{�ۃn���С����D.+��и+�_�ߟ�����</���I�N�/X�-����p���
n�X'�Kip�lP3��oU�ڠ��?��,g��ac8|wW�!��\�[ �rk7���l����*��߈��u��畴	�|��=�\�$y�-������	gȌ��x�v����v-��t�PɌ�O|�R�]��r�V�^�
�_�6�(>1MO���g8M�^�J�i'�V�
߷W4���!�T)��}B�����^h#���c)�"+# 8�({݋9~Q�6��Ӆ?��'H��S5��c���P�/��4������Uz#��a�m.�7���h9�i�ӲY�Cf���X�]�]�Ƀ[��Dֲ_��}����yv��E��b�0^`��^�����CYA�Q�f�ЯJݳT������� 1�]�a.�^)Y����J�W�'�br(g(�O�I�&i�Epf��!��Ɉ(�]�hˑ�Vk���ƚX�*����}��^�2��CA���A+1���F���J���P��O'4�X4"�M�?Ʒ��V�%jsh~ҍ�����BͿYH7��ԟ���`���E���ɸ�mg�8���?��x�/[;M�-᫚?��� ��w&�iY�Lo�����������nY'�/�W���I��⏍^�Զ��T�A�a�G��	l��0�2���5o
�铪�Y���(��ګk�|�F�sl��K��i��N���R��,�����~Eѵxd����g<��-��m��@������X?��_r��L��G��s��|r�F ��?�X3���:+�iT7���akQ�>(���.��~]^�n2S�vk�O���<e�5�Ė��|&�7A���IQ�:ux���{�L(k�����tS�܁�($�k�l>�آBS�v ~7��R
�� �\	<��a�՟�����H��e����9c��G7�l(����Skj� Z-\v�KQ[{�{��b�d�Klz�u�����aߦ��+6ܿٱ���^� P�8ݣ��X#��+v%�[�x��UX|����I�0(oI�e��������0E0�H����.��vѕ_�`ڊd��2�?!ň��vF���@� �,��s0	�3�TǠx7��Gz��	�K�6�9CX�a��펀
(���x�f�dy���(��W���[rq�t�{�z����=Ȕ�����_HE{����n�/+;_]>��Yъ���e����}Y`.��vW��ΐ��ݟp��B�07_�ĳ�["��>o�7�J�0��pܯ ���
!�^����|[[���fPh��ʇ
�[WRn�<�lAթ�ZbNh;r���X��u�Aܑ���h�f~msGD�J����-J~Y�oL�@2�K���k�0�@�H�"-�Oh@�G7d^��eCzͽkfa��I?�'hK��Rp�1RS���\'2���j�H���(�c/��,�(�_cの�sB�P�����,�qT�B[}��"�Y�wnTa3r9���*��u�{�~�!I�٬AZ��G$��ٻ��ZQ8�������*�?�u�yo��/��%��y]�jk�{��I� +z�TB����Я�������	o��2�0FYl�a�mdC$�8R������[��8{>Dly)KDo�I�K~�TRX�W�l�|"����ц�����Al�uu���ay�4tel�F��lvI?h���7� �gx����P������pz,����bT�W�����`�r�$�x���
���n�ic�9�j���8U���ɗ�<��y��$��kE��,COH�)�5��^�+�t@���g{�)�DE��W��g��+Hz�)��(�&ZL(K*o�+4�m��;x�3*/LtD��<7��1L�'	��&�č8�@�{��_"]��'�/Y�b�s.)o9��5���K����_����*�ʠژ�a�.jЄ@%�֐�ܥ�M�1�h1��c�qș���=N���HX��1�!`��w�1��qn�Ց�:��i~44�����M��)�(��w3�d+ԥ��r���Ї��|D
ys3%i��h Tqp@-f�6V~���,��֠��qaMh�/]?���x��o3]iW�G>vX=:���\��P�gD?r��د���Ʈ��
m�o���Y
���*+_@�C�Tx\\&�t�=F��(�6ϒ��k"p����g'/�F+W2Dq��Z����L�z�S|{�a����e4��v�L7��a,��[l���P��o2}�G��%�	ArUª�|yE�͢��5g�G�w�pC�&�j�ߴ��k�W��5q��fZF\�y���8���LfX�6��Z�D�<Q@�����<�z������;<�G'��\����s��E�k�)�`fU�R��r;�'�I·a����@�G�5lذg�oM�k�
71�=�i���.>��c!�(H	c&J�ki�,x3���(C-�om:ݰ��mw�6��Z}�9��g�L����CAsL���g��n��.׈2�DP[��ύ^�����lLI�Z��3_��pWDe�&�1��*�X�0��T�I�݋��l�:�K��oһ�� ���a? /��x�4�{�r4�C�ꃋ$����BW�����-���z"갅�yA�g��+��25-x!;�6ぉ��O�3���C�
p�$K��Ģl��� ���Oj��)���#J��b�*��5�b|⴩~8��#^�:g���|2�c1��9�s�B���ؚ�5T���
f�CHY4�q�Z�9MI�ms2p��ı��� _F��+Lz��\_@�XRS���`�\�l?O�MM�6��Er��X�F4��w<�ȾH��q��Mnǔ��Q1��O��>r˟����f�OqN�y�H$�ϵ��A�w�%��{�C��*���#Y2B������y���$S&G򏌍��WJ5�9�%X��86�����cb�6�����)zZ�"5U(֕��wŐ��]#]�z���k�TfF�HڟR'K�;:z#��u �N�Pš��4*M����{6]��cW�-���,1�Q�"�e���%�$1�JU �7�	���ơ���rb��LX���q=����r`-�+&eI���;�-�S�hVf�T����t���f'��� v-_9����
���}�����_~���Aݑ'c�rM����-��V��1�]��D N���2-� 6EGL�����}_w����Y��Y_��2��੆����NnkaK[T��S���Se�����lC}�Ғx���Jg���Jk��(M��5{�������Sc�ɨQ�t�S����K��'H��I!I�/٬|�]�r3��w@%:���I� Bxh�$*�h� Gpr���׿Dt	�~a��8�����Hnpj�/��ǘ�K�}L|�%mFv���-�W'��L'�~���"����PR�o�