��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\����q�?��e�I8�b�Ǽ$��"����ׯ1�V0������j�*Y��#��W(��p�/>z�<�D��N�x��#�EZ��mr�B ��rw�^T��e8��WIGE�TiUW�Xo�%�gv�Zrq�m�5�4u&W��l�}>���1B*R��C�6e<��Rb�J���WNǡ��\6�y	�:���Ђ)�-��gjm�κ�Ţ�$�[��`�>')�m�3�	��Z,4n���$��l��ׅ�wK���t����dA��>λ�� �Wh���~�6��0���#���!	5��WO%���˅�kL��%;��]�uRC9i\�o��ef<��l��/���m3أ�*$���o-���2Czsġw������ o�����Ʈ8V+"��g��_��^�����&�E�>L���8L(�ǿ�CA�r*ŔG��JV��2���ڶ�l�p�U�����:�������m�(|�W�37s�;��VT�������P#}E�3~/�D�޽zUD���%�.3�Y���苆���F���|���ݪ�F'DV(<��熪�#M��ﾛ�V��Z`J���O�5T�8��lp"�R�[<�&zH��w�)�hB��~'���~�)i`��
I��7��U���p�x ���^��ǰ�W�Lp.G�O�N�s�ˁg2ݣ��3��B?v�SB�	���7-I�(p��J��u�P���RU��#�$Z�t��'5��{�c���̨��6F9Y@J23�ї��,���̍E���}%��6���C��g�lMR���;�쮞i�z���3��9�^���?�0p _�|���ۋ�J�B����;���ȹ�G�3E\�$]Boo���[�pO�j{T��J��"8�X��K��C9.s,J����T]l�nm�����M-���w
y�a3G�+��UQ�7���ů�y7}vvDI���]��?D���[�]Y��<��8ե|3���<�W�2��>ƍ�Qbz]����z�ݩ�B�LW6��(��h7�-7ʽ�xph��XB�n�"�ԝ����{�V�Ț:���y��M��MJ�x�ޜqX���`�g�."�rh������F7:Ɵa[^:�_��6`�b�3�|��)�R��=_(K���\j��;`Є� {���0�K�����DU�/<h絺L*�@^xT�Go�\�&�̅�;n��� 2���ٌ/e�h���$7(aB�x��r'�sW�>������7e��j])�U�6�g"����:�^�{�$V�ФΕ̩:<Z�������QQ{@(�)�䮰���_b�pEq�z��P�֊�A��Z�qg��<t���A87��mߑ����6ٲ��h9|_<��.5Sϐ�`T��z�E��#�K��s�XDQ�<�����9�l2K �̠�I[@�O�e� 1)TJ�����0t�N�	<v6��2�vj;�^m�ݥEB��K��O#
���Sd��,31l?39��S�OTfǩ��+(&��{&Z�O�V lZ�b;u�SC��>O�ۭ
������*��kn�v���\�"w�J�r�����#��CJ`�JM��GR��6�0]"5$ѻ�\yi�6��ӿ#���{!Fحfn���J�/$�9���sH�v�}��1�2�[��d| 94�����*q������R� �4,�b#���;z�������|�I�:ǝx;aB8)��V�-v��jCӘX|#��y`�Xu)�z��X*&Ҧ�U�h��S�+5���-I��`�c�����&\\�oO�N21�M�����=�53�5��K��]!�]B_˻��W �:��Au������T��W�^�]�>�H/M�k�$�����sĳ��@N=�|���|&�:�6ei��|&�7Du�*� �w�W��'X�٩R�(}���y�x3t�|�"z:5.���R�L���]���Oj�٩tWP\d��w�#F+�d�yP/'������x��/$l�a�΀�����v^�7�c=d݃橕�"#�B͹|Y�UQ��U�y#��cS���7����V�u��M�1�N�/le����	_T���9ֱ���/q����*5���[�f��a�bC�l	Q���h���3�RT͟��'�G����֞��˥I,�vMd;�O�A��F����H�8֝���[��p
���+���_�r��0Bl�3P�+mKsE^c e�O9_��2b�ԉ��u蕽��*���t}�ǈ-�Q���h����B�4{_�b1�|��M�{%�.[K��68]ɻ����~��*�0���я��jI�y�5������s�ς��_Q"��Q�F ���ݵ��?��a��D�[o���K{�8���6%�V�`@G��_*p��BlD�GTғ�
��m�Rw�`y��`;U$�e%�!�
�S��������-v��@Y�*�/}�������6, ��H?��JK�!\Yw�d��Ҙl�K f�8 ��6�������FB&#���@����d������Է�.2����]�-�+��*�E�m�2grZq�l:/����9���Q{>agh����(R���i�FwH�\8vy`C����?Q�	F�L� 5��w(6�Q^f�q�D]z\l���e�r�A!�O��W�h�Y9[��M�{���qKKG��a����謰PA�u� ����4���������J�����yՈ��(oޚ�:X\��З�x�|^z�?ٴD������er���lB�?5ʽѭ T�s���Uf�&rա邛H��M��B�����W�ҧl�u�>��T��L��P��`)�Xxsd�����0������Fh� �Ж�/K4y��2�L�"�17�����`���MY{�{�K;3��?��8[���*ǫ������S΢!T1ޖk6����+�1�(��[NA(7�Fg� �0]�l�%{9���a��n�	bݲ �h{�n姘%��1����)d.D1���v$�1�BN'�G�~D���햌��2F&:4Ԭ5E��������?O\�:�x���`�{�uo�g��S�y}?+\J�2x�1Y~-+U�:Zm=�~W�O����x���(���"z�;�ڰ5�ý��rF��CY�L(�v�5=��Il� �C����N����(v��ژ��N��>���J������=��p'vL�rcqx�ӟH���z��r���%��������"���\S��j�9�O���A�U��R�v�~+��QRb�T��<���(�;�@�d^�e��=8,u]�~1i�b�"���E���|s[���r�#՛RNC��P����Q�
ү0�|��K��߂��=�ү�����}�x2#�O����UL�
�<J�*h�]��*�P�Sm��X���Q9���$�y��_�	9�ژ��	�F�dP�+�'��Eܶm�9��:�1�8�f@���N5����]��}p��./�H���BW��	BҎt���!:�ҳ�|ͭ��*5Z���n�Z�<�̞�mKh��1P���7�f.��W��g����1F�j�
f.�}��2�Ě?'��(訜�!J�W앖ظ�AɹfP�LWJ6�$�ik���c�׶0L�����/tPh���ð\��e#�:�:�k�1I�YS��-��tkv�K�K�����f&�%�S�"���BhAh� ��43z}f�|U�	�&c(�?��NIX��e=է�I��l�9SM��U�	 ��V��,x4�*������_���s�齱�qR'=�޽�y��y�F�+Sk��W~D`���ݘP�P��B�04D7���4f�v�ɏ��zJ��S�z�>ng��Bz�Č����v*�D��x)�E#��r���2$D�T��ܰ�Lz�D���W�����e�K��K��sn��C�K���ŗ���|fA�&�����R�Q��&��b��xӼ��lz�j\�,z���.q�x ���[h��j%�T��h��b٣�;�i�?��b�)�49-�����↻&]i�3�.�_	ɒ��߉��_����H�簢�4��1(�}��_�3������f�ֱ�)�r�@�?-6��5�8v�*�[���^�a�B�%qIh�p����ȓ�Mp�܍�����0t֭<���S���%�,Ȳ	S�p??u��W�`���Ͼ����;̆��-ҁip�x��Ё@ی\�gE�}�vPg>�I3�(��<�B����{�s������O�C�]���Z�qwC7U�7Ա�&2X�ؕ�F9�yӾ]�E�����,/�~w%­$7`�vǁ�8��;��]��Y�n'�CU�
��'�� �/�?��Q2}���@w�a(���%r'zG��cQ��-��Ƙ݄�A�i�'�*�A��s�Fɛ�����F�FO��c���._����'q������~\���km�m$34��m�.��4��Ȕ/q(��e��z�N���o��$ID�V��Ū�?�?[KPa��:Z�o]-�x��$�ܤ�l�N%lm���mC�����V�.�4r��k�'�?��u{��툳y'�ՎH����vț֤���F���*~�߅N���4��G�L~����nޡ�C4�S�<�B��&�ӛ�V�C����]�������'5@�@��[ƀ��.���*]D�z��;l �.���*����c�?5�����G�����7q�Z��H���k ��|�B�f�m ��y���'���ⴗN�� �N@�+q��tLt�-���� �:TVB�SNF�B�U'��w����֌���g��B���c)�����D��A5��m�HW$ג��JWhc!�C��6o��]Ua���H�!�q|h��F�\p�ggl����.F�I��`pB+�{�CC���R���q��`C3�7|�����+#�-��7ױ�q��@�X�Ѿ�v�ї�a�N³�>�
:����v�\����Ĵ��O�vETe<��R��=�6�,
�@_ٌ�Ѳ�Rw�)��t+�c\��[��ɐkD5�F|�2��|^�T(7�go�Ǣ?�c�:7�^��%�v_�r�F�.7�M���ަZ|�hZ,����VRWόc���Q֫7d��47�6�����^�
����W;w��4�#/��h�ؿPO��|�3�pgZ�M�#
�G�(���D$����y�4.5�)+�b�\�~3rFU��U����)��r�b6{���
͡�?�IV���/4��}-,��r�~ң�<���J�����\���E)��zZ�����ïv�˲ 됫�����q�M6P��/�=g�2�@��N�4޿E��xvR�ߒ��'�4K4A@ne3�Ʒv���q4˛����}d(4���냺�;h��E�$�!�0@ӾD�T�]��/��Ǭv�Փ�����zK�)%~Ձ�`O4M��Jn�t(���G[�U����5�n��|��Y��(�,1���o�">���}'}p�_�p�.3m:4�Xݏʉ���q�.?<�!>�sTo��4N�E��"��
`)��H
n��~�D�rS������y����S<��&#����p�n2a�+ws�+����w�O��=ġ���9.e�N����a��oq����Nѷ��-r��Zn�S�����G`�1_�{Ә7�c�h��*�p�٦���'�\C�)/����$ulr�������0�}��(j��D{���m���I}��3;ؓ�hyD�ȇ�|/`�@��Q�v���%V���"֬I^�8�`7T����&��UP�!���/�lh��:��������0�
�)�܅��Y��F��2*$p��tr�g�b�Ⱦ�-��a�m��fZȥ��.K<X�.�Qai'Z9hc�߽kc�𩃲�� ���!q3!:K�����m��.����)�ˆ� �e�R�E�"c��ڄ"�٭h�<"�J��]���N�y�|^>0S���"��D,Onb�~���K���{EuG��T�Z�>;<�x��}������=Q���_H��sCF��n��b�NJ�����3]�� W�i/E�jHMa�:�����Q�B���*��^u� {�-؛�#ӱG*B`�9�������J���G]�2�JP��
��3��BZyW�����"Ɖb�U��,�5_5��H�+���d��	Jl�ڐӤ�0ju���������2����8i�\�}�����6�p#����L*L�n��E���	�7�:�h���f�!\�v�CD�f@�?�t!�P,E�s�@)�	�Y���e�jL$�ۄ�U��/���޷=����M�"DS��;�Bb�r���mz�w��޹� &�����(F<l~ܧ6S$hLc*y}nuݛ��e�.Y�x����,���CZ�u���A�Z�檌��hKM��7���J�5���4'C��D^�ZmQc� B��"~�$�	��c5�����	K�$t5R$(�yKHR�̇��D���R =cJ��q+�����(����W�sF"����P�f#�l�#d�F\�gX� np,~{.��h�ѱ�yՂ�6���.B��g�ڬɈ��-����,|wp�# �w\��<i�>n�pnd���n?y�BEf�x
����m�R�M 9��6�g��j��yDO�dS�^|a��P&��Eا`x��
���hqZo�^@��P���{	�>����Z����9�p�@��]�����+��2�Pu6��ux>V�ZF��q�� I��-ψc����+�ͳ�%`���9����\'ت�x�ѕR){ԣ��vԿ���@�f��4r=�>T��TcZ�WS`UZ��sd��7��D�,�՟$oء=p�������.��$�Vigs��8��+t�	A�ۯ�U��m�>��qI���c�P��~�~���0��˒Xrs���P�9l�;	u��[ͫz�lHT�/�V��Ie���d-���7�^\]�QF�Ɍ3��SKc��HV=�S�"ػ;Oz�S�#�52���h�)9�	�Q��2��:ҷ�0U��H��ګ>��J����Dr�eɝ÷$�-�I{�#��6F4����k#y�N���b)�'if:��쀦��Gڈ.cERz�;���9��F>e���w�u#>�e;��lE��C��X�����ἐ��q�O`=���	�b'�J��W\jrd���D'7�K' �3�UCO�h��ٺ�US����K7�@�M�-*�23-�T��t5��J�1 O޶D^�P@�s�U�A�u�\������#���J��;y
����01�/�1#tu�B|�'[���v)�d�-�����g4���F_Nc��%��Y��M�[��6N�l�����,�dʵ��5�z=,���}�#S�1�,xP!����D��BTlq��0�iC�M�`�vor�VP`����%��͕v�	�P��ҧA8����Eލ%�n��a���@�Ǐ_C㊋���_[�ہ�pO��V��G⼽��y����a,K9��e�j����H7"+4;�2�6�_L<-����`����D���Πj�胙4�vkPy�8'u�y�7�2�t��c��؊ޙ��a=4�!E�d��*B��۶�(\+�w���s:.U[Ct�O2��y�M��,r�#�̇�f�&��)�R�B�e2��R�}9UTn�%���L�[�?�4��5�<���h�"�@C������!1K�2|V�b�Q��)�Kt��(��&��j,��oNXrb'X%:s}}����U����K
u���yw������h�8�&�֢)�����}�⟞��#�p/�tDâcF[K�`x 7q\�-_�n��X5�T�神����AD�#�9i d�����Ҏ�J�z���+�P�s����Ӷ��1A�D<J�VW�K��/��Jr@��i
�5�������rP��mJ�K�b�����h���b�ƑG~������x�=��n(���ee�\T�V��m���s���r	V�Ğ2�L��6h���<��:Q�N_tZ)},:V�_�-�!��A�̙ɯ�S���lO�j �V&h�4�������A��&0���y,�N'\�(���S��:��'�ݨV8F}zE͂�cc���-��c��g���<���m=�P*q(����;\�4W�'����k.BprP2�Н�����g[QI��H&�o�����0	��ΰ�&�^���^����8!�5�(d�#�;+챱�h%p�P��UK��v4{Y���ZQ˲�0��R��)}��
T����U."�W������P�/��e�ƨ+��e�Q�2j��c���.�H���~���8��8b���QۨB�c��Z��#��L<�����R� uc�5ظ��-_F�/4fn�D5( �2��چ�8&�I�~�6���_5�>ǈ��p��,���BQ y-�Ҝ}m�K�P�c(�~ �Ǟks�8m���E��;Y+�&˔��7��H t����6VM��:C{����z��ۿ�t��ڽ+y�F�����)�r���V����+��)�h�������VT"�)�?��t\�,�r���.���H��g/�C�s�n�x���
�'���5�A��5O�0,;�ڪ(�o�9Ӷ`�:8��5Y�V���K��.W��c#hu�Aa����]�z(�p|���j	�bً�4�
��k�=n�$���mʴ*e���M��D�¿9��?�du����ɷ���&5�rT@
���;�+���{��b�<5��4(=U�	����T�@�?#}9<� ~�3��w���ނ��ylP�~N�Ǎ�e/|2�d�i�::�6 ��(
5`v@� �ÜU���ttc%a���)�����0����|�p9_�b�G����e�K��7�e�;���F�� 0���#·���zh�Ł�6��@�;�L�CR<T��!
k|C	 eѾ�Z���A+h����7܋�z-jy��l��ar�2;"<�=��:?}�0�#���>���E�a�ȣH�(��A�I9��r�Dy���NsiBG���j��ȡd�����ۼp�@�Nm��`�v���F ���~��߻��B:�0�М�re��cb��v���q