��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_����m�e"kxu�Uٲ"#oB2�-g�j��h�p� M T�(�P�+M��&�[���+ۓmU��a�Z6Y�X�I*j�4E�#ل�!��0z=�^j���-�՗���:�$���_-CS��'�+;�iu�u�t���h�D���}�Ϣ��3ϧfQ��Yy��[f3�[aag�x/g_W�}�}Xw���8]ҝ�s������!#��&jo���J�㎰�:��������{+wv(_Kʈ���q��')V||���dt�	1�*��p#���W���퇉C�*E�r"k�3`��{q&�v����1I�ܮ�Q��!^t0�o�̮�EjK�� v9�"|�ByU$,����i'���0��cM�ޑ�>��n�5���=��6������Z�Lׯ�S� ���y���s�Q�����
b���o�N?�]�I�a?�s"�Y�UX�׬<�|�P#~�������{x�1���x��5k�X8z���m=tnBe)�a�xX����DM)	��]��+O�����`���mq7�j��������Ogc󣦞@,�,�Zp��g�^�\_L$4�k	H	o���23�Tɑ5�.�P,�>�GS����$��s�8V�KMm���%�U!<��.3�Sھ-���f�g��Ś�vlN/@=`�w�_H������"T
��=<%�����4$�D#��!����eݚE�|N�U���Є���E�?2�]J[l�K�8��h�D�-`��]������Vn�[A9����y�B��~��o��8B�Q�з�3ר��R��09z�Z'�r �ǈ7�v�3x:�c�}K�8lU_�y��~}����Z�R!���	Ԍ=5��G�Ւ�C� 3,l�w�q�F�F+7���ޯ�r�b$t�U)��K�4L��z`�����r�+B���f�����&���d.Ơ����/C;֐+���G��z�CL��
-?E�LGQ��
9k�9d�bӆn���x�~gG��^%�Ɨ���/JOFz��}���wND-�hQ���x�=O�T �<�t�iul�oѪ!����^��=�* �� �j��KŎv/[�)�Z�g���'�hTp��4�Wr�U���a�@���W�YO0�K"�r��f��B�l��F�d>f��~�tra�0��ԄH�]\�o�:��eK=��atbN�l�k�h��dw0����kv(Z�8cF1�n��s ��8 Z�h��}F�l� :I]\$����������ˬo��7�랻]�i�43H�,k��-P�����(
i�}�x]0�Ks�L_VWJ�W����`8����{-����,���q^x����9����:�9�⏦�^]$3����ٺ�(/�O��rEI0^A0v�W�ٯ�t��G@���{gQ�&�d������'~X�NcA�{W/�I%��x.m�����/��˴��zj�aL�w���M��z�d�C�tj������.�:I�Ƌ��<��}Y�U{���V)EnӍ|�[n���^�p�G %��@`����,�i�g�!�yY1���]����{*PZ���	�"�{��Tмj6��7�eM�{~6׎*���%k�/q^�b9$�9��>��2H�B�O'��9L���J���Y��,���m����
|���#��m�f���Z��˼c�;4��]�	h�涗��9��ec����A��ϭ�e�'�g�aWp�����
�/	&�@�
>���X���☾F(�1b
���R�'���Â����X50QF�$!��Cv�Y�bHb��NE@�Z�]�]O<���@�����rL��	�oF"b�/�{�1���:��7}0���Q���7��We��p?ɶ���lvp~oŊ��íb��T���,��]ĩ>����<��&[Q����2�S��G��?�c.�U������>%·.�1�R�)��_�%bo�V�J���kԑ�V��@�UG�y��i/�^q%T'/\�ML����h\�����:A3:�_��C>K~��6��EL+����QI�x��mWv�����pB�B׫�1� �G4+�2/z`K"��e5��쵍,��[2y&��^+��C������Z�z��VQ*��9�#��)k��dmͶ�C>�򈚉��COD-�^���l[��O��蹅�II�i���#�l�Ĝ�����V�	�VS�<���q�\����J�I�M�� �AI;�
��V�K�������Hn�� �����=�i�l$�ftY6��� ��F��G]Uݥ4�l$�O_�XoSv�pd轸���t�QQ�A1BA��0�K6��l6�U4��ӧ� ZB��U�xi��#m̆�mG3��?�:f�a�ɶqQ7�օ���������"��*R�*�Ǒ��h���~�Z>LT���U){��g��Q=�ԃ�<߆Q�y�/T-���*�>�'��l(�Oޟ�߿�C`f�V��;,s���J;��o��!v�*l6XI��� ���^ڔ��~�y3���u��\��V�$Y���I�<d&�+Y��f���~ ⏺?��_Y�"�I�:�� �
��-�
�Y��}' ���Al�tewi�\\K�+�m�����>a����-��������M�g����a��ZP���3�qW=��첵:��=;�ҹ��p9��}�
��E2��S��@I
iR���bE���'$*iN�.'$��̸) �2���P���^�[�I��� ��cw_i)�3}l�xcJ�`��AU�����ĺr,Q���Y�������Z��i��-)m�*���F<V�!����#�#����i���ʆ+8�87�h
O���Ѡ�d� ��~H