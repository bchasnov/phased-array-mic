��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8SjfSު�U�.Փ�"o��d��R]��;�۽(�O1b�c��V@�����Or�}��%KOK.�3��k�����q2��i�
Q��H�_X�N��6��f��=�>!�g?%���i�/�#��V�y��+��"�s��T�TB{�����j��IzR�v�>�aت;�qgg�$���%�S��oBrU�UC!�w��[�kps���zh�P�$Ĉ����SZh�+��ݚ�?� qD¾�w�9�b�'(��A	�@6�b�]c�J���.�]��v��&�H"��'�߲Uͽ�oN�8�䜌����<ò��H�i����h�$����P�w�7c��|)��l\�K��z�7�1K����~r6�*�N����,?�p�ކ(�I�{]��*,k�@)zg�E�yAmf�Η�Ў� ��4
A ���*EWXM���&(�X=��#jd�J�Sw�r�� q_s{l�ќ{xP�x�p+�����wD��w�G�|z�!�) ���;*b�|���|ՠ��%c���o�ӣu���kw6�/��U�&A,�o��Sd���b�p�����\�$!��c�/F��b�� �݌�`R�Gf��u)b��l���R�s\a�Q��z���S�G�Ő�D�cܥ�/�x���=�3�fU�!p�g�3��&����:�P����	ǎzT���Ń�Lh��q����;y��zx.�s���JJA�`.�ˡ��� �D��C��[d&)=���U���/�1�%=�0y���;�i��6��O���e��eo�زrֶ����IYrH��`�+�d�T򰼯�ȉ]m]s1�"�:e* 1Ҩ��\��������S5T	'�'��FI[����s<� 5.�,֣kM����������8��^���Ew��Z�'?3S���cjn�֧ĥF��e(B`U�,��w�5ǲ���"�/�p;l���a�u�Í�i�}�g!��T��o˱̥w|d�:ǳu����v����в�ҵ���&htg����%����$${R��x�v=�g�͝���\xt�.�;�4]��Sl8i�E�7!n�����'_2����ȗ$1H�z��M�������@ø�s���oFin�N�__������MI�)������̤��D�m���ݑ� ��*dU�N�XP��߭�b��Y��=���4E8��Q��s� ��qG���ds
m��޹9'�Z݈�y쨌9ڡ[~�5��Æt��4Hu�p�=Q�������m�V�ɉ[ؔ|�&��6����a%���&���Y���Gƺܞk��T�6hr]]�\�Jׂ�L�0���������7�o�rf��1��U����?t�rBzB��[�Ɓq�w(�H�495�*�3���0��0�%���R�f�X���hW���mKU�B�X�}������D�ݍh-�8��3)�*'�� :} �6����[�i�{i�Wj7�T� ��J ��_�m�f<�;j������4�		(Q����}7�����)��yQ����[܂���@��oQ=��.��{F"'+�_Ew���Fۍ@�S���o%Y��Y#�-��Q%̳Z�}z��>�]�Cނ��"� ��9wh��ɹ�e�+�T����O��1�jb�Ε��x����� �X�����I������PQXKՙ�j~�����y�9]G�0������tym���^(ޘMr�����¹%�Ul
2s�ב��׈A�=�'.Y�f��>W���
�>���X��y����xg�0�1��O	`\�O�q�iv���v�7�4J�~�F�AɌ,�:f^��~�c���V���o*�LD�����ȴ�t�k��5PP��Һ�q��H%��h2��^}�Z s�%Sm4ȚN�C��(p�]�����F���Z�` /��X9c�����H�p�M��P���&G��S[&���?�!R�z�aϘvftv�u4���5�_&Ǳ&IR
���O����B�C:��4�z�7?^�'����o��\���|��\�� �HF58yv%�dY�T����g�`C�&k����� @��f�G������ι�j�W��(M�Q��y_ Eo4��F�148!5�R�V-Y"l�'�B���RQ���!��)��{^��E���S�1�	�A5�{[�M*��ʩ�tw�U]<F~��sq�.A49��y�Uk:�d����U9 ���=�XlTᳪ��D"�N�����=�n�%�mb%� ^��k��,�#������2��yߏXݢթ�ǭR��q�8���`�AS�X�A*R�r���������hW"f��Y��cSj9�����A4�'��F�\i��S�Pܔ/����y�/;5yf�eM`�(f��q4>s�Jf���n�P�C�6�> $�%�j*�+�su�Әp̡����CH�Ͱ�����Dʨ��o�͑[�V-iI?t��u�k^t��j�D_�Ӵ�z/��@B�Lr��Q�e�C�:w�(Jyb��d�m陈Qq$�/Z��lEȵ��H.j����\�?q�Z�5_�f�y#�T\&���ڮ,z��j�^��4r���
.{:�z5�HOgD�k�AC�T|	�e��c��v٣��Nd��x�9z6�]���� �v���8Jԉ�1q�<��w����@g	�"�!�ٳO]A=�?�	�۫/������B������	�b�5�B���)��P5M�w�~�$qI�1*�W��������r4�S��Acf������nʾ����Z/I��s� �/!��E�V'DWcC�^}��i��L�1��/���Q+��Yܳ���U_7�9�a���:j��]����#���]�+'�S����,$w�����w@��)�	����F�DUR
Η�#a�!ы7(a
�ضi?���ܳ�e�kNX�����XH�"�\��C�TQ7�����)��Є>Y]�������{�J���H߬X�J�隑�7/�_�n��oF�����¾�=�/�b H�>|��kB[�,����M�^.�I V�F�Ǹ|����U�b� �P�?�;rC����|U�ϋ*�X��R�G�\��g�Y �}�6�o�9��@�*�Y٥�c!0�>a%'�+��J�T�dRr�Oe�)"K��HT���K�d<��;�,�)���_�tlTe6OTO�����ׯ<8��L��|�I�9i�H�Vmw��% �.R�B ���?��H$���-H�	~����ѣ����[�Z�&r �vN3̐���3��n���$�ZV�!r���sH��r��9d/�@�� ��(U ��>�ղ=>��nj�����J���r���k���L�Xno�������_����n���$!������
�Y�ӊP��M.@���^����p狍\�)��-(&�Ȇ�$�)�GV�+��ɮ�!K�N/U���f+(��]�$��=���s��=���U���bHI	 �h�Q���@�<J���&�O#����C�?�m9p�`	�f�������j�Il�_���^��KƫѠu%n0�SUYa���g����\̔�G�����l7qH��9��F�� ��lv5���*b�t���[u��!���M��jp�b+C��3 ߮G���qimL;&b�G��_���U�n�]�4g���EO��l�Xܶ��H�#�і�y�s��hs�����^~}��1��m�y4���1�2Y�4��`��um���N4��o̘Uv&�)�gU����Rŭ��4�k#E?�p���9K�&1d���wG��*��TZ���T}y�J	M�,�6d���~�oyh��
�e�]+�VIK�M~�=�N�	��L�(�o#���;v+��M"b���7�K�C�%�X�|�g�df�E���4KҌڙt���u����F����W��|�ֲ��Y�ӆj�=ݳ���)���`�r�����9U32�,|=���C�q��, bXpխ���>�.�6��
%٫_f��?����OӳW ��<�=�z��Š��t��Ƥ��ni� z%SW�1�ԥ�X�:E��͎m0�t����C2�Ⱦ���5���V�C���C�{�IO�۪VT$Po���'�}i<����� ���lߞ����L�^�X��0b*���t��i i�z�:#kK����q���������T�%�ל2�SuC��dj\�Ł�q��q��d�|�W����P=�]vt��x���G��P����|���h�N�Ķ���w�N	w���m�c����<�]	�o�+�1��Pj �~���m�>N0m�<^s��=�'��Fqr�ůd#T_��sx���}�_9�p���ر]	�/E�P�9~��"�߇�j�: (=��u;Z��Y�'�w�0�҂�f���śe��G�ȦN	��h��!V��Ʉ\��E�F}W9Q��R�/�3(#U�+�d�ٯ�i��Uo	=S���_�DE��.�� ���]�?�zS����8tD�$�V��Y�Z��;Y���$҂���N�
�t��u&��Ͻ���ɛ�P��-@��0�Ce5���YD� �_�"� �D�o3~�9I��S���-��[��<Ӊ @�B5H�2��O*6�(�
����{a����Rڙ�e`C�]hEp�����e�����/�&���LC�S�^�:O����oM.��p�g�X{�w�A���D�[�T\�럜Qk
���1C�H�H����5nlT�� ��ϚϣٚJ>�Yx��I��D�w�� h��%�$���K�)ut86�f}B��TY�%n@������|QI�R�"4Q�dHZo�*w`�9�U�ƚZ�U��H(�7�בL��F�S��3�í�k�6� YɏК
���W��������>���+Z����+��΂z]{��/��?�JO��0��0�%�]�s@[���-:VZ^�b(�ZDcpf�JОR�sb2l�?�Mf ���0����1e��ή�(��F4��ݵ!h���Nq�=h%B'�f��F)s��ng��h���MPzG�+��q��u�>�v�Uj�����R��������:�+�wxx�#����űI|a���d}�O ���׍�LZo�&�n��~e��_�Sk��!��.%�.暪8^^������؈冟�wq�v�$�knYQ��MN���3*$d�\�b7��H[�-9b�ZH��ݻ���]sF9��Ӎ�Ć1QY���y�~�8V2������kω���f�yªp{g>��/}��5�n��B��]�cu�1��������@�|~�6��.�;-nI��I%��_��E�{��L-�XvG�+5w�03%�Y��(�+��� F��~�;n�!Jz�ln�(6��<'��R�&!��A<�Ӆ��Bηj���4��
R�'E+�?w
ep���sU"t��o�R�~�s�ʶ�34���c������Y~�rN��ȏ"��� ק�4���q~�k�N��5Q�9ѫ�6�Ux���lY0�T;?���f�Ω�����n��0GOa�Q��M��l�s�Ow��T�s޼AaSDk'}ܚ�txBw�#��=�8�6 h� ѓ1Q�Ø%E��2%��Xt#[�)�s�������C��A�G{����ObwU-�H����μ�D�'c����2e��C��Kz1㧫b�"�E+�zCXrY>����^O�*����)�֒Z��f!�? G·�.�U�k�o~R�n�q_�p#�����ӕy�8�b�bkuވY#�eQ?��@�uq2��n�DZyl��($�ӍH�B	.��	�ڋG��%��+Z�iFý�9YN��p3应-xG{`�K ��n��ӣ.��ځ�kg>I?]�{C:�A�#̵�'��I苏��U�3��c��{��w�%�T���;�2�&�ٝ�|�ns������Obv��I�z����s�52���P�#�q�2���=�?O����hU���KW�+/�@�`l�p�����ci�g�	lI��^�f�wZ���5�@	pk3q����� �O&�ƺ�a��q_�W4==�;	x���<��Dл�1���_��g$���^��H�"�������p�٫�:��<	�g��H�oZ��w��2[�L��7C�/�u*�FY�XZ�d�!��r�A�/,����*v�>�� � [S������Χ70���P�F��Ҫ��5V�߆�B ��K[�~}��8�P��J��`�ȥ�jc0�4p�V�5&�H*�����Ʌfݐ�
���4�AA����i:������� HP�E���8X�e�ɡ�� VsCx�]ߘw�&8��ؖ�6���W3'7�&���;���S�1�������!�����������3�
���������gm�ݲ��Y+cs��[#X���y��o��b��_�s��jzAt��,I5P�/�vii	7�_s���u���1�	��j�����uM�&GE+�����NjDT;$�0���hٞ�N������l��⧰$�sZ�h���H�pl7JF�qY���GTk��0�+��Mj8��rd��/	�Cǐ�o���S/gO$x{�*r�Y�A"c��(� �d��D�����˄>�M[���m�����O�
���H˵�w�i�g]XjL�,�Bp[8U@�@�9��FY���Pc�n9vP��*�Xn!I��k1iHs�c��B����~��B?��Et����E�5�&�����Y_p�f��H��R����XV	�X����m�cK�9ї|6C�f_|���.�Q:I�N�T����Iwmr	�m���@ޱ����"-=�����Ɔ����7��j%$��/�NO�t��̆3��ٶ��xG�H���[��3����^%����)�A�ynt�w�-�/$��CP��.y�z_)Z~�����";|�v
�c]_���1���P�L��	����	#"�1�xE�>�d���,�'���+_8�RӈYIEN������枒�{�~&�Ȃ:�!��`-:���J��Y^$�B�K-3���+O6.����!G6$�m��c����v*����d�ۆu��!���$q2��sq��lN3���}Jx��{�>��p/�X[���e�7FI)�L�=I�U{���e��)�s�ŦE�ڂ�Vr26�ڊ�1�6��̽K��Dä��ހ5\Qq�!n�]���4癛�Gwa��0�}�R�)�����W�����������V/i�g׉�04���0 `ܜ펌��Fr^����Χ��	�f��g��	�pN)�t�/��崎�����ӕH��lܛ����#����u�#$�IU����� H_,�����5��5�;�����ĸ[���?=�A�4r�-�Y{������=�8.��w�R����MTQ�`h��(8<�Kꞝ�pϘY�;�y~GB0Pn��9B�[S�O
N?�o��Uh�bZu�Y3�MZTǘ�DZ�d`ղ� ��ע�F:i��=���b�T5k����~���p��ܤS.�)5��7��D&x_�Z�܇&����$��o���V������Ymcu�s�- eh	~��� .
Z��~[l�^6l�bX8`��a[�$AY^�sP	K=���]_֒QR\�x~Y��4(��j����g��{�P�0���P!+����}�f�_�h�IJ��렡DzÁ���݌�JQ�n�io����,4X�Q�}��5Ԣ��nZ�9�4{�A`�����?�:  O��	2�����,��a����G�W�,��[��`�Sq䜫�TA�"�, ����X��n�n1U�ĜC#�D�7�A�T������U�$�:?��o�D������p���OQu|Z���N�P9����Г)n���5j|�t��|ƧN*�C�+��)]n���s* ��*5vY8"fB�7NY=�m��	
~��Ou�֏��Jփ:خ���b�ݘmժD=�ڔ1��~m��9¯V-��'a��m���+8�º�|Dra���e~}X�?	�<Gw-�E�>�,�g�_���� ǲ@8	�����ː��l6�(����U&ʆ5_+�u�N�"���>�'i/}���\���}�Y�")��y�]�ڢ`dIL)��&�<4R�ٸ��ϰϮk��<{�҇��Z�$'7�
UI%��w}�*C�օ5S��^�h�B�,c���a�2rx��-z�������M����h�����#7 z�<<�N3�O���kh��Qk�������v��D6��cI!9ٙd��.�2��0w�c��᷇F��5��'�e�})��ǬzI6*�R_�����t�z� Qm2�"s4(�[v�M��U4����.�����s1I��̚8:Q��?�~���H�9j�sev�p^�6'��@�:&�G~H�U�+�f�}uw�ý��Ɍq��G������%qC;��LD�s��Cv��H����|�u�Ej�׋?��Фf���=7>�>_�m��i�$y|�TT�0�0p ���$q���ލ&�?���fZ�?"TK�u�1  �:�%��ݯ�_m�R��WsI:�8g��c��Ƃ*��vJɀ��ٕ���r��r�a�a����r�^L�L�#�K͑��p�~γŻ�+�\.���&��R6����5v<H��������Е����o��v���'2
��cZ}���t�t�z��'D�p���b{�RuZ_�g���Yս�Q���ݴ��=2����kM�sn� �W��i��8�t*�9	�ŉf}b v4�CRj�LK?�&���/�	 �z��	qv���YS�̒���C��71��q;=C�kMU�	�����l�*�G��'�����D{y{e����%����K����)�\g9Q�!�k�N��J�J�f!.��!���Y�!=*W��a��Х���?׵wE� >�e4�`0[��|���\Iè�T�q�	����P��`�%������c*�W�&��h�@*�)ڣ��Ѹ��oҢ����ģ��e$<���swJ�G��5�f�L.M�L���ز��l1��h{fN�K�S������>E�|hj"�z^D��7�'��
�֩t��P�SvfIhg
��I��"�W<�������a��I�jB����H���B�n�7p��ܭ���x>,�Hޯ��1v�=v�c�]�1���ax�;/H$�����Kh����a�ϝyL}�����0@D|Z�Ķ��`�,��Zy������:Z���M�=��БԄ�깡X��~�F�9#��"g�f`�~�R�x�ב�'v�F�rvu��ҩÝ��?� �� ^y
��?|Y��B����1�GZv|hk�:�r��߆���ln<�M�tG�\K�r�q�߱!w�5w$�2��x��S�O���R=`ǠZށS��ߦ�_4�q���2T0
�!�!�qx)*>T��m�0�P�� [�gQo����n�nА�5��N�t[}���~�p��
i ���4�o`�T�CQ�\J�l����YOM_Ozʪ(�/��2��&���,p$����s+���o��&�i}ɫ5�i�8"Q�~� �݀��L�ލ�Zw	6j�r�+1-2��mr!AH�KG.9L@w��s뭏�9��N����o�J�Ub�Z�6�� �*�}�"ۣj�<x�8�%4�9��Z�v�>d�Dr��-n���jC��e.��f�
;�@I�>�M��!=��U�D؍��u-�<�����jj�E�Ct��6���[�i�
N�WJ�uy@L�	��n'�z�Z3=��#eUZ�4k�L՚���PR�9!u�
�����)�k��o?T��1A��/��#P\a�����,P��ԅ����38��P9yy0i˹���U���-�J �'��X����S�qU�K��D!C3C�g��^���'*�wx,�j5F�#~`��j�̵�ppr��vc�^�ꍔQ��Um�i�)�>�3�5`�����׽o;��k��ρy���R����Q���J��yc�0�z����})}�`�
'A���5��@�ݣ��}�4-��vH�D*�=�i��� m�q����v	�4e�%������5��b�ﮭ�b��W7����`������P/PnƀZ��#�[ڦ��m�z6��F�X9*'F%C=�k/��i�b8_	����oo�Zu��k4��O�,w��ۡ(pR�LWOr� ��Y��Bo�,��>$���,&��z`�QM��w։6�{�f�h+�,^Ps�� �6�Tc'�(F���>�۰ߣ��"ߎ���,\�:��J��a%�����l8_(gBeu��j�d��������2I�-��&^R��$�3k"t!���-+`���p���%��4ziYw����p���7�H�[��.����.j@#t������@��q8�.��v�S��n\�^�9^d�-����z��Ē�'����{�mָA6E���zn�k�-��ʊ�?��ڂb��"�����hlöQ\a��hO���E�Zʓt~����:�!@W���� @��j� /H�En�H�B�A�*ybϼK�����$�<"���lv����A��R�p<~/:�v�u�Qo�a�`*𓩺	�4'Ţd
��ݜ����+�٭��o)\O<�4��É���}v|}�&�u�hgƪ`/T�-l���g�pH���=����)��x(�R����3����� �߲&�'���VRAr=�e��ʎ��'�1F���b���i�;�'3mVFP��_X�{���⪵?���]��hB!�����h��������+�/�dS��P���h�)�R��y^�de|� �o?\dRڛ4E3 n$�K7��-���{��f�C���U�%a����qA��$�us�K��'V�®VJ/1q�P=n XH�H73��C-q�_
��z��P,uX�(rN �DAl��տ�)(d��z�(�K�֍!����-�:\�#�ǷN�r����r����5hσ�e�V�����<�A�����p�O�r�]���4���#A���d^+%�w�ؤ*���ϩ�Ny)����r�Ga��a�������.X��{�k��w.� A=L����c�O�#<��b�ɰ(��F��mVc�el�/���<+�y]��y��%^�zG��K��N���Rz5B������*=ps��k�<� 5�)�7Ր�x�|u�4�m	Mao�K|��I�;�Ul�]LZ2./|��N �|cԶo#w������ �*}�s�>�Ƭ�c��@q��F;��X�:	&m�L]&P��ˤ�%���x?MP�U_8r�
�#������4�x��h\ǂ�8��p20@w��2��QSB�����T?͗R*Fqj�`s��?2 ڔ�ڙs��ۥX�)
;blݛ+}"�ܱ�v��(B�
�O�餰��lӐx�̰��T�ٝ��EhfW�	�^6��^���з��ř����j����SL��`}���m/�H�?
��4ęE��sN*���dŖ`�>��Qܧ1����\��jLg�_4c/���j	ó-�Q�0bbF�mr..w^���7)�č���ʳ�/:Qq� h��p��f���Zv
�Uw�z� ��\����戾В��\7ѱ�?ݶwff��9�
r�=���ۜ��Ql����;sd�99�3��l����2�{�x
2�[[���Z2�B��p�|�P��or1r`���'@q[�݈u{�%����k��e]��� �rOg/����#���ݝ4�\��X�<�zc����T%����T������W����Ҫ|�� �/�#\� ��S�t�c��86H4g}�
'.�a������h2_������i.�@�����9_yhc�@���#�7��9a%��J��'��'�P�]�m&G�ڵ-�ӆxe��;�41G��]��R%�����GqI�r���Z�k~3����^�#��Xn;^i�DH�dC��b�66��<&��K�ۢ�Ju��=�6P��}A�>�J�7��� zݾ�\V���viA}��@YٮJ��I�r�:4X���wy�ڐN8���:8��C���R�,�������2�ڑ7NG��$	g�g��l���(S��tYFwј�RT]�Ұ!��=#!9�J���wՐ�Q��X��V���y5�S	/3X~�ʹ�����\�����Y��_~D.꺇|�R&$7T$W\�a���j.u~P��xVHA�'|���c��U�(S��!�א\�Ó#n�}��f!����@Qq�?�4芗9S��uK��r�eË�-}�v (i�2|�}0�2��ʝ�<�����#��m�sY��[�G�IQ�[�hŏ�ǃ�F�	�ӂ�l���
��F���׾�yp7{�b���
��U�b�̏DȉԾ��E/a�*9��Ք��?3��ݓ�vQzF.'���$��ԝG�������[G��"�Ϲ�R�FˇD��U�-7T��[G�m�,���D�y���z�V-@\C�_d��[à�KS_|1 X�V6Xޓl��D�29���XP�L))�˂_(�)ě��l��)�����C���#9��Y�'��H�1,�%��~(�v�E�c6��6վ@��A�����em��v_�t:t���E�����	��{RJK�8���T��M�+���c��4��F^��u���Y.:��o�qI���Yͬ��g��۸�-�Ǯ��Df���r*���0���͑�4xS�ʝ=��a��z8 �A{��=��?$h�b�\Օ���8��g<�	5O��8:Z��Vњn�J�s�*��mĐ^��@�sҳQ!��$�JYE�_Z�Y H���xu���i�Z��@�!���em�_�����v��n^n���J
s�||���Ͷ/�I-��������� �ޏ��R�6�8[V�-i4V������$[��M�������M��ū�CUo��e�~ʴI���=�8��l�V;�`g�� ��-�`M�=و�� u@N�Mm��4�>3��J��}FO�}n�bS�����<يg`��`c�K-�e���S}]�滃�uc�A�-X�no��D��~jTk���.��2��jԜ*p�J/R�����s�\#�ZL�<�[U2"Ų�m��+�	�
B�Μ3!^�Ұ�^�Դ���.PA�L�u�U>�UI՞깡䚀�dP�k��jѦE�г?��	6Yt��+��ra�R�A�[�+\~ζ�Zp�����1�m���l���cx�=w�m]����Ƣ&����k�m��}�R<J��\����m�w��+^���u��2�ef�C�i��eo#U��-���o@�*[�՞�T)��p��l>L�o�����7Q�#[I����B��&���fN�"��ԁ6} >ԅ��aT�Ǌ�T�Hj"ʭ��q�� ��1ڄe\n'��۩������۰�q;B'�l���~��+CnkeC�u�r1gn���H~��B��}2�����;�V9������_�C���}\=��p���ǮGJ����Q�Tj�����e�L�r���`{��5	�>4h/�)�_%��/�u��WQ������U��T�B�S6+3/���v��-�>��k�K��-�y���x��)J�m�w�5�W�7����zG;�VŦ �����Y`�*��b���m��<�B`��3���G�� ��7	g�8C՛�M���k����a۲!�`I�G]^ɿ��޽`��\*3�  ���6�ѹE�9 v+10��s�y���dO$g��v��@���įRe���wNX��Y�MIٹ�;��
#�(R(�L�[�O_���	������:yV�3�g�{K���+-�l������U��*�wj���~�ͧ99�(��y��������A�ృ(������QW�G��Ⓝ��&�~����hߩsC}��=������Qh�u�GH�n�I�;A�7��"��u5K���~-�ڂ�2qI+�Uw-��v��㬼�N�-�,�L�Ĵd���Zm��%E���PuO�W��0���+ps�VS ��Q�翉���3xpZ�s)�H^�]W�T'����d��"���n7]C$ߠ�����R��Y5�ۋ�-����(c	F�ڛ����aQ���A���=,A|J� *�RC��~`��^�j��1 ���@.Т
ә%�շ��b�9�@Z�H&��/�#�ʊ��n���׹�˃�t�p�}ʋ}��͘���iu