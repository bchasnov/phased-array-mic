��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����Mڨ��˳0��`q�M�'���2&��Ȯ�W�4��д��|�6�K!b�'mY�`��L����T�7r~��<7�֬�a�wb<y�C�
e�E.��A��hӈJ���3����]c�w�W:C��Gvq�� ��&��� �/9�Rj�ơ����dGl\jc��{ś�'�N<�xBG�ZT�=ԣ.+����.�Y�@�=˼�_�����?6:�N��σ���;9}?��W(�ADd��pyy1ޕ��Ajϐ=��~x��f������ 򉰳�:׊җ�&-l�u���K��ݡ��L��(�G��Z��m�dE;�*�ߕ�0�ߥ�ͳ8�U@�7�滾��J-���:�1��S�N�{X��� ���+�s��p��Wu[�M
,��\�ܯX�|���/)�YE�m�d�s8�����:��I�t���d��L,pc ys��W�^3�nr�i��$7�"r�.K�X6� �s��yG{��\Y�Xl����>+b���%��!r�l#�D���2��ƌDiC8�J�b�Ē�`]�g�[���68 �k��PK"� Y?Ա(�z�W("�bqLd�s��m����"�0L��]	Ũc�����C���LU�(?�a�)m�^'p�`���P�/�h�׮{=��#�e��K�b�:Re3Q�ܹ�����Bh��^��7��,cR3���/�\�I6�%nhFl� �!Fhu���Z�G���rh��u��E�����S%���7�%1ы�z�G�'�]U�NdFG�6I�1o��U	���&$Js���Uw)�.^|�;�Kr�շ�gM;�s�-�H�����
H����dz��8�&YY�R��Ê=n?Q\����Y2�P����@G�����~�k�7+��&2CEh0�z��%���`u�p#��݄� �W��Õ�9|���Txës�Α���(_,B9�iCm���#��`%r!Ua�ᐆ�	(Dՙ�� O����I���LT,�m	�'m(
b^ش�P�"�V"���E�Յ)�WPK����:�!#S@b�;LQ�(q�/B�{x�=��fD�2Tw�{����2�m��nY�����>�j�i�#u�Ϗ��0VC�5zsKm�K�Ǥ��b�s4��w�jSlJ*1�}T��;���e�=z�B��V<_s�|Fw��]�Wp�����BӇ���B�VfMk�%#����<�[w-�<�%�I���г�a;��~�
�bUa��ʴG�XeIB\��t�>T8d����v�7�P}̗���r:K�Ŝ��q���GG�Ϭ���i������Y_̜e&��
�	��:͸��Х1�.�`3Fܝg�Ѝ�ל�Q��mm'���CxV?��i�+�Jf�o:�SU����!=�HO�^.�5���E@��Pno������E�����6���Gއ�b�"s�ϫ����k6�%X�QO7��2r��xe�U� �-��TGau��;�,8�	�P<�V���]|�-{�/�1����4Շ���x��e(w�ph�=�pȽ�#���5�V���̌ߚ�%��w@8�q{����"
�U�mP�9� {F���̌�~�v�E��S�_����w�Q�V/M�����8p�2}�5��c��Z����|���,.�%&�����:��6k��U9�v;�n1��^u8/y~x)������R~�����C$\r%�8�~��!��0�-�~[�����av��U�sG�����v����<��������֡c:���;)}�
��6�Ծ�'�	��%n��Q�;;���g���>{kT�M�Χ���)��-���l�B.׸-�͸�$ �O��BB<D\�{�`"1��ca��U(�C��Pڏ�ʘ	���^e���w���$ƍ�FE7у�I�n�{�0V�Ex�L��o�,I���$Ë#5�n���ܼMh��I���{DΞ����3��=�,�.�����;`0�k��0�h#$�l���vffgM�����~��X-1z��P���H[K�=�!b�Hދ�{��� ��m��=Iߔ_8^�پ�q�t7Ǆ��"��\���#Cm8�$��&,(�M���l+�p[�������1�O޽sstH�L��v	;�|�I��>��k򖾘n`�p��#�FI��w�5A�?�W�d�� lX���>h�?n����2VQв��'� �v���FGi䠺x"W���a��M�S$�
C�f4`�Y�n��r��y��k�&���y{J
��`y�-�@�7Y*�CzJa���qn��E��aJ�Ϣ�"j�z���-3�Y����?-^�`��f��rp��@O1m�H������q��O��j(|J������٭���p����Q�vf�����q���N�-w�i/��L��h�����k}1�~� �z�_��?�&�,�sf�Q6|��{�����$"y���.��d���ӣ��h� � Ns��� 7�?�(\�;���B^[q��S˒���H��(-��X`������U������7q��"�d���Yt���)��E�� �-�䛨�k��%���ن�3j�F�V}��$���b�Z������D�,R`N��U?ǵkT6�:+�W25k+>tT�L��r���T
�F��\��0��X��.L�h�9Ć���ױ��ɉY�N�]��/�s>Z��v��\�\۰�V�;)?���o��vɄ�L����^�
4�Ċ�	u(|�~�R��r�"��ڄV�K[Z��w�cڷ�37���c��e&Xul���_����o�����d��r��rv�se�����<�!�>��̇&Y��uD$Rjq�4���=~���d&�e�\	�"�o�0Y���7�Ư�F�
ށ�=P=?%/���>�5�~����<|$<��\������a�������ׄ��+x�m!U"�"�J��X\H+b��aSxS�4b3鹠�̞F#i��C`o��]4<�b��$k�v�N�A\��D�M�O���:v�`*o�B���\���s�vs�^����A��W�c���)u��a��EHD~�:���������$�E��_�2''����MP����6�(v39į��&Yݠ�B�9�I=q}3{�h��*���Z��|w����xpcQ�-|����h#* ��f{@��HZ��<VW��D$��!��A��0+���q�d��^�.�U���8�2CI�Bb�ы͟m�V��	ȩ��`�dA�d#��Z����E׮u��^�Y�G+�|n����}MA����p�kk�&��@3��3�x�í#7��EA)��@��ߠ�n.��^���!�?��Csm:��/�6R�TYW��(��%�����a_U V��0��&�?��/M��FS��O�30��s�5��&) �=��{"��9b�7��^s��y��� ��멘��h°I^�C�gQ���)x`~�t|=X[T]C����%a�(�T��d�ɷ�A��*μdX�n]��w�_�-PZx�G5��+����O���E�;3Đ ._;MV.���!]�A�⪁��7��>��d��@�P�xf$}� �T����� ��Ơ�g��G��K=o��kظU�>�+��W�N��P����3�^��آw��g�R����N�H6�_
��
��'�dx@zJ�^�d)\:�e��<nf��EC���,dd��U�/<����= ��d>�&�}}�r]�}%V��\���ʆ�=32��:�C� S����z���X�iK�08)�K�8�Ϛ|eXTYR�O:�![�u��x�C�{�<#�8X� >��)Tt�4��ʶ�ܮ�D\���U�ϩ�_W��4��+�^g�d,7nM@gW�yM#�^=k搛�4F�����w�6��(샧�ΝA�d<o.x�	Q�ENg����iT���逸�c9�����u�����6��Q-�i���1� ���@��Ȯ�c����
����߃����;\�i�F�C���vlR���A:��_��J�[�V�:E"s8&vh��lՀ~1&aןj�Z/�=o�}}�8�c��Y�Y�J��耙(��\ӫ�G^[+3�R0B���v���¿'�.)nM��^my#0.�ݎE���o����x�Zڠ\
���6�%�3W��F�x���hۃ�'W*<�:������ݠ�"��p�����+A�yז3j�pV&��A��o:��ͯl�������@���V��7ri �����p�ϣ�:0�̾j��
IF�bH�Ў_���/T*8pb�d�N�}^�?��S�-���.>m����p�vOz�L�O�8g7N���l�!-HID�91��W�r3�c�6q�tu�ݞ�����A�p�5F�9#�Y��Y���cD$C���콘,�P\5���h�7�sz�@R�ެ\�]��uŵE���\A��W#mx[�KL�[frӔss�I7U��@۷�%��^�'{�Qr�c?�����U|�7��PN�$X���ŅXI�s��|P�٨i���\�&�}{����N��K�������2AR���oP
4h+�ɭ�?P������3� PaZ��)�'c�9�!w�a�C�vmƂY�䵨�Q'M\y�B�^���o�o{�lr?��YF�N]$���w�18HC&�Z��\����V����l��� �ޚ�f@d�D�o�k�cU���8�1Nu�?���m�Y��1�õ�"��t��!e��l�!T�iE9�ٔ9�`д7��p���|�f�2�c}/�g�uL)���'
,s��Ԗ�E��F�n<�	pV%�wx��*ɮ�5&~�d�|���@�̌Y=�e+cq`�sn�f-R��
�l��9�9��0��w��^�_����x�!64<��)q�"����O�A�ץ���r�?��R�ad̴��^C������	9"
��x���pOL��!&�U���U�q��T<� {��1���>02,���_E��3@� n+ ��6�;GA��5ڱ���ڲ��L�~��Ĥ�oI9v�̦α��z�B�&[-T��$�ƾ07bV��e�(�����)�[)g��85g!֐������t��N�����͒�� �KLAI�n
^A>q�*hX�ȖP�4͵���Z"�%��
����t���1L�K�����p&	��e	�Dt���ٽUf"�����Qk���,�`�QWm�������9�`��K��k>{&Xj����O�a�Iz��iK��uNaeqJ��B'r�_t3̝]'C��$I .��J�8>2 �M��Xj�6�����	��g]�\%��lZ@�Z�v�=ul�(t��*�W�EO���tW����1Y�iS��?��>ػ#��^ąe�j�ُ����2b+y�����௜0��_��DMA������ip��$��Y��x�j�� ��n韒���} U �129�cm��ȶ���o�9� $SMh�`v�7���\�P���?��ά8w_���.r�t�����؟:3@��jB�
�La�3P%��x�K�a��I�l���࠸Y��9�ޓMQ����O0�c�Ge����>K�<b�X�4d�
vŌ�v#:D�E=*FN8���Rx�Ϟn�I��դ��84�$__{���6�ฒH��/_հ�<����2c56�y.=��D�=�K�~��YG0�<�-���x����J	b�YS��#�8�;:vl���}`R�<��������>�!�x뛻���A�P���iS|=u��fCS��A��W�5: m)�����)ĊSV�_�"�^�g�K�eWR7#��0�������C�[h*CN�*L��r.@��)��Qs
?�p����{Ǆ�C (`\���L��ȞDpW֡�8��v[� ��ߩߦ����8+�?���ۂ���r�\����)o��8;0�Z�����{p�v��*
F��6�"PN_�/���2E4nCG9!K�h���#ʼ���"��=#���9�~꤭pa��C�r5h�v���>5�����%��0b(�dI�R�ޔ�X���hj���X���@|�V_��x�z�o/�xӼoq��?�lH��_;��:�,ل8r��s�`�=���&OK��X5k "0R&+BH�x._F�^�P��v�����e����g��ѕ-4�֩��W7S,"m�����f�l���s��T7-H�ϾKZ^E�����0�P��G�(CrM�H�p�����TF{zո�[�6�ō��S���Q#G��2z|���V�	X��aRFp�*�p�Q�m���8�49r��z;Ίއq��b������t�'dj�ٞ������^�y܄�#y��x-\���Ÿ%C��Ue�c�"�,�td���/��SP�W�ɘ������j�]�)��^O�`�L�UJ���=���6���|�����=)#W:��U��Ev`Z����9_�߃K���j�ڙ�D��6�lpx���mGQ�V�Y�����~rG�o�i�\�{��������g��w�3��kĻAKJ�t�����I�Y�?c���T:P�O�I�w�'6�T{?v�#M��pj֣o��$-�5kf�t��b���~����u�\���e�L���+����t�+eF�(:�&ˇs����y8l�*��5��
]9��� 3�B�r�"�yGK��4��K�E�i�Ԋ�fnݧ�.���dZ���K�dV�d��ZUZ��A�P���WI�1�&3D[B�(�_iR�T�S��<�<��r	VZp�.5ؗ]1�Ƒfl�`���y)Z��f$3��$~c���o�����Z�^R,:Ӑ�� �RҰ}�N��+��Tp�a��p��Dns�l�ΨW�,�?������A[�Q��f�ox���T��(��61�m��ȂtD��\�������0�;�`8�Q:��l�L98�P���~��+nd������_h��Z+�<��h:B��j[���L���s�Vj���%xLF�И�QȒ&�Mq:��!�!`B�T�/l������