��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\����q�?��e�I8�b�Ǽ$��"����ׯ1�V0����#x:�@:&��X�b�Q����-5��t˱�)�'�*2�G@����>Iq�5!Ϥ<ؾ\���L4_�9u��!�Ay��6��[\���EM�O���?�C�����О�4�\�&�X�A\H���z2��v��F�����Xʊ�l0���;���_GH���\>������eH�|�HH�b�R'�y���Grb^{$��hJpwմb}.�,m���}uA����:�W٬o����2��v���V0��/]5.+��(�����D�1�-d���2�Op\-"��UDCP����q�0��Ȱ����y��n)9h�x&��-P�mG�&���)#̴:�?O�p�Y��$�0@s�{�����A&>�W�^��V���أ����v�~�*絈#+�$��#���B�^R��e$�BE�ԇc~�}���i�ю����u�G��C�l�a,��"�O��?3=���a��	:�<jp}�k|5��p��T�\~"`4��J,��`���	�̈�xg��t�"�$<L_�XW�g�Ŷ�f�X�ܒ<Q�v���{S��F|�o۶���P��P,�]���e���uecQ"Ϸ�>X�Xl3����mjV���֫�x���%�
�p	��1<k��	A��x�}�Q��B$��BNٲ�\��>�Ƶ����V,7�^TV��C���!���:���B�B�d��~ ���X� �̋���1�
��yZ���6>�e�E�0ߦm��'k��#�ޝ]�z�@\YQD��Y�R�&)�r����$���K�lK�|���tAa�6�f�VO��'���taӣԨ:CG�n�p�]�͹<���3�I�qZ��%X��J��"�c<�j$V��n��y��Fҡj"�ۃy.�8ۺ]u�&<	i�(���R�N�\��ٍg���4Q����s�f�1�����~Õ��[q�md[��RTwW��V��-Xx*c��OC�k~��d�ρ���f���`��2BgS&0f�I�޹��n�P��+}�^V��5�o��s�	�Tio�ThB?��
�k4s[��-���3��iN{bR��տ;�,�@�	�OL*�� ]��>gk��ۊ!���5����{�+���1�^��iX��1��S���-���_6]��Cw?3���RJ����T����2WD:��R���x��6�i���IˌZ�_������RܜP��@�-='�/\P�W\�pb6��!\!�Q�[N7E�MI�������y�E@���Q-v~F�c]+�)}���)l@��o��]��d-.�*��	r�k ���:�c��`sdZ�)�+h�k�{��8�h�B���:���v��$�? �4r�{�QʀW s�
1��b�c��i��U���>wl����z��54��@-�l�3G�Jޔ���]wי�z	�~P���H0/T��D|�7CV[s�¬_�z��w�k �)�$ܳp��e�%�N�ϓ�?����6,�A}U�
 � �V��D(��zB; �,`���g C�Y1���<ǟ�X7 �`��tyѶ������q|"Y�Cg�Z�;C(9�����1Ⱥ�X��:I�^�okŋ�'�ߎ�p�Ca.&�`5r5XR���23��<�i����u�2`
]��s�y~u�
)M����Q��&Q녤x.�������Y%`�q�Ɖ*dm�E�Z5�j�ȇ�M�d!�҆DMu��w�9r�_DW��e1ɔ3���7�A��ɼ��<�H-��� >��������|{Pc�2~Ŭ��83}?#5��B��E%ŏ���<��K�9Ze�?hX�2�y�5^^���w�MD��]Ws�3p��{�K�m)pk\�'�w��;Fe	�:�k�!}��%/���2�LH��֍d��r�l}��$%�9`�x���hP+{���2���� 0�i��M�i��K�L!���i:�N+�y?�f�V����:�ox�I͌p�T��uǡ���9�'�7T���Cm��6��Eě nv%2�}A�� ��Q:�U;̽�f��\����Y��|��X����=�ū� }C�:5�����k������b��l�8_ө<1�P�S�9oY�ï~�ca�^�G8!������P9�����״�o��v?k⇉�6"�`�⤴`��(��۹OZ������7[N�1�E���4Y2�$i֪���אb��4��b7��mC���C_O1���4k����t�l��k����xv^5Gߗ5|�&��GUK}K��������Ӟ^<}���`7{`��a~0��6��	G��R��H�؄#��Ǹ]#fP6�����a��YƎ@]�l�wk��׈As"H8o�%k��`eW��S^�}�ģ�Ȅ��VX��6����NG��<��	�&���t��3e������o�N_5�m�A1�f�;n��!Ž�T���2e���(@k���u���XDd-�l֥C�M|���[�x��,8s�ti��\�����3���ZR�š�!���O�Mx�G��řt�3�z�,�_&�L�Vt���mݮ�'^��Vē��M#Td��-�º�g�|���)�6����#���ԧfu����vTS��)����	U
)N���n�"� Y�3�LRۘ�V��ϊ�!8������ΊڄʋI(�ܕ�ќC������v*���xG���At�i��0Y��=6��9r��z¾���Az�(;y� ,���x�g�8ܝY1u���>�9��_{��K�X������^+/��P0�z�?ؿ<��J��*�6�fM.�_�q`zK�v�&�F���)��M5*���e\޷��C�']@c�h��Mօ�d���˼�F�P����K@TPP���e�Kr��f�̧�=��K�V�}�}����>k�ă�+��+c�=��ا��8m�-l��G:d>ÇѶ�$���.)��3s�P���p´��hG��I%Uꌛ�}��_��{��s��0;]rǨdEϴD�$T/7d)r�W3I��8Q��	�a;�|Yi�T�YV����qA�w3��� ��`��l��w�6���������L)�$��ª0��S˛]������h���We��Oڠ@1fy{���6��d�V%;�����3	X�ߛ��3f�#�������b2�1J��V��O�����v���'�.5��g��Ć�&S���Ǧ������݁�a����c���#������Vv��,˫0�˼PL@b~5b���#3�r�q�Ѝ��\<��jGWP�����I�d���a���P�-���j�fHm�+����!fD� ڞ�l�����6X^_Z�"P�4g��r������\6���-���@ 1=����[B���U���L���6B�μ��%q��~�0�eD"L�Ĥ��(h�Qqc_u����,�āy���|v�w\�\۽��Un�2G����W_�(��q���T��nW��d+��a=a]sV������o��;|3�AƸ��S*�����0ɎWT�$�X%K�w"F�w�,ݗ�!z	���i�����h�d[���*�e�&�
�)g�x�r�>f#��T�M�?:f�?����<`餽|�a�^W���yؽ̮���,
����"�D�2�NN�qx�(ZL��|젣G��)r��h��1ZO��ƕt11S1g}���﮷���a�A��v���5G1���)�)�w�Б�98�-�����˧h.<�# �,3�g�$}� I�k{�b�>鉼�!�j+����P�( �3֏>���`���,�_�	��_ 1�����E�J�/Rl�:_�����o$�N�&��G3`B�5\�xB���h����P���vQ8+����2�js���>m�&D�0Q)�e����%�R�^G}�ڧ�
g���]���^� �,�ڞ%O�.^�_R���yJ���� ���P�l�Ҡ�'�UxPe��v����X��;��n��#���՝ ��RlK�,�c���a�Ġ���f�"�[�-�ޛfdz_©�d��a��o5�ʿ҃�As���A���d��ua�wlOB�흴����7-~�����+Ύ�Y��%@6g���]rT���V����R�ٳ���.�"�`�)�Q�����,y��W��%��� ��3QX�PT.��g�è�E�ۉ�Y�)?G�믽��Hnc�Cu�E*Ä�d�m��LvWe?J����z�L@��a1�ƺ�`�w�ӖOAޅ+�c�0��߬)����ē���>���⩍OȘ��Fi}.z>�W���W�Yu�̝�s�?h���b���z�dꥹu�M��i��a T�nl5���hq�7mƽ��o �'-X��1[��U��X���`�=Z4�T"|[������B�F�h>?��s��t%��|�A�'��Uӽ��@�G\e6Fɹ7��L�2:Aً�h>¹�[|��&�.�SQ������y�D,8���o�^0�\~p\Pi�K��)���'>u{�jn`$��(|��	�˺	l�[������
pI�_͹���B��6)�wMH��e�y-����8H�/qs��I��2y��!o�j٩�l4�g �J��G�.��4�B(�i�ժ�of��&�#.���+"�L
��
nq�uF��+PKs�8�ܛx�OO��?��Y��u�<���Mk �T�3m��ѩ��˙��)qh&G��Y�{��L���4q�Rm#�kH���:�oos-�bH�%ӧƢ*p�g�YO~"ݻu$��x� �Ґ�
s����ſ�f�V�q��:DN�n�TyWM��;����I�K9��uNߧt0)�G*!��)\]��O#����}�3�E�~����s��>�%�m�j3y���r?R�іz��P���s�q�Q�9l�7G ��*_2�>x8�~7K��l�<��|�$P-<�Pv>:�������j@rY�:-tR�{P_����|�+7r=-Gݘ#�	�|ϧ�q�;������y*��/���5>�9
��g8�x���������
���Ʋc�D�6D�2��7BX���Kc���X��a������ʕ[,�s�'�#�(eS.N)��C���kA�����g���	�j����qQV0E��Ql���c8^�^ԁ�L�� "�v�_>�݉I��p�TX�|��"˔��**�3}��H�s��iE*���� Kٳ0�YϏz�|�������P#�TmщF�TJ��nguV{FGp��帄C�N�j�=祕O�כ�>���5e"�_���K� ~�(�I��{��uӍx��%@Q����M�+�q�Q0.�c��z��E�O{\z1r"	J�-�v����"�����\�%�H� ����i}�p��8�������XT!�Y�Up���º�t�L�3jPyM���{Ę]��<O���xt.;F�C{XҪ��L�]���'Pd���(�����H���� ��H&ة;=�Ez9���~y���G?�����1�����*�t�Br�+� ��N��cr��ɞb�i��{����}��N�=���cCY|���j {g�Uҋ���oXЋ��dqܹ��q�g*���gO��*Us�ԇ7�?�&4�#hLy}#��s۟D�86����A�<����^���ߥKH�N�&�/�e)Z�BKm��6�$'�+��+��F�C0��B�Ћ�~}:ռ�b�# ]o���RU�u��0��i�VI7ԇ0�& ��K!�7}��bB�'$?��8<�3�~!�I^�&���s6p�MMl� ��� `�� �a���Vn!�R;|�'���>/�a.�a�-Z����µpb�9� ���d�d>ƐX�%R�~�l}�K�g�{E��vށ?:�]�j�����R���7T��z�;/(��]Rmdh܂�c�8��i���� ��h�&�-?�a��u;F�.,�W��֏�κx��_)[Ñ�խ��%��Sw���拚����UFW��4�'�C�Q&\�J=5��f#�F\��e���c!���%�M@���*��o�W�բ�y�LzhQ�Ԙ��\�f(�����%bl�O�A����@]کb�M2q���R	�y��e�l�5sI���HN�"^W%=)�K%��*Q�}3[S76X���N��MhL�		_��)W28T�74��?3w�e�*�d�X��h0��
�c���U�G�TU���]���f_�W��5Q�I�\u��B�1��me���@���OH�+0"�J���uo �h�0���jT1@�})Ë�$e+�Y
�.�������{-�U��ŽK�k�p�nC�X�Nl<��*�*<w�������F�T4�k�q�
��m5F������g`��~4%�e���tv������IKK��.9�nKXD�N� �^�\]�h��f�H�$,79�4,&62����k�}��=��\c���?��&.�6C�x`��RJj6u�$h��ɗ3�hx��	�{\�
X\�mظ�i�Dmh�7\��X�VJ�M�7C�kr7�]�C��G��.�Gbr��2X���Ei�)����r&0����d��|���y�-�;���F4��gȶ��"Z�?���9k��� a���ПLl�Dϩ6��~+��Q0e��'�)�W �{<D��6a%U��xJ�~�'�c�?6�$Fx���<j�x�ɖqY 
�9��F\��`���mt��*�d��g�(�u4�&%�����uͥ�ָ�H@���❪�	Q)!V��94v_�ux���&;!yKU�vM�����Įߺ��-n�:�d�IC�&V �x7��g�A�B)z�,@��#D�vLD�~A �R�xi��Hv�2wɛu�:L��f�3����<2���D.��"ǉ��;Q3���;E�`Z��G|))�ˣ�~����{v�.��tA"���~�Q0���X[35��S������۔@�q��[�^����PML.+iF����yz��v���/�?��9r���#2E���'��SI��|>S�$�2r���-��uG=�K�V�)Wzٟ�h��TK �Fn��E��D�yF[�}׈�٠胊��!���o������ip��<��t��6�!!���~�]8~���t�J�L��^��[�/���#Ğ`��F<.�Hټ�a?�sd��5��o~�ds^� \P}����)+^/"�E��oy�J?o��qX���[E�Llv�JM�x��Vv��vWD?�H)�]u�	�3Tn�҉�I�#&t��Y<���%V!�vj�,��U�4����Y���&ҷ"%��p��XY���#Z �&�
8��c	�e4��>���+i[�kOK{��A�D��FXvN��<�7��WȂ*�tM�ݢ�
�P���e7I�kg3͇*8"�H��4X�_'v�x�Z' ��؜k^�'�������uA�8ʃ@R����p}��3%��U���5�|ǫOVb�(A(p��W0WHl�jځ�	��a���T<��Z�ȡڗ)$�DV��СeJ�Vh��*ec5��!�%���nzwn�<�k���d\#�1�z���k$�3�����W�+�on��cw�����4ڳ��m��+G0sD,����Z.1�kt�_^5��L���'\el�k�:xe��-$�'68��l!���ճ�u�$�j�)�?
��K 1���� ���H��W1�C��w�/6VT1��,�fq	��bY��'��ߙ\F�W�
]w2N���w�{c��������`8�*+:k��ׄG��Z�8��К���JQ�Қ3OԸ���Y��E���X֖�Lۜ�2IX���X�h�vLּ-�hqD�7�F�	��.�n�&?��:I�N��$8� ����ex�I �L��*�S�({�O��4S�S.E���/�x���vd�"��B���2���w)yxPq�sj��y�~��~V��j�W�zĴR0��+�6ڒ����Sf����+9H���^O�}z>$\<KΜk��
���!4ŪxҦ���"׷���p7����0�̶��m�8�G��(Q>��A��]�`U��d�6���D�]Д_��^��h��J\�j4����|\�>�^f��Z�M�n&ӈcK���R�N�ږ9�fY=��.�[�=T�g��z=`��T���]�iX���?���9�$8ٙ��[�gϵ�ȖNI+��Ƈ��R��m�]1��v��y��~�g�ʐd��P�7lWĸ��3j�WG˹u����>"*���f��,�K������"
��~p�����_�
]�1�u��Ei<�f��@����\N7���Q��KA��Ś��B�K����3�h}���"�u�D��&{�#�S:�Lr�:)_/Hv2����_n�ja����*���
q�b�D�,^�� z�g���I2�U�dvK���A�����'l�e��I8��� /��=�'���:r�/�'s4����Jh'G�#�v��+0N�Sz��ec8�����tn�h��g��e�*uɁ[Ve7��yy"� x����m�M
p�t;uuFW�+��'�m"9 �����(�feW�n��{e%�D�{�{z��^PNqn��6�w����^��G�دN���F�u�qx����'qgZ�\�\���_�<��~_�l�����J�P�SR�p��/���0Z��(������KVT	Y���$�	���N9�.e���\����?�F�⩑���AL̈́�#!v����c����ܩ�P�M�&o�<���.�O�E�fiV�^X!��x�;�lH���]h|l[��3������r(�s������ZS����ݺf3�����`PϮ�:	�9rZ��K�[ VR��2��fHr�PKˣ��o��t
�,9>g|���t���:qI�Y�R!�����H�B�qa���T~=�7o�=[�c�Aў#s�"ϝ�2�u�x&}�@{0@�����0?Dxb� ��h�G`��Y����K����0����Q�T�:�W�=lHΛ�p1�8�[�n�B)7'5��efX]z���pApbQ?!�K�6�#+\X!p{t�GH�h�2VŲ��R@YgrL�As9�Iּ���q��X�|J�P�l��4!p����x,t. !�9�jʧ�T|]��$�V�p��Uw3sM$��`T�|�9��w��8w2B�O2�{1b�bH�W�yC�Q���oƇa1��XL��ouA�ρ��OD�<s�'��1.��8B��쵔)*��GY�i	^�X��W���;8) K��I�H����z�oO�C0����pK,N�� ��4 ߤ��+��4���9fiT.=��1E3�̹�u�?�5�k	E�M�$�v*��=5m%��5 &���9��X��s�A��}���~���ny��%/|�T�t۽ب$�#qJ�Y���p��Ӑ�;�l�</~O3a�!�T��s�p�پ{�4I�d��H=`:��;]�%K!��(UJ���IK�Mk�︚ن�@�:���-�ܽ�s�u,� ��O.a���a4�y|�;�~��zmL�b%�z*?�C1'�~����K�"D'Pj�rt���(�� ��پ���e��ܐ(�� 6������u}���}���0�=?N�g���� :���G�K���R�q���4C/KO3���[���3��֌y�YeF������N�Ձ��Q�*jb���	J郘2Rf߈�5dn<,��zAȊɤ���jVȽ0�"��B�R�ݽ=^am�2���1_z��^�9���V�-�(Q@�u?�nj�~2��*���X���W�ʦ㎔�4$Vu�%�<����:����B���} u��ɢ�XǺ�B����<1C�n<�O��/���0��d���JĴ9p���jL�Z8x� (>���7W���Di���f���!�Q�A_���Y���d�A\�a3�+ �ھ����m�7P����r�d���!�X����5��<�..Ɇ��H�OǷg�-tZ�+���5��E��KU���Åϧ�IwuU'�}.��ݲ�i�	�5��\��$ܣ:Y�is�xZ�q��ޫj�)�`H슾um�<k[>�GapF�*��F_@�^�c
|"`�XS�h���v�E����~�P�������˨��~�E[F�l����l��4a��S�qLf�^"�b�� �̘ʠ��X��!P��id�j���)N��/_�:�x#��V)��Q�����)�jc�IMoB��c7N�8�J�wGYL����Ҡ}<XM�+`��;��_�̓�<��:���KY�u'I�5�~#E֋������L�j�|?S<��o��h�����r%Q����Z��S��Z�l0�b5�4����@Ƕ�E��a��CQ��;���`s�E��*��2]���y�&�������Z����Dv�_yY %W�JY� Bw)�,�@ͣ�g�����;�` �4�f̫};xe�f�,ZHi�����	�P��9���RDm-�g��c���۬ƫ�&p
Ϥ(d���t:���#��� �}���S| a�k_�x�r'i�@,����q�p5�]\�Ě|{�a���N���$���,�%�x@��&��]~�4,�aM?�����_\�D��Fp�����Ŷc�dN�Mz�E�&s�*U��g�)I���d�|�r;Q50�/�,�����b�q�Z��Z�?�P��)���2'd���t|������Bc�qmbĢ��v���(���񲰢%[싕w���=�Pu�͈��%�^�C,٭�ap��s�� ���ى��)*�v7X����8�6~԰�'�>�
��2.�|�����k)Rb-'����z�sΪ�.?0S�B�!ѿ��9�+�p.�����g�K����}�-!��hk
j38B��{��]F��`�.���E�����Ju$�+�<�z���,��&�d�#��{RCJ�F��Q�3^����p�5͇���I�`��T'�}c9�=_�������,`lP�&vH�O?͉����`��<)��"W�\��R"�m�&�o�g#<�#x-�h+����v��\h*VWV�#�M@b�ǂ��
F�SA��k��v�.L�1���6��=��$.B����P/���y,
E6�"��k� L2HAs�d$Qg�$�̬��Ŧ�b�Z���>�V�L�s�2�r˚ds~�#	��C�Օi�����h�'
7[P��%��e�KƘhe0g6�����1E�l�NΨL��QD���'��ގ��Rft�́W�\�MN�B�������\��ˇ���ͬ��;q�P&���d��|]��â�F?7$ao+��*����e;6�Z���H���^LaK��.?b:����Ǡt�ő�MFDl��A%��L|I��L�	׶]�]� �XAa�h�3�&=�M�6��=�[�AY�,��_��N�f0���Ƃ�tw��;=ǆ�3ɪ��Kۦ��xO�%	�&O�>�/���\)�
b=��/7��z���ů�૽[���O3ۘ_s�$�$k�t:X�RO���9Dǻь�͡�'�"��1����J�!��t��K�QN'mGR�[�w�/�V�g�YM	�Cq��ڔ3]����o�O!�Ru�ȍ�z��q����G@!ۢD+p�11�U�2����6�r�)��
:8������!K�i�O� ����ٳ@�����;,E�U������ۢk�	)<ʡ�U�w�J�|�w&�K�⣮���#������j��d�˖�/+�j䬋�|�S��94d�5�r<��L�
k��<��T���ؒ8����0���A�n�V���H*}{�zw�v U��q@xن��CcA��/%��P��z�*o���Kì��吱�߱�9��Ǣ��&n�Κ�FWh��� Pz�S�Y3������aL�?; (7G��[b���>�:�`*������πъ����֋g�.���J�$�S�%R�oNp�6�}�b3�AP�OQ
��S�R���c��ʔ�-���I��������,R��P:+�gݠ�j6ӊ��]�j������LT#_M�$���%�+u�dH���ɜ��Ӎ�(D.܇C�P����t��'J �=v�ɹ5���e�Z�}�����$������ޏ�l��XN�F���'c&~S��||T��4gx!e�������^��d\�M����Ҧ:��Y^����
h�X_�]��?Z6�jB�������?���X��Y�#�A���1�ֿZ�*�<ީk�h;7������_���9�1o�U�g����Z����Y/P�bף2���z�5��G��>a�8/��D:Q�K����:sʂ�����M=6�	��򆢕�0��m{�$������Mf#�"��V�5�Yqc���	3o����*F򫔤�/��nQ�Pw�	�<ժ�̢����N"��	��~);��)�����Ry ?o���ŸG!ն�4����C)����dױ�5Ց��E��Ub§��D��?�X�i�q'aR�c��&�Ԙ҃�sp-���|�Y�#�35����Ԑ�2��-�9t`��&�<S�	o��[�Z��o�QTG�(��Lk1�Q�O�	Vac��5S�\%��J�~�c�0՚�� �L/v?o�1�s�0��8e_�8b]J\@�M΂)}��oNۑk`�Z٧O�H�$N��.�H�BɼJm�V�Qo��@avq[�J��	L/�8�����.ʗ��]�4S�,ey���P'�Ȫ���C������a����/�{��bysAc�}�U\x��>��U�B���t��yd�l���<�:���H+���>�9���za_��U�M �K�C��\�U���#B%��?W<��+�?ul�ЌB(�X�c�}L��V�@5Cas�S��AB�I�fiL[���{+..?��F��ݩx���y���T���ٻ���
�[T|Nk�|d�ߥj9�<��22�jtHr�\ˍ#����<������t̀��?~ldDx����_���[ej�˫ȧ%8��ȳߤm�T�++�r��(����b2�HI�xB��5>���F$3p�0Ҹ�v�2ү̞y��\'��h�n��t�͠Ӛ�8w뙂�e-z�}�9\��YY�3�t���J=�쳸�و5.x�PI�㐓%�Z=l��5��$����@�q������>���ü��.#��/.)��h��qL]����j�v�]��Ì���qBp�8�����#1��P C���5�������U����}SR^�l��xV�n��W#eު��0H�+���/�wV$@��'��t��A��z�n��+���7��U\������wu|��t�G�֎P�ȓ�J���&@�A_��V��>�e���n�F��(���$���z}�ֆ��P[�VcUQ2�pL��,�uqP_'+X�f;�S�^��M"���E`O����<��
l9�U���=2~4�2��f�"�1˘KH��4��i�i��}����_���v�<�N@у��6s�.[qߎ;KX�<���~��@���~S���f�s!1a=f#�$ꭨ͠7�e6Q?T�,ҏ�M�%����/���]��A<5���ir�mam�'C+�D��T��,�&���.��5�j�x���ژ��y���M�]��"{of�t.�2�Z=yG���T��ϲ���[M#|V��䓋^@[�=��e��Q�?���d̡s�>#����}��nLr���#�/.�T#\�\�R0p�[蠒.|�x�����P�Q�zvG�X�`H�
a�p~���Dk�~�����s���ŷ�~�����ae���ŃS7�9�a�����9��ܚSB����+�\����8����o�/`�.6��Ji7���<��$��rpI�����[9*�z^>@`�n΄}�p����y<]ufos��h�B�����6hu
�ii� ~;�?-�_��|c���<�B���R��⏗���Z �~S;�l[���n|�Y�!�k%��0\C[���*�:��/��3b�>>�D	BY���Y��7�K2����ƛK��8 ���������A�Qea�/U���"0��Zg���Z�y?��WhL���:#�������-�,����۫��.�z�Ȱ�L#1���Y4K�(����3;t}��w}�Ҏ^ۆ���>�d�FF�<���4|x��Ck��l��A���?��RN��N��Z�>�:�����Oj.d) �8Ʌ��:s�0W;#u���LҐ�1p:)5W�Cc��"���=H���oX���LA^��3|���?k��ε��͂�1D���o(��M�GK_,\v�������\���VO�.f��k�a������>:G=�)�'�>��=��.^�#��G�@$<D-9��4�f�HDF7����'�©�-B��2:t䝷Q��b'�����|C�q�����̍e���j|�h�������̕)�M��������xc�B}�h��i7�v<Ѡ��ۇ��ᮐ%��J�u�z.�bW#-_S�r�R�����������~���>����_Y���āс@�M��W� d>�`4WB��"�B�_uk�G��	y��|B�-����0G]�Q���^@�
As���ET�$��G���_���G#x��R7�H��ڳs�v�0��c�(��2����x�m2Tj�^<�S��O;��"����{W7��N�-{�"_� ��֊)�H��|����j��i&�ɝ�(��b�֥1Y}�
6�;�*���PѽYmpT��/xL�޾E�������U�8/�2�;Ss�?�h�L�ZF�+�hD5��#b���J��$�
���
�M#_��-|�b�붞��_�6���Ә���d^�[TdXC���	N�U+(�@`0��ܗ,���{��E��?>�O��ӗ��g���2t�������IY��$u��EU~gY �T�|j篻*AnN��C��)D���0�5|�s~ 4A�FJ��STz��$-ۇ��#+3�O�iRO8}��R�8D��3h��P��
,Y7�X0�)IW�"+J��FƝ:C����`1 �ƛt^����0L�Y���e�iC�@a�P\�চ�|HIM�j����.�;�+�6�w�&��9�;���<�%�T��t7���Ib�z�HM1���*S�Ƅ7��Ǿ&�?vy�;}R���&,��tT56�#��8��L�xU6zꞢ�m%��.����U#��4Zw=\� @�%�ǭ`��m(?P��αL�$���[�Mc��k���	:\i���Ot\L�	/�~�[f����h�:�4�eJ]����)rV%;jh�/[��xۏTa��Dj1.�
}��s�Hqp"�BZp�;֔D�BJ���T+&$

�������[�6���g���Џ �d
/!�6!�!vWp��S�Ċ��VY���fw)��t�w��d�ʐHå+Е����9���0N�
R_2�:/D�)�����C.H����ĚЊ7�46����.q_h�z��}�Ck[�91�c�cR�K4���e�l�����,������S�9�l`��e�)�1\L�$���_i��5-p�T�OWJ�"p=��Ա3���WfX�j�ѻ���Y�-G��Z���W����G�+�&Z��y�QJiJˆt}}=�w�Z��w`�T�7�`�)]���_���,���V����9�����蛃��i��p�����o$��r��Ws�k�Z����]�8���o�������Cz��.v'e(�.�$e��v�I~��`�{�a�`���'���*���Er�Ƒn���E ��4gV��ԙ3�J~a�j/:G�M�t��NZ��)���?�'#k�C
h��E������q_ͳg^k��*h'� ��7s���a���֪�'�X�v[)e�	�\m\C�^(�7�Vq�ֲZ�SJ�L�oy�{�r�fn�]��aos���X�lT�T\Ll�.܊�g:Pd-�����|�K�b�N��Oqi����1�nv[��	f�֘3������@�h�ڟ��h��z��+f�l.f�V$F+%�LE��r,4l�c';E�z���tފ��~S	��p��[hn5TTo�,ۗqN�d�~naCw��2ۨ%�Bb��&�a�R��M��8�|�|�vkEW�'�	��-%AI��*��? ���#!��}2&Y�
����
|��8Y+Z=G8e���-?�ԑ&*�cT�"?L���$��,&K�87(��t� ��X��ϡ�0�����o��ہ��O���P�z�T/ci��IS�{|IgN�QE���_�};���b�y��"��Ye���q[gZi�L櫳�������E�/��y�p�⬟�����\����Hd���HQv'�4誨��Ҟ\���s�M�ł>X�� J�΄�lo���Bd�RD�%Eo���-=����Bݝth�=s�7oAW�N5�/G(a�r�*D��EW5�Pl!f������}y��y�<��%��|��R不y�\�4�[. �b;�dD�P�^��8�C��IC��5$�5�df������@��N�� 3S��Mxӫ�s�m�2������]a5�e~4���7]q�g�`�⭰]~�V�mw�%�trG0T�T	�
0Sd4Udq���71���{�������� �L���~��?�y��ӳ�8�'ֿ���y?��₟�`�'��o�?�@��O���P닚92�x\f��U���b���jJ����-,����q ���}G���0z�����lho�<�N����H�O����{���-xE�����Ψ�o���I���KW!�P�}}��M�̋;��iW|:����{>Jj�}5k���|��L#���t�d����S?�4v����@�E^�h+ _���u׎dS�L�e���KCWn/Ng���a�d��ֹ�J��{:�����lP������3fG���U6J�c�d�au��8c�NN�F<R���gnpN%�"	�&��Tk���$l@���D��!
W >Hқ���ǚ��!�nv�����4����Ƿ��O���3f����<z�T`���` �$�%V���uoN*7R�+z �L�g9D��Lu�Ȫ�-���_���y�8��0J3�$�?y�
v�}`QV4����C5 �B;��(���#�!^���'��I�vp�QN�P�A�&���4��Dl����K*��F*��g�pȽ�)Y���}�� `5���!y�&(f�����ܼO�k��~I*t�r��Ĉ�_^��~ۏ�Wy]��Q+����G�c��r4m�z<�=�猕yW˒���*3F`.
!���`��7x`���������:U�sףq���(47�F⬴in�0�ʥ��#*�K� �K�U ]w2i�9������{�Һ��?nފ�s�6O~���	=�!D�>��~|s�^IU�0a���*u�z�Z)����B-&�̜_�\�ۤ!~�S��B6<`\�ƽ5�Л|���d��
IY��*��cp�jX��9W�2�&�>rG↯*{�_06Q��@�{�T�7��?����ǽ���*c�([u(,�ۭ�.L��d�a�^���f>�Ayҏ�7�o4��4�]T��`8��&�p��}+p�B��E��E^d�5c�Қ<�E.�`� �-�^��V��)������|���OA�Ko,x?�E��q�y��Ν��+�l�����0I�y�x�
WZc���8C�|�E&�G�){���|�ˉ/��*vIΩe��h�|�α�TcpbR��-��B�E��JF���S�.��]��URH˒S���d0xQ9WĢ֔�����I�:�.ώ�㜔�4�i�6M��Z�qz i7���x���[�lM�:��]D�W������M��Pp}W&�؏�Z�*0�=�����q	��<���A ���!���,)z\�r�( yT�`S������� ��m��id���y�KH��7S�9��,����Wb[c�ZX�S��Z�R�a�
Z'��������pD�}kl�U#3θ�v`���L��'d&�be�&�\�&��ف���Q�}���Ac��PK<����\p��ǋ��Z�2��'cBP��ML�9��Q�>+_PS��m?�ɟ)�� ���}������g,�fT(�Z�&�|"�����,yνp_d)�����7�+nd�/�9>|�4�w�o�@�"2�����̖�PK��3��r�.�$hS޽B��b��.7�/\_z����T$�%n�Mxh\�2�%�y��
�ⶥ�K���y��PՆ,4s�P�X��k$���Qk���܁�ꖒ���9����e�b���85�u�c��{Q���<��$د�xw��ޡ�/PӮ�����H<K��bݡ]ؤ�]s'��\=�nC,��u?�b��dk�P=Q�Y�b��R�%�)d�1G���M-J�����!�����T�$"�����w�z�Z/���2|�N?��J�p,�p�*K/'[�fB.��k�)��>���;�f,��M�JfC�r(V�8{d�$�Þ)�K�Yn+2�3��+�Bm���G��_�����8�\i�đMc�S�F=PZ!��d�:���?�-�8꠨~uח� ���c�+��k�]{~�Ex�+�/����9��?W�V�Z��"uƒ%A��7�k~U�^��Z�0�|J��{юk�aP 󗚗6y�LϑS�	�!�@�8:"�;X�Uk���o��r�e�f2\+�ss���JY'ϭ�5	��-�
����_K���)>�(H�o:��:�|�`5�Zd��MO n�Q�Ь�X5�����B���{A�A����Ѓ�8�\"�逮11��zR|���̟�d�����FwV-����p@���P�%�}y��p��-(C��q���o��d[3���ա��Q���(A�|%�����_�����.��w�>$�eS�2Uo�6qu� �ڪ�n��q�!u��<���f�.�`�8�e���D�E�M��7G~Rh�?��>;�'�C�&;eXLY�nL�QҪ����B*S�� _�Ehc^�L����� 
�b�* ��3-�F�Z,6�I�Ϥ��ְ�O_k�16Cv����v̳]��x�}��{	���Ś��/�$�srTQI�NtQ���n���e�U��fu��9�]��?�Y�3P���[H͡�(�uc}�WD<�WX�ji�s9)W:(h��Z�8�-sguV[C09�C���w�����P���9d��TS<x�� �a�X�"1k��1�X𠲗�����9�4��@l����Z���>R��^��d���P칈�H�i����[��Y�c�
�!����K�:8�p+���cӒ�3ǧ�V��GX��f�w��y�ָ��;�r)�ҩ�����rp��^QP��L)j8��}���ҶAo܉ā�p��U��m�S�S2s%�A2v9�O0�l*��dm�.!�z��J��{���2Y�[Ƕ�Ƭ޳�9���t��;s̪N3��X���ɧ@9��7]�o�'�m]M�q�c VS�4 �yg��'�vvtE^�mjH������MQp�l['j]uP�'�^��Pd�f���t�Ã�x�m�,�c!���'ESs}ܵ��;�Y�a;����T�6u���ߋ��-&�&�Ƽ9_�ѯ8Q^�1�*��C���-[?�������l/���7��Yܼq��+�E�z�/��̙���Q¥�8�$��3�o� ���DC�o���z�џ���F��J��d������������<� ���ԭԗ�&��/쏏��ҹ�1�{K�+�:3�QySϰ3��������w��K�`��$>w􊆂��Q%�?F�����4>�?ʃ�.������r��L'�yZ�w�����N$���6ӛ�*JǼ�Z#cS���� u42��v����LR5�,g���U��5��g�������S*e,2���{3W�ԁ3�%�u(B��P-��
8"�s�`��:�$^�?n�#�-ٛ�����\��b�+��h�Qd����~�:8����A	�ΕEEnz�����5�9cG����x�m	WM��?Ay�,�?CJ�$s�u���i�qG������iG3�>�xh��z��ǙA�%0j�� }"�Ƭ+�6��o�|#���%�[��<B �
&Wهr�ֲ���A.��_ ՗��v����a��3P��?��ưOR�Π5Ћ<�Fd���i����!��F_
�S��ʂ}CjO��J�����kRp=?���ٷj��]�����j�H����ԩ Z�l�d���4tm����@�A���-ˌZ��#_��O�V8e�_d�ZPZr�9,���<�N~�˵N�������T��4�O�\�N��<�hb�;7{� ��}� ��լyQC
���P��H��(c�{X�0Რ���0���9���P�M-� 1		_�#G�ι�[~��}��d���qh����G^�T-+�܊�+����;��Y���(�P�Ox� �R�u�	Y3�ͪ����D��8nۛĝTӮ=�-X��R�͚L
I�0�/B�áJ��6?n�*�8C�*N���`w��`c3�nx���I���?:c�/��1�B�gZ�B� �_��v!���G�z��m��S����i)q{�#lR+~�W�#a3z"Y�5b�{��w>���e>2�Z��v��`�<�_0w�� n��=!���_4��EP�g4x5�[�ΓF�@_�/k�F3�ɏ��$`
��x�� Q@v�VϘ�{��Fy�EU�Yx'�J��k��NAYf �h���\�i����{��(��Jo���� �P���C�g�k!i3"�1�{P����2�M�Fe�x�ل? ���tp6VeK_]� Y�X�uz��z-�]Ms�<Ͽ��f�a*�8\3ɋ��RX-u�N����L�_�_J�����O�J�8��b��ՠ�^6�p��Hr��Kn�(i	 i�K��g�!��fґ'�c��t�$7���߮ě�9jH���)��ΖP�z�	_[��k�w�� o���<�y'|���8���<�͋�t�=�?y�J�У�(3���P��yl�WO���c�nkH�v��q���$8��6�Y𦕙�Lj���ķ�,ŭ� [8|�1�g6���u'i���u���k� OR�<ܽ�E�ans�Hd���oR�X�_��x{-�����n�/[+��	Y��L�"���	^��r^c�l����t���\�z%� Vk Da�!��ue� 2qI�㪐�r�xy�S��gcj��nĝذ�04�[�г�"ʔ�1VE�I{�yҗ��rSY��7� �m��U�w#�GK@\@�jH�?f�� @T�P�'��"Y��,�t�.��N��2���6����K���V�hHwQ�;x�A�+�)��8����%���[�=�>$۴M�V�[���dJ��^`n��W��x����p"����s&����W�Zx�R��"��MK�l��#zqԝ�u��f��	�x�Ӑ ���PO�s]!��(��h��Ȧof4���^DY¥��=��C��]dy��0�'�}��?�v<��H�L��#���2�&�vM���@�$�����KY�����֧Ѳ���"�#q���4��|}��H���LrB~dn���!���h� ���(q��)�j���I+�n�'[C!l����xN'ڟ�Y����A�#;�畦����[�Vnu+��;p^
���V�[S���?���:�AZogX�Y7r̝�;��<$]b�w=U�]]�bsPE�F d
�>�d��!`��;@o��
��z(?{��8-ᄂހ���׬��1������[[��r7ئM��� \���Kab���F������d�f��}Iz�6Z���tI���
!TJR8~�:�bҔK+KwGt�.�0��R���|F���iz�3ǘ&��9H�&d=nK���-9a�or�Mj���R���\��Ӓ��@��@K��Mp�X���
�*��6�i�/R�*DU� $��fj�%5+���1k�١[�9U�R0���.���br^E}��G���z�(���V��{���ў��x]E^��L«o,Y�;:c�	�խ$�c���$�{�h��nb�MA����;���c��G��Y �8��W�a�5~������2�q�*�i�^=��]�Bl�g�F��4 ��xq�h�"rB�[�����8����0Ema�Ԓ~Xm��7��Y��u�qvUx�$ʄ����.kx����ȫǰ@�E�>���e,�V� |������#��L����	�˯L��9��E�Z�,hݹ��1�ڐ�@G�>>O8�F��kߒ�Q�B}�v�OcY�>��|6�/�q ��Є8,e��r=����16i4�L��[���*}6�B�h �k+���_`8��8��"�O��)Z����_5f���chĒ�(;b,/�8�P��R����Dӄ�NJ6���5ˢ��Q�qҴ9`�;oGFw�,'-5I�K���	z��Ͷ����J�$��<���`��	p߅�o��U
��ւ9�9W��k~�{tU,���_��b��f!sAL;zG���/tV`�e��J�+uc�	�B�P��%�4SZ�Uc���
=/�w�_�-^��f�5:q�.>���(�d*������dhΜd�<�F݌x:$P,�����¾l�~��-'�~&YF���'I�^�kFxJ�t	�G��Y��x������0���fK�9�x�B���c�	��n��~0�yW�	\�K�㞾�:^�&�4TS#/'T���п�j:�x\�G��I��(~�~i'z�Ʂ�T�al��H�I�m4>΄�0���0�ݕ�������2ĥ���`@-q�j<��8�?w��fF��a��v��|P��'3��1�A%�E�O� �Y��@$�xd��h�4��5?8j'�������bU~x����}Qxu���ju<�SA������p9<m�S�rF ��zh��Ո��V�B�Z%տ���N{�)y�~a�˛�����يXJ�6�l��6�'?$��(�(��X��8!������(��D�ә�YX���p-�\���T��+�Tc^'7��[E����r��ך�c�S{I]4�N�?��x�!'��E}DN�l��>>���>+��4@=�A��ڏ�G�$��&�]r#G�e���8}�C��qtduc�1��T`���o�� ���Q\"=42�>�Ӯ�&����R��ٔ||�,�A��ģ|�����[Jak�**Fw�S��j�k����5��R���8��SD�W�L�#ڐ�9n��� �M`���6=�g���uj��Ϥj*A�r��J����=��͵��S�I���Wh�^G)|d�4`.���ĵ�TⓀ�Q�ݬ�Oa/@�zG���Mg�/�A2�gٰ���\X�i����<#��N@��׈�'WX I�w�04��~�����U�G�5���@3M�=�L��=��g���7�=l�� ����&Z��\}*G�׫cE�]*=I#Y0|!6=K7DQ�^���B��<S��tb�|X:�&��>��@�*j��4�����.��]���=��.�DZLPz�zcR���Z�*5�Չ:6�e5�P�bvc��#��ڰO{3���١{����ZU�p��ǋq�T�9�m����W'�+�w���¾�F!6�f��Ԏ�{R.p��)���V��!�N�Q��F!�
iia"�-&bz����8����-d�I��]Y�"�d���lRE�!0J`�O
a���(�BT��V4CG�"L=p��VVJ\��O����]6��sF)�-��:m��Z�0��Hx`�4T�s��ܥth`gD�uU���׀�<�)����S��ܬ�2��O�*��(OQ%�(�;��ZSP��Д��I�9��}N	Nq����^3TC�R�n38���-g�UN�m�z���t����݇��-�=W�1ycM���!*b��!/��ˠ�I�Ǣ`����R n��S�w�.R��_t��n��3ڦ�k=��~-�D�䮇.ɛ��+��i� �z��t�(���T�L��\�*%)��0)ǝo���K�5S���]���س���B��L��걯�u�����Dm��M�hX�F5V9�$�Y�ߠ�˕T�>��v�n���8Rh~u���n~>w:�,t#̈́l﫦�8�6���:�^(,���`Z����2�-��c��L�)�h�7��\���� d�ْ#&рkɳs��Pxa���׎��H	���2���X�;�UjdB�RD*7��4���dZk�5Z�X7u"���s�P�!�M��5�^���`ν��4 ��MU�����Y#��k�s����z��kP]-Ǖ�=��k2�0�tyZ%�ͮ@Z,�h��o�>�rg\L0���!���j�y���J!�}��5k��(�#TN[�<.z����
�s�͂�^��tI���)C�<��=��&i���	��o����� ,]��t���O�E�M��YEVf��"(���9��������2o��S�����o�!�ΘW-�����*�L�=��t����4���-�p~�+�̟��GT8���c��c5_B�4�u�-���^��,�i�lr��	)���������w>��P�Oط|��5%