��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���2�U�z�[B`�#�� 3�����E��R�=R��1��TH�G��N�����` �۠���<q��c}�޼Y%�(�"�sڙ�AӛXG�{|��AT��x�PL(�]������r�@�h=n�O�^����	�{K�*�q�a�T�FV���:`��Q�օ�H�m�Z<A�=p�Y3������ϭ�;�jHz�#D(-������Γ�Qk��c����{p������y�q�K�Ʌ&�o՗Vy��P�N�*��}f�G��g��&�W��$�R
����a��㯅�Z^<9:�G��S�kUZ($�%��]&�A��Q_�+�\�~�4�Z�:��iI��`I���E�G�&d;���;u�A���|����"n���П�d��D��+Bӏ�}��r4:җ��	���OR
Oj��u�h�b���ۣ�m���و)�j��4�jX��0�K� ��郉T���I*	 �u�6�t>'u�d�s���X�C�����9 ���?|7Ù�z����7B�5������Ï`�6����4�f�ܐ�����$�~ma�T` �P�*���3@2���5�����e�����>��tVW��oI�K�K�;����A
�f���+W[�@�#��}w}����M��y2�͐�D����3�`1��Cc(� ���L��ׄkO�QCo����0@r=5��ΏJ���E��C���12�K�1_	]�Gp�G��:��DS����٩�b�J���s�vnD�� 蟌Y���W�T|m��jb�b�FF�L�`���x(=
2��V|�y��Y�B�y}��8b����;��f��s��:�س�B����!L����Xp ������q�nm+��W�~w��O �j�V�Ip'p'7^{dp;�I*�}ރeʠ3���!��
�x���3��mmЙ�T♝��F�vE��`�q�+��\��;y��-��`��D9����g9ya�)jL$B����яB��
���lѕ��q��QM�2�9o��:��C%�PJ�������t�}�ݬ�|73�;�� ����g�5D4�B���yUٚ\�ָ�.�G��3|X ��ة
���q�h��Q��D�������!]J���II�h����:+>���Ů�����Р#6��Z�V�����EJ�Vn
Q��$c�m%��	[�ԙ� ��ԜM���J?�ւ����tީ��{ۗ���h�,�m�oLΠo�t�]�JU�&�;����^2ڮ����>ꐉ�J@���B�$���R2��4ƥR�M</���:���{2�<�_�	Q2p[�35Z�7Q��+Ux���@L{TZ'̘̿�d����X&��#����1�)b�~#���y��]�{��0���C�h�����`�@���p�fE��-�z3�F$�T�N����0q�TB��3���i(�U�v��]��Y�*�������22K�"���7�
�%�O�����l."]3��B����v%��M�Nܿ<t�_�Ϧ�4qk<O��m	��K�u�۔��2v-6�`D���X&ȋ<�q�cs���]�Ɔ���nt!�O\�7�[vIFB_Iaʜ�y�Ui��S��X:��%?OT#�>3Z��b���W��Q��� �-L7$�����1ؒ��f@\|Fܴ:	VUZW?��'U.
P�٧߅ڰW��ٻnw+�~e�Y�V��q����;.����#3B��A�/,�!���0�Io���:?�bǬ�d���'�h<�yiӢ�ͳe�s�hV<(�M��]!t����1�,PU�Eb Ԑ�Yiݒ����Zd)Dҙs�Yk:�i��LvR�;��,S��X��_�]��h��_8^h̡��)���Y�L�N�Ѓtz �fH�e�H-�{u0�$�+��-����Ї	�i�����b��:�&�aH�i+n�mJ�]����\��߉t{	���k�>�HfE���^ϗ�D����2���F� ������?B���4�����tl3Rv[�	@s賅�U!�"g�Ĉ��d#e�����W���P��8H�:��E�N�a����蜷v^�<�
�b���䐲&'�_����z�*p��=q�rt���n�?ֿ���~k�W�Բ[AO��)���o7�Ym�a��Lvu]�����@�Y�1504=H�T�����僦��fXI�"t����O�kAŹ̓`���_"��	��?��76�g_�E��I7#5���?)^`.����t;��D���B#��м2�N�=��v�4�Y}6�7�[{J�W����P��(N��B�hg%c�����t׮�QQy�E����惒�xbd�Ie8��9���^�*0}�h9x吔pϷ�&��s���V��R{4��ά>��#��Ǡ��Y3�&�2MiNv�`�i����ߩ�u�]ؓd�J��h��ϜM�E��ܠ7�o�o�p-�8�s��.�L��Y��R��;y��w]�H�S�\.r��0M�U�_B ���I��;����XI����+�
#�,�x�oN���)�6�o�݌��=I���p��6k߂�W枮��9_Щ�ŭJ��n�/����PN{��}�G< =@���y~e_�!�� ·["�dA_��@�����]����֪���
^A���+~��8�}���\��
6�_��&*�A,�6*�4]����{g��$�D����2��kAs�K=϶0l�� %��ȷ��*��.�I$-E_�����4�FbdL�\���Ɯ�rص�S�N�R��n�S�:
�/��]'�5�r�61(a�<�Fon�A�q��9B�˯�Y�h5��@�7��e��U2u�҅Y�[�j�y�[�_����+��'ѹT�	�ZVB��a�+j�ի-��F���9t)K$�Xp;��,4��	�� �Hڜ�,l�y�j�%e ����ڙX�G�����8��
~;J�����&#4�um�"jP�-Y������Dl��&`�GZ5�çe��'/Ag4����9�
��t- pi4��I���/�1z];1lm{M��/�Z�.}��J�/�Dz��Ϸ��
.JOM#��fb�K�� |%��2`�+���ޟ0�<8��R���)�Ȑ�R
�_�z�anW�K}��w��l`�\{��J��rC�'�f9��	��d %Zᘍ��wC�4Ԏ�s/�MW"nB�k2�2��\��y㹐��ͷT�[�> � �Ƣ�|)�T���~�8���M�wL|��e|��D�J͒����Bj�2�F�� �0�e�q�ПYTfg�4f�/�1j��}�2JE�w�}��X�7���/_ ���]��*	�ʮU@�s��V?�0��x-�Q�1�{xP���PUI*y^���#:��^-ϓr�AZ�`7#W�[����u#�j*�=<����>)��Xtc���G�Z��O�pw�N�D,VG���B����+Ԫ�,�c�|��?1'�XsE6�'����o+�Ϫ BC_���������ilz��P�p�7�r'�6����)�z·�-4��G��U=v_��oy�"J�ܓL<9i�}9S����l`��_w .��줦G�	z�cG߂���ݹ�R���K�ML*�
u��8YsI�)z��� @��ۿ�	йO�]�/��`�.��$�|e�t��,5�AR�mK��4cFv��g\BVڮ�kyW��
��6a��:Uiu�E,�[v�悫7���_�d�CъX����{�7m�UE��o�EV�K�'/n�&�L��ۯb���LNG�v�8T`sǁ�)*՚x������zV ���_��`η_%���b>��T^��3�E�����X"X.�.���v������B(N�.N�16��V?M�m�{&���[d�*�@(u�u�0���B�J�.rP}�V�+/vT0'���UD��lA�h��A�<,��7��1_��X�� �Ƨ�`��m���s��Q��B!1�o.�=e��bv��:���U��	u���R]���Hi���\�S��&�ǧy��h��� Q,�Txh��<�#�%�}s��،���}n�7�M5=y�۵���o0�V�<�I�:㺽2�i����g��(�:k�y4�#�&u�P\.�o���/	� �ގj7z�2n70��CT�dk�\;+h����!��)��/���Cu���%��6(;1r^��KR�R���<�C���f�~����y�d����Xk9�I[��x��k����K�Zn�i!q��oM�;����y�׊ٿ�#v�yf�~7�b��!����[���-�e��yI�̘�V9@���E�c65��� !��~��*����գ*V�_�4MH�C#�G�M����7�J�ۿ��u����ɉ�f��Gs~�U�#+Qu3��Ѵ�^p�y��YGNh9&��"^���B�G�
1�[��J�@@�8�Ȗ��ݛ��KJ��l\�~�-B���<�V|�����~@'EǫY8w7F�kN���&�D� �A�&��\&=��`1D�劅(���s���WDm_*�bh� a�\V�}��-WUl��2�Q~%9�!��?��`q��Vuc���x�n��2�O����Y���*��nT��)^C!���[�*����.�1��Y��L!�|��'�H��o�GI>�!<������=��ס�� �(�6  ���]->FUv�;
�<��v����C	zόd������7u�t֖��t��X/��V���[s�ӕ�#�]�JT	����+I��W*h]f��7���*�je�h����m���
�E|"<�:�t�ʔ���Bź��f��4`�-98����O��"?�?(��}l#����\!PfX*����Ig����bZ5d}칮��W>�!������_��b
|j�����yJ���*W�u{��9Nq݄?HA
� bz��kΪ&��9��A�B���w�֊�7!/��ƠP�,�����5��B,_ݮS!���2�
��4Rw4 uԍ��f��L�z�v��,Lt �l��$Ai���9^��%W[�d�&;���!�;K�m��"��O�b%/���ڼ�.���d�P'`�@S/���CZC�҄��^ޮ`o�Q�m��S�a���� g�%搛c$Z� �J��X��jy�Io��Cm��3&����KK� �)x�M��P�흅��-\���uo��?<��+ 	W���Z�:�J�K�a`�u�,���Nm X�<�Sb��:��&�M&T)A��S������8+7�p���T+�i�jRzT_C�8�W26Dm�h�Hf�l\���ص�-h݌�����;��]��he�%�T@�0���9�ݼ!�)nXKnekHq���$"�&��Z�Z�X&[������Zkx=�wP��ro����͎��#˸8������U��%�*_�gnF_B���'Uջ�$;r�ٔ�)]���,�i�dm�(��ϛ�ҙ�s1u�{���S�������t����T|ɐ��܊u�RD%��c��âu�<���6Cެ �Y!v�>/���	ٙp7ށ����0��`�����3�&k���k |�6�_�o�WcYX�����Ka|>�<��I��1K�\ϗ{�na�O���[m��P��D�@;No������Z�t�bT����C58*E��Y��	�,�R����D+��R\Uё�_mNe6>V	3X��,�D�����c����D���
?'�O���T�j�"��e��a��O���Y��9@/R��������Om�d�B_e���/��^YL�Z��BfGL�����&cG�A������F�����+mG6JT=ժ���T��s�p���X&�E�K��R8:NΘ�\��X�J��w������iz���ҭ�˙l� �\�������D�P�a$	�S�!x�r39!�T���ò�_ɵ�\��T)_h�'p|�uZu�'��";�`*��N �@ �h.�8�����I����
n��'�j��-�a��z��I���/��9,��A��Ooo�D��gX1�ȑI�|K����z��f�ג ���3J��>�Wby*�Q�����0����]����P5%���洷���g�dӇ,�����%Bi��������̛Oӹ|���;�.}����7;g�jQ/˽��{XM���"�PB]��b<F~5*g��P,Yu�� Dĭ��<l2����O�����l���6�Êd=��*�yv�D�}b�C��ޞ��`"R�Hqt=R���M,��p��;���z�����2�*�71�:��H6�8Mb^O�����5=F��T<5��F]�eP<�T��~��1m�fa����5�F B��\C΀0�!����[B���5�@o���'�94暽�.���=�!(�e[!�oGHt�	�R^<��6���N��A����kk��Ǫ�l�?�@��d��w��d|{y��<��^	[��_%w��V-��)���z�C���EY��QRm�b��/�6�qj��Ok��q���lG� |���y��(�0{��k����t�H�n 9X��Sda����~���"���KƧ~/���q.:*�wL����x�|=(6�vCB˳w�~�����m��@l��4��x��?-�0Ey�ܿ�#	��{`l'�m#�،�0���I���M��F�0�GF�|4W؎?�������Q�k�Q0��D��Q[&�5b��>�����E�3�%��O�ª!�������1&O5���JD�r�M/Q�Fł��*���=���G��"졘���n�f9(-�?h���۔�$	��`��M~]Ի� *d���[k̈́�-�`s�y@�y�Lv^@�����[㒽q�K�R�Wp����Ǡ�dsw�f|cFC��f�<z�CK6���I~U�W��+]}�~=��?ۏ�-Ũ�t3	e�3R)���0��5/�@rz��P������@KA	'uk������zܘ�0�*;`łzk�Yr��x5����?��4b�]�o���#s��Ć��7���2g҃��g"�ѯ!(����_oi꥞0��"3�N�#���
�>�?������8�{�HJ�lU�	��oMW/�_��G 2�+E|(;�\.
9,��v-�:F�4�E�7l����n�B�׋T�Б�\(�Bwe\�x\��*�p�nn��d��t�L�� G�B<�p�,�Y�G�2�0um"<�,�p��T���I�v߬��o\�q�r���.9�D易8����Ԙ�׹W4ĭT�{��@�B��<��u���Ӧ�$*��w1���@d5}�G�H���
֣���XCV	�]�}���q	΁0ay��ߠ{Aצ�?��Q*�}^�/r�&��,3:�n���O�P��u���߯[�vD1Xn�acw�� �� VNQ�S�b�V�T-pf�l`:GR��B�x�,	����%�0)4��5(��6��s��fԭ׀/7X�h--�L�%^��7�(#�^?I�?i�ZJ��!���"����y+-�Gxh�.���GF9���;ěL*v�4�J�$��I��b��S3&�wJ��|����X_,����ny�ǀ���9%��i*�㵩e�oÿ��uС9��c�t��l--�a�v�_
+��J�g;��mA<�F��8>?:M9���x��?X�����l��!��Z~�B���ծ��w�ڛY@��d.�H�4])$��X Hh�ؗ=�8��]�X��3z��cZ��F����P޿�-�p�&��$���Q`渢���Y�3Ǣ3[����N�@���H(;�%�H3h���GɹĒDPB��D�*�����	���0�<�¡�^������;@'ip��6\�i^ĻR���)},�� W�O'�u
0f���(���=�_�b�>�.|�2�
�'-�ܙ�;���0����+���]��m�(��-����9��N؊;r9t���<r-�r����_�j����
��F�U�؄�L.Q����~_���FB)��8�L_��ҔT��w��h��A�$B�/C�`~`�'�m¶XV-��i��a��H;c1|lT4���AL��e��X=�-FVD�7E�G�s.�9�����1!�׌dÆBU3e�8���t[4w�>Vƙ Ђ�ʯLI���%B�>�R�p�PZ�`�^��L�V4�@\AN�g�Q c�Ц�\�*.�
>�jɣBf�D�A�2��`q����b��Y�}�T�l�)E;��_� �j+z�N9��������\���/f-j��Q���ȷ��]�E&��B�E��)�u�S[)��6�?���@���XvI�Z2� ��@ů�-�GÃ�Y�Ȯ�}�aA�h/�UI�s��&?ku���5Y�ʌtrD�{�)�ۂ�zX�,A
���I��Ut� 9��;�1g�I(��Wg;CO��yF�}K�Ҙ��I}���Dl������]ʨ�����+�h����1a!{WNx�i�=�A�/~���{��~����^}�+���_!.��!��Lxy�q��/0�5� �
8M�ӿ^*>u~�զ�l�����O۬�^S���x�ZZ�Xg�'�|V�K��J��B���u?��D���
l~��V����CX���OGht����g��ORc����!���E�v�ƶG�h� ��R"%l;���K��CwF{�Z�(܁��g�vb1�ӕ��8M��3sz:H�G�el��%lF�˘mɴ�d7fƠFPO|��fDؤh�KRj$��j����� wKQK�,��r4?����<��g��f�x�������H 5@�>�vF�G�`��1�'��,�q�"�~�"v���7̴Pگn�{�r�Q�GhO
�,W*�P�^�A���8�{4�MUX��Zo�A��"��c�}��Q�J��>'�t�)��e^���4ß�e�Wzk�#&�1)�����S��\e�|�"B<}@��Z��|Y��NR~wl�U�w������>�l�t���y��Εjð3����N����,�pZOO�ϲX-Y�����5�|>� �.��8�S�)i���Iicp�o��P�gd-����V#md$X��`�C9'�M��<pO�o}���1���K��ki���#�q��<e��z|�[:>�õ܃Lo�K巩G����[�(s��<�!?�4CØ�<	z۸0��I��%��}�L<t���=AOk�=Y�8��H����Z�#;�`ƶ��̯�5H���ck�������\�A��(Ƃ ��\������ad�)��[e5󈰛_n#��U���09��t����҃=Is��cȲ�"���iu����cc������@)2�I�	;5Ҋ���<}0|��ݒ�鱿�B��$��}7^&l��i���W���]����/�Cc���-$kwo]��Dy�j�9��۪�H��/��̰��9j��r���T��lT��9�+?��8�c��,h��3�o�[r8A(b�m2
(�<�+ߛ��&��E�m���<��gB�n��/���5�0%=�&��KM�R��!b['�"�-�����2�!�{���+y�&�  >���C)� ���W��]r<���n��Q9�M��z�]�@V����ޣ��|����|'2�Ef�J3�aG�3�1�Б��T��G �|�~��\As :X��P��D�yLs[b���:�f�ǫ���u����_�����2a�ҧg;p��3��0���Ԏ	���̑/���M2����e��q!ʕ';�I�rm'\֘h�J�M(�sd�cq��k�ͲL�A{J�쬤��*��Ȃ�n�@�������=�%<b�S��,��}F��iɢp�|��U�Mz��W:�}����l�Xӱ� `� �*��w��l�*�ӛq�T���evfx:�3�ڝ�����E��;����8�6�ydʍ��D96x#RN�q���\e	��~����(�����1��{�����؏�xV�p�� ���o�a�,8�;�g�E���5�)����Q���Ջ!�b;��e4��||�����Y��{�=v�d�r�Z������~��pJ9���H)K`E��t�1��+'�#����헺h�-�Xb����g6�c2�MsIÕ������������'��5��%��[�à"/��xe5�}�e�+/9�@oDX�q'���(��?9�o�)\Q?W�FkW�N���h-���%�_|���zdE�Pt|L������1��we��MZ�I���XA��t���6�v}���Df-��V�z��≇�7p���k��fL�W�3�:��_�kH��K��H�����C2��Q(�3�6,����~�?oX�[u����KM�v����u]u��҈��䆛��1���	k�U�S$3۴�O#xԍ���l��#V�������|돃�<&��Mf��9�^�t�.J��G�+�nޮ���3��UרT[<t�D�����8+!f�RF�ˑ2t�*2r ����ў<#�dG���3��5���p���e���o~U��E�Y�Sc��y��]���ڸ�)���8�}��d�t��wC���e����#XL��������w\>�{~��XT�o�ݗy=�R��நb���vԪ��/&`��c��ǅ/V_�!����>4V
iY����3~U0�v̀��L}K̗i����?�79�6jXK��)ϑ���;d���)S �X�1��6�������O�?È�����:��?���f��apg��[�����W��N�g�e�;����hx��`b汐�xW�r�91 �R[j��f���Ok�������㗮EW�k;���z�q��Ds���2%���x%d��>Sc�8tJd�f���j'����YID�XE��3�N r��;b�%w��ٶ���>�2<�?������@�k��2k<��iP��Rp9t9Rc���Uh��t�J���m�{���Xq��δz�fD�0+��҉LJ��w)aW��`'*�܎{�˚�-$�C?B,B�|�]5`-OV�����tъ�IT}#=��o�9S8�nQrW�<!�g����O��3l��.�*~�;w�a��83]�#�r��v������^�2.�K�%>���&ބ~g�Sx�c\�d6K��P���o���-�O�����M1����-Ԇ$�B&.7L�ؚ�[�#'}{�s����|�-��rT4X�`IiCk�1sj �!������]U�q��Q�/��}*�,(�ן?����~���S����W��Ho): �:>SVҷ����E`V�(~M�3
�7��Z�n�[�Q%!�̶`�A�ѓ<��q^������0N�L�2d�� �O#��	�M����e�i��l�񽍬�H��05�!�3$M���=��B�q��i��l�Դ�>�܁o�ìNR�>�^-��2ksFo��,2��]'��'�3��g�L�
>�v
p�����Zx}Fc��ZZ�{fOm:7�j�B[�� 1����t��a2'�l��Ϡ����8��]W<�ˊ$�x�k2�*B}�թ�h��Nɮ��S���}!�b�0P�E`74>a�����$��y�lL`��g����lw��J��Bc�LBYP"ჯU����w�ev��p�+C�hHӛt�|�UY)L���֧T���	���k��e�8φ6����FcPi�F�����%؀x��4��4C��V"k��뵺��X3�r��.k�lS7F�(���63�r���㛝��zi�65��)\V�#�Y�'�e��u���F�,)3uH��k�?,�Қ�f���������� ��aq���V$� !��y�&B�f��	;:1K�ck�%&1���>�b-��Gr<C%���-���9j���~�O�U?Y�����F��-vܵg�ף��B��q�G|[Q���;� ِqwJ�ˁ�8���sV<�XŔy���4�w�Q��삆x�xQc�Φ7��
���}�&̼4���i��������L�F�ᝢ&vG�<s̽��ɦi?-���*bC�麖 bȼ��]�~��6�1�{�e)[�𨚉�I= ��P�Qz�w�͉#mPj��&!���(m���e�������i���Ħ�4�ts�P�!,���v��P�Eg�kBo�=�jf(Q|��/9��P)���|�n�i��q^ՎVy���~c�N�j`x="i�t���w�֩�0��fQ����2�����Qp��A�(�i�E����
�[.(��3����tϥ�;��M�qE0��X��>�G���=i��6���,[W��f��!(��{���:H!�x�[=�u3��GB�;��!_�lYO��=8E/WS���dQww�+}f"�*��W���P��c2UxC_�^a ��esU���
��|�ec�}m�z\;1Ef�p|ArR��&��)μ��W��@��s�ZQ�΋7b$���5ȕw>��sUc7��dډ��Hzsa�r�P'V6�x����⫨��M;�+��������m�v�����X���@��F�UC���3�x
� 9�M�RsG~ʎCP6t;1xڢym;�a�.��B��<��
��-�+�	������E3���! ���m���y�����]j5m@�ǅ=s#M�Eʰ�L�I���Ao���TfZb�m��*�����D���s��2�i?����x��մ��l� ق ��0	B��r�O��w�\����5��|�����(�|�(�Z���}2���,���
+��:L�cz4厎q�K8�@Z��/�%�u�&���*�uθ�o�1Bi�h��l�� O�����"4w��77߫����2m �w���3aJ;���~�|�vc��q�.�������Rw�ᦢ��/Tm��w�ؤ��K����9M&X���v�� !��S��gF�"%�
]�0�n�>��
g��*��t�T'�N$���P����2�	]V�d�*�;p f8˒�qj߅m���H�4,_��`�����"l��L�^�r¥�SS�O�uy��Ԁ�Y��=ι��+i�s���CԮ'�Oi�^ ZP��U��!E�!�(-| �Z��|��ĩ>ee������{]�"�H	��:�|�����������Ǹ������P±���<ٙ�^!�+�?��������?gأ�|���C��\#�_��sRe���]C!�M:�˼���_L���D���~����2v������6У�'��0��+4�����h9l. �߿�Ϳn��QK=������{X���jXoW�W��*��S0���+��F}aA�*���E{aL��=%e�]Df���ۖ��N�,�,B�sa���M��m��Ci�D���ɐ��F����[8r@{ܗG6��י�"�[��v�˂�����{��z�N��w&$�~V��<ͱ��>ev���_�!ϻ8¤i3iWb:�J��t~�
���+��Y_G􍬻Nnϟ(�K_�v6�3�3����gJ��\��C���-�m�Ե]�#լ����iy��C����������
K������n���	��h�eԲF,Kj���R��X�BB'ł���P���'�oW�44:d���+ %{~eZoܵ�kg
��t"3��_�������g�����ܽ�%V�܏�M�����,��5��p�Ů�<*�|Qpd?p����l�&�4OEj�>���>�vG�P�����̳��@~��ta:l�+�����d���	�g.��"�-�ⓩ�fpG۳�#�����5�Q�u`�;�"_I��F3:I��6�|u~��8%����k�8�ޟVA�0!��#^3g�M)q��O�1�W�����
kO'20���6�hnioC�|�vh1����*�Vݿv��H��$E��/�Ev�G�8� �4JU���P�|ps�b��Qf�)ik$�/مXW��I+ϴ<gE��kϐ(<��v�RMw��ڀ�Zd-׻�v+����)h��\��b{�at�}<�Ο&�y�l� L��M���B�T��H��i�ҸG��%��w$K�����X�ܑ]�uN/�m���bx7MH���^g E��IFPh<���k���J�qj����PN��!iVq,������A�D�-�Z�9KŔX+�PίL4ں��j�Z�u�n��<C[D�����B��$��/�Y|�tY�j)��a(���0uo]�`������	��sX9�p3q��!�:�iϥ����:�������]����r\ӻ���)}�
�yEJ�~I�!ڐ��J<tAy+&7K�D��tU��==�p��e])���g�,�3�|�2�,���ϲk��C�wYr�ͮ!/����8����ց�Hq�-e5��j��]�.�kJV�(��*�6!��4�#�{��!H���f�O_�Hm w6.�E� �ݡjn�A�nO�����7���{^>�K�\����\�"��F� n�1)�[M��B�ə����B�a�rwL�HLHڳ���]�L+��/�\��@�1�Py��F�΁���#��"�E�L�­�BK�t
����o���(iJ0�2;�M�R�DL ��$�7Y�+����_�ͣ��)3z��F���������.Ia���F��/w�4����`��1�e���.�h��M�6�w5"t#�N�)�@M���-�&t�P}6�R�D�>�Ȋ:T�6�{��2�H*�1qZ(��<&>H�|��V?��?�(���;7,�r�L��m@��Ji���c;���&5'�-F�>��yiu�%8(�`�8冠�*�חa�ڻD���c���(���S�O���|��7J{�e�9D��2����/K��c�(��5�43~m��'OB$eXY`f$�X��ȈK���{�Zi�4s�P�HWM'EH��<������������O@��Х[�|M���\���)��JN�6t����~jX�{^\���y�6�w�$my�M������b�u9��}h�L�$y���뗱�r�;$���<��v�l�2������v�t�Y����z%�m��/���b�u�z�O��Y{���;e�@��ߢ^���bЕ�����L~�[pJ�In��ם�^~���WU�"9�䟉D�����º��%ݹ�1c��zz���q`��H��R;���Vː��47L2�a�X��S؟��Q.��K�~s�J�lߤ�x���u}͹�G`2�l8|ǆ��~�)���xF�a���I
޹�{���>GW��࠱������6��^�Ӟ�7r�8���t�z��ռD�>x��^��%�)�2�)T��ۇ-��+^wЦ#��s��Wo�=w��t���]������[��n��U�<���s���qȫ-_��f��n	�����_�yO�lZ�?��D�U���J��&���9g�t����%���H1wx��?*�0#-[~Mz�l��3��\A{�pΐ��|u^���뛑DU��8@�>�D��y�c�b��`aC#"���� ��ؖ�x�d�;qk�φq������mQهm�f�a�֠h��P�c�� 7�r!�C�r�$k�7�gM���Lny�
+��	�X a�����2����4��M�C/�d�g���fc�O��yb�_��7�G�d.�`^����P*��1�{	�<k!����]��`� a���6P��m�_ N� �%�Q���[�l�
2%�;��vm6��`(�'�E�b�U��#@�:n!t��V��X� ���/������ֆ��m�X/?�M42�C�[>�A]M�
��/|�Lr�hl��$9l�ԭ�oTg��D4�b?�L�!f1z@���P8ʤPu2n��i����Ie�$XIg0g{���zf4�|1\-H0�z(P�/�*�\
{�����v�UP�1KDW�xdCu�4� c��l��������!�o�a�=Еx�RB�e���8Vd�b �=��ɟ{�tK9+<��y#���N���'���?0X�P�oQ��ܓp���Sk�T����m}��j; $�B�Y
�o�	M@�~��x#�S�^$\�n�"{AA��s��h��[����鸞>a�������S��sU�b?�JUK.��Z���nq���eX^�!�ϡ7X=�x����B��Jg]J�d/U�����Q��S��rR�<��k|4\){�I�������БC��(5�D~��,nj���4��.�Hϕx.�lN�	�]�a��
��a%��'�S�3W�/�Y�1Eۄ�,}�l?���{��9h�!��Q�<>j)%�S��g\�F����h	F��lc���bc�VI��zC\�����8��ϣ�s���X�(yAi�b@<2S��uLrL��a���?�Qr���s�Ĭ�����i��\E�ı�b�[�%�]��������j�y',�w��;�B��k"3�IJ�)?�bKՔ- ��àtN�N)3��O�!Z�t�khZaD6�9���3`���N�p�F�N�g5�v�I���N�k��ȷ�i�ߛ��;����ޟX�cL"��\W�� Z�=��Q)W`������58�Y���x�S|��00���v�ɜ�"��n&��To ���G���`��h��v�Y의 ��CPOT�4Si�n
�.�^�Pt�?y�I����0�Z��`�s��L`t<��.�2"�L���e������MYMۡ'{4��';o���Ęv�L�����oe�?kR�	���](�� ��o+�*Mq
��8L�Ll)B#sPc�. ���-��0�&�)�Z ����	�Ö1㜌y��[;��P�!p��a��U���ǵ;��Hk7�����P�-ְ�pR�@����5	Z*��Y��;�"�D]�{��3w���1��'28��N�Y�1q���GQjі'���
���l��U��]�Q����S��G�1�A�%��&FZ,k5�RS�X�8CLi6�?<������iw˛w"�[�/X;�D	�zm��6\JqG�;��䭸g�d	ot
(9`��9o�K
�~X��r*�ߝ��Bܻ�>�����Y2%��m�cw��Rgt�X�EŮ�H����X�����N��I�ep���쬰�>]�)o�`x������<�H�ݲ�^u�V�!S}>|E������x8�0���ѡ��.n"�O6Gf��P-�f�j�ڙ`�2��^Ok������M'l>9�ڒ��m�8��~]����đ�vY���Z��V�&��(Eԉ�k͙c$�KTa֮��_������#�m������N�������a͟�̈́�#��\�>��^��g�@�I@�%;r/��
�*it�Ȃ÷�L{�����v�0�OZC~�@t�K�{b౞���)12ܯ�LU�\�^��{�Q�tr gQWLc:��?v������Yz�5�����(�RﰝI��@�^Ɲ��q\Gf
��8{���_����tz�/���H����&�[�u���Hn/ܐ�p#�t��
�Z�[�̮�r������t�Fq�!H1���7�d�.�au��JC�ƠU����^Z��JW�}��^r�D�I��kD<�̊&�X��2�k�dl��K��n�R���BT���Q@�� c?������,Z�a�DA)>�-�ĉ�ID�+ۣ�p^�#	&?G��5r�hp^�)�#ݥ����:����f S-�#_ �$!'���cB��ªaؙW�Y�UV(Q�u�o���եf�`��id6!��&�{9�FЧ���X����P�#�.��Eߑ������t�}c��(��������Ev4�q�U�f8G�c��� ��� {��\�wU��P׋�!�A�������c����f���0��%,x�+Iêt2�y�n���Ƙ�֣�.��8Cy4M����e� ����#kMH�N���d=����,���3��^	`�V��I�}���á��`��hk1;��w|?3GϺFM"y�݋�2?�"ƹ' =�c�ݍq��4���9���Y��;�ck�9��X���Zj��BP��ӂݖ�Rwhq���޶���F�0h����ա,%U�z�� Z��{��䆜�،�(�DA�,�$�ΜT���9iK/�2�P�2r���+��.R
���E�L`"�%n�#߰֙����d�i�}�����cO;��qde�ޏ(K���bbj��b�	�(�P�7F�6o׎��r1u�.�-�.|�i��X�aq��z��Y��]Y. �B1@�*ޑE��k�;�,D�Zg��R�G��W!�Wm͙����p��vI���9�Pv˱)s�����K,��\O��k�"�zm ��y8K�OI�f�1�Ĕ��C�g��Rn��G�E��Y٦��H�H��ݑ	w�&`&�9^����@U���<��^	��^	�)5v�y�A8,�"s�F��>��z&�]�{Z�2oa��!pﾞ��g�o{S�,������W\�F�I~��Y�/�6vF��P�e.#s,2�@�D�9G�~���`��5��� ���cCVR�<�$k�D�-2q�ĝ���/"�_%>_�㮲)_$v��H�](ُ��￰�s~9W���".��Y�V�k�AU�����j:�:q��)j�`F�.�9 ?�Б�ݘ��a��@W�6�[�c�!���E�I1*Q��Ҭ����2��E�`���M�����G�w]�eoj���S�o�fL[C/b�sN `��r�����#�*{��������L���f3iS��X��ܖvﺛoC���Ϯ��1�0�$����(���*a>elV� J���`�/-�$ ��4/�G��#���s<y�HUJ3��<�t���	>�y?�20�w��K��K�-��#��2D��9�EG��3�X�X>�0�6W_0��>o���jE��?��:˥�t�9���0��Q=ˈ&S0������Y$�S��(S����73!�4�ۋ����T-�Kw��$�B�*��sʫ��o�
V ���
�W�{�A�a�m��a��jC,ͣ�Kݎ�k	��Щ� �����9>��ʕnQw��R<�8�m��&W�����Bnx�Y�T����J�iF��xWZ�ߗ�h�eGr颽��jQߛ�'����;������Q���Oz7̄9Iky.�5!�_�|�f %���w����,�B���X�y�gNEu�t v)�apz�(|�7�}aX�����LpwI�Y�o�q�#!��PW��v��ba
����Y� �b�Z�������#@@>��%	�����M�FM@e *N�t93㇏'���yX��p�}-�9-7`(4���r����eǞ{��ih����r(ҳ��n�0�3����Tu���L̪3I�������X�[x�<�z��k^/�Yȯ��F�9!?�r���|��� .;�X��$H�U1� 9��!6/�²<�8o5���m��Z*n�"�f�W����l/z�����=27��Ua�MR�ly'��j?�2Ol}.kf��1��|��K�C�Gv��%YT1�h�x�@$Ϛ��DF@t�)DF�Mcʈ:���/Ph	QqP��,uv}�8���I �����P��a�G����
�T^z���:#9>���E&])�/��E��V�(�1:��O^cP�����+���Y��L9�����G�ιJc͌&掝��9�2_��ŭ�y�X~a�Okfio�{N��_�ykX��y���S,u�o�����0���i��Ċt8��dD�R�P���)�������7v�- ��ƑǗ��Y��9�8M��B[�"�Tx×�2D��ٶ�8q��j�X3�иݝ���B�d��;��T��s�әǠ�3���W2�"O��33���Y��<���Z�
͌Vf���ф�u�q�{v�s�=���,zw��M2U���h[Zks�]��#]�!(�|��%�D h������: ﮟ'o�+��� �c&Qz��hx�Cg��g֓�G6�=�ƶ�̧��w�C,�J	)�ؙ�1�~2�"�ru��p���R�$���3Ȅ^ƞ�c�ʿ�)ɳ�X'�&Ҽ/��ѯ*�5���݆[�UYG��ْݒ+��Jު�\G��݀|W�����L��wkR����۟�ƈc�B���暶�x4%�v����%��@Bjșq����iܯ3��ud�����џ�NcmK+�֔Y�����ƫNs��Gp>'��0���#Iն��{��pk\��E.82J��?�	��s��(&Ӄv7�u,���{c`9�=t��2�g.�n�>`�0�FP�!Yw6�I�u��]�(!��m�uu��o���RU~��۴;�C�1N<~����׆ĝ�v_���X�|򧳞e��[���}OS�����������O�-���Af�������|�O�f�����rz�0���� ||,�o��9���3A�?��%���h�t�!H�W��f�QT�P�m�W_{����#{9JE�ս�S�/�(��c�N,�em]�F�q6��W����!r�<�#��=Q��gv�M0;�m&}[��1p�(���^�n���`�HN�T�wtU/u�{ce5K����Y+�1v�v޻�OZ*���,2͏<����0��zS0A�CHB�[���f��W�-D�[�Y����2����;�"D�O�
7ECs&��������	�_�]�~c��qgU,g?�@5�s5>o,���T�(�ݞx�.�51���s�����7j?�~u���@������ZO��;�lhٻ�ξ7?�o�*pz���I	&���:3�Tu�������_MJe����;��=+�mU�F��݂@�bȐdc ��� ���<�}��)61y�=���+T��R������a�K�C���<��f������E���x:{g��o�'0��yJ5r.b�	e��3�@�@<�$��w�8Bǭ�R�Y)�� �=#��@K��l0�HE;+8�1&�4c�D(m�QV�1�C�=�L���穣��Z�M��!�ť���U	E�)y���c��i��/*�����C��ъ����'}����E�ݼV���ox�ч茸��uvj~��g� NU2^�\V�kr5�7��L�K�y�"��2��3�w�l����`�)AKs~b���v�ؽ��2A���a"���Ù��*P>�sO�rԊ�d��� d×��kA��i=�:�+���.���E_��B�d�`�������*,�(n��4%�3�ۘ�i�_�,uf0cn������:5x1h[�S��Djn��5]U#?���-5�|Y��������ȩɖ���v���V�Դ#�3�-̦��X)Jmg��H}hY˥���*�F�r�����w�u��D�|�'�,��.؉��Mq�(�V"�U������>�����ɣ$�0��S���Q�m��\7���-��l}��VD��_4mڻ:��ry�KWh�Qk�n�Q�����'LW���f�v��L9�%D��}�ۖ-�塜
�uE��|��Ĵ�q�A���A�[�j}�����6�u�Nh_^<汤jj+��a�-��5�j���A$�p��z^ml��e(/���NUh�Ic>$T��YMo�}]�ӏ/P.�{�+��b�4����١��Ri��W������ޡ���,�A��'{��iU�z$�=�i�G�M;���8cҠ;��4Q����d5�}z�t��˽��L�A<��j=�q��O{nj�
ʰ���}ص����Q%�{�m�0�6܇�U�m(CH${_!�����,���9���>�<�����J�NDB�~�ZLU�������8���j<g�M�YM���v�\2`D����6j��1U�vҕ�)��}�~��+�`N?jb�17�88�Z�l��8����G��!(����yj�Ve2+ 1 ���%�G��9��y�>䟾���⸺׺5+����me�y ����ϗx�Rn�~�S�	�M�9�_x8���J}��Q���+엊��nP��BXH�1���D��
�	Ҽ:'���Ԃ�qIx��v��xLk�g�Ct4���r�|�� �	�}�P|y�I�{�c�@�L��I�.�9<2�K�ɾs�eY�9����ā��a����'�v���#l�1=�Y�e��d3'wN<�k)?�sё�t2���|\;E�+��u�#6�]y�G�
`�k �����%°X���{�,ϴ����"TA�A�����u��<���ĥ�"gN�YXe娗��
�W?�mfXP�LD/�nP��q`ADe���}0��1�����6�Ā�_E�⩓�P�6�10x�pfE��u:#�8�U)���� ���T��}�tZ^i�#a;�(�E6����˺;�oB;]��DH���_��.��C@`�F��L�I�3A��ҋ���L�}5>��̓�S7���h��<�ZuF�+]��?s�w[�ꪣ� �Q٩[�������O�O�wQ�1=��)�����w�\#/1�z���ʷ$���ۉ��7�
T�6�4Ӭ�JO�f��6_�����w�͊�"��
�g�GDwK0�9{w�=))/W(-��i��l5�|��e��M$ͅ�����{�m�h���_��/�D����X0+謹Ó�'��Ec�fX7Ċ��D;�> ��ϡ�z#XM��4�"l�G�z�A:��>5��L�cf���d���pxG�BA��Sk? K�^/3xJ&�`!��?�_-��-;7	�����@�K-�4 ��%�jC�E�P�lnhts~!Νs�$���%�<�������S)(��z1Zar�p�v23� U#�X���Fr!h��;�Тϴ�i5��{)��N�s+��M珩��þft�>������ѭ+*���	�i�p.<��
��<*znN���=9���5�ׁ
�vN�@=�f�T�%����V�����.N�ƹ޿�p9;�6Q9;3���m���͔�t�?A<8�L����J��I}�� ��UZ5k]�E:D�Q��s���o���:�Þ�T%6�ʏj��W��B�O5a�l�]�������j����,��h��f�>���T�*���h�s;j_���R;ڔ²̄�mp�`��՝���|����O�/�!����dŤ��B$O��'����F���Iк������"�M}۵�k������)xi���^5���!t�%�BC��j%VI��l�1"ك��TJfU��&4V��s�|�.�4ƍ����^�e+.2��E�.-���j�P{����G.�]�
����p���EQ���w���(U�c$��4��M�h��+���?��Wt�'z��`�z�ttir��Tn�P�S��DQҶlTۆ#�t�LX)������R��"��j��)(}$X?{�\֛P]bSˉb6�ҒQy˄�� �Yc�yО�0|��C�(S���XO�0Y5�MX7��k*oskh��+�����S�
��f�RC�;2�v:��J'K�#�����q� ������s���N�S�ې��<��σ�� �W�w���9DMt��	8�1�H� A�%!��_94 vq�1f��TSu�)��摣yP-��U�FvI��&�_R�B����p����
��g+O�c_{��s9����a�Z�ݧ���W'lw�KP��X�b��!G���R�0���B {���2�n�V�A��d�.��'�?]e{�&��H�#�6;f�a>��
<dKS�Eq$Ղ�5i���;��\<���$�aS���s�	1A�z'���V.V������}�}�75�G�]E�Y����$:Ch�����s��N�_�s�B� �L�+D���x��j��7P�	{g������+�g��(��ݿ��M�k��:~�Y�����(0E1�#'ꚡs���GT����S���֡$d�eԘf7�A�}|J['8�{��������@���u�Bn�X��1
M�����&v��e����f�`i�0v����CE]h�nf�v��q]��n`���g͇ ��p�ˊi�T���b�������=c��J�$�m	��^^a���=�X7.z=㲿����S�<R���x^����	��2I>��K�4!I}�
˧�t�u����5�H�K���a�M*q������Izz��ɔo࿍��,Ǚb9Sf�Z$�+��I�w��d�%�TT��,}hU/=UL+��+z*S����hţr��:[�B���j��O���jB��%�|̌���E,�a�e��iq���.K٣V�z��I��Mp��U|��"�)\�pZ5�yB�h7y?��w�7͘[����yƋ?�lN��-�������d;/�9�a��Me�#��M�^�U���n�.ǋ��QYj��jJ������y%�i�BA�����j��A�Ї���V��0,6�p�c���,!����i'J@'�m��"����LA�T�KҤ2�
�=U�J-p�N�1s���UJJQ7,��G�~��y9.s�嵓qZ���0wg���|��r���,B��.��}\�����[Kp�]��.���>JZ�NOn��)�{��e\�ߔ����%m%�̿���dV1��xv�܅Z�,�ȇ7�Ny���ڰF�hz�_%�HL��܂0T�RՏ��k��̲�]�&������%��md�k�B?�*��J�Կ�w��S�H�M����N�A%fvz�e���/z�K�JY>����P�^�v��/�Y�ƶ��
n��nC ,w���~��/nUe�B`0=�Y�B8TO�� ׫*�h���&���O�{�i�*��̃��
@�C��TJc������"e�r��͌v_7�IvҰ����]�8rd�F��(��撽� Q���)�7�s���f]@I�S׺r1s�U�in���z�mÃ永���84'"��^�����|���(�����8���t��_d��{�{��.Jf	�}�-tIۗ����=�P��T;�hō��s���u���[p�����L��Q��7x�|2G�?¡��Y@��wB��_�}�K�HkR�D� �jz쿁x̿�P��i��O�����e{�j��0�ʤab/��|��?t�	_��득���]�Nt�1�t�7�7�:����\��bSg{�~!|S��CL�=�!�e�� CD�o3��f�.��9{��5���/�S@n���bm7jlB 7�B|����a��>0jC%0�|�b_�D��lp(�;y��tG���:�ܽg������p@���Q7���Zn	� �"�Ws���3��=L�ϫM�"g%���_�`l��2F��$�moQ'�+ԩHB���R=l"����%/>���0ᣵ�����`�m=�T��}\	��o!Yh��\50Qi0`�$�mB��ܾ�P���] �/���e���� ����}5=X/%���l����m/}��>Q��`|�r���3Ktq�R��
�a�>�M�-�K���`_��1���Z2MuFT�o�$�+����ސo,���J��K (#��m�h��C�`���D0<�v��W����s��m���o��"���w�.5E��g���.M��L<�JŮ�88OhՂ�M�^%�7|:�#,�`��3�p����B� ]W���ޮ����t��d@U��E�ٜ�+�R��V?[j��\�e�z�~�ܩ�����?���i�ʚc8�v�r~�h��K�$�pn���Q�mhq��7MgK��BgϣP�N̉�e��߷�Q�i("K�\�h��F�����=MDd��|�}�)�3ϗ,R�&�c󋵕k�f{��i^����q~q�Q;�o�n�\`T��x1��'R-�V�TR&~ض7�4�A2�x��F��,�1AH��TO���:v��]�!�n��N��F���p��!�F6N�IS�����]�W0��z1@�<�`"@9H�5���͜ �ҏČ�Z��������B���(B��{����Pvu�C������P��M�Z!��BSZ[X��Q1����Wp��:�vz�mR��0�|��PPܑ���-M��<ܲs~��f� �--��t�U�O�h*QJ�LM
�{D�~��e��޺�7S꽗���*���f��0��^��D��|�p��T@h78���q�9����;�h��e�Amo۫|���UI�}��G(��q�0i�h�AO�@�8��}�r�Nf���hrqM_�p���ߊ�ۋNo*A�q�#�E��C4��%̃S���<��|���[��Jt�-�k�:+'^L-�Q�t�� ��Yh���x)��E�����d�n{:8��-�����n����K�!6{GͶ�a�Yw�Ӎ��]��jBg��p0�,����rH�� �*X�����E"���>l�õ���-�b�xBIoS�^���{�t���i�`��)����˥P��ڔ;�v�F{�t���A'H��U(S��9:��2�+�3p��x4:���ʸF�Hr}�;J\w.�J�/��-���@��Q<4����|�����֋P���'9з����
�G���\<��?����$g��Gg�3�#($M�<�9�������Bva������]e_} �$͵>S�
�������HG>��V
���qI�6O�FAG`<m�S�ڻև�@�/�f�Ӵ�F��aCn������UQ�L���(-�ݹ�|k�yDp�Tv3^��<���s�gv��:�ߣ�Bz���KE��$ekػ��-�Z���L%!m��rU�R�aA,��2&ΊD�[ݚ��[��m\^�������$��r|M�ؿչV�@�����m��֘P����A������t�1�i�<��?Db��L.e��Γ܇1*Lo��M�4v�G0�o1�Q�┛h@��f�_�"���B�(QRu\V��!�T���Xc<st�컍ndaׂ"Q�|
��t^o[���$��츿��]-�
H��y��N/S��cɚ4a�tk�]q�]��,63��2ȿ�,.�Ʉ��\��Ey�f�ۓ
��\�>�W�y�"�?�Y"4p��˙�-�����0��ѩĈݺ�q�n��oML�6. ������pf�����QPD�@ʾl�0��x��L��::�,��VZ�Y9j^.z\h�S�򱰹u�;b��?ņ�|P�c�3��?����nu
z�n�=�G��ec*h���*uޤA�I{ٻ�c���2e_�,[��n�/�nG}��,����;��5�y�6��%�Z��xf����!LN:f���*x���ӆn� N���Y��aM���s��!d^��ły�c�;����e�'�lx��m$�.������˄�8	�N��	ڃ��1���n�eN�'⤨W�ԁ,���z;�'�LCoZ���o�ü����&��*>n��4��/#�
�r�֊�����aw^���].49J�Q����Ulܦ��%_�
A�kq����`��qK��K�m�b�yQ�o�Ј��ش�-b�#D�hT�,XƲz�e�8-Y��6;��@�T!��40�5��|m��g٨`����fD��ތ$%�P�l��Vې���7�R�Ws�K�E✹� `({�����#�KI�\t;�4l�"ݕ6�ʁ��X�?>Be;D��� ���hGi^x��"�zJ��1��G�VNj�"]�U�HV�����iv��w����7�@j�Pپr�^��.�pa�3�{����x�L�=iUwD�H����(ݥ����n���~z�*?�H������s/���>��Y����N~V�5�ݐ(t��衷ķ ��@ vb�:f�5�`\t*&C[Zu�F׉���K�I{�?(��[1�K�l2ޔ�e�O����@��ë�Zv��V���\7������Z�W�W�j��i�|[CZ�Le"�>z~c-� ����L�'<
���B�Ì{�ǜ���b7
��Bh���p�MS\F �zcb`����Θ�xc�>�1���J�G�jǲ?�	���z \ t�з2l�`-���o�,�w1��0��9F�j8�L�]�r2L֓7���'"t�F�{׃�)���I�Cw�/2�v81��k ������ N��l����3`9~G�q�в ��U�d��4Ó�f;���+@�1�\��T�̒QP���ЎXq�P�h6�w�3�=�2܂�+!=�$Fѹj��$����ƴ��C��>�[vG>}�v�HK!ޛBIM����A&���R�hd��4Q(�&��n�lO���B��<p3��� 6��iB!�1��?�D�\�]p���m���c�D�����KR�]}��w��2�t�c>5��*qE���\3��6����f��&[�l<��2���w��K!9X���a�Q&I~�t��|�EZ�-A=3����y1�AAj���B��kl�:��Ʊ�>������h+�G�}�O�ᄆ��8��?'���4�EJG���f&KJ}�5����҄,�</n�?A`85��c���a1*'OW��Q�D���H�