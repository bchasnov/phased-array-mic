��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|n�\&���Nh��pAbi��k2���]R���5>`�a/.GsbX*�h��uٝpMb����NADd���!�~y^��17_u�a�ʫ�$å���PF�?�髱usX�����~�/;x�@e���'�&j��f&#!Փ��<����yY��Q=�r����f:��^�SKO����28��;LWV�ACӽ�0�%_��tNN���!�2�?K���=���*�u�h��E���� �%�M���-��a�:h���J�cQ�Ѩ�<|��y=��r4*<]K�\0!!ZCK����S�+�E��q�
��� �UjA��eL��Q
aH�����@fL^��6�3�9˲
ޥq�=��܆*��q�Nʥ�XA�{�i�z��t�[s��j��*�P�����U;%K���1���	c���������w	&���Φ>�b�	�f��r�\������a��D'�3ޔ�mnX�c��
@.������ ����lM�� ��)V� �Ԟ�o3f��B�S�����,��$>��E���`���C��\�)M_�����K����%��R�Je1�u�2���EpD�F#�*��Q��-��ߘg�%��8y�7a�#��!�%���~M�Wq�d8�um3����X_�v�n��	�^�h����	c���3�z�P��W>|��)����^�[>�eO3Y8
��J�"�G:2��d��X�F��.���ƛ�!�z�_�l��{�W&���y�WF��\��i���@I!��=-�l��tk~C�\�]�x_>��k�����5�zG�"���F�ߣ7$�o}(M#5�k鼤�Y8��JeE������:Τ��UCR�� w��geO>�إF�d�/l�'�N����
��+�f� �~7ᇝ�;_ޠظ:��*��*��"<K
N����"���60������l�������EC][�I/B��6����w�X�ev^ø8��&6�PI�poQ��R���w����*�q�d������R�5c�����}��M�.�Lp=�������������l�˻>�t<����+K�����&C�8
>����Z��ԣ��x�R5�;ưx��;����n�;�n�ЙA�i|OzN�H�G��.ݫs��z��������Vm��G��,�ω�R��G�w�������/��ҵ�����E���1�\ޥ�'��0V�zN�J�T�b�3�)){�2+�z�i"d�s��)`!eYS �gc�D��bkW�v`�|ʡ������wH�!�GSL:]5�vO6�.?�y�V���{�͞V�������-�ޛ�&�W�s�����qoW\/�%bѭ8P..�5�M%��A��5��A���xa��6I�����_��T䤯�I��-N��<WTY�8e���7dg�X���n�^O��&Z���n��ۚ�����Ҹ͌XT�H8��7������|��즼|ǂ������P���GI	����q�jL��d-aS}1�01+���m�ߴ���|I�B�i�_ᎏ�&#{{�3 ����2�v�(������k��`D9��O.�g�+��l����k��\N$��B�r�L ������v�*�@&��w9�FH���"22��#�A�ߒ����}�,�@��^��W�ƀ��r���ކ���d����h�5OFgk��K��=!Z���^Ӥ�o�'e�_?<�ȍk*��|�����n��=�bW�A�Q�x��r��G�|��B>c��|�A�����=@����|�J.�l��C_��2c��o�q��!m���]����S'�P.
��������J�Ձ�S�>]���S����pTa��#`�Y:aP��:��ؐ��w��]9�5K�u�-�u�	>�5�h���@;�j��8����o �<0v��S,�G�?�F�� gtLd`+�1Rݥ�m�kBd3���е!Ycvk^'�3"J���2��/�X����K�`\���qJ=S�&4|�y�=�ךW�.R5�wqI�od/�+	�a�+li�`�is\�\� �p�bKK�x��'?��{����ը�]����81:��M�Xh�3��������:	�ak�H"��t�DÑ���+��5Ÿ-�?�cQY�0�w�� ��@�^J-N���b?��]1�5p��Mc�f�x��)g���wO�K��[��������)�+�����lV���E�|A�Z�-�dM<)�d�m�XI�0`�7���C�5N-bFh�"T&�+�>�������fМ��� �ٔ�"�6 CmT�e��.���W>�X}tH��	��]�V�q �X��z��J�@�B���0��F�ό����Q(ŵ�vٓ�HX`�5��tw�G:��gO)��sv����G��Дh������9�V/��1��u?MY%%����&��X㏌�������4G���_�uY�%.u�V��^�<�QZ7G����r�"� �Z�"�����|�ހ8����.5^���H����_�q�Ҙ��0-Lz�N��qއ���|�$c_�ȣ���%«\�Ϫ�r����:ύ"�U�d��ew9"L�4̇���zYۜX�Ү�f&1�c���.�l�p�',�jJ��R5=b�y4��6(w�N�'�yⲗ����2�2��yQ����ea����!)�+(�6����Ȉv%hӥTu�'B?Z[Dl�5[L� iUE��_Em��uΈ�kf� �X|�����M�o	��򺅈��5���P�?x�L�HC7�ec҄�;��?0	�O��X!孟��=˂�h��;�@��Z}�IZ�:�^���NZ{^�A���:�F�z�B6��3B�����ɋ1"D�����܀s񮇎���z:�&��_$����DX�,��f9R��n��G+�C�g�t�ʧ��1(z1�u�}�3�vF�rS	��D/�D�/�x�����ͣI�1��J�������=߄ �e�&i�Iy��}۬R�+��Z�k�4�p����h����$�z�U�Y���2h��Si�!2[p���\C��Yu�gY RUOY&ڱ��ܿ� 4����pl9K�P��>�����T@$iu�z���V8{[fҘ��UiLl
/�䋴?��#��(d��g$������q���}�ɟg�9_TC˻N������n0���Gm䳢�#k$��t"��?ê�-Y�k�G_����K݇e�ֹv�a9��e��@1��"�\�g��4�*�[�F��)�amk�Ah%v���9�ȬT��B��	=.8���n���G]<ֽ�'uy���h�<���2�G�%��LR��,��ۮ9�*"��dlxztYv��%�}�2��Ғ:f�{�3��L����o�Xc��>d2On�*b�7��E�A����OX��e���p��J8��$'e�7A9n���J��F�a������3�wC���j_����ے q���+�x��0#���Q�z�0R#�I�@�p���Q"Bf��Q�rrB�s�N�Y��K*��ɧ�O�i��."������/4}j��*Ϩ��.��_�Hni`!�B8:kK�C�T���8~l�?���QTh�G����_ؘPK�qS�M�Q>*d^I�	g�o������(�t_Y�p27Y���K�n�˵��/��57�X����C��B��q�\V��"PtB��Y��_0�=LRkG�4��B�?#�?�>v�1�w�~�wh�qĝ�n/�%5Ն*���W���/dT�/_-i�E��DK�n�O�0sj9�8���0�k߮q�gS��B�j�K��Vi�afV���`W+I�_�����"�F��Q�wz���{c��?���PC|�	�j�e���޸��Nwv$��r��\�[��髷^��W��^5-�P����>�`;��}
���HǇEq������K����
��T @�)~�Қ��g��s�K	�P~�i���ɳ��)L}��[t���y��h:���.�"�jI&��n�>l�|��L�p�=l�}�%yV#��"b�JK�z|�j����Q^7!w��#�ř�#g�0%��$��{%~�(5��J��*Ι��ʪ%�5�d�M�7^�_ៜu��1���Z�|�b�G�bkD��A����& _f���N�.��+ߝE{��H��� ��~su?�L��=47��}C�`�X5:{Q����.��~�*l�}�fv�O�L����򃙘����a��O_- lȊ�f41P^�Q��54�aB�Wĕi��~d�6���lL�~}=��QU�j����[V����{3raj��xc;�#���	�h'�����;ӰNR�=K�����dxL�x�o�0�ռ�c6j���9*�0��l	���_�j-���p_������z<���)h�z��6Ԫ�4�Hy��hc���ܓ�g���F�X@0���]���۳��ŋ'����8��]��T�A��4Ym(̓��4��f�h;�����1�j�J�E��:�"T3:|��;�	ޥ�,ᶣ�#�|���ЩV�d�z]br|�`������a�����9�'A&��O�e	Z9��{��� �Nr�Gr�����"i� ���[|��+X ���V���l�T_�[���j�9l���80��F-�ln�Cp!059� ʻ��*!Q�=�b��,��q4	xz;�>q!�8˱��w�J)[�k�h�3ؚ}}�ϡ�u�JɌSj�2C���m|,^��Mm̱l �)�?�6b�L+����<`���4ɏ9�֥υM��ŗ),���SX�?�j�D`�_֟jn�"4��2����[�޶�~�s�Z���xg�@��)��٠��Rq ˾��i��	���	�Z��-�ߍ�Z�����v[A�s�� S���*��7��h�d�L#	9�f4g/���H[$NŁ?��VB���U&��C���n���H ��?����A{N&�� H?	�r	S���>���vg�2�����*�L���i�\�$ڏ�n���Q���Œ��C������?�$t�~��@VWR~rkך:�n��SM[�|`	
��eK�n���U�@M����X�4�����܅�7�<�ךD�5���[k���*���L����Y)Q������^��H�&��G��RUЧ��ǹ��'z�ܷZ�|�}��B�<��+a� vHv�a�$��e�%ywhtQ����n�$��x�1k��=�����SLk���+���ez�����[���P�ܑ�7���GO�>��z��X�
g�V9cU
UU��B�:5���t2�4��Q��z��*@�o�~��x����f؅��������=jQ��^����`�j�����dX�x�(µ�ճC�r'�.�S}�t���:�+�{-�+���9�K�b*v+q�<�fFѫ98o��1�+PC��0�B�؋���>��p��v��Z_� V�^��ep�'�	𔌤_	����2�D�m>BRW���;5/��y;�[ڷa]+G��_����6��v��N����\4UTa�_�Ӂ�"�2�pFuX�@o�_�.}�sJ���&����)D�uiw�E;�D%H������>�h4<	����x�_r��6m<[�}�/n�0��8tv��dF���j��`f�
��%�'U������5�Zq����R�+��D��.6v�_���}*^�N*r��A(
~�/k|�$�^Aҏ�[6Z���Q��|e�:-�mC�zJ+j��2��pU.�2d�FE�olG��9�ޘ���*�Çn��1gs����^Zsry=*�)0�a�i��h�뮒P�*�� Rh��,����w����Ĺ�;+�hx���[�����҈���ݗ�d���5+��g��#�v�~�.8��=Q��|��#~y�վ�����;�~�ڔ�~*�<�?���b?��F��q�n�R�d�M�ܥ�,�S6��� �F0�(�`< �"'�:��e��vw���6�p�9X�Q6�4�w���U�Y⤉���}�1W��uQ¶�D���*!�X^+����P^��+�Ѭa��D�j����`Fl�Fe�MG<�U:� �$�W��.~�����Z^��5SVK������rpm\��=��(�Z�mH3KS��`�:i�U�L8��!4y�	���� �44橙����{/�Ҙ�*L�񝄝��k�Ⱥy��|g��1���m�����̝�殀�^�)3�̅��(��[����!x�l�Y+�F�gR��z�����S�W�����E��.�6���ɽ9�BS+��>����T�Bػ؆��d���h0:����4X�U��2�y���e�u�h#meH�y�Z�UyU�0R��i<`aY4r��K{(�Q�T���#e��]SK�٫MZo[4�yt�	�}����e��7ߙ�����h�nw���l���ܐȫ.49�U��aUB�].F��V%�W�����C��:Z���%�ǲ�=�5�1�g�����ڒ���A�@Q�}�u݅ƑU�7�,��|��pVI�2�St�������خ����i��Ser#	)v�G���ü�m�)	?:���)���rSa� �����H�'�z)�9��4�Ȭb�6���0?#���~�O����z���*��/a\�$�w�-l���e��r4�8�C���m�� �Ť�L�[ʆcrh
���!�J�+�嵩��e>Ja�ӷt����f~A�i���H�C\m)���y^���߱�񻕌�{�������s.�H���4�`�w������֪2r:�GL!���U!k���f�a�cm�p���G����@���������P������ o���~���x�W��$��)#��+��9�B����3��>���y�0-����I�����v�i\��C+7�W�R��n�"�U=�ݙbC�)(��e�at�q�������C?X(�
k��4o.t��(��jq���N^�Y�z�[N�ƲO���+���UKY|�;����=�x�b���B�����&���^�����Q�����k���i�h�1Gy2T�/ߛL��Y�V�@�P��k=�u	[����{w���2hm�+��JGA�oy#�Ǵ��0�xx�ث�~f@"����ʎ��:^.B�0>-��̗^S2��h"Sy�}�e�<��x�u�� n�X��C����Kù�ʓ�)*oe��n�jV��)股��)��y�h��O(I�����u����3Ə`@�$Ň}�����K�TgɊ�K������YL��S
P����z���5X+�[�KV��@|4��-��um�I@�q7ж�kIrg�}V���u�C6N!�N���5�!�0'y^/�3/�7r�&��F�B�=(��6�1�m���5�QH���n�{�%��HhgK ���"{Q���%u^V�mN��j���$��^��q���_�09�j�Y�M��v�I�bXg�!cy�ܲ��f�d��J$& �~u��7خ*eH��i�s�L�)l�r�������O�L�G*�d�WA�aM��j�Ջn��vF�kM�
�]8п��d�6D�$���.ǡ^?��|B���R��=���Js��I�h��j�菐�wN	�?S�ߝOb���bK0� ���3��Bn�m$��U���W�J�t��[��&���hk�,=�٬)B:�a�O���`G,�,Og�#���/��>3m�����S��OJ�����1��*�Kl�B��N_��J8�X�P����!'n�F�#�|p�|# (Rx������fzU��L<�2�:+�>��͑~�, ���Og�
�R�]�9����Q%r�Ǒ=�e�0+Z��	�fq��8�7/�hw�/��z�d����*��\Nܴ�7%�ۅ�n�rcބ�%m������'�GH�Qt�[���v�.���Q���Ih��sАz�!Ғ�ހx�N`�B.�ʜH�x`w��6Ec/��v����J1uQ:�Sy�2g�Z�㷦Q��wM�^�� ����}fE����mC�Q�������i�r؛o�z�m�r�¢O�G��@��ƥ]�H״N�B�Pǵ�MX���]{������"���
00Û�����>鄖jb�m����Z^ѧ	�u�xa �*G�w�%�LGޑC���z`���a�U¼_��w#��j��3�@bW�{D�]�6"�;K�ݏ.#.v�+B(ta�⠋Ƣ��$����䤳LE�K���.���U�����M��`�jC�n�@����?���-�X��AgS�ɛWo��,���| �1��mZ�Iꋬ�1Rϛ>_�O��-U�1��_gF�P��f�B͡EP�^l����t�BhZ�z�0 �L��@��+�����L�hr���`�� I���K~B��>G�L�?:-W���at�B��&���Zc5�}�
|����yy�)j�zrYT=�=c�ƃ�&�[�l2��){��a!Ơ��Ew���9z#r����m�q+��שg�Ҭ�$�[1!4��� �*����3�O���\�
B� �pK�H�~��(����$K�V�[Lu�C�Ţg�b~N�8�=}9=����&Y�Ѩ�V\���V�1N��4�ڍcU��ܬ��~$K0�Mc�5/�s�.C��sw��g��v�G��#��=�8�e��$�7������e��e,�*�����u��s�9��{�(М�.o\���5j�r"l�I/_�?�`��c�k�IB>��a&��1�E�����(ٌ�mS� /H�$��G���}p���5�rv�C�!rp�׏j�Nˬ�8�cM�}{��G��ܚ�<�Vj��^�Y2z��)��;!��o~K�_7'���^Tw��@1ȿ��|	�N�	�o����`�~��~1\_CGz#R��C\�����y���l�XM����Snb'��m�
(}��&odY��,) ����;�"魦}�;�<x����)���/�T�y���p�E0l�;�H��Ǣ��}G�(&8 aA�m?=A՝%R3"e������62C�:y~6C�i;VDJɢ�A���z*��ݏ�����܈Ra�
)��y����U��S�u�$�G!����|ɟY��`�S�d����Ϲ@��#��?{&_�r�cN�����oW�v��xI��KW����)�o�s��5�e�h���w����}˛�*W&�/�M���D�ꇐ�:������M�����@���ht��n`/�ݚ�72ı�ق�ۻ2@�g���g�3
���I��R�I�M�&�%RL^I`aBr��K��|H��8�R~��I�>�JFi���<�r8�0F����S}a�?�Z���U�R��e��ȣ��-���\ʻCi����U��4n���yP�)�G�)�<�z�����#��]Db��Ӽ�'��pd?.� *��ma�.S�&P��Z����B�������*�,xV��7����� ƃ�7�6i
�1��;�>f�cf�ay`,9Qv%������;��\�$��z��VF�@;�SA�����?~�C�����3oj���.<����2���-��ΰc�Э��^�˸5�I��>�0��5��:6f��^��!D��B)�8�_�	�e����g�9q>�D8vI���(z}L��w�Ğ} �7M
)���Stc��y��'pxh#,59r��yU���Xۗ����V�y{v�$4��D���裉m�����f�;e퓎�	����5k�񷇰��<10�?�M
 �+�f"�`�f��3�d4a��0:����,�/�d`�u�LcKt��F?�_8n[�>m��K����΃ N=��u ��3�G�A��b=y����Mb^��h����x(����Wg����瀎 y��,M�[��ħ�V4�)�Zʕ�$�tbz�L��] d�8���_'jkL;�y^� �l�C�Р���*M(D]�J�R����֡��8h��������Q����:ц�M:)	?��^����O�%"**f%l�ղ��Eɸ��h�YC��͛5@�lrR��\7�!?r�ґAܽ2p�H���Pg8HvF�2��s����_���J�3~�b8�� �I�:JY�h>q�T&��mi�����o?����u�5���O7������æ�c�G5&��O��v �2�?bJH�wr�W�H��+���7YAo�m�^���P�2$]�hc}�r������B�\�����ʰ��$vD�Q�,<i�>K�5W�!bw�DN62N��`��db�0�3�H�Ѻ� ��?����ݨnL]�2ɕx��-ɔiMb'v49�Wv#���As&i`b��*K:�1~���|E5$J)�ĩ�p%���{����Ny��pSrˠ��C��=��]���,��_�^u	�9�ː�9��@4P4O<Db�J�k>ІY@��@u�"�`� ����ճ��AL��%IR5ݠ�Ne�� ���1���Y"p��[���N���.��R`)����ԟ�C�-c@�`Ɵd%�^u�9j�V����OM���u�M�f+��F���/|P�V3�$G�J!+��.�c��hf����n��r�F��$#�KK�����:�M|R\��Z@ �:��L>����Tev�� ��,�������74����6���hO�+>� ��z6�g�y_5H��_��2����6�l�t��"�ҥ̽ ��ݿ�B�@�;��QG�r�aj˾~�k�NFn���sf���)p��N�0i����L65�6����I
��Ll�Ӿ񧺓m~7g9P�9�̩�8x�J�y���,��F��5D�u��� ��V[:���6e���#�SჄ:���$@�7G!C�VL�pJ��׊C�J���f��k*�u-g	f�3e�|�00���;=>���O�h|��OB�#�����W�/�r/�NA���=��*Ȟ��~$�FJ���^�"w�h�,�@#��K�ħkp�ș��n��W�us�m8ڮGn#���	�G�s�Bӡ��{!S-`	3�lGU���F�(�t%�lW���*�
=N���z���� L��H3��i���%
`��y ğ4�q�x,�5�'{]O�m�*�ہ��#v��ޚ���7��ߴ�����(r����XV�0����yf��N(_���[�R&v��o�^H8���L��1]��� �|p 9��9��zQoP�(o!ɭT+}��\��3h�B�2�rg�"$��|���r,�9.EX:a�9~��%��X8�V>�摣�����ŭ^�V�fAjn债������FR6:q��,X#��T;�_N��?��.0��RLֹ�g:���%�$�P�=�i�s:��P�Ȭd/��x������"s�b/`r#aT ;�8�{�R0�@ܝ���i�����o���'bY�D�MGw� !�c��z�56V(���M8HC���/v�MQ��[��7λ��`!���ƶ��^���P�P��@�2ƣ�)}0湳L��a���� ��T���x�vf<-�TD�'�n�����ճN@��� �<����բ�]���P)_&��J��20,�|��UE��A9\׵�[�'h5t�%�2�֮��};&�J�'��*zk��5��=�Uo���k��J�B����1��)��m[g:b���/�Y!����e��:��[~�������M��^F��kZ�nu%e�E��x�����_|��?Vko�TjJ'!���h��}�$�*1z�vQQ�6�*K�\Ɠ���z�K��2��JS0��K�.,'H�ܴ��H⢻ֵ3��3�:�����ubSC�N�GE��w�s
	�\��MK>��(�ps�+�+1*�ƕ��sU�����������{�5�ȫ_�Y(9��k�ciQn|cϏKz2��OM|p�ڻv/��kW�)�\��5o�'k�W�� %7S�%&��w�)o6\��ה��֖@X��	8k���6�ȵ$�lŢ:���P{��P3X��;�W��{���T��L��?1x�	���<3UXK��bOu�u�P4�Xu��ZO�ab���=�o]��)E	��k���me�~ڍ^�"��ԣ�d��g�"{9�ǎ�f�2�Z���.l_�����h�"�w�0�Xj��>&-�M�NU(d����[��ި6��Od�D��C�aGs��#�9�P�N6ֳ���ǎZ�\n�yDGU��8��@5��Q��x��N��m�v���6)[�Y
}t��ג��\�}c�G���yo}�J(@继�֦�a[����
C���Q�w�����lH��6���^�T�����Ҵ7>\�t�/�p��,�k�9_��(�IhDT܎٤���}b�0Y�.^�V��4?���b��h,�p��rS��:�o/�B���,�(��E���U+��[��)g��ۤ������.�^�ץ�4V^��,�	���}�8��P��[��9.��� �q?�K/�����<�O�&ʯ�����7]�i�N��ǝɕ�ͮ�NM�+�js����]*-1�q��K:�Q��)��ˈ�����ʊ*3�0�Lf�P�vs�D;jj�ɵ�G!_<�RB�=��CM�:�v�ޱrҚ�6Gn����q���o�@̬�$J{W})-�S����E��T�L��5\��h$ ���3����kJ�U)�����>�?_�y�����*}�]����S��җE�4H<��٠QO�����P�>�6��V�O��դ�h=�ٳ���ns�#�D��.��ܤX� ����ߤ����:�0SƑ������ L���Tk��4��OV�
߱�^3���oC,* AA�t߱�_��A�vbʮa�=\��w��w�xC~�<Y�ozC�H��;
�?H9b�k|�d�� �2�
���w��{\C���cx���\D��ĸ$�̙��J��p�zC�Ȥ���RrՍe���Q8�Rev6�x�dϦ��'G�-B��D��(�b�=��v�v��j����b@��<��� �#��ƫ���Sr~f��/�g��x���e%�l����l�xᙑ�������5>��fV�^s���@/�_D:)�חĂ06��J�R�t�)Ї�;��m�:�8y#�sW4.`�K��IH��c�J"%7�[��%�eu����&�"z=T�bBх&��P	�z�F2��M3��� �������x�`�-�$4�7T>��l�h�W��g���k�K��1")������'Xv�Q$%���*YL�j����+��9FDXQ���"g5���H��nY���v�n���L��]\ڸ ]��8gpp�a"���c{S
��y��"B_ȁ.�C��"_5�hz�!��蚙@�&E��N0L�U��x�G�VRdw���
�����7�F �[�\m�u'Y�����IW�s�v�%L��z���&�/��v|���Ew���i���鼱6�����o���q˓y:�Z�u��o���B2Bk�����$)[��\%jp�R]t���$��x&�H���>��T|���]VQ g%;H-;r�Oܠ�˰����lm�<�	".�q5e��M���5GN-c:��L-_��m����B�|������/�zŠ���ҭz��;�0V"�H��gA��A'��N�ۮ�~U�7T�TpdgZ	�靋�����ī�p#���N�yHm����e��k��_A~4p�����-3�io�����Lc�zi����YLf��ӆU��y��d��R-~��r�kf������s�!� �x�H���3�O�04\���i�a��b��+�� �a�#�C��r�c�n�3L#n���%q)����C�����0����7@��̂��(��;<��]lw,n�^C��T��o�n�
,c\+���l�AXOW�P��&���k��a(=ϐ����_Kn���c�b����L/�p!��-R�2�A���$����W�^Ar��g�Gu�7e۳ �E� Z�M�{��\/�����a���2�C'�c��(JZ
c�pv��&Q�CPhl�6��ට"�^�5�ҙ� ��f�o�T)�?���)��8C�YZ!����R�b���<� ���A�_�R�U�l\isת��d$:^mSh��諮�7�/ ��-s��8���Rz��2ea�������Q6�\嶲ʭ��a���:�Gŭ�뜸�P�O��6��1<T}�r�Թ5����0M�HP�Sߩ�b���)��H��1�K�lq���n�~Xm[2�H@3[�ݤ�ۉt�$���+�Ur]�@����H��R3��<����k�o$���N��z���X��D��������@T��"BQq�~O�>C��c�E��Ae� ���&����� ]�W�f5g-�|��j �́8��Y��{W�^��R���k���}���Y�.�6�qUwY_��G2X�9�]����]M�$�!t�pL�ÕJ�F �F����f�uܕ��)xg"7���Xd��J��HU��݃�P퐚k[p�n�i�[��}�b�S\ַ?K���Tzw֝(k����l<?}��-��߲X�݌���C9uZEϻ�Ċ&��X܄*��t,P;@W��5g`vèɬiA�ݲ����F��e�<��lo� �[q+DDD1c�W� 8��O�9����;mw�u��Zk�����=?��jⱽ�8$��'��[_���E�kL�����H.f�9FQ�@K-��������N�f'���]۪niG����� ;<ȸB�\P���(U���Ҕo�d�]5�b]f�~0���\�j��lr'��Np�pEZ��Q�~�	~U��[��֖=)���i?�ST�����Y8@��c� E�2�ɒWN��"0ӕ���8���u���ɘ�^��n�r�j&���r�H��S��es^�0�@�[2v���ǾbA�+s�4�� ��{�@dT��۷�Q�5���g��