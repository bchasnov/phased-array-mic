��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�k�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������"0F��}�h'��8��<���9���-�j����,W�_/�H: 2���x���CH�^�g�&{�}�$�����$�B��.}b��t��nI�cm'���M�F`˲������+����o�O�=�{�4�=@9�o7��RD���w���bk�F�}vl�dP�XoI�*�Q�kM'��, �������[`�em�d�%���M(Xb���.�y'���<��	١��,Hl� ���
އ/B��ފ��6��/P�I��G�'���ΦŸ�F�;2,��}ʁ*+��u�{�_�@[U�ɡ�>�?�f��T��vEG�'8R��S��h�#N8��El�7���O���bk׊�<�!z@���O���w�_oӻ�ذ�X�jgojI8╮� JqF��:O�b�!UL�P���d��J۹��?�뜄�:�n�jft��"�l��EL�E�E�b�c�;Dq���.�*Ѡ��d�==2�U5�l|�'��q�Up�_��(�	�j�o�~~�_	��#�P1�f�*S��,6��K����W���I|��<���<~�&΀��J���ؒ(�W�� W�Kyp��R�{C�܆�3ӎ"�|O��<�uz�[@g�8pN�@���`��AC�H`:��Gz��9o �-�m=]�D�0Op�nCaޔ,�1e�<~��!����(({(�Ϣp#��f�h�`� �����_D���KKs��%�L"��aخ̎iNi��~���9T��Rc�ϼJ<AN��E��^N*?)ё�,��ܒ��U�1��W�HL��r_����2$��Z�ˠ�'@tS��������s����/�hF��_~t��d!|'���\�}���y��32P��l[��~\i���Ų^�����W3���@� Rvs�Fe0���[u��:JXĪY^�OM/ �#�>���e�M%Jl7�p��]9�{�|���YJv��t�pQ�L�Wp��_�D#�NU�NJ!�|�����Ȉ$��A�?HR$xovI�)�q����1�?:X��~Pd� ĭ?Z���f;��Vo�py���Z����zh�����X�٦3_ј��~0�G	ѣ��03�	��a��Ѳj�$��K�E	_p���D%=�������8FE�����w2�,����O�j������,
�@�P'����5����f� ���N��]h\�4����+��]��m/�"Zc�n���81Vԭm��u�-��6M��M����o`���J.��[bxf��
mU�}�`tA�JJ֣�
Vˈd�"�x:�K��:��bN��;�DܾF|�<W�ɜ�Ѳ���^�-� ���1��bC>���9�������U��ۉ���L-X�FX�'����I+��G�++�hK���~�n�^�3kUc�?����5�r���x"��;���~�B���E!��ڼ7[U�%h���2�:���j�>z_��H�M�F��Zi�v�b�I����[�k�L ��*7�m�v��pL�3Tm�q.���/ya2Dw�lu�诋��m�)x�<��{�1�0x���L��+k���طH�|#��"�q�)���VF�˿������M	��x7}B�B�X,�A�*l��0
�������G��oe
�/���c���,���as�:s�r_ᔲ�%�s9?�SI)��hobҐ�J)�IT��︸ 4�5�Q���O��v5�|G/�h���[���T�^�u6�L~��G��l���K�H�y�1&"�~�˻�I�B�t�4�	��f��2i����������Ny���ح�/�������d��
�:��p�J}�m922O@�#(l\p̒�h�RJ��
?��䉽(*�;�q|I_̉�󼹦�G�c�ћ��Q�<Yn�Z�����-*mߌ��:�a�Ƌ(3f���!�pEQo¾��:c����#i���VQH�Qu�b�2�������5��nB$�����d�4� qx� �����\� �����ĉ��a��Ӵ�,J�\m�.�I4���$W��zSR<���[�|���й!+p�7�8)�*��)ӱ���^��cxq�K�4(.����j�~���w�iQ���!��6�7��MP�a2�zzI�A��R:�� �9���k�)�-s|B�������G�7�sc٭����-��0���>��Km��P2:��S*�b�$n���o0�C��,ߢ����[:ax��g��1|��iC�s �4���E�rU>�}({�ƴ.����J�,�9T�F�@�4
�.�\*���H�H+W��ċ�(KÀ���'S@���+��W ޲cyK'���%�Yg���2���	O|x��L�b^���?�;v�2ł���0ah;����\ޤjw�n�[�X^4rH]o9�n�#`zK3��nK�ʖ�Ɏ�G�Ʈb2+@������V�R��'>|��UN��
����̖L[g��2@�+7hzv[�#p:���k�V.��#�>��c�P���X⧷��@$_��c�?�����j�ؔ�����fOS�0ڭk`Q��y&�"Ԙ��Z�ܞ���N��yD�O-S~"u�6�i%o'��g=|\x/��%����X�03�K�7����Ma��s>쒢��JM�� S�Uu�>�-H�O�
p�֬�rq-w�I�,r�5l#�V�#4�bz�����ݗ5*G���r+��H,���6Q�
�#��������;Ň%�*?�p��n�Pz�M'2��*�x����'�ѿPd���mf�`�H��:�"�S�p�@�/j��b�W�vwr�P���������I�S�@��HO�2jτowọ� �Oɟ��NY&�OP�*���A-M����� _n��bL���H������L�q�IɎLBw�^��C�= ����vMY�0�N5B~�z�%9a�.��)�eT�Z+}\zO.S�.:�.ߘ�m�_l��C({�q���`B~{�&���{�;/p��򆔫��GUT%�u$h�i[c;�r�u��J����j4�T
^߷�������Ք+�������6���|�~#�~Y6k�+j��
���R��D]�d������6��r0��"�$k�.�y��v~���bH�V�V
��\I��]��R/��/�>3 ��¨��4��o�h�}
E�03�����
�v{�*�L5K��2S��Z��
����gk&�������|���ok}r�����Qv��l��=�x �$(�&~)��]u#3�|�o�n"��%���,^-i<U�H��s��!�]��Q�B��¼AL���)���ǝ�(�b^)�a�nK!�Z`@��h���1J}��"Rn�n�ݧfջ��_o���TP��~�1����SGuv�k�8�g3P��s�G�b$zA~ܒ��o�-��Ƥ�-Æ��u6��K`~Om,Q	J}�`.)r��x&d�<��*�_f�t���2��P��Da��������iΟ%�2���Ű�����'��II�����1�fIݡs���(r�ݴ�94��۔����ѷ�FnKOy.:��o��]�i;h5m�.���*��jMM�;���λV,�Lت���)�zT1�i��Ė�o�WHtnrk��9|S6�k��-���d��e#L�HZ`�D/Gԣ�e"�K���m�����5��P��9��q�i�6*����n(a�G[��Q�J�k��Mn�)��q2�aR�Z�㯉�&�ȡq��_�9� oqr�Z���J�K��1�eA����:��{�v�h�|޶!x_��}ʩ��0��pӟ`YV	Ѹ5� ����V��{�y� L�M���&O�_f��W/�^�����N���eT��P�qx_VF_�b�����`�vH��X�S:���W� %�L[��V]�DI�����B�9
9���24=4��Ae����b�}_��B}���Ó��K��l�^3�+��-�����@��KD�ڮ��*��	&�gE���&���/�'ZPF�������E�`ð&12�k�L��j�دF�:GZ-�q�O:�%yC��h�tm���+���*�#�{'��PR�f�����ں�;a���+�ذ�f������ܷ�.V���w���N��V��)~���㩽v���ㄍ_�c���Q)v�Y����x#��8%�ƻ���|�M;�
+=��C͓�T���7X����ɞn�ã($�^g�Ӛ,�Be���>i`�+)�a>�Ƞ8��80$K\��i+d[�K����"�
�S##,�����+l;|��?�0���Bc;�|������ �@�>� �4;�:���Bq 	��1����V�=�Ш��HG�%܂�Ѧ�<J<ܒ���(Jlʦ(#��"����T��]�78�Q�U��Ot�O}_�T٘��q������vrw������`և؅�~�˕�c�g���A��B�����U�U�Z���O?�e�RE*�	�d,�5�K=М_�a��mZ��B �v���`��Y���~�K��PƉ��W��F)*y/���?y{c� ��C��'HX���b�j�C�;�.~���� !��N�TE��+j��N���>G���|���xS�1\����}��4q����ںԣ�#z:Q��}��;��qGrhh$^\��*�Vk�_�ϛ_�B���I_e�5f�N#�=}�G���^<&�v� T[��5������{�ySt��?�0&�-q�W�/���B�W!��RhZ����^��\��5~�FD�HG�y  x���7� VU�&z��9b�����C�����p[NV�Z�l�E|����n��`-���A.{�Ýi#:t��&�#
W	fh�����{���8�n���n!��Ė}�K�̃�߈����_W]����-w��B'�ؘo�֮�僁�<�F	��W����~.{��P��h�bH2��/�Yn)���!	k{F��5*	ÿ5������g�[�z���d˛�B�k/��v��������vƋx�wn�v���1κ����1g�GN�Nn�i�=��:"@����E�c�dm`V�����T:ԯ�k�)�z:^�E�U�vҽ6:�J2g�k� ��j ��b�������'�`�r)ȑ��Q���fOr���W�Ԓb��Er^t5&�AD4���?:���vH�P8{J�xw��|'J6eL���VZ��]~�&X�XPq�>|�Q`Đg���w���WF�����ӣ��y�hM)������*M7��3�U���oq�9������E�A��a.+�w�%m AJu�җ���m�FYn��f@$���bX�\�������/���M(�{8�d�Rg�h��$W&m���Q&q���; ���8'b磥T��Nb�����u$[�/����n�!��N�]R�K�{�#����f�>s�/�W��P�{�jc����5���f�۽�0�ĭ��h$�q���]���q#��&�4��'*g��%eĠ%[�+�����9[ ?4HHh�@f?��>�@r൓"���"R@5,n��lp��qp���mm^h��=�_�/��F��C�A�����=��`��>��#�-��'��V��|=�<�l�"]��/U}@u��/�6��>E#2�f��S����c�{��h ��|N��Vߵ'q��Z^�sn;)M�'w G��)��&����䓍��D���?ſ�4����!M!+2�}�������8��x���`. 3��^�CD���mX�o](��T~$�T�S��A_Qȴ�Ut����	��U�	k� U:��bQK}�HI�^�"�����/�?@�Z� �Pޥ�=c�yX�6�F�Ahg�#�A�BZ�D*,F^�ff��-켷��)����������F�cx��8�%�d�zα�����;Lk�)����0K$�)�2R��P����O���	w����=�2��1�/��/��d,G����a���� �y���ƞP��P�*�][n3/��z�:o>�nB�k/;z���e����ꤰH���e�D�xl�Dg��U�64�כ�zrڄ���4�Kӭ����ѹ��F�9�h�hD;�g6�P�
�:d����d�T�v�G�O�����1�rU�XTD�>#��#f� �*K��$2���_���; �sˏ�M�_�X�x3���W-���."��G��!"�|�|��tă]m+-��9�~���Ig�[�)�>h��S�S���"�=�B�I~�M^�X�+�CU�'��CI�i(s�D/4T���~k��f�,�.+�0y�*�*�G�L��c���('S܁�Bg-�P�ֲ�/�B��I��}�7~Jnl�A.�'v ��A�5���`�]8Gt�JlҢ��|.-�N�"�&���맀�������0Rl�Ȭ���V�a}�R�� �ki�?$6Q!p��틪�Ό=h ]�8�46�V���LC*{��I$���[�X����l0_"��Pƣ��!�H@tO���y���`������\�62��Y�G$�,C݄�l�V�n��z>d��Z=e�nmh �ѧ}�A%/N��G���KQe�s"��d��1w�x�&�����A��;c�����df��g����~g��r���؂��{ǌ��o�-1�2��C]${��`�瞉�3��r{�(���/ߎq���K"5�t�v�D�%e����қKRE���Ҭ��M�G�I���1���m�|�
d�<.'h՝��^�lΦ@��E�^�B�+�)�}�Js�}17����������7"�L�m��Jx
�E�����.�c���fE�Z�<��q�����u)^���A�q#&���>m��4j� ����9�Z'��;[S'��Q��I��٭a�$-�L<�qtF��A��|_�S
�P�L}���r��y����N�>^�\�Lo'@��Y��:����@�@g�����^@)���i��xP�R����fA��/dU5��e���r�"��2I?� �EW{���Pxld�M�@�Ɔ�z���1�j߸����!������r�}=�߿�k"-����}Fρe(6a$a��Bv�&�%J=�t�}��q��G{x��%U�����lz`�¤�quL��_C��\=*ᄊ�\�`"xrT�e���
:���XL>�1���w��}Q+'h��n��<�D�`[�M�"dZ�[��U}��:��?{����ռ��Z_���)Ɣ#z�O�"5�eRk���'� .w!� ����C�C�/ߋ�?e���X�8]�7��v�#�0E���;Q����u��j��G*;�1��w��6ρMRƕ�~tr*2�-�L�#�,�f׍Z��_�'���/V�{�xX�ou�!�huu�Qm�Cъ-w�����e5��S!��c̐���(4����`�&ڑ�W�O���d�y� �5u���K/%���Mv��r�:	a~<�G��Gߞ� �F��Ŧ����.vU��³ ��*��)(�Uޓ��2�~4��G�4�|h��9�H�\?�P�c܎u&x�I$������ט��D,���q�Yna�D52vrj�S���c���Z܂W��6��9i��] ��?��ǂ�ҷ����w3�P��S��E���6�Z2�F��D�|�J�k�TF��\��� ���4�bu���vI���n�J�P��e�
kb垇��Ug�9�˓�CLǀ����i�5h�1�#��D�q�ľo���~�Z��t�ڶ���<���7y��q}Q��#���g�?;;y4i�<M��7�@�m=�
�K�đ����V�N�7�+7q5\@xנ4@�Y��EV�����.p��c�(�6g����l�S���w��I�;~�KZ;�v�'s�7덍()��8POS�Mp\����%)�k�m�3R�H�`�'W�|�a͇�1�I?f(�����jc)������P�8-3��iX���(���J��ˀ�>XE�ڌ��87,�XH�݋7.�������OVx� Da��Y��DB��Al�e�x��YY���G΀H�k�?�{-ީ{�Տ(��/$�u	Bh:���˭OF�2h�Ǳ#�pLe���3�O'�g�����[�|����^��@�Г���S�]�����F���v�N�����h�U{�HR,��E?�:��ZP�"24����{@_Y/L�Kڑp��)���'��b�w�I�L��]c�"rr<E�Ŋ�P���SH��R��$�/$��Ɩt�,l�K*�M��SkJj�?��v\�uõp���:{$>�hT>�-�/�Km@�h�!������C�\�����N`�ŧ��@�q�(T�aHE�ݘҽ'��{���,m�0߯��j��.[>�z�4�\�����4P\㰋#.5O9�l��ą�Z��O}�4��RWY�ʦ�!�[��7�yɚJ/�#-rTld�#Sp8*]Ϧ�wnU��%a�'�����J��x:F��c���#ȶt�C�vke˾(�,�Ԥ��K��P6���EuT� {�_�>Z��gs�|1L�� �D篰�S�q��2Z&�<S��N�E���c-�y��EY�'-JNy�мH���E�Ӫ,�	�&e��<t*D!ı�q���~�WG@C���D��u���x6�-.����ZmN�ݓ�=i'��B���gQ������HiY��	G��(��Ca�xD���?��(}�ڴ�_Q���%gv5A�� �%�G���7��~�1:B�*Wt�&�쏮���R'3aG�Lam�3�������~��j�E"Ys�����[뽵{�w{��1�u��P�Z�������~	VX��;R!N�#m�dƿ�m�� ��ݗ��\�,M!��H��O@�y�Ҫ(���BOzd��o���#xƥ��Ë��L�ȁA�d�f��U3��LnϟSޱY	�KZ0}|��h�.5ԙ���͝RYJ(-�@�,d�ڋC�`�J30��n�O �9�2a��MҀ:�_������%��z����N�^���:5v����dDP�����`��JԞBl�QY0 
�/9*euz�Ɏ;/����iָ1P]��ו�IB�"��z:p��'�!�u���ZN�g������L_\0s����&��N��a�-IezM;��C�Y�D��g�EIij��}��H�M��׏���)�~Hefˬ��}�V{�(��^p��r��{��Og �= ��=P,���2��e����������Lݎj��B\��p���q:嬉��W��Y���hyc��������ݦV�Mb6
%�t�T]�$U��5A�]"�OA�#�دs��_\ω�:���(���Wh��P�|'��ke�$W���b���gr���!�8��xn���yEGjI�Ǟ�8�p��O�2�e7���"_{�2¥�����-7U�3)o���}�W���LF��!9h��^������"��awmߒ��T�|��rG�M� %v晁��zRr�
��r�e�L�/c�0[ۊL�����8�wT��{?�[�r95 �� �>~��8���)�����/��x�����Bnb��PT`Dßl���~,Mt� '���X�.��Ku���l��ZmO!��I�a��}���9�o�ɦd��׭x$��m�i���R��A�A��$�Lʃxː[�����֮�`*#�־/�yݿ|���ه�R����؃�Z�����$�W�Hio�_�2��텀�ԩ	�4=k�7���0�p���'�&H{��:�������rɦ�~�0Ŝ�?�A�<3. �r6
�3gK���o����LYd� ����DCAE�|�u!o{��*É!�K=�����o�s�}�W��|��(�
�j���3:�_z%Y���f����\]����b�I�&���,�Hm��Ϛ�,AOUFQ3���#�֔ ��u_�1߻Ŝ{ڶ��d��`�����)�@5�=��?�ͨ&9;> �������5�������B7�9�Z�t9�x����ַ���z=�v���p}�w����x�#HNӡ~��q�h�Dd����d��s�7XƴD��Tإ�
Z��N��u�k�9,b'�2���4.����l)�B@�፫]�{� � �S��qұ�޸ޅ0�qf��<P�B�V�
utg��P�o��	2+�3È�<�����d�P_����X+�3����3�s��5�kFmtF��{�q����f��0�C�R���%�I��nZ֒�����)C��p^� OΥ�=e'k���>ͤr.�|6xd�'��Ű�֚:>�m�87��i�m�F�	��>|����f�
�8D
���?*ѥ<�	!�`����7m�T����#��j)S��$�&@��]r��=a�8'*{#:q8#3>-_��t�Ս������Pu��P̜�LHJj+�����
ә����ŹW�y��<�H�+nq��C�~��J{�7L�3���������3�k��H�xI�����N����@ߦ�WhL�>]8������.��-���/]���A�׊J��nB����S���S�	g��F���5��Xlgu�;����CO�%H�uV��������Y�{�&Xt�C4�{<�Ra%s�cO�w��7Dg��\7��@6�C�c2F���������0`FJ[b	�m�p���O�0����л�Fӽ�H4{r4�bu�~�4S�W��ۃ.4�Z�P6G�^�n,���m:8�V>o�ny8�C��{����ӹa�S~��c��[}��$�GEEft�C����j�v[��A��&�3��6�q�#��^0i46U�'��Џ�Ӆ�f�b��a��V �^�׿g��ݸ문�9���}nK�@A�$�?�D�?>~h���
��S� m��|��+�m&�B��p_3��h�B{�xA�M��Sŗ��m�*ߎA/;M��C��d��D�7�I�Q_�!&��]�A ��r(��&��$F#�`¾�߲'<���rBK�j�c.Դ�/�x`L@P֮������2�x�&�ٟ�Sp��X�k�B�}�n�Q�=��P���ڭ�1��gR=�ѼO�&U ��	~>'|w�u9p�D�-.�s�cg�2����4���04�=UDX���'9���d|q�3��3�_ToD�8-0�J}[�f~���VD�(�KTf��S~!u9�*G���P�J�Ԣ5�D�M�!�Hp��('�;����G���3[)����4��"�PK:CH�=�f8Q��릂��u�c���F'I�2ݐg}	thv�h$���"�K(�2�Y�vF>ϒ����f�I�R4�d��Ē�X��;�1����]��g�_r��� ��к�}����m#[�ex|@y�<<��MqJ��G�`�fH��L-X��#3�7�oZUyd��mZ�R��w�F���p�ro'�r�8�<$7����J����]r}�KxK{��nSD�mA������K�}j�[�/���}�p�T�&�������]����bJ,x��@���m��g"��=���2���܃�Gj0,<ꥣ�TJ�o�י�<|��oojpR<��<u@(���K"�_9��,4'�