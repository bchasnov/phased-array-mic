��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ���L�����I&V~u~[rR�C�XT���o����۟�V/]�@�!ӁUټ��)����؊������I�Xa-�w�H}�T0�me��|_��������M��)��H�BK���G֓�r`6��Lg�6�ދ��׌�ŵ�G�0�2�!�J��c]Mw(�C�����Af=�Эh�c��I+ݎ���O�� ��^1��0s���=9�߸K�V}9��^��*!�S�����p�QtVx]�����S`�)|e�_R ���bd���_63Y��UgN��l��"l�����I�Gɏ0�4��<vT�5���m�༇�µ�U��H��z�4�n]����-R������ބ��I>��L�� 4):E���V!����Q##^W`(�
�P�CI[q���Y�ӕ��Cp�5뿳�p�3� �agD oa��EčgF:K�=/��R��MV�ٳ P�"�:����Zk�Y �{��W��ϗ��ݟ)m�F0�XFk5 ����V�ӹ���:>�H�A_!��K�� pxH���КϿ''���H���%��?H�} VL�Wj��	[��WUt��6(2�"��M�2��d�)��*>\o�䝮6g̍�u&���;AV�{joНgl�z�-{@��oߕ�����W�S���i�f��5+��l�u�Q�vdy�-u��D�d�~�W��QX,_�_�IZ��E�]���v,Ik�5R̅<	�{�B�v�ū݄8��Nf�x�L��_��amY�A�A"���g�.��0U�8W�Y5sgVu�e��s,�	Ә�׹�+�YŅԘ�(g�Ӟ�Le�oӄSm�D��7���y����e��󆟤ۦ�^�شf�ȹ��Ek��������ڣ=��1�5#���Ef� �q��B`������+�#��n�$x��dא��ֿZ*+?��ȣQ a�@�����DX-�ߚ�6"�NS��"������ɏ(JW�Q8Y�Tv��LBb���J>��r�6��XSn|�c�`'�	�'f|���D��Y�� �5 ���^��}��<D ��O/_�i4�٥%6���I.��~�0�<y2��7�`��Jh1�e|�A�$Fì�6��T	���¼��n;W��qJ���&���<=�{$�?n������IDw	�^
�,MCIo�-lKeI��E�${��D �����>���hc׀T���C߉�u�t�F�Q���5�2f9�9G�u�dG�E<�7�0$ٚ>�N���r��EL90����i��"te�8ZT����c��H`���B����Ff�?;-N�S�`R�H�|p�̧?��"��9�N(�~b1� oo��� {߹[��sPõ��_�s'8d��Ai�/�G2kc<�L"��<b^s�����Zߘg�iwR����`wO�ʨK/LkOZ��4{��؞�T1�и�+H�|	�O^���d������FK&6+� �ǿ��6�B���N!�X0��7GdP��jg�Σ�4�+�]�Ӽ�4g�;�V�pR%Ch�ѹ�x��J�1O�xB	�LmԻ���Ɛ�t��ly��8��2b<FO[h���x�r�E.c�X�e�q E16Xi�	
�|����$U�ZW#�K�|Q���'������P�㵧Zz�j�oFc~ҟ�$A�_D��1�z���&SoƁ�6�]�6T�ހ g��$�L��FR
'Oْm��Ȳ��@�ݕ+���l��e3��<�RH
�M���;Ŭ��;M���o���ȅc�Y��uv�=;���}�y�]q1����~a���%R�(|����몥�7���V��Nh��[K�ppMݼ]ՔZ�`��Y9���p|�|#'{/�o���V�] g�>��y�JUn�01�7��+K�Gr{����s-}e�Bv��d�i���|��� tJ���}�鵸��nh4I5�M��3���/�>��� B�	/FF�r����C��ܱ��j�+�� 6��<�(l@�<�e����鄅V!9��1e<��8���� �+V�{����4-�V�WA�Ð�L�G�hY����g� ��O�]�"[3�@J�@�0ȶ��S��E��\%�Ƥ��L0qQ���n?[QrY�����2l��t�� �|�$��Aw9|�ODR���RƂ
�Dw��O��ܑ*B��n`)rޙHn����L�t0x�� /�9,�L�y����#x?*^��)T��b�SsWع��`�!ɨw�'�£:�gf�9+v�]�
��K\�0j���,���fj�?ó�H7U5i��Q���"�f��G�� �./�> �Y��
,7-/�(��S��Gz�a������Z��p��-MEr�~C@�g����zv>?E=`��F��pT�>EF�
 f�A���&ݬSI�\��LE�e��_#l�P��T�����+.��hq�F���tD(ڪ���苚P6�
�6=�ǭ�"���%�M� !!-�<�f�r���eKc�!q����b����E����SB���L�.�E]�'"���ʐE����ab��@�9�/��ҧJS(��B"��w)R�q���F�7b��Px�ן��3�)�ӔR�J�#��tF��������2�"�u?!t��j8@&�X������A  Q�ϔ� ��cx.�������%ě��_�}�����J<j	<��y�a��8V��*UqI��D�خ���!��झ���׵���OL8�H.�v�����N�Z��}����;���in���C��S���3�p�yO��g�m]�P]%:9j6�۫������u>�X1 �X��t�CO��04�-grq�o�d���V8���]��{r�9ͅ��s��ЍG�!0�>A����*��jު�TVq7
�FO/�\� ė R4�����^�v�������M��%Z��t,8��֜L��Y��#HW���NՆi�d7n��-lG��������<�u�۱q{�����z��t �vDP<�R�7�/���0���¿��T��!v/c��f�2�?!:�!��*�y����β|�>�1�in<�J�gR��P��H��b�-�gև��%
�����9O�V�p�buJq��6�g�E�yT����A��lser�|��-ߙ�c m��X,R�Ύ����r���ս>ސG�-f3���)��7-0�!=C�~�0Nb��I�B/1S�+]�g�!�@��.x�Ҧ�;J��=v�!�J��N��Ӥ�Nb�a��֊�H�;�r@T�wń-v�pW�)����0�����&��j�E[���"��9,)�5��w�M��H��)C��� ���):6�H� �fVꉳ���dL0�"�?EI�&5Q/��