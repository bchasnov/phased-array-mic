��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\����q�?��e�I8�b�Ǽ$��"����ׯ1�V0����1���=��7̓�'��S�F�ˤ�EN�V�>�� /�C%���!;@3�ɒV���7�/��f��t(�RV����U�~FZ1��A�0I��j��C;`!�Lo�CcU��ۖ�K��G�P�P����/�s3����;z]�0�!M˟�N�w*�!�����l�]1fV�0�?�*�Ұ� ���B��h�y��gz��P�3�6�3D���$��\PRH�.�t-DQ����:��q��ǿ��\�dS`����Ǜ/��\��>�?))$��O�k��L��]��p��&$Vܐ4h;
�k�Ҟ���#��00#�`�HǍ��W��H�R��Lq�
�����i5�n�cަ;6Fv7�������������(C��o�E�8~I�I{�EW0�V�xߘh4c=���az���!ݮ\*qi�݌A��69�f�7�k|�\�G��I�6L]o�ir'Y^�=Z'����Un���nN���T��	6���|�`~���"�g�x������v��x D�$��f��6'uD�v���(��u�B�`nΤ�w���w{òKa6ϴy1G!�nN
4W0�j9A"���A��,
�G�RB�!��C"*{D�I4�@@i����B�8~kS���@� ƈ��e�.�N=���pN,t�^Q����=���Q��2zеַ��n��4�68�Z9?l��������L�E�s)O����Q��C1	�,l=i7��NsTC]8����c���N��S0=IBˤս{��Dy|Z�1��Gm�Rd��t�����Z�
�(Ym�	O�t<fJ�M��Co�����, _����ǌ~R��Y���Qr=7$}A'�9��Z��o���b�%�J�wK�PY�r*ݵ��P�@s=|�d���sѢ�mUz��H���3KV��n�^k�Q^	u[���i�B�5iH��DDؕ�/V��	܍��T@h�=�Y[�K_�B�䩖M٥T�1�a�
2Y��&�؏��kQ����ƙ��3�d��?d��W��ψ�#ˉ�YN/m����摾ϊ��g�>ҺCK�7.����� w�W��CTQ����h��₄��q֊u��Z�G���<y�b��w w���=�J�v{I.J�������!�� � Q����JJ�\$��a��P_8���h�{��f��Fжj��ڴ�4��VU����q���{���iO��%�+����,�E1Kሞ�)�JI~��'v�4��ղ|B��r��v�_���|?����fC�Yg�o�O�sX�r�d�MPZy��=Q;�t���*�ݞ\_�,��R��/�D���ˤ�Vg�IG���.���c׵��\�E�c�"��Q���jA���Q��� _Q#�� Fr?
[�p�lF|u=/0
H^���r�_Kt��5������z۠�d^U:�t���*6Vq��zɗ"/Q�Qɏj�����ur�N�FY�D�p�@�?�,_�g���VF)$�rгb[�b�,���U�ɻu.8���sNPEGj���ЀO'^��o�N�M�^/Q����ݛڂ
��Q�8X���1��}�I���Hm�L5�q�Ox�j��[ׂ���D��\� ����ڌ<Όs�@1+Vm�:3J���ĝ���5�C;й�~��&�umW����P#[p�g	�"��CtGZ�p�i���Ʈ�;�� ���~j��c�n'�2LPr!�Da]�L�P6�b���ox��A0l��>&����p�#!x�퇩7���Sڷ����)"��PbY�� j�ߔ}p���Gg��.
���rmW���o>�zk�J������؇�0���v��@2B����.�M`l�Z{��� �Bw��x�t�� ?����+��:������D��;�;K)���Q������^�9;��CI!����,s'Q��]���^	���{�
Q4�wv����Y�EF�o�4��0<M�"�ډ�۽F��@��"	&%g���/�aPM{��s
+j�@˕a"����|����f���&t�(X��:!�_���Z�/P��C�.:Ɩ/&p����|X�4U�b8�7��+��?5�8��HZe@ogr�e�	��H\Ȳk{���b�q����64��Z��_;�P%�e@p�Fi��ѐQ{ �K��� K�%���i�Y�o�C���D��x����u�m���twQ�$��Fn��0�I�FQ�� g=�7��_5L�yG)xIlQm�➥��5\"��[�@�d�A�c�l��h(�A=3��-r,�������Qw��;4o��*NK���Z���ے����ꬭ��Fc9�gP�t���O;���B'w9�S��K��㾤�'H��x�H��Pam��� b�/+ts��E@��֪D$�}�6K��]���|�e:�7�З��I��9�M�y�QL�K>�խ�����W����`6-��q�Y����]k�ya����L�Os�!����8� ��f��p-8!��CNq�\[HS�*:>��6O�x��*�Ua���"������^#pr�*�F	U~�~+�3g��S4�ώ��m����]k�.^��䴸9'(��7�N��c�J�Q�;���0u,�����z�|`8��8�Vkx���s�V+3��S�C3g_�B�]��2L�K���R6�_Omg��pn�SrJ�x����m��f��)Eۤ�bΒ��v4Q���#U�ߖ�SKRa�̐��4�����7Ū�=�g�>S�ƣI�}�A�����	N!;�}��~������Ϡ� ���e8�kEZv["u��V�HF����1�qK����@v{��$}��[�#��{��k��W����|Fn�1E��!���$T��i�����ʭħڤlI�¿8>-��қJq���t���n�n�*������~'�&��_S�7����J�DUz�;5�]i�j׈Xʮ_�72V4��6�&�D晴��8W�3D�����p�����L�����'��u[�A���W�\.;q�u��!)��Ӫ���N���j!7��}�T��68/-�����55��q	^N$�uP��'Zp��Kx�m|y�r9;r��y�t����Ӝ�W�۫�k���5�2^Y�s��l�B�q7�1�'�80�VE��RF�}�m2�"��+��UȖG��3������Q}�'����=6���g�h�
�T�������s��-��o�+,ւ8 ��I�s�2�q8g��J��H=1�e|���4�$�;���ې v��|��I��xZ[�R�~=��	�"�	r�����5�"���G�n����v$���"!l�bA����[T��F��9�~�U)q��ifݕ�n 2./��c��4�W�*�:Js�;����n�{K^f����]6T$��<G�#R�b����y��`����ȕ��S�c���c����j Y �9���yoM�QUs����I2[e�}��~`ϻu�(��(�!Hb�+�i��[�~X��������u�#L�{h��rd�����=�V�Zb� ߫1�5��,|y�"���e���%Ǟ�J?�xC�a��Dl���{���� ����A�ʉ��}�\)�A�JW�k�uG�Pm��H�ҙ*50J�	��!�{�Gs����ud����-�FpN2�RSi�_b��a���M�O��������I�I/O�#�1~����{j��&�� ���M�աh�D�e�;R�z\��ډ�6���-yj	3���D~�E���@ƕ��=���3����B���{]6�-��:5��vy�N�u������GIxl�r�{�����f���h.i4ߪC�:����N��%�<{�DPs�KX� =�<W7��+'S*3�.�DVY=X��g�E$��R�&���79`���
"��	kCJv"u8z�"�H��.~(��s2t_��YP�����<��Ĺ��҆��j�'����DX���f�Zϭj��9��/�&�ݛ�@ǳR�sI�iWùNn�y�v�n��ޅ�>ϴL�3|Y	:b�*,d��9�k��YDe���`�bۣ��Őј0�+��~��M��-�un|01;��'�f��F�ޑ��*~�i��Y�/?�V���0�1��[>��'��/�J�{L��G� �@��m�� <�(@��K�g��2���wQd�$��˃�J.	t��y ��]s�Ի�r+�aΣ��V�wĒR�k�4+��K�h�p�-"�����D�?ܩ���F�V(�Wm_�6Bs��������s5������c̤�m�Z���P;s�= Eq���i�1WXQ����DL��-�Nz���çt#MC�\���O%��'^H������㬀?�@w�ݏ�-u��0�v #�t)O�e{���4L�� ���eq���rZ�	v��'�T�C.�@,�u+�<G�q��m�t��lI2ok�a�Kr�V��= ����$�	�'�e�V �������j)mb����Ҷ�Zt{��n[{Q��]��2��_oc�y�PU���/�R	�,
l��x��e��c)�I��}��_p7z^�拘ٶ�a��G�S���Cp��.Gh4���jL3k�'��,�(?�bQ��xw��u�{n����	6D<5������"��>�R�W0�3W1dtz�*
��	�*�3;���K|A�����)�tp-�����Z�l[̾�����֩�n���!҂���b�H�D�`ؙ��nij�n�q�@�3U?���x;��X܂(�w�Jw@���?۝��0㝅�R�8�#��t�1��~��V����F�U ������ޢɰ E��p[W�}��g&*PƘ���YE�=�L��`��La��hT��.ĀK��L֕�L�3��9��j�x(�b%靟5O	��BeW&�U>���8Ϗ�"�&�d�a�]�:.aP��"�l&��^kԩouĘ�vD]��'�7��#L* ��;k�)�H;��v�[���	�C�TY�F���1ܦCqQ��Sg��+�k%��9F��4�:UfcpY5�Bl�pe��ݔ��q�1��c��_e��30�Z����K��T�^�>�+���� w��~�)��w"�U�>�tbbl�.xQ5N	\�q~���ג���,�;r��-
A�V�3���ȟO�8�\p�h'$ش\��<�%ƷM�:�7��#aî������ݛ/_C�z}��YY[w��j��v��.�����BM`0���Z�MB$"	��t���H��u�h�OX��;����y��I+�Ѿ�,�d�o���w^Qt��o�����p�t:k�+)k�x�*�=L�Zh�&�<w�\����.L��V�#B�<��t�
�M�@� ��5K���B�����(�x��7@��Ji'�͈�A�~�=c-���Ҥ&Y��E�X VB�
"J���RS��2��Z�0i{�>�C93���g���n��Y����'xV��7�gxkT����P!�on2\$���z��ٺAO�<f���]�i�o���C�92p�����/[��4ض$e�Dڈba�Aڸv{���@��$�Q�Smh��
E�*�ė�bq���v.q<en��Q�C��6w^���Zƙ�tm#�l.�O�������5��qD��b͖��<~X���`I!O�Rť��]�u"f�;�T�iN����g!:ΰU��'�GФ����` ��x�t�gr�߈��ok��q]�{e-��I7Dq�V@��Z���tXo��D���	0Y3��X�%�G�fII���Ӿ\Aߝ@;�uD���@(��y��j��fD� �"pG���!���f3��9�H��|t��J7�ɶuEDjF˟,Ɩ�jk�2��$8j`�"f��v1iQY��IOYu���\�8
�ToP���y^�X������?YZ�&i���3�~���޽� !�?b�����mz��tX�]�C3����Y`G��?B������O�����?AY��Ƅ����,���U�괇0;��U�FJ!rT xz�����	`w�"��;?P�v#RmV�t��1����d������
��n��U?��h�b�֍�׿���E���p�S6�q@))a�[2�,���q�.Dx�2������9
]��}nJo��7Zd+���0�V�uG9�f��jG?)�gn�_��^�pV�Tz�ق���a�D�m~��I�G��+�:�,�Ǆnܽ~%������~B0�+���YM0�c���h��Sw&��V�\S��5��q~Q<�C�{��s���g��ZL�J�����sE�hY�Gu�vl�lp�}4$�G=�0�\��ǚ���r��m�+*	L�W���.m�L�i��M�������R�ՏՒu:F�S��B]j�GL\i�C�Q 	m���������km��3&�wy2�� ��n��#�|��ş����~v�x<YA���Uߊ9i�OH��X�[^fg������5SG�5;'=���x�Adt��evl?��?K"�v��BSZ�H7Q�e��0�U5���,�r�(�ƥ*���9��a�oE[ fF?��e?�[I#��S�:��ۛ�=X&�����7���1�+�����a����� Na����)T؏�kPz@����������|$�l�:����{V!�Q\�XK����S궪����*�	O4�k{}��_I� D������d�T���d��׫��ԌAO��)�:.w�).=mS6���C�l�4��~Í+G��3�8�Z ���ej���(��{Q:PF"g\i��_��f��	D����5/�y��n˶��fj]/�l��������0X0�m�s/Ob]=����źXҥ6ϢA):��\�2+T'�&�����z�i��|IB����:k��^%�R�N%w�
R{�f��#�@��/��ۛ�ϱ3~tJ:*K�5|c࿩Ak�='������;��}�3�ȯ�o�CT|v�,OT���E�;��B���$���w9�  g�27�՟1v�Т�b��N�
d���C�0I��wԦ����t�Nj�Ք�)8�Oi�ԣ�ћ�S��%���9}�%'6����'>n��[}�.��r���Cz�oH��$�VN�3 �Js��J+
�*l�o )+�����/������j$7yKc�{���b$Μ� D]v��(��.���-���k���>�cw��m�c����"��St�c�X��C�"l��7d��O!��/,�N.G2�m�h*i{�]����z�z~lc�:��.\ź���hS�qs���]��z�>��/�8�������X���
F�%gp�]9�G���gS|S�U	�_�E���o�����tM5x� �$A6]H=�]���| 
�$J�}FS��&�9���6S	�^!ʌ%�������)�c��6��4z�n���Rw�nT�p�X��'J5"G񷒭�q r�4�WMX���s^K κ���%�z��eM�E���Mӭ�*}�	}`*+�}?u,�	�L�ʖI���R���>x4eh40F����E�K�6�ŗSϒ0�/8g��������!��*��'�k�٢��H1̮���`O�M$|]�L��K���n|f��jIc�ƉT���  bU���Vo����7�AQ�����X"����$�68���>=$C��x��6��&-o����A��"���ۂ?0r���H�w��y�t�M�K'��($�V�9b�]��]�Y��s����L�ٲ�d���6��[y�f��m GM�����o���n8 N�����"���y��K��I߀X��C�:N㊵�k�Q��e�R%GѝR�����,�K1�[D��Pyy�����
'>��ҝ�)�?�]����>�S!�l��d.�������3��G`U/��C�<5P��6y�yڧ�n�/���¬ZgJ����~��Qkt�Z���%H��7���~w�-���*�?;0�m�Dxn���)�I�����;I2���o��{�>$Z˜pR����C��Vu�=�aV"5���@ep�����'s}���P����]��Z��?�~`zdJ�}����@���\�0^���K��5`���/=��(���)�S�<'�/�R�~2�z�R�� ���Jos�~�v@ �.�:�l�X�0���{�4ҕ���$�z�X����B.�Y�;W�����ڛF!������k�fX��(��l���!�킁&i�ޏ�Ϋֻᘅ8����c�������eܭn�A�x�����'�v88O��h�KY�$j{C���0*F_��x��{���.�z 1��\�<�>�U��o�b��DW:��9���F���h����"�����Bc/�衫�hk�ň�mm�e��q="�z����N[6�r�&6��=k��Sj�����0��ڰ���钦�xJO�ل����j��\3?e���M�A+C� �φ �+�?�a�^�qDS����z����p�ǘ�9���n�|�7�:�X�����b�+^N����E�ÆN�3ٿ�b�6��@� ��˴ٹJ ���j���K�:�tDp�����iD�<Z�7v�h���4��4(���ճ��l;	)�mʍ%�==�9�bS����LT�#t�v��$����)�P!��k֍6�[51������/5>PJ̰E�b��t�1�'�ɲ2�'��v�&�w#B����\��u(��.�K�1�8�"�_�⥮M�;SA}�P@a�*_z?!B�Ѣ��l��"�E�F��
������u_��!$���@j^�D|�m󞃕���1���-��d#����F�T5����d�1��zɟ"7�;�S�V�߭�}+�#1I��n+��Q�+@��(�|���N�'��ҽs��\��+Z��8�[�������g��ȎoDಯ��&�'A ����5�Tş�߽I3���"�
��@V�`��pD���SޮU�����,U��U����~�!��[�/��-凰Q{�fv���a��^�d|a�S�Z��k���t�Z��Io�K�o�v��� �p�)o�>�d
f�A�z�Ʊ��c^�I�
܄�}���|]�=�
��T�;j��,i���=i��(����(6itԤ95�)���_ ���=ӛ�,��
������c�>��:s>YN���7�"�'=K���T�>��!���)ϺFe�C�++%8�lX1G��ކ���vR�E`	E��j�T��4�F��Z^Z���F�w��t���� �'(8꿩��{`Vu�Նպ$p5=�N�˘�-�<��S	��%,c3>���?P�w��lܔJӦH���p�g�h*�\�|�i����"�<+h����f��{�ygk����F��+qi�V`y�EΓ�!o���-}`�F�Z�����[��h�	��A<~�<i��~��ص�)�3�@��#��1�a��ӮݶnկYݩbU��M�[�[}S�X�B��_ �Ih#R�����?�ߴ�⭌�%Y��q:c�ᯣ��H�َ��eޘ�w1�h���~Փ����I�ӭ��guMA���1I�8���D�ں4\�t3�d����@y���9&=%|S�2t�`^���މY�k�)�������A�t�jN���Q���u=0@������������<�m���:�y�$$�������ڔL�-�Y����_�=!6���F��K�T�޼251X�#E�U�:�ٍ*�^���{�Q;�@��_ʇs��O���x�3�����2����QW}[�����,{��ne�O���������f�'��sg�N��{Ƅ{�������lk'  M5�Q���]��=�mw9���&�Fn��|��>�y%A.�"4p��tc��/���&JT_��,B#�ݥ�����)e#.��/����d�o�'�F�4InS,ř8�X�q1nL&�7��6�	-w��1�X�HR�$�۞u,�u���IM�`�$(<���H���M�i�����L+��-����9�t�JVۑ��ƶ�uW�駧�
�0V���Ҝ��@~�vR��iC�5�� @<���;�go�z�+]B}���Va�%JB�o�8
�GD�9g>���D�H-]~�,������aFs�7��!o�;E��z@���bzM�*2:��Hz07��Mp�Wl���_����U%���%��K�F�v	c�-�c���� 춆p�{)e�G'�6���<?I�i����>w߇��~Z�.y��q:uPz��Ѹ>Þ�O�Ma����ˮ�0pn1����<O.?�k��s�S�����Kg��g��r�4j�� �5�य़9&52X�7�ñI��+,�:5OSI_�������j_Du?��g�68f���H��;�� 2бg��G���q��������cA]���AQ%X��	���V��q����O���4W�A���c`���pΑ�����p����+G"E�����E4Z�	�eV}M"�e��\�;}���exL���l�qHy{+iq%�=�|`z�$5���`�{���1k�	5�݈D��ՓJh�Mo����!)��x+�������|�f"����W�bL�qc�p��@%}�b`�}��;8L@�=�'���x�T��C��4YF���KG�"�V�x���Z?��#��j�h�N���b��O� �k_$��h�� �c/
UV3?#"��{m�kܙދ���8�å�'~�(��is�'m��m�|ݷ�Y類�=�v>��$���!)=W�:��n��qiuw����r���^��
?����s�#�}�@�������$M�݂.G��4��h��/����V(ۏ:9�Ja�g����h#4.�H\3z�?δx��ޝ҂�y�:�z
Xi�!����gz��5m�w����WH ��اg�,O� ���q=5uz�+` �C��e�=̕�ζ�v��g�c���oֱ�VL��C����KTs�Yi �1I�;E����#�R�ያ�]o�c��>#fĝ!e�ŷ7�B(յ�f�cf1�D9�9?��g1]\ށtz�?�?�������sX�[�w�{�^�`�Ԇ�+A��I�d">|1�>�"y!�.�<��Y{�{x�H+�Ġ�\46~��n��$��7�h#T�<CF�/p�Cy'�m�}
�G�SH�3(�M
S������Bp��3qe���2��@v:�a���JWX��VzNv��]Z(��*&ӰF��hvM!\Ap�/��1�&��*S��B�����r�_AQ]�ak���J�38��2Bꘊ��@}�:|M��n}W�.0�Al���V�ߒW�l�c�v٘s��կ�:�B,�X	}<�$*����S���@ �ӑ����ߒVu���䍿V=	�q�o��WG���2�K�M)NЙ�.�+q�J��m.�S0k��}M $�y*@�G���	�Գ��fnV9���C*�/�d���c-́*H�����_h������l�<娤�3������!{4�WSkf�rq�>���*�.xf(K����临��f�?�[�,�eȔy���I,<�������h8:�t���۾]�2
��b�؋�,�-1yȮ/Щ9�������T������W�D\����Q�%�e%)����R�1�G={0��R�i��.uR^U�}��L~�{�qi��ˑ�,.tu��fÜ���l�omKS��|��|�����8�I?I&��"7�Z<?�(�vJ6
��A�~� �]V66j�p�&�����L�xdXW6e�ŗ�z,���+6���S����_�{�t�`'31T�_x'l�D{��~"]�?�{� 97Y@�j��WHXsځT�ϐ tw���M��T�j���(&��4OYa L��kV�����	��W�St����MI�f�u�{��c�|�{�m��S/�"<O:��p�\>�6j��� %LZj�?���VX塚��R��&/.-ΐ[���������pi��(��SI���35����a�D�;��B��4�PE ��f����IEH�v��V��|t��}�z���j\��B;�f܁��ȗ���9&p�4`^7�B,��(�<�	@�p�
���b����5�d����n)�er+�#�d�B
g�Ir43��h�H������@�M���G�eA-�D�5�`\�����P��L(���Ñ1j�B��I���7�A�_��bW,?�$����S����&��� .8"E�uG>rF6Րj�(�V� �1��X�"�R�*G��$m��Y�ґ0�y��Ċ�#L�'ĳF�AB�2��	 ��n����|)�5�{==9�B'��vN͑���I����|E���և���KW�����Ȇ4�5/��7���Apͥ6p����XJ�2.���Ë��$��V�,"%y3��&9W
NR�U�I�$�nVa���d�4�E09B7<�"w����2��/B�4beS�;���$����ij
�F���(2���h�قF�3�?��kx�Nv�Q.X�P�ͭ��!=�1�����4��"�Q9KyQbƭ�Y�[���NX�A��Z׹dT�9P������B�Y$vws7R�g7h��.�Vt�����U�����G�.�<� ��=�̿�C`�~IS� _��%�Z(7]��}�*μMciV���^��Xs���'Nٖ�Ͻ�Z V<�ZZ}�<���[pK-f;�KQ�!�\��`q�ګ.�"W*�K�=8Qt��-�8e�0>���y��y���Y�t<�o:ǣ^�Ӳ�B+{��%j戫���)��?��WqK��{V��3�>q�E�� ��ryd.�9Q�&�͢C�Rȯ,�a:u�R|�:k"Z�+���r��2� � �d˝��V�t�=�1���U��S��m��'�T�]q��$��_s�з-��	�2�e�j�`]��������BO($MmQ�	�A�T�i��~��������v8#�a�<L���v��\�6�L��t��3��UX�o�a'^�Ǯ���iV��b�Ad�E��;*�"L�q�<��,�#;R/Q�к0gP���6�K���1�����U,����{��qeٺ]n�N��TUݜ�4X�u#4�{BJd��m�J ��������n�Q[~#Ud��%���'�����zAT�8#no̸��r	}�������!܁p��TG��yY[��̺���%a���,C<E���Y�?lu
d�6Ot��0��&�p�A+�D\�5z~�+�T�S�A�eI�__s[���i�N��"V�K���~�O^�o�鬠j��2�;��pe���B3����=��S-�D�@�ꌄ��(�Sw�J���O�l=4>�~�5Sr�86i�x����O:��#�͟mL'������ޡ�yuA�[��>L��)(S�2Uo�$��%50���26aK��笼�Q*dKw���O���d��_��j��������*�\o�_��b��v��kY�)�.� ��D��BD؀�	T��f�Pʴ�
1��d�Pw��
~.��dR�ϵg�����&,�+4�paj
i��C=�өA�/����w@$���*!��2�5��!����^�b�����ȝ�6f��ژ}�E�P<�R���o�����wb�\�;�eZ����_VM�� |9�i�$�o�8`���e�A�~�%���l+��p���FAd�;[�>ڛ(�٢�9�\r_S�R#�r�y`*�]�_�q|��'ҝ��CImx��ٱR�s�d6"�Td��Lz^���cK�ד��7�|+ĪY��:*6X{o����>N|�����[N�G�~���dG(�3W��E���_���ZC�e9j�~�����8�K�;%�2��e����/�`Rlzӑ����(C���l*X/ž��\q�o�^���I\:�z����J0��,�=��a�Ks*<y};��E?�����!���,��rU^��&s�G�(���m��ݥ�(tQ��voy��� |�5�q>���䙃e��:�Ƹlnxُ5;�H*�����<H{S7),�ɪlO\sl��f���J�p�'�1�w4�]y��#����,��@2*@P=7�.� �12�A�%����T�N����c|ɦG6.�P�i`U%}P�T��_	���y:Hj"� zHu�&�	�	�������Ӣ��K�W����	��
��d�i���w�n�8!�G?�~*?Ç/�-��͕�T{C�άI/��P�Nu�=�X):K�L�`_�F�1�_|����UlĤ{A��=���g^� p���,0ɢ[�e��aɳ&i����V.i:��?�3ӹ:DWA��
jx�fd����ꐡ�14q�ɷ�6���B$9\s(e�e�"����=#�Nರ�d��T��Kq2�=5X���������h0/P}6��ż��Z���Y��Ly��Ye���%�	���f�Bǚ�nX������ �6��ec�P�o�/��.�P �!��B�Ʉ�RN)d�_e!��<a�����®��/��ߴ���2:�b��׵{G;���%O�N�^�O���� ���YiL�6j�>|KFU|j�!|v��4�~�ᙩA6�a�^�����"��-%��F�:Bod-R|?	a��h����<�}g�����b��S)q�C壜�&Ԕ�8}[`)��k�Deg��Z�A�_�E-������dɺ����Ub���/Yl�@7��4�����Z]iT� ���F�&�
�4�"�s��7�ݱf�z���<��Ǧ��ЉNؒ`{õ��]�5<ˢ��R3�hk�x�~r��bb�d���Y�����ɥ F�YGlǆ�t�}c�K��t��4���m�I� ��c�ӏ���b�tFKeY���.(��������߅��E��a����p�����q%�*�����޷n���IaiU���d};�rb�c����Y�4&�U���?�xFɢ�H2��Y�Ơ�=8�2��n�z�n�-Ȳ�.�<�ޘ
������������|�6�
�3!��{�K��@
����h`w�j�b���t����j! ��h��艔w$c�����ŉ���㭧�s��鲈n�]K��4g�]����r���1�Z���+R���T`��o�qO@f��֎�w1@0�i�El&�2��!�8W0h�׳�Ԛ�-�~c3B���ecΚ ��d��S�?
��>Q�/
#B��v�@��(��r��u����)!E�ϒ�TL��I��e-�����e�."��I��5�(���˗Z	2��x���;ۑ�J�"��.r:+�}�`��8��O�#a��㤏��5]S��&ޭ�O��E�t,t ��/m��'�˦>@`G��d��\��lH����ܷZ;;�Y��򉧢�t��H��y�8�&6�r�5j��/B��As<E�`���#��o	��ގ�}�#G������:�I���'\�Ly-�_�(=��8�cr�ż]w�'����X#OLh�QҖ�2"<;����7�u��K�0+0R���ķ��Ҿ�zD���LP\���sk����(�R�Ne��g�c4k�G.�#F >{W�$�>� M�UgpK���*�0�0�n��	{i|���.p�MG���M|h�{�r���qhɼ�6s�����D#@�~F&'jmeq�g�߈��{�}æg�Λ��_�[�$�2��}	V�'G&�%��3���?���%�K�J��D��Ŋ���7���*ϵK%�B�����0 ��a�АU�^�]f0(�QX�D��nG1@d�#�*�:�J��
�������;����L�&�؋S�_��<̈́����R����Zz$W�ZD�9Y7��-�i���>pR[��v�q�kC����J��`މ,g ���]G��Ҭo�
ؙ��\bF���uC�ɧX��"�{YT5�Vo�D�� �j��i�*³��ؾ�����V����^����膍ef����?0�*�*��{�v�0L�H8�.�o˷���Z9x[��U�[��VqǠ����N��z7�>twD�Z��.�aZ�%�	��;����:.��S���������xh����|H{v�W�;g�ԥ~9�}�i��Xs�pW�Ub�P��؛���+��i�~��ogꞭ�S��!ɟ�#�"���,N/�A�@'ˢ�������3`�+/����K.�z��/h���K� 	?V����.G�v̅����-=����o����Y��k�sV�������m�2	EW�<l�*���O3���ue�WH�XI-l���<*ڳ�?�0O �Ú�l�a�]�� ��Z� ��z�i�oV�߀�@3�s52�	�^�Iv�� |�x!(_��xW�(6���P��^QZ����<]��A�Qo��s�+^{|ْ$zƓ&��(��k�k�|)B[���*��a�m���?k���1M%�?q��T@R�P��#�:"7f��6�7����`�kg�i���Y����B�Z�H3ρ�=�QQ���A�]5A:��u����.J��R0}�ٶdhWI���@�a��	P�A|�@���k=�,�"`$�3����lp	<�Ř�ׇ���6{D���wXѣO�T�O��U���w{^�J�C����8������-����Z�;!��R6��<[�|�4�q�e&��(�p�H5!n������Go��Ai&�t6���3'�[P�]tza�O,CPD�Z�X���n}ϟ�"nc���k;�a!�y��L����j5�f����Ď`epOW����|��9YxAR .uA�Pe�"?R�����>D�A镀]��5U!�u'`C�eMw���h�p����B�)M%V���X��W-��nݐ�2�G
i��;mKy���R����#(��]����
��� k~~�{�u\}S��	*o ?_S�q ���?��i
C�B�{Z�L�u��Ke��ov۶�"�"�r�*F�v���CH��86����4b<�%Ŷ�5�X�K)�����N�V����	��������̉�4����Հ%��t���wn�#;<��J���&KwǊރ�n�c��.�5��l\�ލ:�5���O�P��9�7�*4�4a�����^Tz#���őB��'��)���4.V����ؼ�M0'����T�	�ܓ�k�Wẗ�?���T�5Mه�;�f�vp��7�1}K�����9*UT���cMA���9��Z+���U�V�tU]��+I��1�A�?y ��R��)Ԯ�U05��J�&D�����ЕD�4O2W?.�wm̾==L{��|���;u���Ǝ��rt����V��"�t�K"����	���oC�,u���m7[ p���-�ɞ��+�����g?� �O�S�;�Iy��s?���w�Hr�\�]�y
:�ONh�y�%��#��� �bޭv�V�܅�\�Ws�"�o���ٞ`�b�_{�nl���-.��E��\:��0�1�Si�c׿b��)�����;�S�7,��������7�l���.�7�]#�
E�`�!L�fye��MUI�Ӗ4{� �\L���!%���h+�S~��O�1)�
M�;�)��(�t���A���iz�j�.1����z�����w|dS=c����Q*T�h���P�N������TEh;�V?0���io��H��e��NR�C関��cN1&��<H��."�`S����r�x,� l��p�u,�Jbc��x�Ir�'��\*`��;+ݸ(�7�)�Iqv���/Ia�]� <D��j�,Krb���s�<�g�;�mH+!S�6H��r�m8\�>ׁ,2N ����W<8$ޫ�ݶ��qF�C�  Ng�܃T	<	�>a�E/̡(iI�C�;�B������+u!(���'[��,Մ�!��gтj��^M�HAy���$sy>}>!���W��t���g���sV�
`���pu��}>������v�)� J��"N�L@z��/�?zv��=/�᠅F�_�F�Mk��������G��N6�j@1���|����{�,0Oɺ�CQ�Y][�W�+�Uu��O�:�l7L-\;M\җ�՗D����_���}2�ԍ�6��tT�6O�"������+$�BtL��
%��!�aݥ��S���#o�Ҹ��=��©a��D�U�)���
�'�Eo�e\���&�:����9�,�3���W��,8QQ���w�g�Ŭ]&:��ε2S��s�'�53<L%vf�
t�������҄�Z&�h���� _��$MLi�+��EvX	��t�%f��%s<�M�q Cm?ޮ�AU�}5h>�[qB֗�F����������)#�͑�Q���BX_� uI�Bi��La�/�>̟�z�u�?���\�`n�g��+�/d�A��p}��=�}G�A"�������qߒ�ڮ��У��=a��+�6�J�7�a�1WX��1�{W���3�9�D�����g�
�
�U��ê	ڼP2a1D�ϵ:zG�o��'�v��:�a�X��%r��������M���K��K�T"�KwGx�u�?������^`�P�7���S{uu�S�,d�An�6&��7��&�S-�摓�қ��E*#[HOc-�9�W��,zml��Ū�Ҋ��ߓ��D�ȟ�3��B{~7�I��vF��{��CE�y��!j���3tW���:�?���R�<�)��?�L2�WGc�̓��S���W!Pq�T[���2X �[���U���Ҭ����M�e��%Lh	���C7+3�F�	�ަA���Fn�NAA���֛u��^8��@���Av�0ׂ���#�~�i�0��xe�؇�v�1ߜ]��������m��DD��32��IQ&K�O�obŏ����H��\�)�w������t���Ji��	�/��*��z�f�,����R�#����y��L���D* j?������#ݒ	�m���7̛xC�g\�M��H�L�����"��춚d�v�!%���̹:s>q���lۡi!9I�T��*4s�����C���q5��e/��;��"
��O��T��L.�����iK��Ɉ��Rgu�hu�{�iZ7܎C߉���C�ʦ-.P�j6؊s�jH��ߕ��g��l��RD>9۾�����Mn
y��y�!�Qb�H��������"���`�~Y�(co��	��"�z&�	gf�E�Z-��Qʵ"��p�G	�*�������us��¼D�X��H����&tJ�C�����s��tN0�AٱX���*��	�CPgL��j3���NiФz�ƠT� ��/2���e��1Y(~��)f)I��c�t;�U�[��6�1|G�|��D�q-wm�&�����8�r����#B�BN���E��MGG
��F�8���N�q��xhQ�J\�!_��X��A#J����P�fl &�T��g�Od}Y�;�f�#����c����e-T]l���ןAT�ZGn�7���Z�ܬ���^����s�
�����j����z����|����d��J�$b���vK���M��(�i��Eϰ���%��4�k(AW��??	dX�ws����<�G�5�F`knn�{�s�)_�P�朿я��j({���j���.y��Z������s���g��*���?�v�uq-�%�2'4!d�ߞ)�v��'	r�19�â�C7�䇱)�85������f�N)c��/�kk�6�3�m7W���	�����~�7��U��v�9�5CC���0��Ef�dR�.��$��㗟K�x�2m�p3@�q� w[�-��X�������>)�p;.�ڏi�	<MHb�A��Uw�HW=k�S���I|����t���G+�w��3,9��'��zM�_O�32cm7��%DN���\!�P��,���v4[8O4�j��l��f�ugXOh|`>�Z��
J�<���ϲ�h�c@t��w3v�I4aZ�4� i�s��Zw��3�$u&�}}�z�Ó��ǌ��\&�%?6�J�r�Uw�=�u��������su+A��b�,5>����$���wE_�}�D"���z{:j>24� �m@�6�"�d\In���:L�n18��x���`�4���$4@j�!+�>aĳ^^� �h�E������g+�Ro���]�+�]+pP)p�/e<aO��մ_lz\�_3 T����C5�MU�,��m��8t��*Z�x��\��ϊ�]�7��&Ҽ�C��-r'�o��׬oU��@"�t�u�Y.ޫf�~{ǁc���G��c���C!� �x�=,>x"���bKS�T$�mƏ��%@%|����.���u�p%����+-Y7�n��a�e(}�D't�Ӱs��uL%���y�yt˧g�TP'3�[0q�l��#$��3�t��3�\����sF�,�_ݡj�W�j�� �`�� ���LW6B�,2dpDw�?�'��+�Վl��6������܏�$/Ɛ�0�� Qd1����e�V�:�U������Ϣ��$8܋ZN�ys���m�y����n"B�����?(ѐ�x���QQ�/_Eg��c��[<!��>�FG�!K"��������K���M��.�@!~/���p����^�zğ?z𘠊�~<&�6����:���Jr�����np!�Ȋov~����a��w4�]F�����+~��' ���<}ً>>��m�u�'<�	�Ѽ$.!3^Qr�E��<���hCl�{������c�	�ofeH�a.�9S7/�)�̓e����d:�M�w8w���ڑ!�	�v]����p��n�[R` y�-�}�*9������9Xtz�W�����ؙ,�0���;%�Q�qZa�ڏ���t��#5bL����D�s	��	�V�d#�c��u�~���8��psϻB2~��9ʋ�'ZwT�����IX�S􄠯����O͎*]�i��x���'�Æ�+iv+ÿ������Y����qvi�C}Y|xЪJb�ZVL�ֽ���=ʐE&�.�p�Zg����#c�9xs13a�N�rC�����ngGG��ۗ����,hv��+>{�$�y8��[�����>7�D��i�,O�jO�e�v�]�v��I
�]�����n|t�n���Mb��d�����0��FսaL���4�u��j�����1����rS�ڿ���D�׆� >�\QE�h�4�t�r��"�>a����������B0X��oL�:	��ˈ&��h�+�hjeѯ_u����3���������1	�ZS*Ú]�O��8��W��~V�������o�ɏ8�F��T�=��iJ���^˰ Hw�x�UcP�[e��5y��3�h��i_����9���3�Z��@�ͼ���|�����U*��MH��IР�:��mR,3��qb#�����]º�!����gL�!���8�8���*m����J�CX����d�\�,�z�~y�{HSBc(j�4��qIq�},��9GHhzZ��١r�\�(�N�5�:\1៭~�ዤ�K+H!���!;��	`��hr���J��A"�,���0T�E��ü}�}eM���>Y��Ќ���7�J;?��LFSm�c M�BؤJ8�ƙ� ��rxl��S�)�-��i��9�~�D&]y�yGT���~Q�ҋ���[�Ji!Y�:6���9��YۛX@'jgԙ�󫢅o���P犬�?���-������H>����a�����/M�q����N�-�R^���>��r0Q^�Cm��m2YY-`���lS��פ8�g:��7�VY��l/�.^f�⮋��]q6xG�3L$��pq�73��r�Õj��m��%��̶�{`zu��f�˂`)��Dj6��0����.t۹=�"w�@还F;�T�o�=��ت������>�&7��y����kVV�	j:6�}=�p�W�����e>!�1�^�m< ���z*�So�D-M�}��+�-R�$8�o�d?@��Zm��M��a���ctI���������mId�z���$y��f3�$���Xc���/���t8(Y-���+50T�N��:���EdS�sy���ݕؕ��'N�,�-��%W�v���n����?}s���]n���9�|�Z����VY��^�6F�Y!��{u��L�Bao��y_"�*��;�5����O2HT�3���Elr�)�	^v�9�����V��Rߺ3����Ͳ��n�"��&Yp0V��~FYY��u{����U�s�`$K�9es̉O�djĊ��+��)����]y���%��t��=�'wh�1��'繯�we(0��Jl�>'sO׼!�i� ��\Ij��8�#a��j��"p�����Rc3��_;
��+�m��U0v��עFǋ�ff#v��y�%��۪vW�Tg�q��܇�&5��;ˍX��_s��>6��!%��]e�yB$;(�}
�P�̟�*����gǺ�����(�~<�X���h��4�e_��j_ϒ���N����I���C�@��-����7�>��@*�����?>�K)%��q�k�:�Gx��G�1R�o�7��h��ֻP���Vd_����L
�"]�C�lb�w�g�xR����ǭ�N
�y5�^�*�^�)4䫳7ݱch��Э!�̞(� L�d
��.N���VR�s�(J6�Rq�s�RMA[���ܽ��'I擿$�]�6#	���C��  �cH���Nֈ�_���=��w0���@n.ƥdQ�0|����Ҹu�� �5Cl䯖�^*�	"{���:
G�7K�v��@������b��Y����f-X��[��5�ZR%�!�ϯ�̄˂�ͨ[K"u�sьV{�����[�-�8�Nb�zb/�I䭡�`SD��w���z�kE,�r����e�$3V�q�Kt�3#ə1�/�@aH����x�Z����ȗ�R�����d�S���PY�찎�A�,V�:O�/Í����U
��7�,v,�B6�A}��A�P���YB����6�k��KV<�橐<��1!̙|!�8V��^[�
�ײ$��3e�W]Y&iw��_�|�s����e+l%��k�C��c�������{e�	�Q{��ǯ$)���·���B�\z���-"ꔓLog�z��e6�\�k��Ú����=���'s�� ��p<&}�b�e8.�ؘ�u�)hHY�C� JΗf$'��؈��Q&�Jr���-��߃oR/_��y���W�5�F����sĉ:m\�	�/U_ؙ	.����9V0��8D��z.q���7_����4%�W��,���x���Pd��dDfs^�n����h��g��Y��L��*@�krJ���N������X?{+���u��	Q�|�Yε��J7b�o�1Hr����՝(��\�2awC)e�k>Ep�1
�-Z�!yVxh�*
�tW���ت��G��1�)��_z���~2'y9���Y�or�3���\|_�J �`�=c��й��@��x�4zG�XOG*!��G��H}a�~DX�1:�y� [%���E�Bt�np�C$�i�[���i��_��I��VNU����eJ�Mrm�g���1H ��oJ�9u���7/?}P�-�d0k}�M,���S�2�'��?��h���ɲ�����tF\���4���AV!:3�ۻ��+J�����3>��j-�'~�8�d�����w��t�q��������cR��No�;�?Awn�s���)eh�7���q�E'���L��r6{���)]�k��.T�&�9]((�mX4m1����瑘��}3ݶ+�G�~��؏��i-k%��"�����9�,���-ᰔ;/�>2�f[/��𽣘�,��\q>|�[A��Ǝ�~{La�r���/ԋr�4o
�����z�	r�� ~�݋�AR��8��u%@f����=�\����,����*m�!~Y�p���טU�vUlK��-�A|��Ex_�7#�`�����N�2����E�:���y�0bSf�R0���t�| ��dQ\Z0����F��;�M�u�	/����$���l��p�d��:Oh����pӿA\�jy�/Hn���p��f��Mk�5��$��� �N&�f�u� #M��`}���zPd� ������NsW|��&ǯ���Ͷ�&r�
5"�x�q�m�u�%ј��tu�����O��Du�� �(�j����P�0L��"�2c$�Ů
�A�j�� ���� n��X��ȅ��"��j�'����J�ezB����m���(��)H̃���K�w�� ��뻗0�ws�љ-$I� cD��AWKx���`Wggb+~�<�2.^=C&X�CW/G|��R1�p�![+�6�]�s��,�Z,�s/y ���ƾZ>w����[��3h����_C;�#�}W��u�Β�]�hB=[#�"Y�9�Gn��*��?&ܗ��I=��aBC�m�.��]�`�	��ڎ0Z����� r ��V!���_�
[V@�j�,�`\ڷ�=��>�Jk�R��c����c�1�ܽ��KmR~�L(HC�ta3�R��7�	��R�f?К�v_����Z5�Ŷ���5�����]l�8��T����'�1�x�Al��p\�&K���|��!��S������v�f�h����;�LJ�E	٩
���gyߤ��O�u%���]k�G-�8���Go�kM���c�����|�DʌW�ܸ�}L� �i����C�ՃS�-��c�@�kd�c�?A�v��� ���TÕ����f~�ó�y�WT�(ak??��ĵ����t�K�.�8hFF�s�5Hd(�����e�ҙ}w�Z�����&|����}S�޶��=�Do�(,�z�-{51����&�Z��ګ�IJ�p�[�6���u�2�f2n�i�G�I���j~%[�G���(������_������b�K,�U��Ƭ�"4��?�	v5�a滅�2=���Ǖ�����'5醿�
B��h�X[W����"����X6���E���5�<(����s�|S,3g�c��n,&����F��z����x�t�D���Ц�H������Q\�IFs9���_�K9�(��?�wM��h�s+{A�P���*׻���`��y#���َ�-�$�{�+�iZY�^���~���F/��I���3z[ڠ�l���}Vjz-k;���g�-��;��b5$�sˢ��G���i�t]꺵��ab���lo�����S%@b�;�]WX/N���_ E�\�Fw����Tw����LƋ4]p,��b��mCCgJ���8)X�j���a�[�4n��^dE�[���2�a��L��d�̼�+��I�%�l�"��"$�{GgO{\:��0T��,Zr~��L?�{�ɵ��z��Ԟ[�^������zw;bù�d��g�ڲIzY�A�K�YTg4#!77����4�Z@�v]�?�aZ#if}1��z��(�xeloI5U�F[J��j����҆2�&q=��L݉���0Ap)kъ�L[k�s�3ؼ�����^�o[����em���haB	1Q�4�!��z/���Qn��#�P�t���LJ%-�5i[X�:D�cw��&��p6}Q�\��׭�ͻ\�R���{�	{���,��"�y�ۆ��;Xzv:�g%�p�/�G��NuW6�����N�8���ž���#�ܟk8f�-N�+[S����CPN�7G�q�φ��|� ��v����#4����bٸ�`�E��ʽ�N<]�	>�M'*��(�j�3�D7M�C�O�jz/ 9�D�*d����|�W��q"���_�{���:ca]�[NJML�2�Q��PU�Ю�N�K�O�.ǁ6���8ss�
���QB	�-Q�`鲙�]�#R+���?7�/$������Vt\; Z�3�N���}Mi(i��\����Zh����
��O����n����1�p���i��jx�h����!�T1���s�������G��5�����[�Ժn�۝0�y͛�U��-��y?7��q��� OB+/�p��砿�R[�w� ��>\(�}%H����9�W�9�ֵK¼�x�JD�b�,!Pu���lx1��ΌƋ��7�3qsPv@��d㞪�=��]띎�3��9�/�[ ��X��9-֞��ܭ�V�ɢ+���D��� ̢��_]S��� �X_��7�,��Z����@!����,�]��kcP}�u��v���0aTP��q@�:E��	N^nl�=4�o�i���R����ʧ��jN��Ŗ��Y��٨�v/�IOm�����T�>Dlfa17ʵBm��1�~m��7,z$�<�	��Ol�5�eė�Ë<�5v����F(/�~r5{� ϒ���Q���[H:`�USn2l�p�]���Ds1��l�I,.D�.�V�� ����2��h�ʫ	��=`���
�$HW��{�Y�a�R�6��H��`�I�W�=}�����%��_����w"!ח�d�5�! ��5=�D06'Ui	7��>q*�R�%&~�����F6����	�brQe�Ќ�OU�R��cQ�(y�֐�Mm9��Q|��۲fS��o��Q:�J#�vP�[~��M�Ţ"v����xz���}��<0ԍct�E2ܸ����dR�����|2�gٗ!����b�Y�A�V�|�\�
d��`Z㷸�*9��@�~�q���DlH��
\�{'�v�64���k}LH4ۢ�S��7'z�S�I�WG�C�?���4�y�g��k�/r��)�����T9�6�U^�C��~M�iM/�=ټ#��T�l���QC��b��^��Ҽ=�xd,��-�� G?�/28�ڨm^���@��J��n�t9� Æ�f��k���� <a�������E?7���9&��v��#�5~A���f�T�.�Ą�#CY�����z�����as
�l���w�"Q�LΣ�(;�Q=� %���I~�|��o��)xE�՗g1M�]�.�u^�Vˈ�2q9�d�D��	��o�)�8��?��2Ptd�U5$?ǀ�@���h�?�t��h>j��q_���V��@�'�!G��k<���Q�E���H�0ory?��ȵ��G~1p�<4�uĂ��a�)צ���^��D���������LShqS�a�� �n<_Jm��v��]�->줁O��=����1@���P�������ӡ'��)�m$/mǬ��g��������<�[��b��\H�]�W�9�h�F�R��t���_ӭ1����b@u?�*��PS!S[��
֚l����n�L�P2��ќ�i��^X!�N@ g*uHG�U>@>��AV{7���8tu';�C9ͦR=|�&EA���T�:9F�f`��#�ا���@w2���ٷ�h��r�
΂/ �n�Ş�[�"�w�/rE��C1�s7RJPw/���G���T슭����ȫ^3ه����R�|цp���o�E(Az�+��1W0`����Ꮼn����L ���O*ͥM��X�&��\���b͂Z7���p����.�F�? ���I�6���N'��B	&��Ton+|���'�%��g*�������X~g��Ʃ�iĐ|"a8]����*>��|����_���HN�������Dj�f҄$�����v*����B�z(�L�s�r����r.L�.�� �c{q�)@y�%4���s0W�"d['���􈮠dI�1�:ؗ1�zM,�<�K�+�Y-��X�J���N����K#�������$H�Ӽ\��G[y_�o����S��x:�i�U�g���M# �e�.Z<�	��W��}(�!�
8T����I���8kO��0��S�z�%Kw�����Ń���@�� >x�H�mq�1��_ӥћ�;������W`Ϯ� xށd9��2P�:�r��ɽK6�<C��6�Z��+�!u���Jg���|=$<2�X���Ǐ�v�Π�lj:h�̸D��i�#f�֔[�����iX�l��&�j�/[�
�'b��qu��w�<�PS)�۲��&^1�#���<�
�q	�����瓬���m�r��p�*>�-�`���` �}�{$��y2��>���~�/��{T�Jm��i �b�	~;��9�	�g��r0�;��u�Z��Ҳ`�ҟ���WGq.Op��S�l^w�]a%�����I����G�z�夡Ϋ�H�+���4�XYHm�ev�Ŀ��U�I8٣���@���Me��G��P(�r�F�i<��(F�+~t4�}���vܕQ���)"7���
��d�)��я��h�u����'n�d5�ܲ�y	�X���:Œd�uEӤT�O^��-���@�B�a{e�(�[C ����J7*�x�*'x~���p���Sc�V_��2Ok����lxq7S�Z�j�8�l�l�W@��M��iuKd�L�u}���ʨZ7�W	7�Z����R��>�^F�	m�G��Tk�@<Q��z�EXT"�!{'�\����js�xmC�������,�dz}�}����v�0y-�+fgA�B�B�%��l��d�m�^_z�s�@���co�~^9�_D�4Ľ%�c5����6鑩O�3l�:��?�}C�um l���W���Ԡ�^���ւL]g�d/K	��@*-d	��-1t��<4y��F�Or`��E[�)����2Wp�t�2HםI��>L,m����P
W{S;�c�Z��ݖ�1��ct��¥���.-n���?�;���y<Ko%�<��3�pdPh@�Ӫ�P4�������^\H�7o�&�5'X���v���7�-����=YO)�sٱ?�Q>��f.�1y�4�
JD�e��?wL�Z�8Bb
�͋BoȾ'Y�-|f����=���G$���>���
���x3:j��iU&���Z�&!�	)������U7��&"crƠ2�s)&��i�
[Z��ʍ���j��KG)�sq��vEtFs�I�tH��p��_��	��}��s3d[Jri,M�Ϝ%��['���`��e��!�����Լ��x�C�խ��ws݅�ٛTm���
���J����
Ҽy�����/���fe�M$���f�>� ���P�'�!�T�/1_�}>�ƺ�[�,�!�SA��MdS��!51B#���$���.��uM�Z�R�p�R�h�8�Thg�2��Ş����*3��]Y�?��"6���ׅRyT���z��`aU��{T`Q��$ǼWMjX�Z��1Ĥ=�MR�I��b��h`]�=H��D��S��q�`��tw�����C�r�g2���8�|��)[|��d>����ӟ�.[4C����I�l�:����(M]<���繐z3�O�;�)S�c�-��J��1*91ńpc��1�|�T,����˝%LQ��3� ��N�6��}�Wƃ_#�j	�HHւsFš�@
|G�ޞ�ԹE�>�R�?��Xٰq�F�6	�B�&�^��<W���w���0�JO��C��-'�d ��6�������ړ%�C��r@#��̿|����04V;i2~���C�+� �{[��;d�ҟa��K��2�5����kG������T�w��N��� �D�x'����y���F^Pv	Cpit6�p���Q1I�d�:�dhv�;A:�|�6bJKa��̈�E=��+�O�R�Ϡ����u"��..�"2��������.�Ѷ�Ejߌm��9_�jA��w��H��Z�}&�L�:�#���~VTz����*�%Eb���7��`X���t�W`d����\GWڗ7x�f�/ь�������fxٖS=o�&O��⇋���,��ާ�qnAG�(��(X���^�-�gJV�&Ĝ8^u� -�n;�-����J�-&�Ԝ:;��÷���b��F�����7M�������56o.6D����6�{?���ve���)���	��N�c֜�8	�r�Ef�8���Qb�$�^�M'�3�(�
���]s�l��WG;=ɷ� wA���n��:M6%��@�U����"
өʚ���_6��,�NZ1Y�F�0������ε61BRS𚰮�f4�h�1�D�V� �DI(=�n=��u�_ݡ�fbxh�K&sʉY��_4/y���(�_�F`,�5�w5��d�D���Z$%���o[dl_^���%�T�	����r1���J�NT�mM�5\3�y���L;+�Zm�)���3���41Iu��<��y����N8�y�?}ǀ�媭�Kt�)���ȅ�����k�j�L)Q���⵻��gj���cĩtR+kN�@Y-`8ſ��r�*K@U��IlP�IF�I�H3��r����������w����J��n��¶ǳ��$4]��	�$��²M&,�p�6�w_r1�
w	��
{��?��i.Ʋ�QUh�6f�u
֎�p�@�sH���(�g������Mg�b��ZŜ�#	eM)s�6��)�$pR�Y�N�`	"�����~}�klޭڷߴZ�X�f{,"e��ߖ�*�Dێ	������O�*�\/�#��1���c��%�'JGp�14PBj�lq@o��.|�����Z�ltb��7qը}�\a>-�{�����൛�Ω�[��c�bϮ[�k ��կ]�P��f�#�`�g�OU}�l�-�{W�G+DN��6?Իp�[���^�\͆�dn�iN�ú�9�U:~�&5���6}�i|��%��b�TJ���al�dF���Biz(�n���[��l�c�Z�_�8g�3	�+���./w�d��D�����~�@�ܤ@�;��dUp�il#'h�9��<��dadM�'8r�C��K�g��q����`~!_�b�	d\R,gu:������-¦,���m�SKY�v�9X���/�T�,|�6H��&�*����E�{�,�9�E���tjH�[�*�C�f��?���Z�M�M��ʣ�d�S��6<i���|K�%#�������->�8�9�EW!ɭ�0Q�Cg6@�`��e4B KsD�'�6w�6�Q���n37N�3AuF�|$�����B�c�$����1N���1l0�#֨2��`����4l
����V~M��W�KS`�����%䝕��_�ʟ.p���)E4�q��q�eFUs�S�1!����(����'nBI����e��.����;�/P�V�tz����^Dg��Ռ��c�9��g?���}:�3�:��Niƾޡ��[�/*�/˘o���r�#=�G�� 	{'ˢ��
����z=���vxI��ƨ5�A`N8~�%H�y��F6ה��*�3������U�X�ڊ��BA�5��R� _��p��H���R�׏��� �{���E�D�$m�����_=Q6��``��(D�R�kV�_dK�)O���࡝w4~������kC�e�?��,8A}����% �i�_��W9����p��t�9��v1����+��Dw�_�R\D��X��i�B�֑�)r|"����32��
P���r��)�����7� �K���s�A�vŚ)�o�}Ķ�\�R.��]��n3H���>����Mf;#��aGf��rZ�/+��KJRgw��8S��8s-�0�?�&��7��Y ��� U_��f҈�`ۉ>
�k֭7>n:����%h����00���炀���aX�1 ��XD�������1N�V�M�b�}ᩧ� 4+X�1+�G�B��ܖ3,z���p�1&\�!����m`�!�&`�1�H�z@Q��_S�Uyȹ�Y������>q��&�ف$o��9~J�}ZZF�:)g!2�yLu�k)Bb�I{+� eϫB�N���+,
A��t�s��(�U�"����X�B�_�<�,�m]�^%�B�� � �#�������m*������/c����h0&��y_#��A�y�o��t�7�n��o���Yn2bC��V�o�ȉ�1�;i���]�S8œ��9휞P��=�p�&b��������^��r��/*'ݎ�E�����I�?x���8%+x𷐊�]K��$��N�:����:�-�ر_�z�t�G^i�,Fw�+�{1�[�!1~�F���5��CF;�)�����@7iz���iBD�bW�7�W=�{�v�����+.����XR����[���5\�8ɓ<�bm��i�a"�)N�LAW�2ү�1,�`խ4��!�Ž��~/����oY�$eW���/Һ�>{�@�˴�X�.�{'q����E^h
��)⊻nX��� ्�{�4��QZ�F��1淋�Z����[b
,�����̯��3t�Pc�H9j�o�"�W��	�0�K�|QM�b9 ���L"L� ��V���4�i��Yx�����7*��eh��=u)������z�����i��pj��X��Lo���p���Ф?��>4�9h�4�C �S6X>|�¤��y��~m>����9<܁i4�h�_g��+��(o�#���g'LVƨ�/A���Uކ�8\zrn�����ſndz{΢4��n�p2����"�[~#�LϮ���_� Un�^}�4����+�E�mZ���|���6o�̉�s~]�(�c��׻(�U�;�X.�����#�{�QWUcc�w��W�����Ĳ�	�9�LK�H\�DɂyKh��G��G�`!l>��)�AP���%n�O�w84��
񶖠�UY�F>�Z�OB߃�X��Ƀfo����7ê��DՈ18�j��Qt�d�d�� V>���P���pͯ�M��V�g9����b�T�oK�akGh*�/��N2���3�W��҃'S�X�H�  � 
f�-SA�'ʪ���#��^
�H/MF�v�Jҽ��1����CѳV�#{:�a��V��V|f�8�V����aȏ蟞Twu�Pt�'C}\^������*�-Cǰ
��%������g+o:�T_c-w�vL#\:0�5����yN:�,�s7�<�R��Di��Ve,���0�'���w�dG�"��A���-c�c���I$�Ac�j�:�!�CV�!ک�e/��
��?���jWw���o[_�'v��C��X���7�r D�՘ GO���n&1�;��6�w�25T>�=ʨ�f)�f�k	$3��������n�WZ�o�_}����8����D������O���.���v̅����=P�&4�դ��!,Fm���r���[ms��$\@����{�$-����;�P�D���n���;�pV���L�?v u�}�M�� ���|�l�h��Ɋ�$�&Ρ���"�``�T��q�r7�U��z..0� 0$4��P	c nO�ɹf���7�p�ijx�N�_\�odX�o �?k=�e)���£ټtئmi�%��ߌ	��]�!=!�C���r�al����]�{�ɧ�Ȅ.X�� �ny�m4�jT"O7��}$<2sA��	>@�˼�%��+�q�i��dNewߣ��_$���<|��ѢW�uR�d��SM�!h���%/�Y���D���c��޲����Z��������-���ۅF"q����AsTs�A��ŀ�&^���#�k<n���1��=�hH��OZ�|��\�}�H��Q
<i����^�)�L�/����o���p@��#s�ϭ�޲�#�~G���CA�9C�\���PL�[!�Z��B��R��I�<������n��#����}�ܚ	(�CP�<��qk}����5?�)D�d�T� ���NS3�G��%w8C�7�ϝ+�m�iQW-"��uf�+��n�Y�g?x��i���!��EM�Ʈ�^]���+�
�C4��0l"#I�Οvh���[��/b��X��%�9��Zu��pק��#���a,�\�d����˒�lR��%�3��4��p��uԯ�(��4\�:�0
|2hpG>�v�<��ݸ����`ѢQ̕2��q):��}� ]�_��q��p��E$?j�7��Z�A7O�V���!H﹯w�L竪�H�y�x����^��y��8K�������i/b����'Z��=F��i�5U{�P$�����k]h��6hj��a�VJ�! Bp=B�ä+!�A>mOz8�Q��F�A�<�n����$����= ��n������3��и�����atU��N}b9�o������V>ĩ���)���H��������j�8	y%nA	�K��NM"N�7�~��#A$>SL�	�%|�hk���Cu���{�Y��¢�g��:���R�tt���@�.��Q�vB�!*�yHݰ1���['k	uDsE�l�K�$˒P��bV�a��nS
F��+^L�$�]��,Y^���T#���dV�`�HL~\t�=�?_�$�5�L�z�$��E���O�Vh�������
���a�RN�BdD�e&���YY�x_�� ��S��4Пsc�6;ӡ�X�����$�j8O$B>�i:����X�s�j�^�;�iDd�3xK��ڙQTӔ��JV������SoMVY��2��Ї��Q_6CFˢ!冲�ۄ�U[/�rݮj���3���������$�%ڴ&�0t���1�����~E���UMR����(��Vp�r뷛-�w� �j�Ha�Ll��10��Ch�H�Ǵʴ.���u�{�G�:���Z�����q�����p�R��f��r�M�m1�HAw�b=�3�u�`<�B�YG@*K.B����Y(� ���Q�AÖF<R�U�bm���lc$�̵S��[�����/̜��T�St#�
�����T~F��b������7|��F��E.P�{�-k`��V޶���"��	?=tcmI��Wf�9$uD�fc$m�E�h���[Pn�!�PPJ�B��ͭC���8���b9�u�O�g�=�8����^.mJ
c���3��``��@���#�Zs��-�p�]?�äO?�.��5��g�4�����7}C{�(P�G��6��IӐV��׌E�bځ�z�CY�k6 �p�M�!�ŋ$��� �~K��N��A��]MD/ɼ�/�Ƹ��y��H4w���ꡗ6�w�`W0�'C�H��#k�j�DŰ���5�� *�m��(�����C������a�v�;�0���7И
K���K��4���} [?Dy�b����������.�:d��{)�zi�2`��w`�(ٲ��Gݔ�;�(���v�<0�%��~��ѓA� 0�'Rpv4\}�,� M�+J-�/iHwu�9�l�������u2�)�#�W��$����d��n��ݛ�]�FXs���+{�.���b��%��/?�雥E�n��}�c
���Uͦ�������e�=���J6,��:�nDRR�f^��h@�!C�s�j0���B���C�">9)5�<��i���!�#��W����ml�+q�"D�ٝ��fFSI�v��-��^wֳKS��~oe����6_�Z1Lf5^D���C�Z��^�W�K��ʇ�W.q�Ҧw���8������&�`вL��f�oOҝ���N�Z{��������L�hN�xՋ"�_��Дb�)n�N ��/ȹf�����~�aG��0ł�r����k���=���)͸\A4ZQ������	���e^����[�lu��d�0?,Cj4�6l������Q*����jD�ͪ)�$��:�^Z��0����6�VP�؂��"rg:>_n��좆K��h"�I��X��)6[o��z���O�i�Ƽ��'Cy�y����6�}�x@A@�Խ,���D�qF8���	�u�}c*zI�Q��EvC��c��#N�~��m���;�+1	�{�]�E�D(�_��;��RیB�]k������@��(FaB�@O����a ��ɱ�y�V>�S"�c�|i@E����9�k�gh�Aے�_t�P�`q�A�	#aGR�/�=:�_�+/lP�����?E�W;ZY��x�슭����Yq�s��Egvޢ^�fX�\�D�Z�ض!%�]��%Axf�`��e�B֭3ܠ�	º>H���V�}����B�G��XI�d����0��?�SH��.��8���i�{�B��)���﷉������Z? &�t�E�"�Wq:�N��4\A�i�Ve2�f��y�u��>y��0)�,[��z=&ꥸ�#^�0��{?'���	6[�U��ʔ.�4V�ۛ����4hPxo�Ū}T���=���VG�*o���FmEl2���Hߤ����M�E`��g�R�B\�B��₪l|z��e/����A%��2�듮�hv�6_�@�T%�,��l��ӇGB �/�?!�$[19�v�GkH_K�[R���J�[�Jy�i'����2 �������bl7W�[�}�V/:���e�D�ߺ8��yu�Fֽ�&���.��H"L[_��\*X��8+��KV�(	��B���~³A��d9��8$mM��bD����O1@��*�a>�kBV�^"�'������x݄s���]�΅���^,����`����h��$�`B�4&���!HW�M]�N% o���n�9M��].J��~$`�T�?D���Eʍ,3�H���멆B6�ԓH�г0Go6�kJ����`76ܢ�L��L�<Y��g�t�����p�3��zT"7m� ���2�5�i�C��0��)�5e2i��؎�������A��8�J<�����ƿ���w����!�*�cT�A8
prk~��8/�����R�B ۆ������>ȹMO�d&�8���U��]��
e��S��Ɏ;w�!�z�rv����85���S:٨D�H�<�K`t��U��j��\�sr��a3v�q�N2��#ÐR�筊 �^��}�/�m���>�������.N.���9�1HtLJw%g����O/������"Vʰ?{X��WMW�IB�B���Y{dkH�\������9I6!�VEb.����!j��$���_����Gʃ�a�x���P�ѳ'\փ�.Z�
&�(
�D -�RUa�?a���k!N���s�M2�?�γz�U����xp(��{��kX�M۬!j�G����/0�*)J���Dq3��,�x��bv�_�`�D�`��^��g2�l1ER�����YkIA�^3:��Nb�|�(��Q�{*~~@/����S5�!Ģ�䰊�32prf��|��2$�ɼϊ��*6�F�b�cS�/%O�*2���<&GM,s�0>���ޚ�Pn
 k�v���YK�,�0�HؗCQ�����5A^�1��ZdX�e�1�xf7bi��qz��AZ�B��&�D�K�Y�� $���H����*��@��J��a*���ࡶ'@��hA���A������\Ұ.����*C6����V�@C��CEC�J�Ɗ��TP�,�9U���,�l���"��G�tAN�-��]�ȝ}>"'���?�
�7��P'|�C�^)�*ҥ���^�0�F�oW��e_{y�ؽ�c�H�?��#V���@����rv�a�4���K���v\��]d��˸ M�7��\��s�ӧ��ku�EW�~�
~W�V�w���nE`@Z�j�|���[OT�����6�yh1�mc��7Ap�KY,qZx*.�FӐ�肳�"g�>�V%fI쾱Q���!���r�R�~�n�;�^���,�R?d)�qTg� Z�E|Ee}Q�ќJ;��`s�$.�A��-j~.τ�椫�1e	��꿆U���`������wS+vw�-F��w�c !��7�Y]3R\B�=%ݦ،�Ӗ�*�5ݙ�վ��gDy��-��i`���
y� �nSf��-�Tn�L�}���c��D[��E��.j�my'c��f4X�;����T�\&\Zy!�R|d�m��?3E�7��<�d�����1��ca<#&Jf4&6�21���������ϋ�R8�C�U���fq���5��g5�ߑJ�zW3=�Z-:���X��{����tG��?� C0��|�J������P��)�'1�a��]Yl�{�M^0�S���bM+�H��-��c�GL�h�RKa%xp�.0 *�5p^_KR�	�P� �lI��$��c�G.P�!�m\b=��%z��dl�4�����T����7�u3ߊ�(�/�&a��'D�?C�'��	@V�O3�f����Z��'�����)�6��r�dΡ"��	rq���ByH���ߞʛ�E˫}��6y�RA�5\�̚�������!�*c����(x�U'��m}�F}��ݩ�Q��8E�V�Q� 5N�k6�uay���A]���I�nRm� i�O�Ag����;��@N\y>c*1I��Ҿ|�{z-d޾ҟ�z�]2D��yЁ�ĩt@x��Yj�ȿ�O���.�&k�Г �weiT7�;#�ld;���cQ��#�n���|ݒ��z�6w����Mz�F��n�m' ��_�k����ۓ�Fz�r9e]!u���L��`U��c�b�Q��k��V�=���l�VK�t�Erg� RۼhG	{�eʆ��3��;�����ȎZܺ����Z���+z�=-F��oA{������|%���s�ŖW��KOJq�!���rƐm�������f��s��׹�V�����b�mu�~��wE{�9}��O��	x�6T�)8h�ꖳ?�0�ip�n�ֶ$��U�}}���_�I9�Yt��A��M��F��+,CF"Ǚ~�r(�ر�47ոx�T��t�NV�e)�� ����G!tO�u{[�|��=�}��ex��)Gtˢ ������*R��q�p{F�g�������7�������a�����b��4�
��]��v;�]���d���r7�����j��s�ʌ�CyI�u%�K2l�T�"n�����P!���y�@2<r��Ӯ)���,Qr�'���y#�c�p�q�>�vS��E
iJ�(�?�̠M��X�h8��pe\ԥX���xF+<�4����+L"�y��t�N�Ӭd$�R��a�7b 5ͥ��t�+j�Q��$'�R<�9i!,��^p ��+�mm��@�6��F��dI3c�#O���x��\�B�&WJ�Ѳ�v�7���(o��!��d���B!$��{���"=3ue�J��g2�ϵ�-���x��e��]�n� �r*�y5��K�<І��t"R5��~���z1HS���wϩ_RMF@y$2-�@�Z#���)~m�DsNR�Y-�ӡV�'ڕ�M�
�^�2��GN�g ����=_�/��	z��x@�C`r}�%��	t@��^i�������Hx*^��I�N����T�_\�3���px� ��|��=��eb�;?'���3�-"��w��C_V{3Ii^7�]޼<wxy�Ʀ�;3��l�ȥ�:��]�VB��1�� vƑ��5p��ҵ�Q5JDF^-�֪+#WtE�M�90f�����xpF�,��f�D=�Y�\'�]W+�yc���{l(�;C��ߜ�1򛰱3��
�iVSxb_���!�B�;�Y�`U��ĺ�[���;o��배���;�̓鳯��ܟ� �nc{٭Y|�,��La