��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��/��Q�w���a5P��B�~�/�'̙���S{���^�qѝz��'�hřD~dVr�F�!5�=��[�\�bYzy��d�(5���*������j M����J����Cw&�u����Dg��>_�,��o��3�9=]�sn��5���A<�-��Y�,���AU�G���̻N�	�Ϩ�g�ϵ�w�Ω�k���R�9HO�o�u�(v�W�T�yVL �q^�Q�0/�����)1�cڵ�E
�W�D�t/�Ș���~x��R�X7�]0|��?ͭ�m׭��e��%\rN���H�i��8A(_�P��0];�ű
�0X�����&�Մ�"<I�L`���`�����:��������ߣ��4�!U'��|�R�F��L�	�|�tW�S&��	�p��%H~7��;P[�u㲥JSiu�t�>:�j {M��KK��O�l^��;��O���������'�B���@�XM�m%�ڄ�x��V/+���0���l��ZQ����N(�s�N��/ǧ�_�����H?��2�{��]x���=�I�9�@�H:��zY�����}�ݒa�$��.��9��Υ�Ĳ�N��$ݣ/ڡWR���D�q����	�qV�WQA�@D�tE��啸&X��X�a��i"�h��V���iO� �li���BvG�A-����Mv���4D�ʴm��}f��m9 t�p�ϙB���y��+LWϑ���%����%m4}�L�vڽ�b_'�|�AI�c:La��k��n&zÏt)�y���C��g=��MB��<?�n���3����:���6��W'�-�����0�(��tT�FLo����L���B�`����A�Y.*n�f$%hzU�����ս�r�������QqUJa��Oح��j�Ff��$Uϵ!��oQ[l�ѡ&h9.����~v�L_������d�>��}����zv�u���D�����$b�J�'����>���.K���m�x�S �i\nP����P���������I�}�D�����$��@�c��� �X��4@����Cw�{^���6��9��z!!���^:��a�L�^�����2�����N�@������ /\�8*˖FYTK���&Y0�^/K�ӻ�e ˴�V��n�=��������C�;o�<��p� ��
�V��#.����A&��!�����h�@쮶�(71�ti줆��+4V���l�:7��?�<b�Dm���1��H0^�@%K�  C�%E��9���{	����:�@9P���Y��s�.|LG+KIߪPŕK���z�ha'�a�|�$_}��딬-&(�U
���'���4.D`�m��	���lY�,1o�!V������~�0���ͪV�Ns�����J��`��o���h�B��Q�v����H5�,�9�*�.���ᅓ�[�W'�,4���V����p1h|���4�����k	?j[0�O�j%�U���<�,S�[�(�"���VO�PP7P���;��|׊F������xK��% h�VK7���0�d`��+f�L������S�����>x�h%�\���fdق7��ר�J�_9�Qؖ���Ʉ�z6�$	���g`ҫ���3|	��<�P3�<��4zkw�f�DO�W�����b��j��T���x�m3��A�e��_�4�enC#t̜d��t�Zs��hI*W�Ii"5������U�������'�V�zKin�(�K��he�)��D�u�=�� �9u��E*��zHu��p��kq!d4k��3��ef��2	&ʠ'* ��?S�������Ң���~|��Ŀ�������G.�!��՝�z�Z� �:���z7��z`.x�"��N	 F�̨�k+e
:C�8�S�'�v�V�Y���v�XF�"3�}���7
��eÅR 1���k�]��s���~��h�׉�^�R��7gj+�.���ԥ�mQ:��
}!UъC��'��M�.��ļ-3P�tR��>��� a�#Q��0�|��^��_��.�k����ю���@+wm�r���|W�˱FͯӇ��u��(�D@�Ws��1&A�F�3���\U���ƣq�g�?�����/��r����8����bK��ݴ��8��Q�u���ײ�^0ţ�#��j�&�3%�v3u�P�:��ڹ��yH�yW���e���Z�uSJ�-*.u�#��wٶ<�5c�$Dg���j�x�x�r-�P�S� ����\��~}�s
<�I݄T��Ca��P���3��١+���2��%�=��|l�O��?�Q��C��1N�U=�O�*�&��5Dm�o�ĹtQ<�����	bkc�o�����('�p�O�Pu:�G�Ѭ�d�~�g0'�����s���Y׍x�L50kG��md�����m$R;^�ק,�
�:���mB��U�c��RR׉՚_�뇡��?�D2%^�X�c�%��B{��S�ױI?�)Oj/"�N�8���qL�g��E��
�m5]�vk5Ma7:7�
*+�Fأ�9���֧���;.���ŲbCZ@жW
j'������S�8�]���W�ײ��G
G�c�� �D���46��� 4��,����-����g[�|ymhƆ�d$P���� ���'U^3oҌ��δtUL���#�{��Ю�JXh��K:E���V��dJ��A޼S_䇎omĀ4G��9�B%�[_I9oh5i<Ĭd�ҟ����7棡���u�~�\�b�w�,��Y��=t1`<� "i���x�	"1�<�l���Sp,%ْv��O�,���'�kT�LŬ��ASi-� ��&�xN5e��<������h9���8J�K¤�6�����[/��-��Vٜ5$����Z ;���а��/z5� ���̖0�0�@�aΑf�!9b�X��'�B����g�敗وÈ�#;lR	��oy�R�`�$2{��,���uMy0��T��|d���x�
r�i*�zdgJ�&�aQ���%N�S���V�c�7���^�.���K�*z��h;LJ��k��\�d����l�P�jm�?�:�߅D~C��%���4���q gq�:'���lA���Qv��_V�:�&4������2bxU9.��9�d�}O�#�x��h��YN�����NǪ��AZA��C%�{�=����󅊂S8.V]a2����Bx� �QA}lm��䶼S ���X��ֶ*jO�I8Lt����^��O�x��m�gǐ\��jr:��X{���9��ݸ��SL���!o���#]�R�+�B�.h�5�{��5���ڣ��&��W~����R���U�!�0k�ZT4��!�v~�c�QMζ�eH
�Ú��$L,����7��[�T: s֮��%�E���_���&&��
�PQ/j��u0��a2��mC�Oy��D�Z�<�M^.��B�$9��eU�#M� {p��Ƭ5�����h5ɢ������vQF� A���8�?��d�����BV:��X��n�!2+:� F��o3*7(9,EM�I��x�����l),�pX��w���A�(gJ����l`N ����V^�R��K�z��ic�b�ƲR���6!%�����(�H�v0H'�����&�!���:���7z�<"4�:��B"�RL�m{�=ɐ�W#�$=�Iڶ� ����x�Jߊ��+e,	����c����!�Y���e�~AٝH;&�PS�&�N-9���|�4�A���y���aSn������&��M��^��
�/qW�N�A��qG���*��7!(d��p��A�7k���EC�i݉?4Yxv���{k�]v��Ev�!-]%��MEw]p��
��e�QжR��Ҽ��#�͕�c{ݛ$�D�tx}Ӆ���đC<��d���^0%�E`��_�v�U���4��I����ҏ.Z* �nK� ��U���=�tG�a����i,	������{��D�]_.R���ږ�Z��G)30��м��=�p���o�#��ȣ��TpDW�8���j~R�6��^�^4!�O\b�T��>Ԫ
@|ZY��}��`G��^���>�dŬ��7@h~�J%G�q3������,������Mي����i���ߦʗl�Lg*�uӼ���,Ol���T��AT��
�T'�%�l>,Q�S�P�?бdUĹg�]D�lNW��������Ho|F��4��+s����mp�X6\�a�\/���9�}�TΑ�{�� �=Rյ55a~尜�ִ�5z5.�"�0aهZ�����E��<
�h�6���E(3��K�x�	�d���dQ�O�������A��a1� � ���W�8M�(`"����J�pŤs�vZ�޲�[��BLor���h2��d)b9�)�ݫ���MO�З����k�[e�	���	��1����Z����8����k�H']1��%�9�=NH�>�n���v)U���I�K��e�����UMR�?���$��vU� ����X�6�'�%[Ε}r[7:���q����(���'Ŷd�J�;�yˆ�%h�������s���*��W
rۍi�֖ ,�b�B�;f!8d`�v��U�緲8^�vU�6�N?���X�<�O�����X�&�.���
+ru�զM�2���`�`��K@a�ھ��n���8�0������5�.7����J�BaAe2�f�|����sa?�XtW�T/P�/5�ꨏ�y> ��%jv�yf���%]?V�3(�ɷe~9-0��H0�7�bu�Ii��O̞A�C#�a�<ly��h�.N�J�P2R6IX�?�:&0١�����Ϋ�='��p�������Z��g8n>�/��lZ���L,��e�$ۢw�?6h�8Ǳn+ڎ�P��Nv��t�\g�Ū��q�6+���rT��,_���+���]S,�Q{7�'K�Ěr�Z��!:�uBla�R�,GuL���
�2gF8;�� e�Y���d�<�S4[�+�|
g�J���H��>
��p�V�pB���ɔC�is'�k���$Z <e�^��؆��@�-�N|�� �������:�4ht(����D���a��{�$�œ	��n�������3�K�V��8�p�̵Yn�
�Fp:"sw�Y�Q���g]���FͰr�-`Ŗ�Վ��/%�m�7��黏_j�^9�Dn�8ֈ~���ħ~���r!�IwtKDY�c�7���&o�#��җ�����C�n#�-��5�{��J��#�A^ul����o�pk�Ӥ��W������ِ���'��0TK$�wت�Ƙ��%Ԟ������v�I����|C��;S4�"�����:P��g+FXj��m�`\b�}b��
��Ͱ�HR�9e�E"��M�v+� ��ǿ]--2g2�W��D��}~�R�kl���!m�����S�x����@�VV�y,}����b����ů|aϝ-x��o�\�;d�<A�4e�3����hr6��}x�!ʂo~�s}�:�?����c��J_�{ΐ�d6�^�Q�x��q�I�cΙ�2f�C�zTH
5[�-N�"�X�����0���T4ܳ�Quͯ,5��i���j]�B����t5B&�n�z�$2�0��H"��P2������^��s��O ���o���ìw�ݛ"7*��0J����&�j�����e��w��!=Q��}'���A��j_Z^�*����e�Rc�"�&J�o��^�æ���q���,5�l�蟌E�\M���&*����l�l�x��6���v{�]�������Ve��`F�*}�p&���_�bl�Drn:�{\bg�l\�PG:�4��%�(�N��p�>�_�H�_��b�| �Q�_\��ԒEӷ�
&5�Ѵ�([�8vӬ��?�q���E֎>B�%x�>��s��+�A�CV�ᵸ�N"�ڠk�=F���q�M���z9H"0R_K��8�b�����Au�<� 'u5�x���e������0�k�¥�~��Q��ӄ%���Tw`N"�{�'s�������z�Y�� I�aՠyFM�])i�+�1����j(���{���8�G�&.�bc� �l[�"��奮��O���8�d*����2-)�WZ]���u�f�Ac���u��Re7��0�ߧ���
y�����T?8�"�Fjl�RS��.5C�xl�51��}��%&O_3?��Q��*��e�mR�@XKp��׮����Z�;+B��>�/�W�2��H�ճ.64?���WW>g�F2[�wy{��m�j��(�&�k��=t���C6�j�m���5--�@���i��ê?u�㿩���y[b��}���9x�/|�����潹s�h����Q7�r��%��OO�R�!�ffb�&>/��/%�6�Ȏ�I0�bfILD(4�6�tP��3Z�y����Y���n��Hv؊�|-��/�m~�T�� ��:cO#p��E�=J(a��S��s�G��1�������9"��/	��ݜq�z��H��;�k�Y���>�e�ѻz��p㣮I/e
i���~�/��W"u���~չО�?o+k�6S�;�i۝nH�A�:�	.��B�BA�;+�4�0��u�$ �X��{�.b`����$�؏0��� 9�H��wG!��
�V@x#a���N�L�Y}Q7@Za_Դ���sql)f=v��/_E�<VIcTX�Ɇ�z+O�� ��*�~�7|��~w^9�%�����C�]�Sv2B�:d�z�"s=e�Qޘ;|�M)������i�5pE�(L�Et�,�l���L�'p�t�=C�+6G�6����Y<��w-��������6rH ;��ͦD.l���m�����l��[�U�p�1��)Y%?�[d����D��l%���(�4ל{/�;P��F[l��E�-0}�-���s��
k��Ԓ�������Ŧ�z|T���S��}k+�R3b*�x�?����)�|WA�uz!#�X��+u�޷@/m5B�����#]<��~W�|T/���V��*�7-�@����WN`z�,q�T��;��yd�mL�^��	����$�|�>�tL㨳��i���kY�%���l�62�w酗�N�P'��~���d$f2Q��5���	]�x{��O,=�&��
�p�CY J�!�4S��x�9��n�++I����8��O�� ��� H2�t�� ���m��<D�!-�p��&-�m�Hye�a�7rt���,Њ_Z��4�����ra����ţ�5cSR��32'�������&r��f�������E�nhԻK��%WGuo"����{�2�n�M�Ύ�(X(!���ʍ��Bdi������Cg��T�r�:�Ɛq�,�ϡ�#�z/}��,�H�CW7���z�X�>�6�R?YNl���Ƌ$��X�R5d��Q�AE{"7���w����̀b�VW	%^�M�F�\�����j�g�������:lwn��>�@u�F�.[ޞ9xg��M^O	�񅅜�O����X�GGӳ��#S�������*������8��z��^�وk�����$=�%�[#:�$��r9o{�8������d�#��~҆�6�V�-4��D	,���6�$7;�?��G��#���I���a�X�\5\�\��
�t��w�c�(�uNk@�HY� ����i��k���nYu�۟���=T��]���ߘ�r�1�H�%�ގGD'*��Mk��� �6�ڵ��Ne�n)k��X�#�ro��#��+����n���~�Kڲ���9c��g���e�����s���9����֍��Z	����кܦe0>�.w���S�X&�����UH>��w;��a���=5�h@v'OȠ{e���)b�u�A�L���>�"�:h��R�B ��J�Cܫ򜱱�Ia��:��x��2�ľ#=_Y��b�ʃG�����]�j�~��[�~N�R�3�|o88����e�0�V�("�!�N#���%�c�"�͘]>��������3-�r�]�\�C�:�Y�et� #~y��(ħgS����,���7�5(�/�f�6��C��s���J�֩w��H-���U_2GcS��l��)���\^Q%q��K�S�K`v�TR4�D�B{�����l�@=�s���Yу$޽}h��獱R8����Z��p�P E�&Gh�������E2{����8i,;�c��JM�9	�@�ه#导Q
��H9 \�3E�K=��I0�pk�� �������$�?��x�>׬j��Y8�@P���sZ{�2N&#h��޿��0���6����P�c�s�������!�Q�.�opCl��Gh�#����L"g��9���}~/c�c�������,+O<C�^#JҾ0�튆C�a�4��E$9�l԰wV�:$+&8U�?'�)Ǎ��C�O�D0?�u�{x��ؚ�#��5��Fqx�DT����.}!z���:�m���Z��%s��?�?��M�H��͉��B��-����!�˵��ϸ-2YB[n�]o�Q$5�;X�5:�����Y9�Ǯ�i���(w�=�=P\�id�ㆰb�.J�'W�}d|����I�h��?\g�x��7#|�y�Dܿ0w~�6T2�Z�[|,`����������� �<��u�Kq��Ć7�����ndz��T$*=Z#٦��.X�d�g-١:���ǉ�|���y󞜲"��yq�%iE�m�x`����գ����J'��� ��B7�!(�0V 	E|�ڱ���o'�	�r<e�Y�j1��ɸZ��)P����5������׎���P���g�}�o�׌D�^X�LzS�r�o\ �<��E���:��N��By�����[�
3��F�U��)(�%�����ӨѰ��I8�}ַ�-o��5N�(z���:��C�Li�H�0M�5���_���p�'���''��5n*'��+	X*�|��o��q�܄��EA��4J�v��/�ۥkzC���ȱ7П����/$톖?h�?����s��i=��ٜ�߃�#��m0�^�D�*`l*Wcb����U_������L�"�e[��b��b�g��QڊI��ܪ���E��> �O�O��`#���.�����B4�z[�`,%�l�\��/9��DO���d���W�f�,:��df�[�A��W|f>@�d�^�%��9�޴�L4d���F��PR����e�F�����g�h� F<ђ�" �����&o�lC<�n��t���=_�QR�|ޣXy]�%<?ٯD�c-f�\E����Kp�����E���/d�r$�'����Э�)��ٱ�;��s�j�+���p�+[�L��~z�������P eOugXS�_�3�?i�j��7U�A�'�2��׉\�1,���g�3��uj��Y�2�^ēKrD���G����^��Mؙ}�d�T�qs���A���u�e�'d:��&Q�2���3;�w8���p�6L$�I7��#T�M"^�|$�����~uz'��o	��}��~?���w���o�7�IS�A���*	dԮ��5�|7��DB�ԡ,��QA�]�u�)�Gt/��w�Jƃ�>�w�;��L��R;����.�\�$�(' )�	��}�̷��?m�a^*.����-0	YX�ذ���t^�Au�*�����̷��8�L�+��x|$�klq���<`3�`�o�tx�%<W��x��M�y͆���a{w^tb�J\C/��b�NX�\�SP�:圊{ߴ�ƃ%� @�	m#\C�^1n�2��<�X�'Ƞw�X��d�t�H�68@��6L�`]t�+�wF{s��j���VP�s�S���I���Y5�G����t�-;���W���5gpFG�H��iw��U-jE���U���zU���}��Nfw��H�8�#���[Q�邵{�{s�U�_6*9�)[�Bi�,�D���O����PN��Z��m��H��`�*�)r�W���0J3�Sk v&-b&���cl;+��sf���T���^��2�q�,?�]؀��X#$fk�y���ߋ$6 @��a@a�` �@gF�m�I�.��qnP����/ज़����+�"D��)YW�J������f�Ջ�lw�!=T�׉������R�*����mer�S#!�Nw�L�S��^b'�z��K�#^�������t��N�������ͅ�8���İ܁fdv�7���,�.�" ��lG������������w�_'�}��r0�(�i�E��r���Mئ�r�����1�'���J���+�D1H�!��+B�3����Qɻ�!���˅kK�i���Y��#\/�t%֛R���?4�G]��%C��C	�ga�f1�?�77�Ų8��гͨ �'�E�V`�� (ͺ������H��{_��T��)�"�Ȭv9�馟��JQ��e
�j��u>}v�3��I]�2rc`��K�܃ftv�]Ak}|q0����V�%�3Q
�2ļ7��� *MQ#@A2%`�����c�X��#7����+�(�כmC&�������L�>�c��]�62�[���fn�b�;��U'�����q�T_����W�R\�b��K@=�~�\��K6��R��{/�;Ks�O@�O����W�>�ԧ�7��{�v�|���]'�=uY'�B�����E��H�g2���Ȇ�q�5��B���<ӕ�G��~|��}�$`]������=����	�O��A��?P,2@�$[�)^N���J>5�VYeo��� �x�ϲp;���	E��n=-��Ը�%�AwR��ͅ��F=�vt���5x��E����g!���+l6`���s���Z[�q�*�P�J�]n{A9���ê��jYh������	��&J�R�턫ɨވ.
nI�!ޜՍם�X}���ҭAG�������2�0��v�8�NK���3��QwƊBړ����n1Dm�_fH?�].*����\�tCo7���1����bR-gx�ȍ���$pF�{nf?����:�@em�T�:q"8���[�ZɜlCB�"�z6���Yx�eǊ�w�Lk=���FcP"x���}!��1f� ��C�u'��V�&���0IJ
�7H��+����F��S����%�R�Y��[��	#5ɨ�)��W�q�%Q�UH��Z2�T���I��s ROQm~o4L���R*$�}f*�	�������S|��,Dq������o��no
�N�u2�w�6��!��cy�j��s�<���n��ZQ�w�[�O��"S�#���P�,	������}?�"# 9=�w����R�{�ήNB�$v���<2!͂	��L�Ӕ5Ϫ�b=�ܪuJ�Ժr܋���ţ? d��*��|61&ִI��t�S�)�1x�{c���'��o����}��K��/�e<(�[҅�'�ED8n͗.�l�cN/@�2$��'���W3{Z����$������uT�h����A�pL�A-��␐�GZ�������490e�cX.�t�bF��X.���\��2�����LR?�D�`�N Q����mX�a;�����::���d4aJ''v+�������r/2� 9��:�"L=n7)Y2i���ǔ4�	Pc�\�\��z�m��$*)�t�fUկ����.UZD@�B�i�c�X��O�Ei���^��N��+1�7D�P:w���1z�;��m��f1����y`S�ڈj� o��r.	��C��ƽ3=���/`P#+�B>����]gº\����]�*%5��b��T�*g�����Ǵ�x�݅�()�C��W{�XOZ��\$��m��I{zaƀ��S3U#j~Z�N�l�$�f��:_K-���J#�:���Lo�V3�'�1�G"�6�+&�[��x9+��D�x}�m�O��>F���0+"gA����	+��h���7ĖX����̩�����ӌ1��]x�`��4�.K'}+bl�U�9�g��ϣ�wp���ˎ�J"av���K�l>�lM�w�9yڱ���jLB�Qu��U\��3��n;�~�>Kz̩���D�a��~�w9U��3=Q�r{�Ȫ���v�?���#�6e{I~�&��]-��F+B�a����wClQ"*̈́E�M��2F���'j�/�*޳ۡ͹�E� �3_��S�ː�r���ay·�g%̱����i,<�J4�_ ��S�Oq?����4O�{�K.n�D�D�V|��y�.�c�F�&ߺI���k��$�9��C<U޴��|���KZh�q���߳2�a`R�"+���(��ޡ	��?�B<��6��?�@K�c]_�]��"�չ5>�v�waΤ�9a��ȑ�fR)����y��XǬ���� ��7�1�	�C*�y��@'��	[~>�k������{�^5*��ؓ��>���c`�q�[&f\6�^8��o�^�fN�Q��*���V��
R[#"�{Nh�p�s�ٓ@��%$�z����I�+����h���?��Z��n��:�kbf����Y��JaP��������Av&1Ӎ����x�m��y���Hk� ��n���J�j�?6qQ x'�b|ֻ>�1�-%�F� KN�IpI���W�h����t�艜�lu*lW0+�(
SP$��e{''X`�V4���B���Ե%�5�90Br�ȘL��l˧��qC|�*��P,����h��C�9q�+uD������^]�p�gj�6*�v�bl8�X�x��}��Sa�k���T���$���`$\΅�=i��g+m���GZ��<:��+L��SW+�`c�܁�J�z�{=�kԄ0��~_~�wz�mPNq}Ἑ�H~`��@��J���)TE
�C܇�C6e�RE�)�;L�%�����ʐ���0��uq]`������A�&(|QO�QvT��`���A��׹�v�$��Z��8�f�S8�a���w� e�CY��w�">��b3��j�먊t��o�)��&N�����O����60C���r��8��e"��U��{�ߺ�z�l.}��z��5���tU
g�hdӃ&��J,�O�<��ʰ����+i��@<s�\��q7���\,QPt�7@l��>�j�0J�A�9�^B�jX�����]I*�+u[�=V'3n�d���$�s��{Bhʦ3V�F4�),T@�7�|��B���O{%@$��s�b>@�* �#e��{LR~��P$5��_�bʽ#�p|]⏫�V�������=k��˺Is�U.Zs����-�>����`<
<����/�!9W��^���ꓽ�)��U?$��`9�u6@]��k�����
��w;<��/�A�̝�$b�܍}�?R���1����w��O}�~�=���N����Y.9i�	���!��[��B@� ������3=�R����?j�w�]���܀�?J�w'�/��r�s��Q�#�7���IL����&0q�:���Y�4�ތ(b��u�7 �U^F��с@� �e8��@uy,�ؐ0N�#[/}� hD���m!~��tj#)y�_F��O���ܼb����kdr	}����Xc��e�	� �C��hG������ܯ�{d>�^�4��l><�۸x5�b4L���$ndg�^M��1�R������(�p�o�?�������� {XaZ�ǲU�Ե][9!��X9����y������Y=�����kc� �9ZO���E͠ʌJ�@��P|*���`�	�4�2�}��P�OqГ\�'��t�%��7�>��XВ�%�@gU԰�ۆIF��!��_)���؇E�K.o��J�QD[w��(��[�7����]ی:�?�|�u��Ȟ��B8����E2s���[M�5���ۻ��ֽ0�<7���3��h>Ķ*�@�S_6�vm���CKv[ﶩpߍ�"��%՗���
�l��á�+V�e[��.�`ƪs�\0 @���nw��E��ȉu��T���dZr�*I��q��� �!,A�{�����|�e���2a|���:��-,�c�:��IS�c��CS=�����mY�h�We6a9"�n�լTH�g�%xM-����� �:��Q^YwR�`���/=SY��E�����s�F��0q��ޯU#6h���_�����VQ����~������!����y͘��#R��q����z�|Z��!�sc;W���[�#�)M�/ܞNx9���)l�<����R|���^��3�I��l��p��o�Y�����t����bk?֧+�3�v��p�����g��B�F�_����h�E�Y��'ήĎI�h����_�ΈB�m໒_r�a��zH�aLcr��m<X��n:U��b��hG����^
�Ҷ����K${t#���H�/^z�x+^��xe`�`-��V��B�aR�/�CՁt��U���%��i^�z�)F6�]�r��ϵ���kA�z�lYf!��n���w�;�i�����䚕n��ڒYU�ۡ#egy�M� �X"�!N��2}�t"�Hi&C5�r�F��@C�/&�p+�%��:�ŝ,����j2ZȖ]��ދ*:IDm��A�������6�00˝�Ǉpږ/*;a��ӎT?=GvC��o�Xs��}�̑X�*6��b�>�Li��߾{{�M8�MAXu3�>�������dKX��M�REB����GZ����JV �Xaĕ�?��A�9�� �p���gvʧ��.�����qI�o����o�}��_���Z.c|CI
��C<��G�ް���;2��ry�|����A�J�\߶4��$��z���R�%BR�,F�g��y�`�&�Zz^��� KO��q;����37ʂC���i|�N�a�X"�;�]���]!� $���P
���¦<�Λ�c.e��רZ�!̻��9�	bL�нK]�)X�i�,�n�:Ѥ���q 6t�����e�A�	ae�h`�v1K�v���Q�0�WА���=Zg�ΚZ5;�f��^�75��R�3����8ۋ�ׄ�F6��8zI��-��B�t�Ϛ#�D��2��b��c�OI�;ـ��7��F�Fi3!��fU�!L%�;��Q��^T�2G����3۽��lZ����=�m��C?����y�bg��k���[��p�)�$�`�{�'���-1�+w6�oD�*)������Ml$�������L���B��=bc�Dp�*�z1�)v��t����r`�B�m�.�l��ũ�U#g-#[��r���k ~��Ԕ����Z�x�ƂZ�Re���0���[n!�4(�����/`��ˍ�9�m(�u�s�lx��.��|ԕ5�`�&fI2�bJ�G!gyM}�D b�:���e۝�QP���H�&�ƽ7��e�:�F!�b�77�1�j�pI����a68�^u�Σ!��>M( �	���Rm�q&�:�O���E��;�|��E��jA�Y��a6S�Wvi8r�T��=���z���W�s�2C���g(1���x��:�+.^7�����)+�x�ٙ#��I�;������7N����pnn�cd��v���,���@�>��1k�E��g�(����~5D�"��R�oo��ե�ǩ2[tD@7u�c�gjpȅ�,�w�B�j�6��g'+A�)A���U[���o�����e����t�I=~�|��=��~@�l�gڭ�F%���ؗH�}m�e�6�Ed�֏5s��D1��y����	A�5)����L�֣
ǟi�p<R��Գ�r.8�H�uL_��%��Q�A~D�]�9�4|�g�8`H茹�PÓ�tlV9�� ��AV@���2�]L��\�<��~*l�N�3�V��w.ɱÍ��3x�_�N�iz6�ܛU�)T�H��"�Q[M�:� ��K2���^�������4�7;B�T���Y-�L^ܺ�	2���Rs7)��4+f���wR3��_���ϸ�s�p�$ 7��;	v�$�����p����% p޼Aq��B�9�P6莸�dz��㼈m�c2�K�,-:>��j��� �/i��A8�3n�p�5`�M�޽� �4��8dNwLF�_�6d��fDf�z�hX�[�ST��M��*�F�֋o�i�?�Y�����[�����X�2/���E,Y�|xev�r��R�X�~,��Bu7+JJ����V�T)�7�cC��_�`p.�m�/�C����h��8�f[�Up�+z~!��'��Z����U��^�ǌF����5�L�g�0�<�2�@�L�eQ
c�4~�Ňa�;K(�8A"��T�-���Xn��ؿ�Ą��=n�/�0Zkt��9���Ǐx�؋�]�9ޑ�LC��ֈf}�"����:it�f��6g<�s��9G���ST4e�p^��3X����wG��/�Yi�q�֪��h_�/��ۿl}�"i_����B�"��.+�3�0�/��l�$V �i���k]��D\����ͫ �Vu/�����"�>�/�U�.���h;����]92�rľ���]�Y��J����0�H��~����^ɵ_1���?Η|Ұ�ֆ�r^�RD�*��ɾ	S�UR�w����W�	��8��6�S�aנ��8ݤ�gC��oޠ�ܱ�qEi���~�&@�g�WK;Z��R��Y�U�-�./cG6�U���m�oC������*�Q�ϕ���{}я�W�u�ݙ�xV���8�<8�XN��H����oD��*S`�`=r�۳-��ZȖ���hu0�8�Mhئ(��1�
����u�9~n}�y����l?�c�l����.}��٬�3�b�����0a|���|�}JR���	��!����٣�\�j���UM��K<���?�K��X���|F�k��@wݧ O��6�m'k��[ĩ�T�����.Ch�k �_
3-�����B���]�0Ho�7��b��wU�"Q[ѽ�q�= g��y�#�[�/�Z�b2�.
���#R ��?͑�=�KݼW$g��:Li����H�Q1��VM�*��� ݸ��	�9��,(�-�K�;�G��C~a����b�y7�����Z���PR�w��\
x�Yj�i���]�*85>�|$_�^ ���V��a#I���>2�m)G��m�;H�M��,u���@�=S�B���H�W��%>Q�t O���ԗ7G,ּ�^��?!B�';E�0a�D�[���)W]��N�˔�xoR�D�i�>P�f�q���`��%��L�[�TNN{3��,âH}��<1����12X}�������¹�|��i��-;�����H�rO��a�ѡgb��o�-[����!#=����K`�^3s�����D6R�V�L��}G�T�ECe͚��<$z��fFz�]�c~�Ѵi}��پ���?O	Vl���3Gi�ZUlK�jRJ��]�,��q���ĐE^��D��:�a �6�{�Z�}����ms8���5��F��y״��sa��Dعzt���Ť<13 '9�7�����G�s�U�|���ݐVI����a���!#�֞���&$�Z���0���"W1^W��B^;;��K��$�=� ��VZ|�.�D0�붋� x㛒��Ѳb�SBE����_�P���4���l;M��"�b����ɩ$#� ���gP2H{߶�2_[�x�s�Aْ)�� �;��
�,~`�W�=�����(�D�1�d��K8B�ʩ����d]+t���5�Č����j޼��[�YS����?ډ�PJ%��m]wX}�P��s}P����!O=%,��_�����E����¿t:"��h�r��1j�����%=}q����۲����p
0�5��Qj�-�d	0#T2ueA�tS�ve'.ha��ʺ+>��&���n�o���ev�jI�u���� � �a�L
�D���
���Cv�C�G�1�S��_FF3��k������e[6��z>*���@x)p�T �FM���3��#V�j=��KQ�l��2�.�ۧ���-	�͟��8�.�yx�O���+ͭ�Vo��A�=�j���(f5�y���p�\��Ab�C�y�b�̾a&��n�W�_@�&��� ���p>f�J����X|��F�7D��T�ᰐu�5��C��	���kq_��P�R(}��	켽C�p�ZŪ
G~����zpKː�����.6�yy�K(�s�������%���U��������$N^�k�k`z$�3��eU�Ʃ�t���4��j�����<�P�x�,s�@9aM&���;qU�.q�I���_�(��~��oDl�a�0�^e3��k۝	�2:Z�H��9���oW�I�>�۬P�g�=ʀZW�UR��Bt���{;�6��I�z8U��n��t y��(�3SDñU(�;bP���Ueh�4è�m��4l������W]��z��D&�����[�F����;��3`I�+ƃz)����Na�^\���˱d`���9�r��O ��=�,����JXPM�����.>���GR8� ���׭��hhq�"r� y�������d>^$���R�9#�q�N-!��"����(���%��A/L�w�3tQ�:�� 5�Lwn����?�|��`�E���Y��Ω�m=�g1նx�ބ`c �� ��yx���mUգ� �\�����ԭ��`%��h� ���.X���+W)�'yP�x�;��6����lK�s��}pM��k����+{!�פ�����821�̻�����?^J��їW� �C��Ʉ$%��]k`7E���$*�DhT����&9���<�e���z��Y2J��sl���B?Z���цѬ��� Z<�O��9�7����(��O	gyѢ�H@���Y��ُ�6�9"d��`Bj:)מR�����%��;>���`��s}.��Lg�~w\N�q�0I���wN�A��Ȑ٤���s^d֎���d�DI&Fw��E]t"�c�?�?��_^�}�Zt�#V�f"nw�En�c!|���}h$0*��0�8��T�lcLF�-�7�������<�7�B�6�Q>��c���p�_	N$���OL�e>a&�TU�cA�ݎ'����`Ig���@��k#�6T.���
�էzcc����(Z�%g?[�F�@��ƭ�<=������B�kT�'�~%�_����1?*j�n�cR��Q}f3*�^���مt)�S�<�M��r^O(�ȓ%��J������	lЅ�	���=�C>M��PM�aI�I��pS��?�:H+���������W3�p=���!���I�͢�O���>�,������G�c��hC~7j�4 ��ȴ�q7.}O_�6T(G�>?Y^����|+�/T�Z� Il���e5��[5�UX`i؀ �%J�d�d��'V:}Q��_�Q$��脞��F�DB��V��O#��C�z�Ot�� ��BU+��;:��4=�yQ��ˉ,�և3�+X�X[[q�6.��p�AM���u�η�w�]��p(T�w����4�3�����H�O�B�)�Fuf0=���C���OK��+��Q�(��@4�w|��ԙ��-�#�r_�G��
�c{\���ɄAlcz}+�N$��I�ō���k�Ol��C)L�WE1x g��K"�v��0���kH�l���N��n��\�2>|�ֵ�j|p�xР��k(K�|�U|�S�1��4����-�`u�%�4����B�c;��sn�l�G�����2�ԆH�����"�Ȉ��W�,w���(ZH$h��_���=9�Mx�C�9�w��*4�����6*�08r��2?>2�\������!]�_�p����IV3.�R��(.�T�h.uZGɽ@#������1|RM�MJ;e�t�G^ţ��D?��S6���ɥ1$�d�-���V
�HjTRks���x��~_����)Y�@@��;,�Z��]�L}�q�D�$k]�'D��93��Æ%œ�}�^n�Qi���	E��[g�^HW.�@~N6����w�� ��%��3��B"���<F�,�'��st�k�T+��<`$�B-�֮&�ݺE���6ٶ�w;|D+�x�wC�:kc2��8h�����NF`��6�zW�$X9���C��+#�O�;x r���$"�����m��ﶡ�)��f�H��j>GN���k�����,h[����j����8&,��Ջ�K6bۊ��;�X�̍��<`���\�sT���xHvra���Rz*�?��W���
�.�E>��D���� �]8�k�#�2UA�|2��s�[vU��
A��iv��S3UG�e�D�����sǖ�3�7�.;-��}��IU��NvD�@P�Yʷ.Tq�FgaI����R�`��K،��gͺ�uϋf[{�����5�i��j��)���EW���8���F<U�Ns+����b�ޟV��󢥁n���Ӕ�J�m�$\;����lw�:�<�pU��PÖ�{�sEI�]ӵ�T�	6^�_n�8���p��i�l�?��OI\���Q�5��G@@�ր�3�u�L�!ts���yCF���c;�ֱ2��D���[mQ�֥H�|�Ҥ�dl�H��(mէ�a�=�$�=1~$�F�s�Q�1��;�Ѧ��%��
d������&�D p��'�����t���5e���95�<f���#x+Q�����<xx��- H'X�!�0Z�%�=l��`I��`�J��^y9��A��J��(��@%kj�f�k��&EY��+�cA�/�{3j7+}3	8%P�b
'8Z.��깸��'�5{׋�ס���,ͽ�߆,������Ii3��@����(&�wd �o:8��i�!���b��QS��Jk��I~V�� �O��BعBw��#W�ﶋf��P��P�7�&����V�>2�t��:$�]O*1bw}�"�'\O�D��/��/�*�Z���H�������D�0 	�Rө�O,�tq������E�q�p/�O��^��:�c�� ѭ})�<�s�ޤ��DP��o��� �%�媹�b�z�����3�����ώ�6ٺڀ�vmHEeu苋���Ǳ�99hS'��]E��6Fam_s�fL��dM11xs}��}��
�pmyU�бJ���PX���5�c��7��ڏ���Z`$c�`����xO�b1�<�k�B���y��W�w���Gq\��O?v�5�k���,��R�'$Xd݉2����-;�藎�z$�}A��j6�ܖ�1�lT5��Y��g Jfrn%�(f�_�hz����8�؝초�����k��ӭ`R�,Wv��7��Udڸ
�ր��k��7+Ø�f֐�D)Aސ�j�傇]A������ʮp(oTγ�Ks��k
!�6/f�T"u;%�O�t���^K�[�?(N;��>�J���]H<��Ɂ,b��ؗ���%�I+<��tP�0�|�t.%ض�.(�A|A������a,�����e���@SP#Y�����C�_2_O�Fź�*$��0�U�R��i�j<3��&�1e]�]\P�
4��F�5�xp���X�q��T�vj#�ppV������u�HgRf�3���X��A��{N?Ty�l���k��\�ru+�ܿ�3�ObΐͿ����jq�yD`FM�{�J��Z���p�b�D��Q� �U� M�,�$��ȇ����g}�X�
�憙ՠ�� d�܁��G�'|ߤ�ӕr�5�rd(�6k�s+�
�dQ0UI��N���BU(}12�t�>o`�I�C���$��[�A�V�=�ѓB�3P�a�GF��Gp&�
(�{[��U%V����6�R���vr���=sZ7�c�<?4|'$�ғ�Q<s���� �3w��j�b	P� ��ܭ ^�x���twe��:Cx3#���0�J� ���+r��s�^+��
~M۫���ª�k�G�A'i����>��0�zl ���y�Y&s8��ど����K�0�)\j��$��J8�ί��K~f�.���#���M|쒠Ɓ��P��4�y
�������f�0s�Ǎg�cn ��=UOSjɼ� ̖'��(,��S���k�-$Z�e�)��A`4���|w��U��{�1�k���Z���H�&���YkB�����⽸������ݎç��
 ��!�l$��qԚl���K�V�����7�<�9��Q˦����m�(P�>�鳴�	�m9:�f���
�����ԊٙhlD�;m'�$8N$	w�����F��߯
���=���?���@��q8>��������T(�[����騳k$(�����.��HF�r1��{����-^��P�C��8���گ� ]�hC�C��L�/f�/y�j%�O�~xA��QQv:ONiP�B�7�)>�*?����e��{VA)`�A7=8�~4ÝT�M]�v����ؘ=��4�ݗx�7� ��Q6|�~/��lh��B��6Zf�]��	�1�b���)6�90:�1�}������wI	���N���+4[�>��y��y�3u��Z�9Uz)`S�@ǒ���p?qp�Q��a���ɛ�B#�$�]#��*���R����D��i!��ErZ A6׽R6�n ��ai�e�	�K����x�l�Z���5VcW������RL���=G���(�T���-Ygm�uP�8|���h)�.���MZo��/�W�#��XW��+�%˿-axa�y�֧(/~r�[�q��#�@���+l��'�].K��f��	�SX!ه����0ڂ�f��UѡtnRJn	�:���<���G_9����%�1Qz��4�<RsUd&��������b&O�
;`d]'U��#�D�� ��vJ7�0�GE���J����𘔕Q.	�6S2:��@�w�\j�xm���L����w&f��.,��!�����rވ�"}�����O�Wr����pŏ����t)���6?$��J�|��x��p��@�����l��eږ��������An�lS�3�g�I%lgK�k�u�j�n�8>c��� ���K/Ļ�]V����	Ȇ��@�9{���˴�#��<�������SW!�l�8���-��z܋lq�`����0`S�CeE:��`���)�x2S������l��ĸ!��8�2Dہ�]�f"!u(��䔭�+��wk�C�@5�di�FR).�������r���]��h������NH|F�g�m*�d!�NŐ�	9���[�X�����ߪ$�P00	=�<�n�r�4�`�]S6��-���\w+?��~�U�B�ȇu s�L�-=l��1�z��4�[�$ua�z;p��CD�o7o3��a�J��M���k|S勲�`k5��t���,�7�;E���Nʤo�a�h���f�rwR��^ �˭f���B9���'�xxxUz�Db���Ao'|���M����A�0��� �̲j���T�{��=pz��R�`������e�1��W?}�^<�@�o��ih�1"�����{�Afp#@��Mg�*�ĺJ��[?j���S�q4�a���W��wE��Ћ����m(U����,����(�n�h�>���_MUl����U8�bKK7o%��D�g�+�Q0��#�a��8�n�2HJ����~���_^x�At�r�k���,T�rk�l+Y�xFɀ��
ƶ���	4Sx��kӸ������Tl5f�e�谝3�_�ad��u�*�s(z�Ǜ�h_,^�K�^<��zvKr��;�{��潹�U~��B�G�<僪���q`8��L�F�ok¨��6EO�(�||��7�$ma[SGE3����k�Q���akT���j�I�$���^��w��be�3�h�
��J
�I?���P60�DAԚ5�2;H[+�(ݰ�03�2\�5�X���h9�kO�Y��p�r*�R��Z��>i�^�8ގ�ګ��x"�Q�}��߅x�����Ql�+g0	��R�#�P'\`Rr�aH���X�NkhsG&e�pf�iBp|5ߑ�6�_Y�?�>F!��$���1}ƒنr:�k� ���:��9ڏ��5�՗��#71)����1��x�;H�@�'�����F2��,�����r����d�ek�S8ˇ I��q �\�v���Y~9��^���Ћ�/K���I�ҽ���M�TR�%Q::�˯�o�N�8��#��_��STW�����گ�V���->j0Ч�&�K���]jS�z�{*���!=i4��L}�}Fhp�R.��,}��6Κ����3f������Fj��.��9��f�e‬�y�^��L"q��y�������m�W#���ɢ�z������0���m��Y����?�Z���~/��w�z_�Wɥv	����Ξ��%�Npm� �|�{y��b�#E���ܩ����7����X5��o��K$�롽��5�{���9��NnPV�d{�o�H&R���"�c;���鈝B����`]v�h��6��G8HT�&�"���D�n�5քwֻ��%]��,Z���WMp��5^"2�k^�dR��'r�2������͠L�y�=A�FQV0�I7,^zWS����a���:��X6]i�Ԕ�Hˁ'�#��0�O��̵�<X�Ƣ�F�K׉�����s;�t�O�aaC�N�ˤ�(9z8Y'`�H�1��,�Mu).X�Z������^�a/�g���WC%`��)S�y�`�Y!�=����/�5�}�6?
�A���N[�I����t���[pa���I�u���>�*�h�W�3`1+��pjE�\�IK��=���U-��F�g�{�ђ��Y����4�R�5�@�2��z��~�[g��O�>S��O��4F��Df#�l���I@�qL������!Gw J���Ϗ~"ieI���v�&�կ���U����*ڨ����ƕ��\m���M�5k.����l�m�s��׺��j��!��[I��ejٛ��&tHI�]�f����	�'��9qG:g�?�/ˤ�^��r���2=jĕ�U���mm��|�2�Hd��?y���Q�M{�xyx,3��Q�jVz<I�Tr]Ϙ\�� �Ba��r%'���HGC�(���$�R����9Q]|��*�����R0���'s�?{梣G���㫊��:!m��qe�0a�s	a�K�!�y���56u˵��ъTm����r&��}�
B��j
�,c�P���p2�D#�S�42����]�rs�w	��y��k��A�~�D�$Z�8j ?��3��If����{'��QL]^�-�����NVZ<4E�5��U�`&n�=�#m��/��d�.3(OX/|��R��d�\�	�P'cr��1�vҰ2~��S�J��Kh|8n���m:jW���te����uk	�A�j��ݒy�B��j��l[���������������o~:Є�4`��0Ҵ&��%`L%ޒ�V�snZ)��tҸJ T�Gj����
��@�v�(PDKF�M�Ǭ$������G��t�n)��N	Es0kH~��'5mWsZ'	[�ᇝlW˺�E*�S!�떾rd=�Fp�2��5TK����M����d��E���o`�W�%v�ԝ�������h�h �hġ'tSG.�6�C�a%�\�q��9BC��U�c%J������q=zduz�e5/
8�������*�����b�`>�p�Iq �8s6�X�X��g��EO��q�Xk/R�����4��p9�t�!_φ���'Wb�81Ed��չ�Ӎ��aBm>ם��+`��zN���e�F�j���ʧ��z�(��7V��p����-	����T�%�ܱ��L�!�S#�U�$�*���J��c���v��`]@��K��v}B�W�	'�T^�h�0lԹ��su�?ù�pѿy���_�jrh���T�j���Ap��<BsM�m����@���gB�7A��K�,�s�i
z]��i��^//��,��C6��D�KT�x��/������ Z"$�i�͔�:��^9ξ��4�R�o��:���M���E��y��dl�� �QH�cۭ��ő����� A�(;ɡ
��`UB��)w"��:��u$�6,P�,��Vf�0!��ʟ"Ơbwc|�"d��0�i��N����٪?�(���%�0E?a���It�8d�s.���iU]G�R���M1&�f-��d�O.ϕB�X�b����Hk���u:��kf�<����Slo��{��غQI��"�'lHX u�-��jKk�@RU�t������ENb���r�W�~n��J���o-�����W���^h����s��%z�]`V�Xxn�Y��8����j�~�+�_aV���̅�������[�S)4�o���23�5��D�d��y-I`*Z;�C�
i|fi���
&�8�g:�P���v��j��l�&���*{���)�Y���8�Q�m�k#ސ�v]�9��&�8G�̪�j�V3��"*e5�q�i��@�f�6�p�ߦ5��xɉ� ���P�B6�o9�����Ą�[	��J�(��S���@�6��z����x�����s��#q��pW�j�+�4�AM�q�?��^�W�Wd}ZHI��ٶ��4.�t������A(��=m��UX�x-#h�:G
�q鿥*��;n��"�t��Yy�sa����ˢ&�Q��-~���p��n��iH>�s��3��AN��RӔx���7��u �F�83��m�p�00�Xx�I&#5&�Κ7|K�p��7ͳc��5s4�Z� [�T�J%�mؐ ����J&���SG��Yd��|��$7��_Fp��M{��򯖕}V�aMQ�d*HZ��?S� �&{������
$.�J��m�R�	?J\H8���4[�} 
����\����ׯ>���ߨ�(A��$P�^���J<Xu9f�wݴ��h!�X���Y<����嘄X�ń��l ��C��K�\�O�սf�K�^�m�����g�b9����:��h�^R>'���Ϣ$W�d��j���{�<��M��l����Oׇ[5Dx ��\y�(�\n��|���)�7�o���?Q��m�?.r�����!@�Q���ޱ�ގy��477��ȝ���$�v�%:�I���` fȺmST�Q�2�8��1�n͖��*�<�g�ƥc+�?n?ʛ�/�X�r�
d|f���������\�9���+Q�g��5�}��AW����vL��nk4���c�t�%sאמ��(
(I&�+��2:�B��/5㑼��I���1�WD�c1���$Pp�f�ǆ�盧�O�O����Ɖ�ɾrn9 �yI��je/�<<wv�&�h�=vo	9�f�"��k �E��o��h֔�dB���㴵�{g"0
�0OњqP<x8<l� z(9}4TA����9�:�v�C��ld$��N�8��!Kbx��]��k9�d��d��Y5*\Di�#�e��b`]ؐ�Z��^"��,��u o0�*j���ϼ������I�ڙ�:���>�(A.8�����Sr��ϴRk{�K{I���BB�����f�①J�pS-�� l��h�#�{0)w
mM�4ҙ��D>��9�)�>"i6^X��t��\Ɛ/���$x�U72�G�dΫ��~�4����Y���-��~���)���i�X�[ ��䱺��$���M�e)u3�����e�K��'�V�AgRB%%e�+�˓��;��]�>^_��a����Z�� ⭷uS&��� ��lHa|�}~��;�C?�{�IR7`g�}�RJS�q�<���bN�i���\�K�#����E�}M������������갎s�=�҅�m���N�f遃bM��� �s�d]���¹w����Z�Q�@oL*ujQ����D��T|�e�E&� �Q\�v�eH/%�R=<�/�?]�4,m���Y�����un��� 9)�f�	YD�*�r�P!;��E�E~J.�̖8
�  ���'j���A�)ƈM&@����;yF۠Wk�������<�����3��-B�<\ԇ��]�j���AI�\��q���I����R��*9ۛM�i��'����(r��ʆ�B����q�[�_�~�be��;'R�	t���R7��!�N��\�[Y���h�m��$��EH������F�:���Y�����F���!-z!a������_�Ь����M�m(���q/Y��_C1΅����CbٗrJK�AD��^�2`��f�x�-��/�����i2t��h��q��X<k��Z�!��=���x/��������v����̌6QN�0o?^���wN����p��X����ywG�����)<���h��k�+�f:��Ȁ�Jwx��릣�icXq貣Z,Dӕ�����ʆ3"N��͚t $�եF��є�1��,�$b��(��h
�iX�'�p������w������Č��%mc^[�������CV��TS}a;�Y�smVTŋ 1c����Ӵ��y���v�%�~m�nk6O��m�
jE�����JΉ�2�eb���s�ؐ�f�z/��`N��O�G��x |�G3����!Pɸ]�~�g*EV�Wy"`������'�Z^N��c�f�#�]�C���"Ưjpv1����@|%���'�o?��W �`W������KmFr�M��mK<�
��\��[.��n�Eȁ��=�|B�?鐤9R����������Ǎ-���A���!8��3�s�ը	�;��9�5��g�Z\A���o{���.<������l�Ԑ�wm��I���zˊL,���$錈L�}�{5׉O�"� _*�Kr͚S��6T$�+E��s�,6�7�$WE�=�����xG꘡�dU_7ٙhM�}��]dP/�w����}~@e��[�t{� �1Y��	�Kfir�s19B�8،���y��M9!P*JR��*�2M��w=�U��T���� ���e�̣��?:Q��,�}]�b�"<I/���U�d�$�?ΚR\=��A PL� +�)�SVk�Q��x-�c�Ca�7r�o�Ki�O��k�PH���L��}���c���QثT^��m@��xtT)9 a�qzH�հ�v���P�97A'ނ!;? ��݃z��`�A�x�Gϰ`w���k�J�,���/�x�6z�(�d0����r�P����<F=e��U�#;�ކ(��g�K8I����gA:sꂛ_�����ٍ'�>9�A5$��r���{����$}�Jt�܏iL�������,�e�Ъv�R����T�-��Hb���I݅�e�@"Ɠ.@�rZ�Cã����f6tP`oTyd`Vx�F�tfj�����(�5	3��,�h��0��}�gQ3x�3�hBgX�����a��8�F���fF2v�S�ʷ��ť=jOn����v�5��T
��\�S���GZ�U_�Y��u�8G�H�`��b<��;�siL٧��E>�G�U,+��>B���h��	Q/32�E�=� ��+n��zi����[C�K�<��	�b��	�S�4#�c=$��s��ڬkȂ'�����n3!����z"J6j,2l�
+3f���*^�D�\�hz�-�1���q���>&6(�E��&m��)�)�?��(���z�G]��8��+S�x�P[�<}�V�/^������_dk� @��	�(ֱ�I�H������I﫤�>��8��ҋkЉ�>�\��j�ڮD��F1gc��!0��W�*�Fចs^	!�-��$_�P��Sɹئ�L(�f6��Az��K�_c�
���A4?�m�$���Ї�:���Ц���K- ��Zܖ6P�c���m���������������V�:��i):_Q_�}�W�����E;A��!�jP��&˝A$��x�<Q�3�f��k��hH�~��+`:�6�0�����(Z�I���#K�b�l�mg��AޕF�	6���_I�y��_�9.���omyKA��;~Ľum��epCJ,�Z��C_�1��F_��ݻ=�LS�uJ}�㶃�]:����_�c3�z4�s�����6 !Ѹ���r>g��;ZQ�j#d=k�R�(��n۽x������9�Q���ǯ�2}Ą$�w2��l�V�Y�'��&��'F�)�`��L)�G�ڨ���~�G���1h�����#^�i*���6F���a���&Z �pn��A�ˏ��Z�m�p�j`�i��v^	�/H�jN{�����δ�՝��Κ&7X�h�W$>��z�uxT�/�
ԭ�
�t�1�\���zø]�"4� �ǎ�o��e+rkV�J5���Q����DE����B_�ΤJr���>����(LN����Iظ�_U�K ������� �?���&�f �Kn"�5W���He�ٳ�v@X�ƒ�leD-�9� ���،�z�{}_?�¶|��6�㠝m�Tg���udi٨p��^�{��5��|,/�{鵦�)���a7���=9=>���3u��̻,�>��-i�����s�H�hk�â����W�����nטHH���'���P&V�����MF,#\���&f����Q�f����.��r���P�41)�ۊ����	�� ��K�'�fFŨ�{��Y�{iK�I�JU@~���;���Nѝ��W����Q	�`�d@��)��&i����܂\�Q�D�Ql2w���,e�5nI͊{�:�up�xn�2��CK����������{�I�~��N;�I����`nP뿼�a!C؆ek�.J�P(�ٳ�igS�j�� �%�a���Fތ}�M�G�\[E���� � "c�x�Շ*�7���Ŝ-�<yVQ�/(����45�&�6��!='���`�O�-�~��{�e77ج����s�ۻ��>f���h�Tn:��(ט��J d�<4^{'�wP�A��L�AY��3��rb34W�1�lvB��v�gL��*�HSַ��<q� �-;4�{��G*����3�N?o�39 @|1�{X�m��
D�8�;��� vy�
]�ӌ-��a�m\�ĭ�_���6ϋx��l~|����{����J�moI!Ҳ�0�rk�8��87M%���Z/�*��s��nF���H�`���f�ѢiZ�[2i,�h�/�y��� ��;�om)�%V�uȰئFV���x��/�y���U�֌B1��镏�<�a1�}����wgPLX�Ϳ1����,��5���q�P:S�1���1��n���H���+��F��u�mMڇ���0<�x��w��g�aG�t�,=���ɶ0��FV�� {��Vs�W�L��{�aX���Eb�D�!�c���8{V7�P�!�e���O	b���α��S���<��\r�Ê�tHm����[����j2�A��v�E�tq�F�*<��V�v#_5��D�?�A�!!ެ�$��$��kj�����5� ��z�v"=\؄s"oG�8z�u�2��3�/۴��ݾ!�&�5�W*��L�lb�x@vV�����U���D�:�)˼��%�^����o�;�����h�K��!s�7���/x��F�,[a=B�O,�y ����&�$@C��b�ߤ[0!u�k3�Z�Ų�-Y�}��#�h�W�
��
�ɽ�{5*�G]�[p�2_��5���?݉4:j����vF���<Hhb���"�����5PFa6Ɔ�PR�k���!y��@�ca��yd@s������$�������I3���p��=�W1T�6�͸><�$ �xv��,��=}2e_T�����H�����I,�{h���g�4T}Z���<�=�M=��NY�l<���_f��D�	�s��5%"�ԓ(��B��H��SW�d�V�߈3�]/�>�K�d<l82q���{��{���^=T��[{���\5�2:X�s�����o�><߇1'��4S�.�]�]V%Z�o[ `F�Xy#�=�x#���5Ȝj����<�w�kw�3��"�����/)�!�B��r�a/�"| ���m�m9��]���r��N9�=	�;"l��}�h���lq����+ɫ�:X%H�R�ȵMa��[ZUM��[U@�B�'�3���R\L7�`�1�i�<	\.��e�����0E���7q8�WU��lC�:8��t�)�&�5�^�	���d�=���6����g�I�����)/�i�,�	|��o�Y5/�%q}��f���I�S*=�	ĞV��Q.��"�D��2+d5��O�i
r7�V0¸;��*TCo�Aw�9�hIV*i�k&�|t2���n���B�����F���EU���{��s�8L���R6�/�Z��U����ŀ��}D�2���_��ֵ��fZ���q�Ͻ���EEɁG$u�{�@k�~�C3�4�iXT]�rP��+v���D2ۙ�/�t/dr2Wo#��b�&RC��1gI³��+Uc5�
��Dn�Au��f# 4B�ǖL�����z���>�V�Ϋڰ�H'90�l?*�l��Pt�S��9 &�44<��Pg/&[a��9�`i����>Y��Z��M�?�2md֣��gT:
vA��g��w@F�:W��B.���	�8AU6�]�2�0ӎ����c�$!Ψd�z˱�ؼ4�W|MKh� 8���m���/H�h��Y�9E|��e��rk��O79X�7/aO��V�z(�ND��lp
q@j��;����+{i=A;>�ݍ��j��ލ:������IMP.���`[w�ٿ����;k�|��i6Ŗo���vh����[�Nt-ho)a�U���3���ҊwkT�F����/���6�ၝ��s�@l�����VD��{Y�V�3��fwx��Te��$Z�P%`��\<6s��&c�l���]B@��H�TK��!Qn���X��,���H*N�E]�j��,���;}_v�U������ڐl �<M��mF����o	�	�Zv��ސ-�)��e�sC�	��8�8�\P��\���,%�Z��?���D�����Ah��n�"�`�����$��|-N*�%Ps@μ�ީ��sc�� 2(,!�4�#�I3�t���cf֏0,�
$��]8�Ӓg���h��\o��G8	1�����̠K�2����r[3ŷ13
�Wh�.Ӗ�'j�;����(FaV,�Ϛ��p���a�`�rk�I\:�)=آ
6�ru��9�G�M��������g�g���g5��m��U\�+���Պ�.֡u�w~�b���pX���&=%\~�'�d*�����g:���Jh+1�d/)���nH��3`r�P� X@I�M�HQ�j���b�Ӆ�$�B��R޸䰔WU^%��j��l�N���ld����W�o��l�&В��H�t9G����=�<	r���T5�@S_�{��ކ�	gpcG�2S�����i��_��2�EI�6p�������N�I��a(���Fq� T jA�u�ʮ�v�Aa�=��8!7���1Ѿ�w �M+ �?9���OW[����mJV��ܱ􉿵�������]��%�O� ��c�k�9�d�,����s(���6�A�^
d��t���`ͫO*ζ�9L1��ήq�_��З������V�b<U��rޒ%ue������j�V�M�K,n��qB��/�=v�uW��#qκ�ſ�* �*� ���L��z�uƁ.hg�~�7��LJ�=lf��Vqr���|��~7C%C��ط�H�C�ؠ& w���?9�HOZeTn�|k�c�5���>I�e�rY�7�hA�C�����Q�Yo��F�P¡���>1A3C�9�n_�8�/gv
�hr�FJ�����}�����X�����7�n�e��Y������A���U�-�Y��u��6o�#'�zk]��ۘ��LM]����$�~i/�mR��K��5�**m 58lq�"�ޑy��xkG�݅W�OT�����A�v^�[��f/$�B�jZ̠-�:����!���=�	�&ڥ%t�����,��8��b-:S��9u���~2¸6%.3f�i�T��_��6^0"+�1b���a�p])gC�2��]Ԫ�fZ�T��y�"�C�z����!��}}�����+�W��j)d@{�u$������t
�oɯ�&�嘍�z���wu��.�o�T��aaQ����k��_H�F�F���d��R���ϜyˋI?��T���x�CJ�C�l$�����GzD���/?N����p�������g��1v��s�D�%_)�Ӳھ^�1l�|MBb�Iit�Ő���@�w�����]���c9K�H���̄,�!����m�~�ç�x�8e��M�d�����CuFɩ>>}�f��R�Ft8o�Y2���P;����h�nk*��>�������^�@ �jGN*���Z���8�A-P�X�؍���{B�,�;����%���l�E��ߕ='���89�L���K����DN�֋HcZ��b�xJ�$(�K���Ze��d���4o]8���[J5*SH鄨�A-��I6c<���2|?��fc�@5��#~���=�V{��l40��|̈¹N��#��<A	�`�)2{b�T��C.��l��]<d�Bd���tlm�'���'Fޏ�{^�X ��+�)��"\�ǘ�W�d��Pv�C4�Xn"��̑,[O��Z["�7~Xa�t���~�+����NNE
�B^$	�~��m?ˉ)��)�)���qRU7.W�keD'z*E_�yĕ��X�Ӿ�H�'\3���Q��,��-�'��Xj��e���q�@��gnL�Ey���_��:��6���|��s�����pd �96�i��D�o��w��(\A�T�
�),UL���D����	FLr���EѲxk��JLaTt!�"��J%��J�]�R�>�����xǧ��_�`�q����t	n�~!���7N)�mS- Ԁ��̖��d(b.�h ���0_�opl�yJ���¤B�����9�����s�ix������V߻���8�d����Za�����%��G��R�K�c��P9h�Z	�8�7���)�X���������?�ѳ�F�R�7���.��P˗6}@�0�$�azrj�v5/@���_6i�^I�t�ŗ�
�x����,����`��ٺy,qx8��5����L�
(�\�P��Jū7d��J]�}�J��'�l���z�(�i(�'{¿��q,Wc������Q�b�͘�Y/���M��ȸ���t��q�v���L8���$�ݺ���$�ȸ0`�i�
Hxp��E�]��!�Z��3�(���@]�&�g��+R��a�PnG/?0�:j�5��x�����Zn�H=�؏���0�Arp�gU6��}7#;���z��aM��i�8WW�S~���2>�[E�a�[5ҭQL{?g��\$��xG+)0GR����wnY��XP(�j^���錌���ܼN6s�m/�f5:��W�%zO��:�өw������)dh(z�U�)��� he�'5��69T��3oWA#ϒ��]����9Ӧ���i��BU���\h�\,�q��I��~o�*�!������+"��GN�b^
x�8
M�j�[iF�����M"��`���}bi�����-Лg��oї����̹DY����߈����.���S�mȇ�dR�9�Tm�UP��Q�����AA�ĺ�|q�$����:O;��-ʉ��T+��$FZ�x2]���J]�#u�S	��$�!��SGng\�:�����2���ic���g��uN�]�2X�B�$��zcf u��V�?�bj<����ۃӁ>I5���R�6t�B��y�MC����*M�3K�r��O��|�[rp�ҧ�lz�>�U��)���iw��\���JQ�vi�Pb1���`QY,�ϐ�E���^$��d��?����(�izD��3KW� ��N��R�듅ZK����#c�rG
�8"�_�?�=0F�28�v%@z�pĝ�օTt��W�zdC����P�"k)�I�3��Uz�pN����W^ﺮ굦���V��<܂����8�n����:��r!��c��F��[�dU�;$����������a�G?m�ژ�c<S�[����mhL-8ӗ>�@Itch��0aG�^.�b�m�ni��<�)��۬�u8r���`��8#�~�S]�����׀[�Q�XB0uÖ|*��,c��ޱ��?'�7��3a�̗I�cI]��`�o��@�z����-��.짬U�����n%+v$S�fd�n�sS� �׌!t�P4��W�^�Z���������timmGP��zG�܂
��B��r��*�5$�w�M�$�5�0�`I�:��^����t���E�Z���!�g����޹3H*'h����)�������w�2�n�Ӳ�J�D�i�La�)~����������~���M]�XV��ߢe禍X�|!'�p���9�^蒥��H�֨��E��i�S�[-�i)��������+]��O�22��}H)�u��V�̆/Щ�:�/!yfPc;]�bd�{��G�ЇhW���'|I�1�伷7bH��tnp������c�����B��zz�@w�{���n�oV맄{V������E���� ����{2�����xY�ܓF�[��v٘����nT"��X�n_1CS�����V�7�h�b��F�C۽ci��a��5l1��9���]��4=�ߣ��JT0{�A�J�Ԉ�`�-�9s~�� b��b�Eϝ�5�"��4��Rr9}zVa��ƺ��W	$�t�@��s{1b����v3�@���Ɖ��y��~~JZUJy��:��㰿JQ�d4�\:�)�ڏ�#�O�ȧ�&�������P[�	���~��F��<�X�� ��������]��]q�C�Ȑ&���_$��U�P5�o�:R�3�w��(HF�a� ��Ol"jq@���n}WNC����>���	�v��� ������:�E�zAqK�����TEs���acG*���@��a�������Y:�?�)A͹CA�ok��;kr��Tf�5 ���8�:��.��pF;������r%U��v��'H����^�<�J�;l��Xr��7ZSq�*B_�����Ҷ�G�_/�i�t��+�p���̗�C��UO+�Ȍ�0���$}ߋ����>X<���^Ї]� ��>!�&��|�� IO�h�l�U���{��w�$
[�۲�6����ߡ>�	�<��"�d�R���:�I
<q��O#-���H!��Ѩ��,���8��kd8@���ҧX+:;���ҩ.��$l�,u��;��]��sk~�<����:mRL�(PM��=s�?I(��-x_��]7F�Km�-�B�'�h�����A�t���ǣ��ބ!���揔����)pP�O=X%��i5*X{�7�ntk���&��J:	O����ŋpTD%3) k'k�hSԦ�����	ֶ���N��/m\�9a���)g��sm��P?]�qOyX�M���&��{�O�����k�E�,�c�F�g����S?�B�z�#gU"�>�����	���>tZx���C�wx�ť����^�F�/f���Y���GO�c� �����C�T�i�������)1��h�\e�|��i��L��A�1TGQ�?z�
a�X�m���Q��ԉ�~Ke!�1yI Q�]��5�n����+�_�T��q|8��^r��@*��C����Dnk�����N�LDF9��L�b-����?��Y��n]��Oi�[���L)B�F�F�~\�F��D�fSY�ا8���$��*�,�.�x�D�lU�n4piކ�~��z�������v��Ou�sl�%)-��b��vf!̩�ԙK�H��*��DK���5i?�^�}�5T4<�@��F�Q��S��,��ü��
uU�Y�����:F�"��OS��2P��a���y���Ѷ���.܊��|t�;ߺY�g�����Z>(��H��	����0� (K�-ZS!Ή�ܲZ��^DC<UÕ�|y���=�z�_=�'��U�Va�ذ�
/�gAUb����\D�#�3b�3V{^��,�l�Q�J���N��s�5�rEK&�K΍̌���U����zpI�$�n���A��$Vi@��ްľ��ۨч����&�9U	���(�X$�h5 c�R�w ��oZ�ڱ�.��@��C�1��
L���H+9�ۅh/����0��;���wjh�i�3�u����&��W�đ�=x&��K$�}����n$د��pM�b�-4˲n�C#}��?js����M�L�>���j߳���~k���3���*�+�@_h>#IrK��6g��PU���<�B�����
��"��6�s����W[)	��S��Z��c"����9�E���N�=��^Ԍc0��`e�M�����2=�Ԧ+;pE�� ���t�%�=D����1#
�b{/�R�$3st� %��Y���RG�j�ų�K������P%E\��2�ă� ��َ2�[�R��и\�KLɪ<q�]��fy4"��}YCi1G���)��|�.1j�R�W�S��L��}7��^�5_+��Y���t��X�e��/��������R����a]�J��迳������SCi��u��q��zk�{x�c^r�	%Qa��gyK^�
I��.@NP���5�;���*�]}񯆚����t\� 		@V�^���<C�������N
��1���B&�/���3㇖̈́�VY��-�?{CfuIK��r1�w���S�.���I���L���[����ǿ�)�0)�"�g�ߔ5r
�A�����d�>��������_��S;~L�H�B�3O�<�%=t�P��*�R\>7ǻ1��>�����]�G������P���x��0+U	����,z�]��X���hB�	y%`F'�7�9���ڟ��+7bk@��̒S ͷo[;d���B6=n�%/M�� &]PPZo�qԈ&m�r��U�H�4G-��o(�����!�@VD�y[��ۚ�� `&��o�#!���x=���x�՟v-�՟�z:.ŋ�n���ѳh�7T:U[~1�2���h1C0��t:�J[�����%s�V����%��;��{0/'W/��;��q
�}|`�ec� �x*�{^���x4�\w�HU��׮Ǧm3O�蒲��*�;��|+��(�.���",��=��e�m�=��]ַ�5�v�S���`Zy7D3�JQ3qĢY��@f�-�������꼡�2f��Gy���y���BN�����<��9�$���OJ��,��{9���1:[HH�GZ	U+W;_-:�l{ϭ�s�}^��[a:��H�t��͈��ج�[����Z��+�ӹ��a��q�?�o�zI?��-��hGo���~L���]�;P;��~ `�Y�]������Xzhhl�~ep���5R�v�z�X�w�T�<qQB��1����ᦆҿ44z�}�/Щ)��u������� #��٘�@�G�P���.�IQ��U����f��T&��J���C�}�#��� �wu�Z+V���p":�̹�s~$�G:\b�IE��R�0��
׋vwq�{1����ܛX����`+�(�6��`��hoo/9��_������T���w�4 Iu�dV��
f�]yf+�+8�����'Y�*}g��yxk�`m\���H�6��I�:Y�u��g��;���=G�n5J#�X�kʯF��"��K\��&�ͧDW2�gc�{�LQt�
���+u��Yab�+ y�}8����Td6��j���Ӡ%������V��s1��w{�óJ�yx��݆
h�߈��ʥ�>����L�?�6X�׽�3���� �F�G�i�[]sbG>���<�.R���ҽ��I��;���[7<�Zx�1�����%P�m~��Qz��J�/����B`_hfP
��c�7���IPȉ�Y�e�IUfU;���t��8�j�$�XXv���<��A�5�|���m���P��3cց2Z��t�7�>ٟ��q���}Qx�o�7pY}�S{��?_<������d�EY.���ua�&�2ԅ����N;]�a��]/�F�9I*���+���1i��ʁ3� <�e�2����W{�r%C4�Z�����< c����G3E� )�r9����2�_���^O#C�e�d$�)�\��'�u]��S�?�X��+���hw�3�ց}f1�т�xDz��j��N�?��ᩏU�x$!�¸��jr0~���G�J������,��j9^��oy����L�ܙ��ƥ�z����f3bmFx�۰8+?CyA��OM�gg�G5r*�.��?WM�ɾ :�H�\1Ad�D��3��6�� hD%��j��Y�p����bА���"-�M�)��p�~�W��1?��X_8�4���D�g��ECA�Jv�����R����Gk�v	Ҳ�rƬ�_���(صW:�BS�"y�C�0ٞ �T�oH{�y#��M�8_@��}��OA�7�8���^�I{�)}�tT�MA"���[;��]H���P�F<c��E� A�ֽ嶝Cf��@:4W
������?����gC�f6�������24�~����<��A�KO|�3@���L�iD$��h#:?PP[�Isg`|��_T�Q!�;�4�EÙ*��1���dp�zmW���2o��8��f����}v<�DlTԯ��NT����ka���d���O���F\�ӲW{��-j�����4���B4c������xAͯ��%�x�'���|�^;�>
�S�,���_�soW;G���|WF�?\���%	U�z�R@FS��>�D�	F\>���[��獑;]G�������'�PM�5R�K �e��xS֦x% =��>������;�,��k� �3�BHf���J��|E�a��M����� w	~M�A�#�'����E6��K�e=D�k�0_��h|��Tr��ĿB�� c�0j��/���E���ON�)I��c"x3�$�B�C�g����q�ݘ��[�}�g0��G8LrM������+�̃�2�`p�.<���s��Q�q��v	?�s��F���%Y�6D���\����~��1��Q ��8� ͐�k\@�J��>H�[Oq�W�1:�,���,�hmd^K8�b��4�.+F}�a��6�t��rn$�*�2G�k{���d�~�2�[�0��>nF߹�q7�C��P�y����q�i��'#&""�]W�6�Rˢ%�q�i+FH��/�y �R��oz�����)�'���Mu����O�(|��2�<�LH+�FOn�k�S�� ޟјq���ݖTz�E�Mh`�bB���攧����A�t2�etհ�0�fu3l�p	��6W�+���HF�g
e^Wu���-x'"�����X�p�I�X��Ņ�D��pYE�8����|K�c?c�N��S���X�Ɛ�ޢ�[�6��3=��u|"I�wP�1n��I�~��38 �<����h�P8~�<��2�~0�Bl�w�RFUj ����5~q��bv6�$A��s�� �k/��{�����ޜ��m:1���M	��sU,y���߰aw��P�]�@L����k;���Y;Qr�hj]�6�����XU�2�a*U�ƀZ��O�������RL�:2�gc��7ݬ\VE��6&�)Cii|�nQ�����
h���$���Jbq�&��n�w���-8_��^o�X+ ��H����h�)�ퟀ�>Ԝ�~��_�E��`�^���o�-�x�`����z��ZZ��Av�"��uښ�[��US���
��د�V������r��Tzsx��2�5�ͬm@w��\����B��
��{)��ܜ�b]V����w?:��Sʇ��l80R�u�%Țryi/'��� �vSk�Vp�:�3f� )W�ì���*m)�D�FN1,j!�焽iW�X��l�W�����! @�������"��_��d�`�C8�[n��/�&���l����G�J�utH?�-�}�}��]���;jO��ݶM��&q���!diJ�	@z�>��K��v�|��Hms�"԰&��!�;�&m��B����"Z��%�]��RӐ�^��Z��>����gD<òu�l�.���I�+��G����4QH�-�G�!S�~OW,-߁	@���ܟC{��bC�D��ȍ(�=��}
��q�,"d���AZih�B�ѻl�@3�����/ʹ&j�'�ş[DHi�K�?Zr0��*��ͼ��f/�����4��j1uWg)]P�G3�:�_�������B�[QBv�{��Dp�d�0H�U�0t�^X+�W.�7��T3�a�$k�S��6�\�t��@�#"��V�w�*&�ۯ��{Sy��������?.N�d�8�h���!���3�G��N�̯3������>��8��CO����=O�O*��,�Ֆ�A�o��Y�D䭱{&�����݆L��N�I����z�A�������`��"kg�J�"�j�
J���eq�9N���~�s�Y�1� �C�՞I��)�:u�=)>+G�wC&��Q*J�u�U?9����a*1٪� �y
�z#.��_r� re��kH6Z����,BzK���J�Ҋ)����ﱲqN~��sg��0�%�b�y�w���~����r�3kPC)*W�e��\�In��a��'P�Ι�:�x'O���S��5�W��r�h�}kxq`\sޖ]��v���<�eȔٵ�>r�ՇH,�8ꋉ�3}#ZM~�RO�ьY������cߴr��'�=�W�AXJ���=ׄn�PGP��py�N=R�����kb��Y�f�?�f㋶���������Nxp (
ޫ�;&T�>�	[���h�p����� ��ÃϗP7�"���X�c��B��0U���#3';�Y�7l,΍Y]<qR�r�)g8_�֪9���L=Y8���dڣ�Z6��]�آy�������%ٓ-%���@����N	!���2�B&�nx�t�8�kTU.KQ�o�eW-����(/6��Q�X��5�֨?Q[Xd����D!8c_��/��}1&�qZKg���_�*9��ô��eg�8	�*2o�XK�7��y0��$5�poT�4�M���܋f0$Y:	#���9]�A����0�a�P�l�]�7��ҷ�߽xƼ�oti���ZK�Aˎ��l��Ie���(<�퉳�uP�q���'��c��Acu���v�-t4[ٲM���ؿ"����Yb���"p��;�F�牺@t8_����MLL���<��]�*�i�!?�(�7�#�r�.���oݝ��� � �Z&��.�:HZEť�ϙk�ȁ�|c�[� k�!ШZZr���I>�":�����$1���I�Һ�)gAr��4E��T��_Le�.=AM�QwW�@o+��Z����:m����Ԟg;ϓ�]J�?kA���`-�s�)����(����̫�g;lӰl-�l؃�!��;h�
����7��<���.���괭�a���s�1���A�ӧ 1�~���d�����qՈ�C�i��*��oE\�o��K�e���H��鰠K�fki������b�����`�cgTj�N-.�����M9ڞ;6�a逌�[ Q�z���[�����/�D"�zO��d���DiwE:��5�0q��?>��EIc)U���D�3y�^Uf5f�Z�PRE؞6�!��\������G�7.	3��W��Bh�����K��z<���U!e���eK&��ox��%�^k��d-�ݲ�a�p��e�����V�Fy��H; �"i5�O��{+պ�g��%���>����XW�zXR�!���t�XX�� P�u�z�oib��Vm��T	�h��0��ީ�|�^?��Lgsn^�Dj�a�W��$3�={f���@�n[���@&bo;��{�YC�NAJ���w��,�R�Y�6
�y�@��pU�*8{LX?M���-���O������35�JO� �#��?�p0O$H�h�b^=yq\��(��O��vAh��������DW��>��L�̔��UӰ��?֙��d\}}�G|�7�0�
U�����7��!��5���W�Rlu�M��q{5��]�f��8&�̵����k|/�G�n%#��/��0��FcŤ<��N��uK� (�S͓,���w��۠r ��G��<�{��,�St�a�G�;�S�A~�Ec��G�v���
0*犞}ug���nK�3o��;T}���ݺG8"�B>�Z(v5c⷗�*���D	��L_�9�����H����G�3җ|�×���:J$����06�Õ��!�%��(vq@�{7�i�EJD�h��,I�����2�NS��YNɮ�ZO��Ei�M4��V��v��v^���#���*	�*�O>��2���L�|$�|t��������iKT]�陼��ڬ�[�
-�v���9-�7:H�L=\���q����_Ņ�z"�F��z��F�]��K	�ďx��5zUڦ�].��tg��F�_�h0�����SdAH�ʿG���:�(B'����7+��dC�ge�ݳ^���u˫
sK���=�0�ګ
WMFx%:U�q��Gm�ޮ���0�d�9tztb�/L�]q^!_�AO1�&��iZ/!�0��"*l�
�^uV��8~�W�ATe�O�=) a�����a��Cp,����1�E�E�bVȤ��A�#_׶aY	�,�}y�xd˱���5��N��3�Tn����j�ƽm<R�?wZʃ�n��u�6�.�c�{���Dwf-�d�1�n�I��o�9/�D6Pbu���`����q*tEI�*�Z�v2�#��t/C������  6���>6mL�3�p��{��qX:��8�����6ǆg)S����7�\��Ig�{9`X���J��te�A���Β)5y$U�NPW�iYQZ�܉�H�<(�6,!z=�NyE�h�c�ۿ☘GD1;0��@T5d�7q��l6B..7>R�i�W�� ҹ.� ��	Y2r�����
���1���1$����6w�&G���G�&e�y�=�,�����Qh�� /� �����D�����7���i'���~y@����*<f)�%�)�:�=�E=#=�|�����@+Ow�UVa�4�/%�S0Φq�mV�n�߂���*��$�Y�2�C��[�e3n����p0]�B�F��T��&�%��8��,��;X� "��u�٧IG]o&t�JKz�:�	��z�k�`�0��2�r�n��wu\O��I�"��ߧ���� ��b(�� ��Y}CR�a�Cp���,��˟L%�y�Uڧz�WÁl�R�X��c�õ��C(���e�r�Y:�k��PO�9A�XYQ�6)s�I)���#�����7��A���I�KM�i����(��A�l�H�hi��D�z� �ܧ��t4>�{�ۆ�Yi*��v�੆���_���32�]20KO�%�0r��.��#��s�Z�W�o�%ʟ�Ё���?{���U
�Ic��R �RZ!2��o[�gǕ*��b�y���3m�2����"\g�Spmsc�A^>޾y�_J������r�d���,wZ����A�i3�A���;�fqm��%���с	�>�:�*�R�3
u��!�5N���+<f�fE��%a�XeF�߲��
��䟩���!8X�)���8���^l���<:�B��b�T9Z�`2�^���4E��-��!���7֩���A~UE2�6kJ��]X55��U�6���U����&J"�wK~ʎv+�
 �*��4 o���v�&�7�+�Xq�:�\i��`�����u�✶�����0���t\6d��A�b�LS�½�<�E��9�!���,r��E�q�d7���&y���9Ǿ�Ģn���Ր�ph�"�8s�5��՚67l�p~�?���<
]�ۺm����N4�R�Ҡ螽f��^��ݷH��E8vǫ�7H\%>��1)/P���!QMةF�5�+����s���z�zT��U!hr�.�U�I1�Jm�A��m|��o?��+���~'&�$�?`��\�����/��f�����В�8��xbl%U��6�!BLy�Qʵ��D!=9�7��������\�O/!�i�ݲx^�7^�����:T̝���Z64�ǰ8Z��G�9Ӯ���@�����:&�#�@�+�y�N����o��6>��Cˌ�B|��T�d����,���ı�yy	�̚��.8������P��q��:=�T�,x��_f��B.�I�0�"�m<�화A^�Uy�X���@yGcY��P�H�c�Zl�v�P{ީ�}KG�vyL�7�N5i�v2?�Ķ�ZԖ��Xp�d-�g?Q�s���#q1!,��ѽ48~�$�m������
���Y}ڃ�_~"Wl��1{�c��\��E}=/����M=�c���X���2��g��
��T�Z�>�Ì�얹��7��#�A}���%�q��I>)�$��,�f�
�G��[�.��}CT���Sd%�ʌI�I�no"M������k�y���ʭ�Y�Պ����Y��ɹ�O���H5�.c��FY||V����v�$�1����p?�Y�_d�?7[ӛ����M_�$�-���<fz��eEr�3H�<�jjvi�}��iz�����`w@��J2���r��s���Ro3�͹p-3�
5�#~La��Kܳ	9�oYI��L�n}.�R	kϬWw�:�&����T�3a?�����c�ɏ?��TJ��dk;�"|-�tmv����ŵ�u�q?ƴ���A��M
�#�WS^b�������i��eCK���k�8���SE���U�9�q6�w�d N~u��b%؂]Wb%#Oe��1�v�~%g�0�K65�ɍ�
�-k�0�D��d�#h8L�?0����3G���e��'HM忇LZ��͢��q�b&��0���Ӻ��>�w�'�a�̨dJ��Ƥ���ߩ�Y.�FݷysJ��o'l$�C��l�}�>'���J�׻������Mo>,�Y�?��?����PX$a��_X�o�A&:����w-��e5���4yA���9f��6;��֝غ��g�f����=�%l�
��t?�<��_���H����6� �$�*��@Q?f�˱\nF�8�
4��ˢ�C� &L�5�7����!���2�ь���5��i��6~7��tгLT"2E���os�0�Ёm-5�ej��b���"\F��X� F$�{�p�'cu��[FX�-����yě��i1�;)�}o|�.c/wv�u�ӂSUK=�ډ�BR�_��V��UJ��k�ҩ-	cD�5�6%OD:iK�&���rH�'7����8t��)��k�J�7^+͞�K������4"M��IE�DR�I���y\ʓk�d�C��񈈀��|�£���&���ny��<;�DJ������V�O�9�'�GW������fGE���q4���+���R.�d5[�����_|���2d��Hղg�i�k\'��t�5^j�Yr�v�|�m�+,�O����o⨗���*_Q}�?3f�8f6�^ �o�ӯ�RkR �IbF�n�F!k�(�7��2��7�W�{TJ���T�vvEw�zS��	"�U�N �����fF�2���X�+l�Q������"��pE�e��zj�šNLP�5�����5h�J��2�B�`4�6S��q�8D,�C^v0��>�4A	=�����^B���9jO����dEwRy��_Xd9��A��OAP��'m���MiQ�b����#��ʝ6l�^�4�I���v���%z7��7 N�m�U|�B���ÉT���ξ��ӧ�!���~��E2"��`���������M2�Ն<;��QC�\ㆭe٢�� �pl�i��%��f?b�DhkL�b2�����%6�X�ЧI���I��c)���~mVXչ�C�lY�^US�V;�^��OvHǶؑ|�X>�H�i!lǃ�3~,](6�xS�w��0X��m�I��â{����#���P	`�i,��]f;}�E�9(@�L�¸���;�Z9kU8�t<��8*�d%}��PF�r#���kZ�vu�����d��I���,�T���\��Gi�X�̖����� �|�X+f�=�;I�i���>[n�������bz�C��!�� g'�OK���;8���_�ࠌ|�S4V�[X���:�=:b+��N���Eiy��8sL�O�
�����frJGU���ǕG��l�#c��[@�|������hU��;�� w�m �A(%=-Y�3°��ʌ�,`P~�6�VgБ0@����e�G��s��H��ă�6���͒��MCN��B&}a?k�Ρ�hVRUɔ�M@���dS�$ ��ws6�yYh�b��G�!���"��`�S+��#��鑾�G��v��W�����窫u��G��1���K�{��B�j!<���-�>s��ؕ�2��N�{(����`{�%��S��%N�e��l���vf%\��2����6�:=��ԭm��7�ު]�u�ǻ~����0H�_��mZ�ib]��,�l��½NЅ�/~b�	3=���iǷ:�8Hn(�P��&5L�%4�6�I3�~`�#"����mQ���g�go#�9O��f�o9�4|��Z��lUsgO���%F���	 ��:�x�4%Y�K�FNQZ��	�}Y�ʙ�s�(�u�!Ă��k�	���eR$���g�ж:�Nn�!�pp@��n�׮�e�~��Ƃ5�]�n�����<�� %if��k�'�͐D8�_��P�����c]�����T�&݈ĉ�6}r;y�4(����D��O�K�f(f��zcd�.	;��/���}�V-o0T�D�߰?uo��[m�_5U�����9X�ǌH�s��CT����;� m���`��O�o����|�+��pZq ��cQn�8�����J$����:��s�d.����,������Z���Bd;�"a�Z�
'}�U�,�C�����NLдY��f�pZ�yW.جȪ����/����;%M� � �h9����؁�I�����VLS;��߁]�B� ���J�?�:�F۪ٯ�۽�s����r�~�b	'3gg���>t�br�5����`}�=^����r�J1�Pf��ٽ1R���Z���@��NtW�����-�s&�r,�s�j@�/�%����c��[�z�( ۳�RI��/���¹�5� �=�<�83˗.>t��H�ԑ��&�߯�L����vW��j�9U��V^���Y�1=��d�τ8q��6���ҡ`�3��?xd��4�e�������6�5��̫��{����9�����k* �	Ǖ������֓��m��u�3�E�v��Y�G���UX��Xg��OA��*)���ԧ�����!�9�<u������x|jӡ	焋��O�9���ǼfN8	���Aj��|bM�q���i���Z[4كn?[Vl��#4c���1��U�����S�H�qs��Zv�r���Ĺ!gH+�D�(�D���"�H�,h�i�"CȰ'Jgl�'�<��^
Wb���U�0��:��ރ��]�s�?�H�L�V�d|����Z1c��0Pp!c#��Í�ʯE�m^߅�R���q�NG�#40�A�!��J��/��{��;�	{�Y�;��5��5kd��0��(y�3��� '�Z�;�km�r2�O�H����g�\P�ı��!�ff&F�66�lF��A��K'��3)0Xr�d��QK����6�Ya�^�R�~]�w� D�T+k1�y@��v�*���%oxv���rr45�q�	�Z�TP�y���ް]��J��{im�G�I0�rW1~�2YNz����&,�5w��3���ɉ�l^��_ҬK=g�$�@�&lW�J�m��=h�$��m��'}j�����W�Ӂe'S�v�x�-�|�6�cq�_�H,�ڝB��}
A˝��xwÂbJ��G�5ȅ��&��g�x�V�TȪFR'�	�~��Ag|�'���r�����MAҾ"��o,��a�S�����RZU2�y��o�=����܇�.Ϙ�$A(�\09��f�r--A�f������g"s]�,yn�1.��[�1*�� �w;����<��0F~\���ԥ��)j�u��Gq>Jȡ��/bn���S]���Izύ���y�@`��F��䂬-�7{��W��j���mnLG��g?V�%ָ֛-�T�E���S��3@#�j��E9��tT0���t_�9%�M�0���ڪ\��