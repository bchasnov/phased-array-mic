��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|�&���ڴzk^�2�C�bR��g�2��@@���³ŜbG
�'0�f���Az��1��@Vs���Z ���R�q1!Ua�V�| �z XxIɭ��I�W�~j 2�P�KEm��E��r5N��s�ٔHQʻ������郿�p��Gi��W"�F�,��F	Jc���zxM�L���W���rK�N�s�[ϗ}]q8eq�6}��y����|�G��3��֔��-yt�0��5E:z�ؒ����c��)t=b�cS�����h:%:Fߠ�-��O�����QV%���v7D ���O�f��dP��&O���cЖvη�.Q���#fq���v��A��2*��D��}���^�}���h� �'��ӹY�Ϙ\�ڍФp�5�/�RD����Zh?�b��]җ�MwA���ّ���,L.G��дy+a?v�w�ӑ>��m�i k"y�n��B��K��c�:UF�wvF�X/�_�GO� w��T�?�V�L��!^{���I�< ���� 6+<���JMD:�Z�Vzo� S��ux�Z�}2{�Z��s/��V��<f_ ��W��Ӭ2{�,�(d�fC.�����opm�j7��JlE������g�k�ߥ=��%�$�Ⱦ�"�������9��ȴJ�[H��ا�?.�*�l?����x��z�"��M�j7�"ar�M�ī��>�$��Mv��7�,�d'+�jaړ�̃X4�!.�֨�~1<!�p���0���u��z����#�����׸����4��E���W��ƈBm��6W1
��o�:�[�8�8A#8��8v�wHA�\Uֺ2y,�>h��ŋ��J��~G���Y!�Z�JuU ���)�%�8��Q�-�M5)T�ҕxq���Km�n���2�ŔT�ye�J��xΏ�PE[Ӂ�t�_zU��u�M �u�;�$���?pw'�e(J��a�)�mX��2Ș� ���3�7��@�������1�y��^�TIfPX�s���S;R�ﻶ��"p Z��k[�"����M�A���������r��ç���!h�~�@�D�%�1�IT&|�:�mօn���{U]�],�9�M�u�q���i4����A�K�p���*����ȣ@�rB���x�o
yQS6���+�����$��^
�|�6�&�r0fHm�#6�Q�ٮ=o��P��x��Ȑ���,t1���'�NC�ڜ8�#�ڐ��_�H9��/�!1#h�v�����G�?�X$���༢}B��@=��ޜy�Z�����>�(]�s�a���9%k�����M[z;^�`��jQ
�*��W�(�35�H�Y�d�SC�'��(l3~*��gi�3�L@5h��#myd���+z�����[����@'zg-��_�Ʋ��D�V��֭s��(���wS�=҇��[^����e�4�毫H<���7.=/�\	Gp�$p�3�aZ}���ei܁����\��[F���~y�X�3�4��٘�dΨ>��{ݐk�R�w�@� iK}���q7c�� ���90R����e���G��y=���y���B����.��B�#��P������6y)�q�.T� ��;@�i���;���C�Nvj��%�TL�qV�%9�QD5��l�m�D�`4�.�HzAZ_�����H���r��Z	 �pŹ�;�X�1��������ʻ'p�A?	k^�v-���G�؆Y�c�Y��]y�k�B�U��������a�I;���{�wʂ-(��}"�ӷ��b`����ځ�H��H�.6��<��?�9�k2~��afr(�����=��K[��"C�ӡ�xy'sw�ŉ�lyݧQ ��H1�s�|��q��_}�~
:e-�c��F�a��e�籔i�W-i"�q-��0?XǏ��P�a	����Ӵ��������
}B��症$$_236�aˣ�;K��7��Q�.yy�`v�,�8ʞ	��&Nf�[J��-0I�\N���=��,M�rխ�T�@?MYK�Fv�$��"���t�-_��1���y����_7�(��[&f�����+3��FxSRUo�w?^SϘ�e�7�bI���a��R�\q�&݇%尪�L�.�$�O��L�=4L��{5�����L;-⥥��*�O�c�x-���Z�c=��Jz��?l�J���i���I�O�G���n�cz�~�ہ�`Ԑ�o��)���f�5����$��[2X��5������3�'�v����D�a0oLmF��jV3O�,L��'�QU"��d�t�t���9Oak���@7'�9�Q�� ��MU��Y�F�x�%4.�_�>_I��T�����a���E��R�Fv��=u�l�6�-9"+��a�}DK����0�%>~��7O	/F����I��o�"�zi*D2�BX�F�6f�( 1E�kũ�8�12b&:�{}^��g�d��n6��q�����'	S5��п7�xڃu��+���-�M�8��[�n1�h;�a��݇��k~�N.���1�)�Q7͡�[�v�`��Ƚ�
<���V�җ�[������ާ�AJ����ՒNA�Y�&w̲i�v�\��A �4T�#���a���A�Q��$��e����Y�h�.^�=({�����:i��+샸���s��yX��#�%�Ŭ�jA;ʏ�y7o~j~�3��(���Y0R�$w\|0�^&Nڭ���Նj��n�<������Wn�Dx��ճg�!_Q�{��("(�m�/��4���y�tL%[:T4l;���V�S��0h�;�c
ME]͜�(�3H�xͤBy,��K3��}���a♨�e	,�Nw�p�gT�J�nѱgڀ��	�ħ7�ƛ�9������u���z�$�MYTh��ؔ�ک��g��PŸ���=|�*���|Aש�Q�������¯�K%�Bv��{�T�����,�c�^�TAʆ��rl_�ycw��|NcU�tӬ��������|z���w��ǯ�30l���[j&���5�ӫ�?��4��ǐճd)�Ʃ��DX+/Q/JqP[e<�x�R�h���V_��8�@��5��u�>��}H%��ֺ3�a���t��?��Y���,�ɫ��P�!�#<j��)9�	MA=��u�����XݚTܚ�Oy#()�Z1Ҵ- �ӊ[��J��p+��-ۻq�g!yE�B�$��w6�7o^�~:��"5{��դG&���q9�bQf�,UGJ���
�
�j*�4��?k�(����oמ������V�(�D,�_\3��W׫JE�>w&��7��� N�d�׿�q�����"�\�y!o5f��ԑl�AC�L� ��Ȓcn�_6�7ժ��؎T�>����:|OFr����l
6L'cr3Y�"������ym~����.\7Tf{)�h�������B�i�zp��U��~G�"`�^i��޷��-\g���6Cn����T.�B�?�-��d�DMV��� ����dX����F�XG32�c��F�ts#�YړޚurV�6)0]�����27~u����XP'�)�4k}m�|�!X�߲1Av�5:�P�M�XK��(���[\��E�q��H����xdQ^�||��7�TU�m�{�'��j3���v���Qh�"��.��CF��.�c-E :�1�F�Gl��Q9�]�W��CT�RU�Y}������+㍜vb��X�
�u��;!�,;">CO��R�P�!QJ`A@��T���16-y'D�=޸�<�ݵ>̡oL,�i��PV6��
s�V1�)��0-���m}'g�m�K�T�!<�9�#G�Ӵ�]�9a�u�TYL1/l��ok���w%k١>P�$^�I)�D�����6�-5�p_�TQC����tt��<���hɚ�'G�.���oᚢ�,+3N�U[V��W���4���g���n�jg�&8V.�9����<��#P�"�h<�L�G��袖ۛ���vY1��
y�4?����|�|�\�d�qcUGK3I��Eb`f�4B��GL��,�7�^f!m�|�7c(��mjJ�8��4 X���z�0]�5�y�m���|g�(�s��7d��%Ä�Y�z��!��4�<Ow�����ݵ:t�Xi�k��FR���ouӷ��d��	|A{f��O��� mҠ�5K�̂��G�k�i�µ�J��`�tA ����O��Rq6+>�����t���@�Q�Ĺ�=9Wx���:���F��z7�m	&�k������w �A*ZB�� ��
���w���b9�e��P�
=��nƢ��P����/���'=,$���Wa���6���+�j����3ޥ_��7�+"G"q	|�;��_�����������o��:�YkH8nx��3�<j�s~?�5R�)��@�����}+_��3��ӵ�U�3�6���!�H�3M����E �Ip0�����ȣ��!�lS':mE�R$��핋å�����rt�/8
���Tgd�b�UW}1G�P���ܻ���A�sN��*���qV^�����~�t��bċ��س,�.~sX�T�9(*��woA�R�FJV$y��hO�=�<Yڱ��F:~�\y�X6�,�l@T�"��ă�W!��l���]�}�Z���h:��S������t�>tm���מ@S]��VvH�"�x;���#<���/r�� �L㾼M����cn����>CF�+���q@���Z2�]�z��~Y�Ի���m���(��6�X�{��R��/D��ߤXh�Sk ��^�m��sT�rC�9�C�>j{��b��� ��/�w5,��}W\k��3���A(jD�O ����.��b��H�ږ�t�y���E�Z^ړM�Sm#�:K����"O�[5�����P���\%%�~��z袔�D���a��,��<�Q��n%R�^`��4eʴaaB�Ǒ������#k9c*`wkW&Y܁��&�;u�{�n�WOe^Z4��Q$�M�k�a���
�T	Ч�$]^������p�|Py��^��=��mX�@@�u���{9G��9>2h�Q�Kƛ�X�w�ׯ@rcr�Ȉ�܍�b�N�S�>������I�kDn	,��Fl��P��`�d#kW�o�t�\I�O���Eir�*8�t#�g� ��B��
~>�jAe"���E��POap\�h�y(�ے��瑇6�+{���EUW�6��\�ǧQBks�~����0��jP�{��
��8���anP��Y�G~�n����D����o+�u��j~o�|s�pyN��86�=mg�)A�#ڕ�==�sЊ�A>4�,]���4D�u�𬻄G0M<.� W�I���檒���� �/�����d�H4�����������c�����Ɨ�=Y�#����
j�=7��>�X���S�����"�E|M���z�,�*k]>vm.a(r���|WIT0��g���:���dF���RX��`�ZcZ����s�[�i��G�������D�Kl�u����^y�^��M�_V�5۫�)ߗ�	�Z�m~3ܻ.d}؆*�'��{�+���26��i�����%l"�:5~1=p]Z�76Zj��B�
����kXs�R�{�9�l��ٲ<� ���%P8D����Pֺ�O!��n�-O��N]�::8�W�5D�&��y%�^�]��Lp2+��םӛ������8.�3,�7��,�����r\{�X���<_����t���A+��M���ě�R3*�����C?]z����#$��ϩ\����c�:�6�\�q�o�4hg�z�ye��a��������7�h$t�M!��*��4�~�;�:Z�b˕ B�j�;�æ�?���\�s�fB>K�tF�K{	�i	WP�x!tס�J�d�K"�j�����>�?��q,�Y�~V���tK�hi�7�rLf�~"V2��~��e��Ϻ5[�(޺�� 
��x���gr���!�B�ȟx���L�F�G��GEdN�ذ6ɋPI��9����k�|��B��7y*ߪa��3�C~�_F[%l�6���i/((�̀�W�O�&{Jۍ����zz?�jL�g<����	����^�s��O;\�
i�+B���8� �S*|�{�:�,����
��ǈI�b�����&��;�@Su�zԾ/D�Ʀw0��wG���o��mC�=����	};	�b}�t�mL�9?��|�-�&!�	�t��mB��n��p�