��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�k�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������H�W޵α���N-�`��6����ݾ�FF��eF4��_}<�ےA�[,�|{�?r+-��]n?���A&Q>�Mx�E��K֎�>v"wTD)3�2C�
!h׮X�L��,�kҥ��o�F�=n�Br�W��N��7j��t"�z�b�^�C�U��IG����ZyWH���?����2�16��'���TY]�Q⒱�?���)~a�����#�/(��:a��)õ]��Gz�4��~�=��N<̰�A�ѭ�'3jO�Q�㷛Ġ��㴖�ldlE ̩�U޵�e�d�ި�8�����٦��8�KUEwyM�8b"I�AP>�E>�g�{a٢�T�E��Q�@�I3�:��;ub���n�|��;{��8���q{Է�_��{q�g�9jxr'�b���`�%���)H�-У�~�~E.v*4Ҏ:#�����VD8���ׇ�;�"U�>f`YCR1���-�ҝ�<ŐU	�����&�TgN>�%�Sﻋs<�V��
g�~�R�Ľ!�S�4c�N5�tZf�hx	��OT/&&�^	\*�ox� �2�Iyֹ7���<��t�ӏ�P�κ�{���|�V[b�m" F�*��'Xp���f���LK��h>4n��@sz6�`YТ Px�F�v���G!��xk,5�F{/��]��a��pC�@X�Ao��� '`����/���]`o;��lx��f)��le�q���H�P+����$l�@�����q�Xj6Λ��7T���`eׁQ���kl�������5��+���W���1?ٯ�D*BƛߖvH�r/�w�o�N�hp����%=2��슎����H�1d����ƅ�t|+~:��HY�W�:��6�|�� M���:���×/����Q�R�����X% 5�7g�~L��B%w�S��O��J���W˧�.���Q�� �ԡ^�x:�6��1N2�iW��O����A�<����U'�\�,��������w1j�[���	�$���Ҙ���mS���N`��u�nUw�ku,��1 L8@��ؚ����}�0�1�]2|�ޏ�ǀ,�5��2I��7�T�m?����Yn ,�g�sF�_��}q��V|4�!�'I��vv�/qb����T	 Q�����>�"U*���Kw.E�? (&���@ \9�Y�\���, y}y���B���:�?�&LY�{Ĭ9��W>�w�c��C��r`��S�P�Z�\?����%�Zoi�:̛��<'?.��l��P��gf�7��p8h�8�s��d��n=�+3@����h���O �(`���Y�ٻA0�Gꢍ�ua�Hx�����^=���=2a�KG���ޗ�5j�'UW�a++i�p
0�Π��Q>
�M$rB�W��-�E���E��*-0��;r Vf�Șp�4r�~8�P�Rq�C��9,�+yP<mpH@:=���p���쪄�`���4j���@�W�^k#$F<oB1˅�g_�ד�q�t3{����ϱ(�R*5�m^�:C�[t�,Ys�Ny�u�^�sXk$������#��'��c+��ysI׋��~��f����&�;A�Q؋v��4