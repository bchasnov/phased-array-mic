��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\����q�?��e�I8�b�Ǽ$��"����ׯ1�V0���DO�B�N�^��y}'x��˗�ʦ{���q 53J;܌���`1�${���}�DV��J�>�J����&����^����O/�-��(ΐJN&D#�2���R
h�tt����>�$�J;�
�o�֬p�t�����S��Y�/jֿv��h���ɠ�?��6��sϿ�����ys�i��KYȲ�8����ƧX��~�;C��k�`��$�������P,ו��믈�F
C�H���|����%�Q��@�n��f��
�D�Y����U^L��~O+�� �s���sP���*�]���h9�`.�Y /��SCp(�˲���o}#v���1����u��SR���֢�;�	�%���w5�i���ŕXx8�&�m"�Tu�W�&j>�rjR�+{5>+��S��ɓ�������\+���싙1ne�!%��ޗD6;��Z��"��۽F0��F{�0�����as�z�>���jC��
�.�ۖ�N˸�D!����.�Aqt"	��:xh�U]nJVP�����Kz;YRu����x�0��$����U�~^�^�ԯ0� M-�Q��Z2s!��R�]1Ӽ����	[�2��5�Qv:�=���;1r,HH"o\�4�=m�:nI�oB�s��¡e����>��{�u7@�c��g$ 7�⭆��œ�a�H
���Y����q���gU3�"�*����?nT7~�n��(}�([��IC1x�9�^�8��o��\�bX��N\	�V�ɰ`���_C���GO��m��
]%7�������i	�����U	�>�8ֹ=�F��d`zΣkɮ�o�24"V�2 !S����q!ջ(�V9�$p[)C���\Jz��Z�"*�HUiN��J:�*���Q��9�N�v�)�j�TDƚw��B�޴���`��Otpu������	°�%	T��aO��.�\�

��]���qT��|��>���S�ᘞS��ͱ���BzwB�]+����ыH��8Pqk��#^��i�d���޾}l<�m�����n=!r��].Js򟅺�����f���]�>����N��F�ˇ�W�͹�!�"HXn�'U�������F��_+�yY���t{��4s��)��k���p���F��|2"�ED
3��t0�F���"�5���5��`cp�$�t���j��R����8����*���/-�x���}G;j$v ?�3b;
&"�;q|�ɂ|�Rf ��V\��HW
��ukx� KB�����g�sI�ƴ��0�4�]���cRe+���Bp�s�ua�t�j@��N3�f=��_�ׅ۔�7!P�1`��h
�-���;�1�	g��ve��{ʢ��ixO't��3����g(vXp�~��(��;�)�M3�����?���׊-��|�����"�_���o\��.�͂-�X�U�g{7J�����Ck�$F@���4"�~���@�e`Oǒ�|�ѰO�{�z���K��^���Ue�렧�馉f�ջ�z�e���'�	���9;LAQ@Ъ����'G���*ET�~��ܗ�U���[�|E-dw���!Y��<��`̎�r7�u�o��E(� N�R�9F�t{m�/4�9����
��i�9yH91�6�����|AZ�iW)K��P�5l�-��;n���W\-��D�}t��JW'�=f�� �G�a�C�q)��O�P�f��`{n4�4)�`�q)/��كޓ5�%"�L䲬�V荻���cן���4=��5�� ������}��&�C�5��Hz�^�S��$|��G_03�Óq؄�)�P��A[l��B5n��d5��VQ*C�+���#���Y`>��V �AU'�r>7�h$�9f���c.BFf��,�s���S���m���5|���R�����r��:��������	���Y��s 8�з+����J�	5Ԋ�W���1/0:}L�@��\� Xu���xә�
:ώ=��k4�����yP�Mʻ��>�7.��	Y���!�0Џ�~�v��_��/�
o����P-�K��5���� Xjs����ɚ
X/�qH�E�h���\]p��'�����p�bn>�*Ͷ�A:#��q{��ŕ$nv�/?�nI�1>�:W�ZcP�@�3\�;/Q�x�&�����o�r�%>Ћ���'�o�ʬ�M�O��H\6r�F8f�:� �%�g�:���/e3(r�,�0�Y�{G�G�^v]��ɛdeL�Ϭ/"�Z�O�i���L��N��,��!Q�1%�Q���� �|���p�F5����H0����MZͶ��R-f"�{rg�N>������y�2�t�]�˒���n�6�Y]���ɜ~c�
F�/p��_���lo��n�%���@�VM�Û!?�ܖ�NvU��b����S�(���@z4����Q"RmU�߄)����I�8!'�2�����<�:�>�ypf�KL��(泡W��l����yˤ�sJR�+X�Ơ!4��0����poC�;��W�|(�\�v��{�*�A�WUl9�Qf|��������S"��=��\�J���1��T����>������G8�� �A5*IF~��{"���T{ ���5,Rl�S[��O�jO)�PM��i�ky$;�ǿAeX&� �Q"��nP;
��zn�=�����8.:���C�n��V�_�����������_=2�	_�hE���� !sP�.%r�� ��y�Fr��,�Ȃ�c:÷�8R��d� ��=1��D
:+el��_E�8�h_���& LR��	���8�L�x��-R��e�/, �2�]��X�5'^�5���׳�߀����]"ǡYܗ�3�I3�2ւ��[�F�都�E��ת��"��l�d�jZػ��d�
L`H+�*9�qj�Tś�D�ҶuM���|�5H,7[َ��C|��:Wf�2�1�n�����k�m^�Q�̘@Ql�����i�~��Zz�O�:>yd9���{�HOtN��3��6X�2)��}�J�R�u	�����=�58ͺӮw4���c:�
0�Ღ�_��s�ە����}ۦ�w�|V��oe;���CR��'��[�C�1��� �s�Q��Y�$u��-�N��������W1�x�/S��e��^��7�#�Ź
�@����WG&���OZ)|��[hKKn.��aA���b�m�&��,���l���n�P�=`Y��]�q���5
_���F�QS�ߜq�%e*�$���M��R��]�i*|�ȀTQ�U�G����e��X��j��a�Q�	e�`��H�@cF��'�=�`��*̀>�G-�9��X��;aH�k���"�}Ҫ��\��t"�'� +�wc~�f�#�T�74Շև�ݸS3 o�y����A��`�b7�\�qS���R�d~'9�P��ԋ(�W�+7>�R;�0{�ہ\f��5vD�0�n�4���
�MY����+9/�����>`jC���2�_[:j��b���:�{F}����uքa	j9 <��0t���e'3�}�<g�R�%���0�T��=oCgH�4�[�N�uc�`-�7 (`z%}�m�����e�G��۩H��?}�u^�~q�z%�4��V73�ᵤ����*_y�Cw}��m~���9n�13�J���U��]ӣ�� �XF�&��Ur�|[�z*�2D�MP�%c9��d�;rV��x�<&tYU���L̢��R{O�z�=q�d�Z��pbC�%(6J"�������f�e��j�|��� #=C�ج��,�U,�G�6�b����u✜X���|N�ϥ6i�Ł:tP8�&�)���@V��A��ϑ�܎�w��O���.�<�ϳO�.ȕJ��&���Z뿜�xK^�?����kl�!.�m��[n�u��Ş ��b���K�Z�:ݻ>�
a�R�j1�y��S����?�	(�Aaq�Q6����o�hj�^:��O٩yx�L��,DpȌ�`��t�A�r��pB/�z�~�?���).��^xtF�f��rRJ��=��2σ��Q<��%X"Lm���\��/�������י���q:?�}g�F߅�zo�h�6���5 1�fΙ����qng)�k��0@�]�'f��]:�IjT�i!�}���{:D�ܷJP�e�/ s�,N�����Xg2�Y=V)�^!�n�ǃ�/���7�(���0z 9_Z�(����d�h3s��k/��+I��&�<��@ʒ��N��'Kbf	гE5�_~V:z����fO�X�$b��J������;L��u���=�x�& t)T�D�!��/b���~#�B����o�#��.�BV5�	4�`�C܀7@SN�B,��)\祤_Xԣ}��X[xA���T�@t�wh�9K��;
��b�l��-N�{�|ȧ�ڀe��$���Kp�N��UF�@���M1��;@�q�B|�?�{��p�u[���>j������x�:t���;i� *��x�����{)�*��¯���`���G�7r�	�m�F��z�`��S�a-oЈO��BH{�!uT�s-�J>�_#��f-�O�;�>�b��7�H�w]��?]�}]U��I��x?=�_7w�9&Q'ϋ�'C�3H��Av�S0	Hy!71)x� ��=Z�]����� L���w����Mٲ����;\�͔B���B7\�I`ƚcq�UOm���H�c��˸9>#���@ID�d�� ���(9�c���~<$O�m�h1�����O� [8k,�����?�}�Z4{�{3�e��%���K�� ~��h�=���#���><�Z��df%2��/�z��՚��a�j�:�|�V��]�\��N�c,q�@R$kx���+��Y�yn�]L�`+Oo��7�F<�p�;���&�E�x�ҵD�KCA(	CϏA����Go]�q�b����@RV�)w��djRY�	�ª�f �-Φ���V�{�b���S��q誫H����l�_D[
��L&9��C��j?.b.�f���8��ѕ��(0]B�=�77@�$�J�4�Gþ�ʵ/��w�bIK�5?�gh��V�h]B3��ﱻ��I �'Ѿ������%kv �e�|�<r�б��m�ؔ���ewf۔���I���܇���|���21(�4M$�<t৭ALo��;���3����9L:�`_`8�>��#q�<9Z;��Ӈ��j�ֆ��l�	?|R���2[nn�T�P����F���i-��.�8q6�t�Zz���C����F������l��vWx���A\z��sT7ݸ��m�e�4�k=c��~#�B��wxo�'�D�,+7O�Q�՛�-4~l��� f;[��y�7��ܴq�ʿ�j�1h�X����K�z�X�	��:���
�Q�Ҝ:	n�Y��}��"���h����y��j��J��i��P�2�JWV+d��k~+]���'�dF^J+��YW���f��i._?f�O6ab�?�"'A�5AO��*s$^��C��H�F\�#�&ԉE������b���cn%"�;�R�l߷��C���Hߘ�s������z�X��l�B�� םn�*N;_@T�p�c�I��������S8�����x�Ā~:z�����'�'�4,��K��g����u��r���ȟ�<��O�Ȁ����$h�LѲ|�+0�{�a�m>���N�Ƞ����y�6'T�Ͻkcm��	n �� ���� 
g3F�OٔP�]`��Q�2�Q��'T�Q�����?�p�L�Z�:e��)��e�<mjzHT86�6R���x�:�8����_-%jv&�S�d�L�
R��D&�K�ߐ�)���g�f(3��(��&)���>e!�z�+Z�n;��L�1�9��S;��u[	�����4�]�[�}�
0�������B��	rh J�^�����w���E֘zoP� t{;I�<��ċr~1��.��h�����Q2���jG�0�?4~<��ambK+Z�	o�৪;ki�=ʇ��u�|�][a������MB%�����]����A�nC`�} 2��Bи%Hq�r& �}*�Η0E)ǟ��$W��럨�f�Mt���E'<~���F�OCQG��n�j����$^Kx���oetH�gy�&�?�)��\�x_á�uELy"z�m85���_+}NP>�l���֨�GaN�55��Q:��������)?SpE�<�,���Rb�-�d�Yq�k��C_w:"Ah��e�o�36�V6�S<��V�V�BnpH��x��Ű��J d�<�D� c�s1��(�7>�Y�ے���!:�,�kon?�;� Wf)v1wF@��B�������4��h��6�	J���Tr�z~x'�,��g����@D؍��Ӯ&c�L6�n��S�
Ĝ0�Ӄ���Q<���8����~�)�4��[����fM?��.���ˢ]j;�v��j�<<���~���:F��	�&y^"�:-t2r|)]K��^W����hypv���F�ϴ����������֨�2�����̄\!Y����E,������e�y��	t,���^��؅o;ـ`bD~��6Gc���2�&��b�Pd�nI�$��S,����N#C;�� [lr��AG�۰d�'����s�1Ζjڦ���8w�|��-<�p���K���a�$b���� ��l`Ll��ID���6`.�UZ����o_2�a�p�kr����br~b,H��,�.�\��y��N�=�ӜTUQ���*����r�m���	~XeSO�ݯ�C)�]� 7��pM�Ft���ᒙ���eE���ģ��� �8�T�8ڛ�q	&�^sM��U,-�t��1�3p�&ȇq*k_~��>B���
?0ɵ�"���pT7O/�M�Vf;ψ��%6b����}2�ĹX(�A��;�E����7C|���;|w�I9��y�+5�o�qw��C���w=�u!Q��M�(@v�y �*ނ���gp�+��~v;�����@N�{Α�wT�� �H�G���j�aKK�HY�a{��y 6���o�d�\�,�������Z��k���|\�^�A9�(�RWhJ�cZ�dP����_D2aR4��9���7���1�gvH��������ˋ���l�?�r���#�S����ۨ@�/I}X��y-���� m�>SA#EFS����+��^g �w��޹з޼��x$A(q %A����@�������0H_A�S��C�2��ExH6��v��cJ4�t��A��W��s&��s��o��lth���/��rτ�ϜP�ܷ�R�&Lfw��C�ق�[�� �Z��K���D���1,L�f2q;�3'w�`�l��kŇ=�<P�9a��%���U�ZrH�9���es!��E����+����۾�7A���f��y��AH�W�Z�$�˹�Gl�Z�l풼X�`�%�r1MF��J6b|�g\�'�Wa��e!��Y�̯މ�	��V�^_�%�U��vFNXl�m��������h��Y����\R�'�g�
5=<5^���x��(�e����D�)$�E�/���7�,�K��a�ʓH8��0�����S�9%C���KVB�����n�UPG���l�E� �I�;���6��j�:���VY&@��A]��./FV���؈�X7�BF <�\�6��d��e0e�����>U����K��"R���F ai��e:!���f�i�U�b�� � �kǹGl�� D���p�����;�vu�b��	4O����,(0Le�Cv  S�7��2[H-�J��!�Q�a7�I �i�.�����1��������f�[�xW�����	lL��K��Zy>���7.R��F�s�,�ʜѶ��i�KL^���bQ��2	s�|���*���DW���u����-뫍�JP��$XF�!O?�J�OŲ�R�{se�����"�D�Uko jN�i�w������3C�*���T7���8W1���qQ�H�kle,~τ�(��w#n@U�B���!�.�� Q��H-K�J���f��q��R$��.r
�ld�p|�-�S���	_N�
��X���yp�:���M�ƨP�<�xs��ֽs�g5£o�#-RK���ۂiP��'�*�݋X>���3�bs@*���َT���h�5E��Ӗq^��'r^�x�d�����{�<��A��2�fږ�W�p���/Z�&�p0��x��cSv�����2i�Zt�ޭq'M;KMiI+o��9�:Z؊O�����I�8yZ[��]�p�Cx~S�����]��-�&B����&Y4�|z*�Y��upn%۔��h;��Is4�n���p����3�^�Yn���iK̓1��"\�p�#`�@��f1�Ή�/[撗T`�uJ)p� Q
fd�N@����~^��O��x8��P��`��jY�I�O�a����{��ݗ��GU} ���z"�׈�������
�7�ZWț*����iAt�� ǁo�L��
���^a��}v���A@B��m�����F��c��7ࢤvҴj~e��O�1]���s���ے/ql��ޣ���;�g��ݝ�2����f� ��2������
m��H��Q��fr�q��Bj���o�<�c����g�|��!�bW�Ep��$�7.x���%9s ����v�͊��ڸ�8����F����Y�(k�����B�eO[U$�@��L�?��1j��� 	+�/ы�C?H?���*
��-M�i+���y~IF���CZE.�f������9��W��6�]ٹX]�eW�e?���=ہ��6�Q�v����[�
�J���Y�5���]:D���J����Xf�Ո�䇍B��O:v���>E�A��.�Gҹ�g��I�|K&;�
�2�Z�Gۺ�a�5B�����h�/D��P*#�K)��y��(��X�1x����t}�6Db�5dݤB�@�c暐ަ�Ћ#F�&��2��[QUR�N#��8���Ώ���3���=������1�JrK�n��q��'hZ�%��G˔t���(�>A����7T����醲ۯ���W����e@#�����g��w���u�r���ȅ�I�������}d���Mof�DY�uKWҭ�����RɁ9�3j���MF�b�t�gK���.W��t�a����g�]�A �G0h'����jX�l���� ����حRu%�I�����Jox$`�����ه�B6�XG�K �t��;�o}�3�NIص��־��$cd�����>���&13nF�6����o�����x���Bi$9��m2��_��ct���
)�f�N*��&;��t�Ĥ��<�4�R!�		^-塯��3-��!��v��8ϻ�KN��c[xge���(O~6�;V�;,7��ޢ��Q�e���v�
�O64��9���.��DG/_}�ӊ���ЫP8d���>Ɂ~a��i�k�O�J�:�R�H�Q����xg�wUPݥ��(��IP^�wM���@��ꡂ�3X���7i;�(���~��
B·Y��	�at(��f��SE����LЋ�>K��L%%�?��/�Q��.!��|�����򣲝6^�ZK�K��nۛ�c��<#r�*�y���ʿ�{X�4O0t'-t��� �yФ��;7��d{�M2s�lz-'N_�H��-%�S�V��Ӆ��nb��:w�&@Τ�\L��� ���С���'ɜ����?n�ߘ��67��qQ����N�)P�P����Ga�N��*!��$�b.?��\bl��Δ�w1��̌��==�+~*6�+h�wj��N�'e;�-��ɴ|6���c����"�X�@��z�E=oHxs�)�!� .w�5�ڨ��q��۫��?���ϡP�Y��A2��&k�����$Å��� KC^�v�fO��3���dm[�9��e֩��)��G8z�����L�=���Ԧ��Һ�M���&cY�-y[��`�p�F:��"y7�>��l�Mn��QGQ�s����<\B��qm�Fc��Z�[��Р	me��7�z��/B*���C��j������{�x��%�%�k`�I��4o�����H8v����ړ�g�s�c�r���������W�l�-�s|��GFb�ł
����r��$YN�"d��1�����"��M���l\�Z��gd��.�u��`K�ݤAa�d֢�v&���s��tb��}��5�r��9׫��T�RvQE|A$w�����_�s�3?�4@�TG��:
�� f8u`έ#�ǰ^���$���}�Ҝ�u�������k��x�F[�f"Y��o� o��/T�?�lP�b�/1�t��6��X��X�Aơ'��se�?vqO{��l�Q{.qG�D��ځTl�4�������P�J�Z`[�6�����'}��	5���Z1��Pl��%[���_~�x&[n������6���|�7ْ�O�b��9���'�]��]����8Z�?Z�'�`�Q|�~.R%���d�m�-R�q�}��o^!J�E몪d۔q�jʻAL^
>�Q�%)g0<-QNۺTx�c�2�kQ�J�!��x��<t�����s0Cd(TiMפ��:k��0Sxm�"Ivm�ĿG��Zu̔D�M����E����w�s���*s�  aDD�&-^��bmw���Q��%7h��LZ��̳�lY�?��F\���M�C����hEA9���f%({�	���g}-��'��L����b~�L�;���g�7��h t?�s�=�?IS�R��.y��<�Z��dG:/��y��À�Iw^��-�b=�h�DI�m�䢡��E�lm	���_q���	b�$�y<u��β40J4��Ic6nY���
��o3 h��Q��Q���B8�s�������kG�mA^ӹ�0�W;�X���jx�lT�)�<v�a��U���i�R�A���
8�\��;s�%��:w�H]"�oگ�t����8ۍ���o�;�e�T�ʭ��%�4�M�ش�O���u"���l=l�ɀ��x���U`L�8�'�H,e&�w��N