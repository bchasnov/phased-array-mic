��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!���"WYj����i� �N�7A!�@<e�]N��?�jj�����W���a�q���#����MP�F�pdoF.8��+:���h1�ԭL��L��[j�1���߀/AP�0,r�F��x�N��>�RziB�M�\�P�ua��B�MɥBe�U�����v��+�R��|BC�:6u��8�B�����趟���*���I�lklry�.T����b��`��qe*@](���R�Ե�3K�i'3��)Kч�˲7�w�b������ᤂ�������]�:#��Ǣ�c��z~���%/�J[��P���&�Ӻ"�|}$ �n���[ߖ��eז5.�8��Pi�!ػb�t(�_��Ė��z�����:l����[��Q+�#�L� �r��V�	�٧3���v���:pZL����R������T�q#�˘�8o�z�d�D��"�+J�(���E��[z������3)�l2rM�Q��&TK���T���4��d��gf����<�;�#��:I�3���^w}��d/������	A\Kf�(�-�^�d��:�Y��#a�5��6��G>���k���?�(j	VB���]�̯˽���]�7c�	2% ��ۉ��<~%k���C���{_TD�����q��T�+`Q1�6oC���XO=��I?�4@�������(; �[�RS�q`�l�ѪT¢�i��l����;}r�sW��l�l0�N����3ն�x��o�d�rr	�r�=z̙�Gz6����&��s[T��c���\�&tj8c<�$}l�z������b"�b�����q�&�Y��#���}��&?k}�LW���Y��vΤz�ZaH�GO�DkY�
~�����hc��뙤�}�h-�"�!���~��!�y6:H�a.~Jޯ�[��!׃!w꫍H�^Y{�0�q\�ƫe �e]I�1���Y��[�%���톒����ڏu}9�1���o�$���}^H����)�~��>Q��u������%Q�:���\����A��Fy�4I�;}��@$��V��G�r޾�f,ƍʐ~z���9��"�)5�|	jk���jD�!�@��j���1�쉘�m
����r����;�����3�d�g`=�}r��N���r���z6A��p�AX'Y�!9.}R����p��vfKw9�F��:ORA�?A�*h=����ލ7R�-�n�
A/}�q/fu�Th���~��� A�~sg�����`)��r�RI�K���Y�L����a�BA��X�:��敔v�C���>�0�5ˆ��e��� l�=�,Ƭ���k}��Mgj q�ӄ�	RT���
|u�ݢ�RQ
*2lx0h�<��ߑD���[*���d�C@v/0�������������m����jNq�����`���h�,�A�����:Ma���iU���<�E)�������/Y<K�6	$A�TXa{5��ݳ�#to�&����������,�<���`�T�Xftc�t:��{"f��Ϟ|�4'7���&�Q��y�1���!�/N'm��EU]G����Bw;����`;h[�����]�'n!�����x�����G�M����hv۝��M��36$��|�}+x&'����D3^ٜe�|-p�	�<�[Н��&dbļY�'�3�n^i�{#�D�	+W����D�a��q�a�̍lIG�y�hS��^4ǤO�%��V����a�)�B�Nen��[��m.
\�K@-2��D�����ZDA����0"����bm��[��=���~��ž��qv�+�������V�<��R��V`�Z��id؏�!i@C�1��3XRaܓ�g�"���J�~�<9�>o����c�;|�*�+sj�����9 ��r֞��}����ܱO�nf�?�]�ʮ�L���>�2h��6����'l{�ǥ��f�ȉ�����k��b���86�̓��|�B��ր��T���ّ2�V(����g�}
UqW�CK�<"�7Ն-^<�Ȳ�X����5�1Ua�	
BR?�S���&}q�lX�A�/�s-
Z�'���f���1v�J&��nZ�}�cZ$�$�;��8X�H˦Ka6a�؂��7#�� 6� j�f>�M��`�<޸���q�n�n����&&�X	#�t31����]��p�8q$A-�������	մX"���[^c����j0(&�`3�.J]�f}�{B8�<�{�t��d8ڏ����S_3M�Y�W���H(w�qF;ӳ8>�Tb_csJܷ��n{�$fD�,Z��3{�M
A�L���@ǽ�<c�`�b1D����[H?$[RƲ8������:�my���W{^D�c�W.�C;��'+I����8�?3N�<؞�������5�!�Pw�D!�9I�1���.b���664����[O�mg� ���X?�:>^H��,��'W�قͽ�C�� 2�iBQY�W@��*��=�������^F�{���wL��Mҷ6G�I����D���1>2��,c�J���l��P������bHS�D�f�vY�k�h��}4=�$crFh����v��D,� H���$*:Y&k?�>����n�`��U���II� �`"���\��S1��8R���H��Y�
����i��E{�#��S�v&ⰾ���v��
@�.X�;!�}h�̓k(�%9���vf������P�Eķ�{j&"���FrJLx�`��>�2��/�,��AŹ#��k�#��i(�l�"�:"�b�_���7> ��c0F �6vS�~)�e�y0�Z�'�S{ьq\	�*��>N6������C� \T��)����^),��)���m�F�(��#��m���b���A�8���J�t�o9���=��x���6����(]���%�h�Ė��K���zl��+ynnfZ=�Q$�K��i�q�AI?���L�PK��ȧ.���U&���L�s4|UՐi�زg��L�{&�X����XDt�դ���pT�
�4LZĚ�#������3b`R�Ι�cQ�"���Q���y%> S<��G_X PEF�!O��!dM�t�-�ྀ�A7��.�2�+="s�[x�h��ط�)
 CSy��2��bL���w%0��w��i�
G엞�`,�Ww����K/8��i��o�E��B���g�Pb-�U��x�Y,	�?Y�r���n�ׇ2n=�����$���>E�
@$��	����:u�z�l�Xr�������"�zz��[���Do>ڒ��]�u@��t8|�5���A��)�4S�"�D��'��ԎRkP�k��Iҿ�g	z��TصX`���MQ�8�VX����O��o?���z��.\��i#��|��g*U�4���1m�D�V��pcl��7��+�j_�n�`��jW�k��ǡ�&7�嬝ȥ���4I�Y^ѥ�~������l	�����v�u��$���X��\l�9�:�Kb�@]/�Z��`9�τ'�Y�#7�w�T��˾�*bf�U�2\�1��	�
��y`߾�j%n�z�'60������+ 3Wj/C���GT��i�򸜙tM]C{	���v�xc��֙7��3�jy2����a�j@e	�����yOJV�e�/�I,���֋ա��� d"�%T�����3S|�"�m����+gf�L��I�8��4�-���S�Z�i��t��d�����S �����f������&hδ���}6��6�.�w!b-@�ei������2��|A���7�]���o,�&�N ]n8t�/(��!4O��E�Vi�9�����ZHn,��U*l5�9��4�h����9>q:��3�d$�xJP:^dJ�r�;-�r��9��/��a[�3���{�hR�J� �?V8�����ϵ���}��iX�Y�Ǭ娤#w13ڿ]�x�'��de�]l\ ��ag�*ϗ�*�@�Ȫ��ښ#���VJ��Tq���V��4�ȃg��+����̈́��G�0��-q��cB;�
�;�쇺xm c��5��5�܄pd 	]@$TN\#��b�$�]�����t�(���%��{�+�=�5v�Xf�9�
m��*�&�o��k2��Lx&A�K��a��g��j<���+�|C����@�����!!8�V��c t�4����n��8�NPz���!<k���p��	7���im�����7?Te&��|>t� p��*)���[L�h��@l�fe����|��������}=�� k8a���X��ۈ���l]�3�
EɟZ7�C{Ώ��?�Z��J�ǡA�V��h:c|
��l�ȅ�XE|]7[��SO��
����I���?���6.�ŊE��(l�8��ٚ��� sn�8�{oJ�J�=v\�P������9�]%j�㜊��E~����a�[�j�9���u��w| ��i�Z��$1�@����,|��uIb�U�`�_U���QLI}�����T�k2)Q�6A���v��}��D��`kN�YE��4壩��k�a��Fi��F�-W1�Aۋ���B���~��ge�7�J4�B�Hf*�7��BJ�^R���4�	�K5T�BƠ9�k��"���6	�Y���Zſ�A'j�	�	��m*)"u����A=�Sq�7i{�Mc���c��C�C�e�њe���i)v	\	�ʍb�`~>�c�J��1x���\>��8V�)U��m(�
i}��F���rq�*���lP�L��'?�ړ��<FM�_�(�l�<���,>F|�w���SΥO�ͺh��n/,�YuM딖��؅h1��F��~�5"p]��k���he\�8�fSB�&wo�X�dxF�X�q��Rr'}�{Qi|[��$�D�b���r�i%�Hx�q�`��O�� e�2�b�x�͵
����������ą�͕���|��Ӣ뎦G��$a����nn�N�!h3���E�l�)̨ 3��\y3�y���(J����=~�!L���Ch��^ؔ\B��D^~����D�=�?g �g㇣�C�KZ7ܦC�#����C엘��2���o� O�Qժr��׎J�!T�̮�,�Vir@k�濁���2I�4L�K�&��� �A���D�F�xҁ���{ז������n�H�?�I���n�,��j�M(nv�U}�M���? �gB�!��{�X}�XWJ(�\���MưK��&���z�� {�W.�X���2h�ER%�]��a�p�\'�t;������kc��漪����N1�-rz����9��ãu߿�Vă���sR��F�tT�m�v��!�O͠T� �!5�j�kE�?�m����7�mDy"ƿ��Eq^�	H��\9 ��e�4����cK)Δ
�T9��,�f�l/;NA���Gmǃ���⶝%�U�� ����
ye|���b�c�:�%�%��{;6aj�G]t/�4���çU7RH�W9�Re�y{���M�JC_�g>vL�����b�0#_l���s|v�}��ʍl�(�A�٫��p�o��`�w�����|�	�`�EF�Q�fT�-?�}��S�+p��j�qA���,6��[�\[vs���8���m�{�"?��Z@���&h]�N|�9<���R� ��Cڅ�3����w�<�,!3�1�{%�&�sow55�j�Kߒ>K�*V�Vu��j�{N����M�m��'$���C��P���T�5o�N�3��=_�.�g��F������
�b|���t7�NŻN��k������^v��TT�������o�2q!͘2����f��ܡ�Q³x"X���ͭ�a�Π���֫�e�1��K{����qa���k�8��yTH=�\م��
�B�y3wޱ�ݟVp�?@)Nt�=G(��C?� �1�pv�w;?H-�1�h�Z��y���~��f�}J����npI�a?�
wF�Kr�[?���uS6���p1��I��g�
�q�9\����v���p���>cG��]�k͍�����q��?W�ȎsQ�]U�~�>�bP��5k��ҭ��E؇��K'��̺S��}��Ef"��[��3�9�^��)���c9l����� �r��/*����u]�S7zW������;0iϲl���ر/�Xm��2�Aq]�q������oT(k��`b��쪶3�ё�_?�^�`R<֒���Y�P��
S��g���`F��~���Jp���\�Ҝ��S�Uy;�B.�� =[�6o:�"4��'z�&\�����+��l�~��Tz�q/.��f�6��VQJ��#�%I�F᧖��?:�Uorh���5��Ϛ���.~/�R��w��d;7o¤~7ړ����Yx,3Ի<�y_����[�Y���6�h=N�uR� �A�� ����\+��s�8�@����_~��~�7"�5Ch���]eqX\DN���g���V
M[�&��ą��Ia�#7�e�`F�cƾ߁2���Lz�7=��B�9q��7z�yfn�w�={!���ϗ%~���[��_x@}���r+)(��x�Bm����Ћ\�k'Xqƞ�v�{E/�3�)�p�Ej�-w7�o��H�lQ�!]�� &�+���]���h�g&�\�a�����\��Nn*���ٟS�Lh������TS6U�Y\�Q1Aj�bZ-��������ͯ�E�2�3���!��Ԫя',�~Ɣ+}ܶ8+$T1���Z>�(�03|CJI>��������H�x���`S/��(*�P7���B��Jdڷ�4�����k��r�T�L'g�uK�F�rO+�Ba4d�^X��6��|\�w�w�/�|��&�7N�Bpý�!a �Mb���9��ĂCϭX��lA�l�f�.0%�C�\!�m+�b9����W��X��G;5��2o����I��������ɭF��K/���Έ�d�mB���1�f�:�{������?	�oJ��������_pM�����W˾>Daur�S�x^�{*�JJAwc)�z�np6_G۟���.�4pN��L�Fa��$}e%bwM���6;@�R'�V@)x��޻~�nkz����� �MA�|���{U�ny��X�l<��L�`gۅ2���yE��u���0�g����٪�XY�eX>�A-��,��X��u��~�^���(���5������{Q�S���`4l�����|R��>d��PG�O��VO?����O3W{��`�����X�c˲�~d�7���
s1��ؙڵ��<A�k�t}B�.�UxK�����X#Q� /�� ���Y����3tr�=��;x���3b�%�%6|�S(���Gwu�=Y���qF�y���8��G�%�^B�>o�լnc��&���Ҏ�R��o	�B��B��}C�_Evr��M�J�b`���������� 3Q��8�1!%�(L�2�M��ƺw�cG�rꈻ��F��EѶx���<�@BM݈˟'L�-�U�ۆ���h�糰���/j�'Ȣ> �y�W=���-W��~k����qw�� �x5������3s���e���O��F}��%��J�j_.�Ů�$G�=���v1��oK_/��?�g�"p��x<�q��.Gvm�z��[k�d���14s<}�=����JM}�z�O^|�����g���� R���k������3n3��#q�o�C�)�y���������PΩ�d�p��x�%A���$����z���Z���M��S	�e��p��[��i��L@�OP��ٖ)�&��;��}y������xMcV�+�G�X�aV;���LB�?��$�58�Հ��� ���ۮ�yv��gH��r�6�`�c��/U ����2�}��=[U�}_g,�tto8<����g��l�HO՜�"��F[��E-鰝�xE<�& ,[�v����a%
����ѻ�#O�zT�ƨ�kkA�&%��۪��9�v���_ߖgj�]_��f7��m��0m6�9�
��I�`��D��4��5���z�O��)�D�3{Z;Z��b�1(~��W��G)���|�PG�"��DML6����Uiz�~�i<5�XM����7`�qN���і����V��":�A,��� ���F�Н��C)�q�
Yt5�o�9���M3*z'#�]H��p�r֋9�L�/c$�k��s����H��(n�%T����
ב������1Q8S���䪥 �V��:?���E����|��J�9D�4����4~d���k�9B�K ij�/}A^
3���r}����wg���
����I�^�R����:��}��sLN{��`@#i���=ȷ���-�Т2�]��*�7� ���Y��,�ϟV�e]�Ͼ��������4�VL{´F���QF��֣*�Q~�kqbb���;���m�9@eM�Ǐ��F
1���6�(Ry�|�	�I���s��'�uh����<�p0�*`�̷)c�lP�o�N�*�8^
Z�q�p�I��V#t� Ŭ$ϱJ`K��;_�������^&����˽���"�x���m��[!�c͔$ߔ&��'��J��~�������p�7��l����x����m9�PP"�b�!Z���yz۫ȿCH���-�7K��k&ydwYM:���p�j֛N9��tb���~8-�g���C����6끀�U!��-���`
ﾸ�iХB�_�I��Ly�&3{�c?�]@<7�s�2�n���%p	t�)���`����*��_^Rg�~��}�[��q3���|�Ċz��Emf�[���V�V|�V
��N��/���HY%w � ׂ?o��BV.hݱëyL��5U�h�
�ӈ���+��ޕvD��iؖ���qz�[��~��.�¿��J�*{�y�x�.r��S�w�#���"]�뿗� �<iR<������6h�^��B8c��Y���?0���|��	�!z;8u[xϥ���H?v�>�@q���L ة��b��8|yL>�ו h.�1BQ�W.Z�i�AlÑ���M~�X�3���3���9���T/��/��re�Q*O�jԺ�~�(q����w(<�d����m��`T��%�������p�g�S-^�0�Һj8�}��:�'����v�Y�Wh��{ǿ�f伩�e~����G������j�����R�Jib��+UWK�#?s�+~�Ы�n"��#���'t�#��K�Io�����?��a���r��lm�Ð1#�!���]��
���6�x*����?;2�灥��Hw�i�7������8#:V�;j�8&�oG �G�&�=^�.wo������w��hŀ�!;x�dy���C�� ���G��3�s���0z�]�=
��)'4���V�K���_�O~$�A�8�输?��ɨ�&������f�Lp \�{�ģ4Q��r(��
&�x���hv���[���K��n�J8��}����۔(�������<zc_��i�#�YMOQ���^��LҦ�n���Y�G-����u�5��(�OVг�K�+PC���cM�m�s��6����"� �5ӅHW"@���[���	�Wj�W�ʰ�����E��G�PeL)�%�?x��p9o�[0�<�����o5Kg�9�(IH*
��XԲ�8�j	)A�P@�C��\nJ��z"��D�+���G���4J1f�~�������Ep�d����u�G���T�E(hE1�k�_��ģ%��ɵώ
zfQ`<&z��f࢛w�H�\�`���a�}�qT������Z;ٰj-���H��-%p����}�+%�t�Cd� �O�B{g�vd>=�eՖ]��t޶��ut��]��C�y(�t1^�����{�n�J���T�5��YLK�KmE�֛mʠ�n�6QA?L�C�cJu�?���O3r� �0n��W%���}{~R_���[�V�*�"(�y��z2����Rr��P4�������ym�K+?ϙ��ں�]�bx�G�0�埡�����i�$�Db�f'���8w���߯��8;���`3�F`V��2#��U�N�����lO��ڕ��8�*5P�x�����]R��?o�n'N}*qs�83I��&}���{�ooր�C_�vN�ST��Zߧ6� �S(p�3{gc%�N�bY�P�U��t��OP�r�E}j�a���c��B�^5�^��+�8�x�1A�3�˱
}���xԳcq��Q�f�����5H��_����+�D�)��ik}#ڊJ�B+��
l����OH��d���5o-���lmz!a�Z���� �j*Q�5hl3�6��Ez��f�	[;�4S����fS4�Y�:���k\���v�줭Ni���[��e��{ԃZ5|`݋.D��ӯ�A-DMե���� �R�����㧃.�ǲ���Y?[q`�&�f��P W�{y("�'��Y��O�( �(��dy<��\�#]���]>0�a8��e���w߳�i�/���ҽ_�U�P��B�w���#�D�"�0Z�N$Tx�kw�U��̡�|�U}����Q�L��=n����O����7F�g�M��	ee|�&���j� ���o�*��5w���`��Ã�z!l~�7pas�MI�۵ɭޭ;&�h�C��Q����Ng�yX�ė[B�@i�Ap��J6���3;��{�@�,e��o�PKn&nz7�.ZҴ?��l�_��:K��)f��̴ x$vJ�c����}�X��#�j��">5�����@(Y�ک�t�@��&�@7&>�;.�R/�
d=�Z� k7S'�)3�@ݢh����y�}��d�Ҁ�΢��\ޭQ	�L]�s�Rk��#ڟ��N�r��l���s�3����E��:�������6~����V��:�3_1�J]i������p.��,Ch��)�%�³u�����V������[+�K�?�����Ԫ�������3��ɩ�ۆ��`1������4�"�單˖�Z!h��ѧg)xX]"B%	0�a; �z~q#��J~Q?�<�^���V�yHv�r�^ITU'�4:8�ᢜ޷g�6)���5�W��[�!������������cDj�Ou�/%�� �e=ށHP[w��@�9�O2bd@���ue�h@U�:R��gB��ri�f��A]n��c�2�i]?0Rx��ua$G�P�ѱ�A�� L����Q(�ُ6L�(�l�X�U�Ɩҟ�)����L߿#��W��KǛ��-:�qxռX�R����:~�W�1�P�;�拶Ƨ<RT������!c��~ϊ_��ЦϬ*��Y��~�D�p�)�=���GZ���Н��>�3�Ħ�����\��FƷ�I��m�n��r�ü\��Ɔ�0!}8����X���^��1?3[��k��UA/۬�-��iBhy�h�L��)m�崟��$P���yn��V�3͸s�)�+��3����E�u�,�)4�{�:H�Ȃ��� Ff�LHo��o����m�RQS)|����5k���UF	�,�yh�pL.���j�O�M�g6�|�%���7�Mpja:{&>���|�w�qp�
�1`��!͵d��x����|����'�kU&nF���B����Yx{u����J��Yx̪��o�~���>�X�#��]�ӡ�4,���߃�?,n� �G�29� �$��9�����^��-�],�{z�7��MG���N��0y�.t�S�t��H�=��@��ojx)`%U���+�g'�ڴ,�k��`C�rc���u�Q���<��I��>zwZ�BC��s�њ��ƣj�#����J�Y���wdm4�W�-ʮF��;,�����B?�s_]���
��HN��Y���5�����nh�ψ
�"�,p�(<G���0����0,�@�,;^髐I&G;@x�L�7%<-T����mu���4↦9�8���B�_���W�|;��4·���~� �Yݜ��(������x�}ĺ{j2�i%̾�=�~苳��QB��8k�V�_}�f�B�uU9��͹�V�ห�E�� @��c�S����u	e�"ݪ��+�y��o)E�$�[3Y��I���Q�v+4s��K�qA�!����/�4�n-�_��1s2��a�#L��߆x{ؘ����������1����}R(�%��h���"5�;HH��~8��4c���A��B-�bBA���*��y��Aj�!��[]aF��!�Mr%h~�$�í�z5+a!aT[����B�s{�_T��M������;��"������h������=�٫5�rQ����sN�Į�Ux���*�}��l�{>8ȯ6W�Wg������[�,ͽ-G��JN���WO�<�+�kh�eq���5��B7K�W>��`�̜��2� ���0��3G{�f���No��ς���2�V��q��~`������:��UH �:�ɮՐ��~�D}�V�2D���k��S��s��&S�(�o��� so�����M1�~#�V۩��Y#
�t���l�@;uf����|w���U���xG��Yo��;���r�M�Y���l�����~Ͼ���b�`җ�,�ra��Pâ��į���H,�S��F����O�B"�{�ŉ�3/a���3�b�v&đ����L(���N��-�V��T��#�F��rb:2�F��S/>7X�=�+LsӧMA�Y���f]#��ӯ)�r�k�Ezn+U�نY� �;qv�K�����^�9#b�o�V��cг .�����*����R�
���?W��}�/�x|�̟���J��ǀ��wS�Y�k�z��
<�V���+L�8�-Kn͸�Dy�X��L�}�eۨu�{����O��;0��L�H1�A/E�#F1nQ�j�ľ�O����S���ԅb�ȗ�qX\��T�s�����W��w2�{��0���Qj&C8lz�{����;W��8��	��}�z|]cO�>Qƨ���*ˢ�#������&Ԋǻ>�niq��CD޾W�E��ޝ:���ef���ZH�p�`= �T�?��˭$r.���d����6�-<�6��~ �gzMJ�����m��ן	�F2 s��o���A�wr�͉.�Y\%g�%��?��Ӊ��~�t��/Xx����V���lt]���\���d�0n��57���-�D��
Y���Il�3ZS���"��1{+84mJ�_��&��HG7�n�U���\��h��c2UK��6�H�D��RC'T�����l`�?6��:�LX���[�Zj,�x>o/���v.kTE�Ϭu�{������
��np��jkY�&��[O%��m-,R�� �K(ʭ�j����91����aĭ#�<�QN�K�qOlϐu��l6&�S=8����Ս�t`�S���0�������3�c0{}�R�݌�/�9�Oe��,n~y�1��2鞭�sq��@����
eW���u
[@x�
a«��%�gAEۃ1��	+��Dƪ8�P�B�"d&��f�5%�-�%�	��ϫ������Dp��,�p�Z��I;�/D|8�9��?D,pb�@��èfvI?`/���r��?F��D�*h^o26��54@M' �܏�ɂc�=�ܦ	� �w��O�l-|>��l[�q;��mW�è+�EΫzq�[~�o�ēƚ�4Nj�J!ح�Fj<�S����z�������^ƻ4R:8�R���-�z��Q8t��b������#�o��d�:���hP/>[˼�H� ��|�������]�s���L��Bf ��57�ʓɬ�?���(o�H��.G-���lOXjg��x��yѲ�QԀ�ǣ�ջ��Y���*�Ѫ�\K���^����c�U�p���+IFL8{�_'tȫ��>�Yd�L!K`�C�v!mP���M�W�Ø�a�o-]��ƴ'�u!WRڬDq��N΍��	ryJ��]D?@��߈��k+��[��d$6`K#�D�4�l[�}>X���_����yv>'2em����,�`��g���l�<�k���Ѣ̀?���_#��s;X�yi�zbЇ�:�=e���y\������Q�\,jZ4&ﲛT��V��"k��#�\B?r��E��,�)�C�Hƫ��g^}Q��J�"�����.h����r�oS"u9���S�L䝺�] �)6�iJI�Qk#���>L�eG�N<`�<�����f<�w�ZN@�6��τ����_�C4�}�'���P���b���O��y��n��8C��i+�E?4g�uY0b�0�8�b~K�7��,�P�_���3�]��N��$�4"ں�d6�&jl}��h���8O�����jg�l�� �W+�g��&�l�Ώ��w
޹-D�J�,{^�P-k�(�VwM�!p�'���>��V	!�cI�[w0|��|5cfq0#߯�|w�G�xQ���ry�bTJS�`�d�X�-Uj0QRB��hRh]6�@M����[=���(���K$����!��s���Ak,����aś
���^���ŝ��O��Ru�����VdD�áI��З�h�S���H5Օ7yM����Aڻ?����?���'w[<z}��R��ZqA��tv�`����W�	tP的8~��EP���FA�%_�a�uE�l�?��$!�/Q ��)��ό�a�ᄢ��;$��4��Z���/͜H�cu*�#�X߷��T�?�O�
ӻ�[��w+{ �$�XV�B�ک�z�W)ɓS�Ѯ�S��5E����3�ص�ź�:���I�2:/#�}nb�<�D5=d�̼�=�kd�k�Ł,�,�74���co��w�04��H�]*�g�l*-D9�F��5������(����.�;ņ钑V�B
w�}���율�����J	s�O�qo����O'�鎙 k8!�i�K��#	r��e+�D����f�XW��m�\�L�8ec:V� ��ʮ��G��<���f��\A�~�I{�ʖ!uQH����g�����"V��z�FH��Ϳ�֠&(�?Ɔ�үB��{Q;�/zyW�`��GI���������XUxpR��w����g�����"�� 1�|�#�J��?՘B�:fom=x��NmldتڤUVm�R�=o[� ?���U���=���+ղF3�#bk�G1Y�tAs�>��ne�����vؘe n�[I�e�N����mE�EYn�9��^[�����0�a/C�K�z\����5?	|H� z�8�7të"�]\���!vFk	�c��U�C�Ldリ��H�;����S4M��"�a�\���µ�
�����EAN�ݫE�uߜ�V����.�
"�mH�)d �Ȍ��H���*�t���}_u� ���%��}oy�xL�yu;��U\n���������~=4U/�%��3g���h�n"��0gj��<C}�M�ٴ�X�QӨ �"l~艤<9O?V�_.C�4�n,�R�bn�U�(ź��K�,4{�;��/gQ��8�#6?�6��萒O�W��[��_��j��r�C�\J���tq�QJ(�2�wP�_�f���9��|M6GL�K�f����|ן�KIWD1������Ҝ�V���虬��/3,�~���ffA���ʜmb���
�}� Ѓ��dzzO�E�P�֎�ԓ�w��f5�c	�Й{p�b�3œ@� �Vl!��z�={���*C��ϡ����C����8��D��̉����o=�I�}
��Vt0���#��Dy��K�M��L*E2�����-�7ɘ�i�2Je�:��g�
�S"6���;�O�Z�{�.�p*�k���@qv���gɀS��q$A({�:5�z��昆���Cuk-Y��D%QȾ�p�������ɽȭ����X��k޷iW�0Է"�b������S�`	��X/N6.H�w"HNrI-��fY�:��I[��C��H�ګ�$�U0��8d┿F���4v�L�DC1G��(���U���e�e����W��l�#���� ��Z,��Ƌf���u��=�i�2�Jg+��5'k�dv�k�ad�+,��AK֥�g�w��)�= ,���.���H��X�� �6�>�}ޠɭ� �����Aџ���!���zQ�&=NZe7I]?}(�4�yz\	�����ϬMR���.q?�rrj���%j]���
#<�w�*�: �x?z
�v�"�ĉ��`SH�66��+��7�w�ǫ�ۿE��<��Y9ѧ=������Ye�.���gdm�|�����x�K�P���fi�h�ު����S����Nu>B�D��u���ϯP������Fl���*@I�|�-2��枿<'�8I��Z`�|��Fu�	�x���ib�|XǶ��r�솔�f^�/��#6OZ�]�ku�r�6_�V"�P�?�WmC��K���~�csm�EZ���L7$t^�ϒ$Dt�M�&g��/`�l��/�T��k���f�q��_niV��{I��̑�]9��4ޝЊ��Ȝ�>=�4�e�<����#2��{���@�p�wϳ0�KG�e�w����Wwٝ����R]y�6��P��b#�4x��؞l00u��Xj��UVሮ�c<B�1z�!�U�.~iY�o�q��{�p@a�n9���H��p�W��Κ�,Ř��!�<d�yyHb�|?̨|r�8~;�W�e�a�,���JI�����������Wѽ1�����u���B��������W��c�,F�ol���M��2u��Xr �\����d&�7tG�d���n0��U����q��N�' �*,���`b�p_�ƃK�|j �����Z�����\ !�(6L��@��m��������
��eHI��C(���&"��3�ڸ�s�`�@��Wj����+������(G��(����B�Y�~�E��k��Ã��@(N��`��j�@b>�e��T�Si*��)ê�6������Sr1�G� Oω5R�q[���?�i �	҈����.4/3��]0V亷��a�A��/i���	l�O.���o�K��h�	�c�(���՗�dJ���[��>m�I&
�{��2�!�^�	|�WP��`hj.���c\��Fbt04hJs���iA�{�R�9gWc>vF;P�$3�@�V;�/�R�9�?�e����)�77��R�l��m�e�@:�`q_5}�m� .�;����R̍���p׬J]���X
h�Pbf�G���j�_9�%��>\�:��P��J�~���S�!��,LS ��h|ou��6j^������LQC3w�7=�y./l��ށ8szP��P`�%j�6Ƚ����,��G`��k���BJ��6o��a�g�!!	�1��C�d8.��x^]����9��IX4�QYB��E[/���������f�c�Q���vW�>�XcV�N�6��<>*b-Yw�����E��3(���#��&u��4ZLq�Ӵ\�R5�"2��TR�k�E��$zb��dBQ�Vb��IU�Ҝ����癬.h� ��}))	J/�h����1����_�!�<�q�T���f�����/�w�}��~��� �ji���D��OjuD�;�X��b��)`uV�:m6���mʮ�΢���4�St}�~�j�Z�+�����r�p��6�o2-��?�0`oqc �Z*1+5j?bS4;��r!�wʗ��h��!=�L�iQ,
�?�O�V��u}~B���*җ��zK,jEk��*�e��������-��x{�t�%���ͼ+��%��nzs�5y�R;Vb��d<&V���}?ƿ��֪�WMwֹ�KY\D�h�*�#�Έ�d�6�[��Ωߴ"3��$3�vYܥ��ވ�PХ7��E��OMB�y|<D�#���-a��np(Na�$g"I�B�(I5���u8�E/#�{�� /X��Fq�e;��+��ͫ3??k�l�q�����9���ʄ�o١�[\�X�>� �b�YW�,A�'�$,�
��G^l�z��2.a�����0�Ţ���i�$���tg�b%3�����V�69�����L��^�+dz0=���h��+Aúg��F7[�%/6��L����}	�Z�ڔ=F�qr�6�7����QQ���Q���G
c^v��Q����O҂����>br�e=ho0t��z��B�)'vI�e��||��&�K�c����y����q����+�T D���v��L�I�:i�(����G�N_�۱˴,>� ��`�!3�����՞���dA�l��Y6e�߈џT�8��S���-����Ƭ��f_F���O����oe^<����ݒ�x0�c�wU;�W��nܽ�ʏ}M�>~�*%��C��c��܁�`N3#*x���}!���%���fdXJ���(F
�8q���r��4�y
����aQm{���-��*Z]�	��j����k�cJ� ����[��x^B�17�U��4i�v�@�TD�++^��~�A�d��
C��f��p ��8�6Μ|	��t������_#Eę3�
��	�@⿉dkW�Ѡ��@*J��|��ht��Ǌ�L�{>��0�1&}�"��)�,����������.�2��=���QSԾ�o�� ���GwjJƊ��`���K�3�H�	�����vm�A���0��i	UV��٫��7D݌ި=��V���ӠQS�"ljd�g��$厷�JA���V� <M|m��l7g�C�@U�6%��?1^v����?�	Ƭ�‼82+|D������8��|����Qew�@D��/�p�N�0[j-(m���VGK Bp&��������C�c�s�N�eby�&����Nɘ���ǝ�<�{W�I�.��M����¨�d��4}��B%����J/#,!q�G%�?45�Ny�3���#EVE/��+����B���(/�\?�gA����3�t,�'^�T�&�[a�q��m�����8�0�2�A���"$%7ΧGb��"b�dWe">�{h���ǹO;��c�c��Ё��q]�z�8D�w������հ��H}ex�e�j9�p�1 ����b�yF5u�a�3lټ M�crl[P*P�Y(V�͔�TMF�eS�G����C/�Yř+���R�d�Ӽ�ӏs-�����q��=]ɂm���xU��!׮D�K�0��}�{�[R��Pt����`Gz~S�]5{�&`p%z�+�c3� �{�X�u�{�e��0B�נ��qd��w,�R���+����W&H�S�"�`<3����F ����]�9j��Ħ=�niE�:�%�e�q��w���08���G�^�R$G�`K�N��΃�=$>�0dE�j��|�O�cp.��hH�JԆ��\�Z4n�(t78���1��0_���S�lqa��M��pG:p�ֺ�A��S���Y���b�yhٖ���?!D:�6�&ӢG=�NT�b�QW%,:��l��A�?ޮ��3�&�6���+�!@�Bl0h��Qg�*�����,��p��.I<ۼ����/ѭ�o����[�ކ��yw21g�� ��<��?��(�����Y�!�#�>8���` ���znb<}���_6���{��	���Z�N�y�Zꄺ&�dUЂΫz�VndЭ1��r} ���t��Ԟ��h!d;He �f���>��m�������P�db����ۼ���_�V��M ՝���LX/��&(K��q�Zf��[�96����'��#)bI[4�2�ˡ��)���~yǲȚ�-v��NRe�u��y��.��ٚ�n�Բ�K���Jj#��U�բ��WSN���B:��e����F'9�9��pu���Bw5��\�wf
�orj�k S銆�ѻ�3� �^�6�!�&Cy?I�&ͽ�1���v�]Q��E�'�����U1� �����j7�f�>��W�i�mb!��	E��\���G)N����̨����2gPX4*K1w��2�Līb�¼?̟�i�"AHx6j�L?� FQ��Kł��£o�4,q�*��q0k��ݸk�U�����_���~[v^��Cʰ�.�v�%c�a�z�ף�f�.#�2~�ȝ
&d���+|��kŢj���U��	" �����F�t��l��Il* ��Kܼ7].lE��������9'p����Z�S��Դ�ةf��[<R�@L�\Nb��f�=M�2����i�&hj�]��x�������J��M5��B��7�/�;+S�� _#�:j�V�I�-��v5@�-6�'A/�t�0mx�̰�ƵS�n!I=���z�m�t�Os���e~�+w��?R1j�$#�R�-}�1�4�V�̤R�8=��}�u~��N��T�����2n�kOL!%*��tIn����^o�ݙ>��n���?idM���3���ҧ�L:@�W����DGX�s��qj�l�\�}��1��5��n�H������f\,�M���7j(Vm���vJ=f�؋a�\3�B������ _?Td2�.��Q�LԜ7q�x�TE��~����o]�'�Be=���h�{�b�pCC�8�M� Bb�d*�P���^�W��p�evH�x@>���QWf�D$�:�/�f�U��������.3�C��n���� �]�-� �X>&Hŉ���#uG�yC� ������%���OI���;�gխf�% ]D'�Zl��÷����'�2�'n��G��=WH��#�>��Cw�\xb+J)�\���г�j����*�2�E���A�ee
X��Á_�{�ҟ��w`M�whJ���2+(�LNǻV�&p��ؠ�u���V���5;�����Gx���^+T�vV��>�����1Rg�9w/�	�!��	���2�,���~~s-��`(�h�5�z�'g>/|ȣI2�
K��n� �B!v��a_���Y�%Ph�~Pl�Bք�GTsAC���ٽ�k��"|�EP4㽑h����m��^�B\�f3}pY�����6��M��(����\�{���雯��2Tnr���70쀋�~�U�u��'��`m~쬽�[&���9�Zfu7Jx�W�*p�;�uϘ�~/�q�3�A&�n��Qԡ������?/�L�9o�A�32�YPy�Gu��C��:�p��<�Xy%����+�ǅ����t�$F���d�<��5wT�5Ðy:Q�*��	�B� bK��q����ʞ:��2
���lӈ�f��d|vV��OH�����|�A+M,V��͊M������ر6e~q�i0���K{̀��h�
Y$�D^��$2#����L���h�s�a���q�[		]�M�j����4F�TX�m����D�?����ko�O*�,pb�-����.��DUo��|�Z��8��W(i`:si���ՙ�K8X��� l��y%jb�t�2܏#����<"c2�� Y�T�&.d�f�/fk�^!���j�9���p��2B/?S��	űܖ�i��'�#���X�զ��k,�%��&9ob��w���f�Ul�{�o�D|��k�>���+�T��[yڥ R.��.�����T|�av� Q�*@:a�5�Di�UՒ��{�6d���%��ц\H)�����m�ܑν�]p%v]���R2?M������0̐]�Fl�@������m3�v��ڮ5���u�P-�KE���4 mj��_�f����X�߱�5���[�@E�'���J��0p4H_V��˿�4����<e��|wݒ�R����~Q�G��c�$�gy���G-m���gq��"qQ�u�=��Z�����������i{we�'R�#(]E�������oW�����S�������Y2i���w��I�@T@�3�i�GN������CE_�����Z͓�f����V��M���-����[�L5�k�9U9�\�}�=&S8�s4�/��������4[��-�tΖ��8��O��7c�������v����v�j^�zf��)��(�ms��0"n�NT��S5U)?
�m���74 %�G*Z���0X��q`��L�I3&��0�.����>���b)�����f�T����#�����Ahj�1:Ե`��RR�ˊ"c��m�&�>�xB�oy]U�oix�sr�ёV���@�;���Xͧ�S #E-}J��)~mXoA[�C��Jlw�^����0k%[����מ�%,��&���=�����b�k��z�`�� @,��P��D+��{ Am��V����A,Q=�G�GT��ߦŵA2�K�t�b���z�T��1(:*F�.�Kb���*^v��=��F�X��b���@n��j��v:]�����1b�S�?bU]1����h��b���2���'p�m��|��ո�c��M�)vJ���G�����Z��y򤭑&V
=�~�0\�b)ư��\8�G��S�y��8�XOng�oP�vao���bL�,��)�ͱ�Y�}��*:��`�e�T����+�(Y'�AeӉI*�k�$�|k,�g;�����;��A��U�~:���Mi5�Qۦ���W�J|��&��W��v�A(�(�6�/lG)�f�0���x��@Su�n�dGw�������s	s�~���8z�6��L۶q��*�'��WIm��W9�vװ���I)>��n�f��/i��b����v�p�i|�9�5�Sa��\3Z�S
���'�ed *>^��jFN	O^�T�4��&cBo��>���_��)h )Vуad�m%�����wڑ��*(2� r���>'Xr�v�7��U�Jd���Q���	ogw����y�Ǜ{Z�x�#�t)���{��.%4��WT�n�h��@�I�$�l�z�����*5�_kN9Ծn��{@S�ѥ�rfa�ԜA`�u���J�����hS
�W	z�~�U����㌰��`�PE�֯%=���`ލ��|��i�=���K���TkG��W;��&�Iu|m����޼@��.�ބP�>S�����Vŵឭ���-3L"�:y�s�m��گ�%%S7��`�T���et�bƀ%g�~�X'��	Ɯ0�W1�g�%�#puI�m5'#|}/6�~Ԕν�5��m�BIY,ֹ��&R�V�2����Y��|�Kҕ(v��\e�����$�-R|��P��.k��}�@�Z���2و��(G�	NwM�jr��f��mu����V.��0�һ��X��"�5䵭�i���@͗�-%�ħ�'�/?L��C;�x�{�%n�����Õ7R���H��Rv�\�A �%�z�:�\����Y������E�����z����;�^ZU#q@N�����r{QL��� �%3�V+=�u�E�z�`_Nt1_��Y����Q�M	.䊺Ϋ�F�,9��W3�:帒t�a�'8;�T��4�(����MK���g��{��$Sƀ vk݂�+>���̎��+=�^��/��X�U�)�{��1���游l��N�ǏI%ٽV����f��'w�Y��h�8q�h�	�����
F�iv߱�
�In�`I°��X��B��GG]�lDY�	�xnL���K1��sQ�ǨZ*�*i��0�Q�؝<V�H6w���.x�T��^��CR�A�E��K?�f(�}'Ι4
��9�6��3���2��m���d����m��=���U�u���D��ҡ�)��B A��g�m��8��l�5��W��T�\|Ik(9�!���r=�vjW���'E9Д�V�hh�ǫ����G��+�<}����R7���_�&ngOg��ܙ�yW�G�Cf�"�oif^���X>�W���tӰ%�S�X��Ц���g�L�G���1uz�\XY��� gr�m8P���Ͼ��D~l�]�q�����vw����yC�oA��"�Rį�?��+#b�H��2�WZ�zH���h�v$���������;3KK�GY�,���t��0 ��n�H�U����T�N��4,n0c�+�;���ӐNq��Ԩ�N���y�v~E���r����p�_%��qcl$�����}����`�M�IIi�;�M��t��o��\�:f��&g-)x>��=^S+u��D py~�j�[��9M�ٵ0g�Q�B��[i������XvX��)������˔���f�E������p��z9�SЪȫ	y@�	��w��!T8z\H��)�G��� ��J��X7�aX~�l��hSRF�K�����n���G��]�V*��Z�_n��5z	�jj࢈��w��c_�{mRl<�;T�@�2���;짓�V�ֳ��R<��Af�NL^�f��	��)y��ϰ�Tc(	�B��2�3��"���(_c�S�x�mw�n�g��,�J�5��u���~�)Cɰ�;��b�⇒`fQ3tm0)~y1�`[=�`��/��'pݵ�A�J�#D&pa�~g #?���Orhʭ�}2��:�9yv~>�D/�w��Z�2~ʰT��Ks����7�����DP��u}IK��L]���q0M��D�QZ������9�ݨ �Ft��f.Y�S��>�c4Bl���Y�3�#�X��{\�Ojs�1�P���d؟�Z��7�ϑC�.!e��w��2F��������&js8�9�%+�B\\q����j��˛����5�0�;��D��h�5��$O>^\x�~�4�v��瀦����,^��Tu�u��0c`�A��C�cH"�g���X]�_��*W�m����Ͼ
b�{yC]��5���镰�Ԓu�c^��1_��!؉K��-(�)��U����������.x�y)o)�0������kHf~u;k*�ңI5�9M�I`ܰ9>v�
=����$̩J�m6N|8���e�j���A���K�vv؞�QX�S����u��Z�~�X���r
z�ie���A�#B�>�9��;߻���R�2���+[���.%�o�Z9
@��K����Z4\�i`)��v)Z�95I����<T"fE� X�����ΖRúH���f�KW�D�u;��>,x�'E�[�������C;�#{�.��@YD�=�9F������wʰ�Ue�z���5u>����?����L!Z��vb��i�G��H�)���a�!�*���h4�����M������*p������e'�;�O7k;�aT�����ϰg'�c)T6�%O���J Er�X�{X�6j(�O*��e�͉�¤1�����ٮ;�3vbd�����x)V��p5/�	DUaR�f�XW���j�fg��!���G*��
������^|Kl:.�w����@a�F5p�{��9�!
˩��~ᄣұ���i��}�4J�+n<�G��_�W<��F�^��9�:l>V0�C���+��łz	��U�V���P�~���6*p�a������Ő�>y�è�rɴ;}�wp�����D8��I�	JF!�j�V�0'r"��ދyT���QVv�v�ڽ4C���/O��[0#�X��mpy"�#���~9?i5�X�_��o���ėK�H�����z������t�E�1�;��<�"&e�(�Z��>�CM/��b7�����/��yZ���'�w�� �^(-T�����݋mc�|P�*��Z?�m�[R�9ďꊔ��M��G[]��&z��9o{���_�Q��q������8Itø�fÞ�(�M6�:�/q����ν��K$��t���,<KRw�XxeJ	���SE����=@�oad��\�����]t�������K4��"����ħVМ�b�z�Pe<�A=�_/��`�� �d��@�E��j�p���	��^<���L��a�98��Ih�G��(n�6����z��&)��n�[xP��_����,�G�l��#�D2�-�����W�7������%�6ߊKag;���նFhz�O>ʪ�}P��n9;u�eF'���Y̫wr��Vf��;�_�a��]�`�ڍ���в�'ᆕ���UG��񓗏)�H���21����w#����o�AOg2��R���Ks�;��� ب�4M�6	+.�u�'��gd�˯��#[���Vo��mEuy=MTa���Ą�wa�Z2��ޞ���o��P.���#<bs��B�4�h3mJ[�t�a���5E�c!ҫϞ�Ĳ�7o�>!о�zᡪ�IT������T�/ �J���l�3_�Wѱ�"�y�x�	M":4AJ� �+�ʧ��2��֫nY�K4�t ����@M?!��F��0��5�)��g�V'��0R%��\5aJ+-�I������2&~����C�����F(�pi6ǵG���-n���UHZ�g�Ǿ�TunrWS��FVX�b1���]�U���;�l>�c��|�^��Y�?s�-�\h&M��������p��6ӯ,	lp{$�Y_��lϭ�����'��%�BڣKif@R':N����OJ#P�b�0f��%����g�(�����J���!H�붒|���9?b���=����`oC��� �ٽ�j��R�fop�z�+�O1}煗�C���/�r ��o] S�z�:ڨi5�L�/	NP�lQi`�r�w�ڒ�'4w��Y��;�V9:� ��\W��|��%*Ψ�~Z�~>'y��9܅ʚ\���ʉd�Q��)w���8f-)�7P0�o� "��OC]0f���6(��!ۉ��{�2�A������ڥ�,,WF��@��|��;�碕��g�v�X��y��Z����<C[H�H%�,���o�*FJtz�q#��d�P��k(N�6"V�^���e�F{���O�a%.����Q%�*T�񥥲XIS�&jG���	qT�&��]>���F��*,$�a�oA�^3�����I����$��}��C�M��9�8�A�(=������CP����׉��_�/�	��F��u��$�&I.�G�D�q-2�'!�!�{��z*/�2ϰw�K�I0�3 �����/��A����2���eX�/l��5������G}��{�_s^�����-mNF� &Xh�sCQ;��?s�u�gmV͏9�P�
�]����֙F�K�@���W2Nhcm��Tz��ڨ�I�,�?���<�����N�XIG�U���k����l�օˤ�Z�_����)�y �&��̬�)����B���:@�DA��N���R�țD�ӰH3�u�T���fw����EW��)���m��6��|1��~�B����Y�-|�SW)!�B�����IALk~�����u�e�O³01s^!~	AN"�$����&^��7��A-�:��{�
]��n���!�����I��� >[%G|��"RV"��+|s'ۼ!�k	�IĦ�P��yU�9T��o>��8<�!����zP����o«���eX`jG�<��I����+AF[�l�o����_����s3�y�3\�~J=�oO�?���� �F�*�~���j��d��E�����i���S)b7X��gѸ���ɥA�i��"P~�8UiZ�!y5~z����N��t���_�� =���&L��edl+�VP����w`&������- "�K��D�wA�V�̦�lw�6j�#5Ǖ!��}�\HQ\m)�ֱ��U�
+�L�-ru�fr� x��T���n�x�,�4J�8FxO�R����,���:��7J��TK;�/�%Z3�fI�ڱ�	�9���v[k)�b&"��T�U ���p��>���3N	8�Ӳ����|aȹ��v�S�԰T`�j��L=�1 �8�{W���w��#�ߋ_����R�N�����HOу7/�}������YQ��~ݯ=FG����U�撿6j��7`z���+zU��1��L-+�b�iƽqȓ��/�%,ڗSw���0�cY�>��D�Ж�į�г���뮢���h<�36��Ğ0��:�Q�஝�elX%[��Vt�Np�:N7\�Ҩn��[`FJ@���E�Jmp:V�T<��(�v�_F.�dzg��c�L�b�sm~���gB�4����'C鯇��򍥄'T\��9(c�p�IwOOM6n���!�^G>n�8T�F���%�GɎ���a�}^XS -�0K��\i���}-�E�֐/�L��-�)�I��<'��4�<Ê�L��dq��bY��<�P��� �d������������$_�❼�_���D�����s�V2��60Ԏ'+0��u�3�UU⃫z�����)��8!�l���	��1�X�x����Ij�_5M�M$��#��8�_�ʰ5Iـ�[:�:�pO!ZPظ����t����H����p�y�D�co�c[ ��ζ0���c:�ڳ�F���Z��^���TX�ѯ�ďL�"�۠\�O��p_��>h�J�)�D?�2.���� YG/캃5�U�)O@%�c:�ڊ�� ,�����z�