��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ��<��T�@d�Gu�!�h�����j~���C��P�Rc���FfxXs�� PC��԰�O����p32iXA�t�"�Q��&?,P#̓�*eA�9T�x��0�8nVHAG8A��J	��c���G܂y��S7AC����&� �?�,�	�B�Ũ��aU�P�̧Θ꾸^�����\�(+��F�I�j�z	�Ϩ��y�g�8!�2���%Q���_�m�$�x���b3,B�6����9�@fZ{�G?֔H���R ���o�;��Hd�����������O��3�m.��]k<�B��I_"Z�L2��:*p:߶����aȈuJ�L�_&�݋�w�����j3�����:6���Ɋ=�����e������0|)
m�N�|[d�)��H���ڵE��Jq�)Tꗓ&�^`kC��O bC������h�j<��+�E�v�)��G�i�SN�p��x��Ǔ,�z1��@��t�ܕ돹S��Iເ��8�^x�)�=��V�fE�s��a�3c�e �ɢ5xE�'�fr&��W`��r�E�m�_R�W�(�|1��hR�%�O��p�ʼvkn��I���T;6�<���d�Gt����d��qkcR��H�5=�E�zD�YX�k���B��&+8�w�}��3V��Cbk�9G��3�����h���7�#���J���j���d�]�O�x�kk�J�1�A_��,�&�:�C����+S+�p�R�^4fN���U81�{^��_!�R�q�Da\��p��{��Ox�o��,ȕ����
J��wܡ�V �p~�P�l�}8���KP��שX���B֬ȼ���_�R_�?Pٷ�x��4TZU
�4E[vS���J(R�v��3��C
�U5џ�����!�tQ��"�Ktf�ʜ���Y�O�����S�ѡf#�;�b���=Wb���� ,�gsZ[�����;`�����&��̾gU��٨P+�4�:���>Շ��)e��Κi�l���]pT�r�E &��v�{�L��ۛ��3M����e�E�g�
1g���}�=�Q��j!s��+��ɗj�%�)����	ӕ�
�qIq�bZ����לb3�+;��A��q���p\�߽���]��<�z>���Iso�Ϙƺ���>��C�Ȫ��\+��hS���v��`2�_�:�96@}jO���2y���\uD�J���h}�bF��f3�?JL򿐭k����k�V ۮɸ�\G����Z5Mۏ�w$C�΄�w�@d�����%h���}��i��K�Q���d���IO� (P)��0(L�� ��Y�>g�oZ�n��6�I��Sv�{?�a������"�' ޜ`��i���&��vEr*�+��樨pĔ��U�x0����~��G��� ]��0V�"��u���OR�8dC���J�(#�v�S�Ci��`��<���!���J7�������>R5�GOAe��)RiU���5�(9	Ϸ\��v���i=�����F���{f�fpX�7״՟{���'���[�+} �×?�kݹ��y���Z�4��&%�E�����]?���ZQ�"�d���b^���
���	����ff��גּ�����V�*`��[�l��z�K8�5l�ʴa<d!T�
"-52�fGL��`n���u�o<A����V&(#��؀���܃z(�M�C�d+Y�[Z���ca���CY@�u�������7�X�`���[#ÖӪ!n|@ ���~�z��Y����<�H�_�Vu ̼���j 7��8�ָ���ܨ'�鄤Z�2eUf0\~"������U��E�TӖcS�U����8��I�:�W�[*�]�	�-p����JMr�����45b�l��
���z�K�t(·���{�e{���CBP�0�Q�ŏ���e�	��h�z������]�o���C�Ȟ[�"m���A5s�`Z8���Xx����E���o�
�<ۂ��}q~���|�~�x�,�da���/�����.x�0`�7��|2/��r�"c�[��&�0�(C�����mv��-d�+��v/��5���`�����M��
�{��O�x�4B�f�i\1 �cW�"^����[����e� !�Ԫ�-G�!�3�ۤs���x�L[���/�c?��Iw��Ҕ��׎vI:�^$]�)��CQ�J�Z\nҞ��� q@E|rQ�{�UH5H�@�D�����r���%E��~�cE@�U�wT����C$�L���[C$.�����;�	p��)1i�ߊ��J�!���:�~� `ozF&��1c��Ҫ�T��	A|i��ډ`_z��&4K�R�{��5.2�5���qWL�����E��C밯"��"��6��.����\�٤1&��v��o@�Qʜ�)����a?��~���9�����W�K�c;�f��qKʛ�������'[�A(Z5�,k�
J�� ������{���]��'g�����Lp��|f�T�w�w��]L6�Hg=��C&WDۢ�M]D�~jY������0�h�N������^�M�D��4�:p��`�d1�5�-]�Xe�¹}�jh�[ݲ�UfcS�Ԋ!�!���ب�X�Q[
�r���QhG���jkH`b69\�w/ X���>��jw��pfSw�"���@�h8��?��ι~�V)y���m٠�H}ԃe���j*�J^sI-�Bf6&g*�jA����,"��&�t@�_�%�_7BC�0,%��0���;W�WǐW`��֭�δZ
�Lӽ��^THtUO�2/V����CX"���� u���H�ZE+�}D:�P�J��q�M���?l���*u��<���z��=���h7r ���K��b�|���_O��b�3_� ó.T�֜js�jx��볰eЪO1�?!�ڥ]&�;�b�Z��Q�C:dW��U�8�|�!%		�q���	^G�x�.����t�u�U�S�0\*�gC����|�/�,'�U2��.m	&�xZ��a�B���������3��(�lm�0�;���F����LL뱑�1n����X'|*�A�����"1@�;S�Y��FP�E������9������.e%1���IRMb���	��)�Oa��O���(Nf%��=.�wɥYv�$��o7*j~M����N�A`�����[��<G�Hռ�pm,?�/��M#�K��;�QH�c�F$�Lz'�)�ˆ_�*�@����ZEO�c���_8�!�6�(|:���A�w�rܞnw�1�P�nE.{�HD�Rq���1�I�9[,��F�oX\�UBi2�W��:�%��=�����2
��U��������i n�Nn��TD�'��9�/��sg�5)��6QcU���Ds��}v�.��[_�\۬]�x�\RVʡ�is���N�gx����U�Ί��\��d���d�_B�02���ABI�~�/�����d�+�%ƃ���!�f��|�8��{���,3�2�'�ߠeS����u&����Uք����L	�,J�ۊ�t���;#���tc������pm���J2�j-S�鶫��dI뼹Еa��7sc<�D�7�Y�~�Z�oɶ"�#��R����6[�3�����:�١L+��8r�e/�P�1)�pVm���[Ѹ��o;d��ؗ�*�DD
�E�z��֩k���x�QH�Bzu�D�Aow�ף��L���8a�iF�aQ����j6���I������Q��Ԍ��n&��f �ҝ�33�A&̎�2%�#��.�Sg�̂a]�N�xn U��G��M؏�s�"�S~琮ô�K0ɹ0���b�A��� ��v\��b6�z`+N�N�R�)�
�ao���B��k��dI!��n2n4�H�T+�r�ZV�ī b�u|�����Bb�|����G����Cc���,E��?Jg�jś�~��[#��,7>�MPN/�̜��U챗0�݉9?�4"ٞf� wd+�����^v��KYF�]k��aǌg��I>�����r�RǪ�ȑz*2��$���<��	���!2��A�w�Ш���L
e�IfV���I����CZ�|N���iݮ�P�<>��lb�Ќ�p���s~�g��a]<j0��i! a��V�8gK����6w��Q����4G}�ի�h�Ë�CT����O��'d�"�ѭ�}�xLv�����eM��1q}lYgn.���F�}��n�^0�]w���zu�4�=U�ι<K�E������`�1�j��"V�۾�u��D_Tj���:�p��3��s(�,f��c���r�JUF?�Gi����Q�d�R�4�ׁL�-1aH�������-x�m1l�^�րq<�׾��+,=��4��g-C���9+~�z�^{�~?^�f����1�a?���:W}��dy#掚���}�:v��U8�q뗬��8�5|�[�.P-Z웞�A45{Y��܊?O}o�b9���Dq*��3�E
wb�Yi�w��M�k'>��~�c�;��/�n�Gùg*�3�I� �y�S_
��|�?Cb!�	z$�\h�C��Zx\9w��/F�xpآ_'kGa���`iK]�F��R[�����IX�kzѪp��eÒ������6 Y�^%
��-҃F�_�A$?tA��:��7�)�rF0ļ5x{���߰�q셆g9-q�lQ�e�Rs���'�/�3�m��wč�Uў���+�]`q�9������v�M��fv�$ r��e�3�� "��U���}�5�r�7����H��mJ��	��o���Pr�0�]Ĩ�Vm(@< �o�]7�p���l7�R������:k͟���,S�-{��	��<D8o[Rc�p����9��P�+�L^����ڴ�z#���utg����T��tx�����bf��iS@E�L��wHV��J�>g#
\\�}�9�m��G���c�]��'g^@[��A�ٜ�T����G�m�q2o�ՉB��ܵ5e�e-�oI���ai�;p��j����֤8�zh[���K־�ݦ���J@_�v�Ծx���Rt.K���s��H� �����#'�=�_�)��������ƺZ�?�cW@��N���<���I���ZD�n�9SB6��;���#�9FI���Ĝ5�6R�H 3�<G״�F��ɩ�6ި�W�t37��� \1hxiꛛ��^�;u��qr�r�e)��|Hwk�v�4�TO����h��5��SY ��
���_�G�X��f�ecV���{�s��]S�|o�$�+	N@�#��k�?���kbm�����+n#b �������T'_O�G.3:zOb���F
̆<&�-���~�	t�8���=�ԈR��������J����P�	�"�\����n�}8���P�E��z\UQ��Q7�&=�'��Z��mr�qFE����.�f�h�Ӄ�ɘ�"�E��B�!�Eă��\���ôDj�����o����U�hf�y����w8���D�s��`�싄ⳉ՟I���Y�;�H�l����Wb2�1Q�7���q��/pD�j`]r�C=����3w��`RD�h0������a��<Ko��WF�<v�8ȑ+�tA?� �9t�7J�s�
�V�v�t��3�ʷb�T�A��V�D	�#�N�ٿ�jJ�(ċ��.WJ���P�!�E wCJ/�,*R}�Z�y�}o=j��
��ޤ�	a)e6�Sbc�;�Wӟ�Y��5T׬�En(Y#|�ȩ,,l��3W厵�!�+��щ��3.�c���2�gD��)�G�[��uk�ӹ��'F���&���ڕ#��d�phm�nEM�_2�p��$���N{�<�G�c����p�"�ţ+HB9�T=Fe��D�W>��Q�(�ub8&\�eō�L��>��e&���f�G2��X����S��,{���o�x���B���Iˋ߶��\�-�LnZ>15�ϋR���9ͧ��*.� .�	��(}Է\����嬲N�����v2cξ��ɻ=���7�X��B0��`���`�� �|*����y��2�-J=�I!���J?� �o胇}�w��4Ƙ4�[t�v�+`R;FlA��W/�{2�E���nE �*�� �P���͎�N��;[���+������JcLp�3�(�f#q/d��mM����u���p���
	��O?[K��t?�mն7
JᏟm��K��Y�C19L��uDM��꯸�LnXuli#���r����s{�X2���D_SPT"z ���5>_��V�n��{g�/�MdY^��jxE��^˧���LC(ǹګ��p)*��<��i2OH�4Y�e��xT��+�X!ݖ��kө6;F��Mt}n*`sT~:����ɔ���Sko��Ϻ$�LPü��@�r���D�Xgk������9CXB�(w�X��m�o"�
='�ϴh�JLg�6��LQّ$g
�EgdJ���&��������yv|mjÙoT�?��x6m3!T�/�]��	��.�7�e
ةS#��D��g�l*��]fhӎb�[��V�`��7�M'��Vn"���mK�L��/=�q{�dP�ui�R��Y�unf�7��J,�E����oy�ɶ�r��b3���^ebһ�R���;l�2}���ض��~�Z� CDں���ԝ��J�&Q.A5�P��0b�w{�Wh����$5�O_2�[��t�>�V-�� ѽ�p'u86�,c_�G��1fU�<yК*�}^���{�P��f�w�E{Av�EM�/������8
l#����9zb��UjI��ep�gp�}9ƭF���-����c[�C�E�J2mD�l>Cی�Cm�q��f-tNWF�?����)_Q��>��_��d���] �?��ݬ�躛���Tbl�h���M��шW|_��OI�9=clܒ�,�-:ǒzev�Oa�g<�q�1�"��;AC���O[�ed�/\� �w��Wu�\�c���+�3�!\��ޫ�c���$����j�ׯw���{���f�h��mg]3�0?��r�ܦ��h^ʄz'�*qxj������>~���:�f�-m[�&���
�j������gR])"	!�ɬ!f?�Kƒ���"�Cmt�̹�c�͏�Yh��w�6~h�9q� YF ����D�8�Cc�e�@���r���|
���Y+�Pqȗ���<��h���1ױ5-�t�)?�;Tʈ�f�j�Ŗ�`G�K]^�IۖQ���~�趼_��g'��f�P�4��k�뙮<� �OVD�b��"e��(o=��a�G��W
(H����X�<�q:�+�a��0O}�p�h-,�r�pF�E?q4�˅;�v�`�I�zZC`W���%�YA�� �҇{���뛅�Ճ��nޑ�9���6ֹnԾa�9ubJ4�ӥ@g�Gc-��=j&G�J`x����D�9�BX�}蛃�������`ܣ��z�Ѡ?o�kE-��n�Z\B�z���W �BL��?x�D��㱋������+���.t�Sn�ĭ,�O�~��d9m��\�a�}�'���e�!�Y��
n�C���)bl���N��"�t��l�1�H��c�nP[�֬���w�hg:i�Dx��������4��)&�f�4�O!�9_��8���7J:��nE�l}�W���?���3�w��S#�ٵž�w�ӿ\���0��[��T(XZ�W1�6d�('��^��CG)�L���@�K��ߵ�A5��xai
�ƿ�:	m��q��H�5�Q���
�wWa��K5O���C*+��uK�$�@�������ª�<�2cr��4b�f�%�Q�G�BJz��<D,���[�j�"��o�W}��;v��Ʀjh��0�L�ZR%�`I`�YR-4i����@'j��9/C:����4�e�}7�Vꐸ[��?�����I�{=h��x�8���}A\�C߷!���b؇��=���Xc%�C�+&�{%eq�Jhv��YP'0�g�pi�?a�n��AI>�?�(���w��;f�C�<�7�u�*�>�<��7k��s�b�]�R\���NF���0�QP��prD�3x�]�c�`���OXE�,{����耘��k`���8tA�B}�I�_��¦�\x���Z�M}=X��C)i>�'
�'����X�\7�؋�͒*#�/hS�y����Kԑaa�d���h|̲?s�.�[��ev�����D�8�[�{:���4\W#���P{US08���TyՐ���
<����a���/�鹌72�Ec)c�$p<�
 ��ě�Ӓ^�E8ϔ3�eY��wC�o\fp�В�NTB5�]I-�$�;�i�5q�U����y��N?b?��!�JRl�Z`��C �r�h����gl��էU�,p�?<��:�c�݁te:�5�(Ƌ&%٩���k�>c"����΢��������?�T��Z�B~9���o ��|cz+�D#��YJ1_�?<fV
-n~8�Ww�Y�5��c�z�����\�f;Hv�2?�l.�؍f��`��b���6�)�!&b�� ��b�`���?�.,�� ��~ū<��6ޑ��#Q�4$-�{��n��e��}�ZN5����l�!���Un�T�5�U���
�f�g�D��J>���vO�y��5�.^�ItM?�:�6ɄmӌY�4s���uw�!Q_`��ӹ�ʛ�\�׹=��R�r�?���@c��nG[��Zs[cＡ���H�c$I�M^�+8T�H94����M*kZ���� ��W��������3�Sɛ�X�����:E!�_t��֜�/����a�����
č3\A�b)� �����n�vRZ�Aq]�|�@C�P�����O-��ٙ˛h��0��F"z�y�P��6J(���r?���IN3V)I]���K?W��oW�F;fU���.����� �6�_Ue�����	��{ȢBk�u�@3���t�|��W���Ix�
�PY���H�@��tO9�E� V ?���ҋ�?699��Fc�6�z�+�h��U��4cbJv/���N�}�M֫d	h6]�O4j�Q����|61_��a�T*�th����%�.skM���b�w�*�@�v���i���M�YR"���*������$pl8%�\ў/`��2p��#�HNVj�Ä�ކk|b�.)�W������b�M�Є���`��f�.�?�jۺ)��!'Vu�׺����طuR�ޙgc�f�!ٍ�F��0ʋ���x�Q6�|:.r�"_�hZ|�Q?!��ϕ�>Ek���wqK@7�N�榟�e�m!Ա���Ap��_a���Z$�-���8��Q���Rf�	�n��^�Ӂ�`��x�#�l~���]B �& |�Y���U��D�7J�����a��,�[-��jf�ٜ�޷�����!Z�M��M��`���ʫ\�_�!�P{|(�1�ωs��r�F��'��?�C�d��s��%�M	�#��v������o�f߲�����3��\�MR� �y��.0�ɸ+�`�O�NTq�c�w�N�O�v_a����#Ȉ��"�}��i��E��	8L��
�A��Q]+�}�`?=g�te ��s�ٖ*%�,���vmür��/����{���4�$,�,;��smZ:KQ]�0  �ْ��G�}�'h:6���)5k���(��~#�T`,��Ba�@~�dX�����ϖ>�I7�k�{����X�l���q̸^��pM��N��&�cP%����x��)nE`f����� ���,�E,�s�cl�ފxH7���Ġ=�������0���ȱ�2�ĄO:��v)�=F�I�>i���;���a��ڔ@��.�} �*���;��>�[�|W���S�p��nD�������q��t|G�+���HƘ/Q۳�m���p���3���B|ѿ�,��Y� }6}D����iQ�~lB��O��e�P���z)a��ݢ�����l�z~s���/�܈�TT<��	��i3�f�/^�3��"6GUR'�0(�c2)�0@��@����O��z���7#��S���;�H����;TX�ֻ�⸶�� M�++k�K��vOeZXYTW5��#L��h�X �=�m:���M�V8J��w��|�H�~񀲓y���~�m|*�R�1@�q��5n���-�ђk��#����r�o-� ��:��(b���uh�H�ْ��$��v���B�S��w�e�
~�2E�3N/MX�a�2�Nlt�\�z�_���;U	�{�$W�OZ(�|d����(�W�zS�ag�(0$��-w8�v�+���H/��XǕ�\T�J���B�����#h�<��G�Q�U���~,
�STM9�lz�MA�I��@~>biǮV����"m����]TɆ��%�Y
��N��{��7�QG���6�9@vI�_��?�~l�\vc<\/"M/5��W_��b!Y*}��g:عJ^:kWԈ��N��v-�$�a�Ɯ������s�D_=P}ݷ'_�Q@�k�r��]����:����iJ���O�Xj�8*�1(�X���w�h�h�J�Q7�����5�4ɈP����<�s �~4Jc$`���h���B�ˑ��'�vT�Zt�cV�d�!s�j'��r�V���yU���rc�<���cQ���`�^����^e:����Wش����m����j�8�x��#���q��k"H5�:H��l�q���uu&M֙�of%�w���t9��j�tĴ��:�((,i�+,Lqޕ>�Y���j~ho?��l9���^��AX֗��� �_��Zx�%
�w�YY]���1�"l}B�9�	����0�{�����⁶���H��4��hG�ͨ�pa�0���ezA&�E�����գ��T]�7V�Pa�:�s�V:u�2� aB�/4�����#�qkWي���2���nZ2d�ޱ�RDW���\���!�C~d��%��[�}ɩv��b0�kp���t8�(+;�(}j���d���q�ۅp;	����o9�'K�q��(-�����Q���b�1���,�v�kN3'+@�OD�6m��|�~�n��
5�Z��7�x]9��@La`P��#:-CNi�N���'���Yy�V�t����{~=ŀ�"s}Q��*��8$q�vV�~��n�&�s;(*���`D�H�敫;��c$*��d���+�uF9������d*�F	����Y��	h����Y�68��<�y��c��s�t�Rq����a�!��X,f�ur�IP�龅?ק���̬�S�M/7wS�k�yD�8�6�_��T�� �G���R�NѼ<�rb�3	�%_�5PC#��8����{�|Nl�l�M��H��[ܴ�%Q(_�ԨV#��2.2*s�k��ಹ�b���QDOտ>Z��������N�t����N`p�ڑ�\�57J?]G���<\��bZf_�^����t�^�i޽i�6��@��ijd����.�Ͼ��*-�1�{�0Vg�Fd�+R���6��$ �/��E8���5�H5`
���� ���D�Y[P	z��U9A�
��+�G�¡��Rȵ*�hZ=�����v�S1�U��I�1��h��p������'q>>萷��N��y�\�@h3x,��D�q6i�{��6ғ���x����"��/ޝ�y(+��bI^��="|��������T�fw���>��1�� wW�ks��Y�$�>1���&��=mΊGU������-�$�,��*��J�s�H'���=⤔I���%G���U��a;@ϨJ=a���,����{̤O��a僱���X@�W�&��Y���ӗ��=NTj
U��^q]�J[�T�X$_�P���E~gδ�
{�����g)u�m:"��.7!n�)�y����y�B�\�5�X������S'^���Բ��<h��hds$��m��7E�g_\�T!h�1�]I����e���,�<�����!��S���s���c��R�؞*5�x���Y���Z�i[b�Oq���`*L��B<���<<l��6�*���H
�8���{z6�)��)�Q�s�6�"A�"�3�<N�	u^���cX)+.��v�^��}h���<�����!�\���lk����X�$��>9���/r��<f��꟦HUȖt�z���۳��ʓ�-�6$j���x��� U�Q�BX���]��}x=D�@��V\��6�!�bq�V������=�2��f��C�9�2�(>]A� B���Jm�-���P�ٯxƾ|@�Z�����2�w��{�5E-�D'��Q�6t�
)��qC��Z��h�p�Aʕ�w���\�A�rңD�[���7\�J��@^d��tŮ�As�R���Aۂ�&�+�T� �%,E6�7Tq�xEs	�������O�4���/o�Ǽy�Q����y�R��J���:��.|�:�Ā������ӫ�tG#+"b\��i�Df�ig���{�D��هH���w�Md��� �%`\�ߟ��^��~[�͂��3Z��R���#�d��s���&����'T�d�؆��y��4^��jʙ&���q��զ����1��� P�9����")>'��V`�C� J��x}R%�k*�>��K����H%�uޫ��[kR<���UhtS���п =�f@�o���*���ɴ�ܕX e!��qՕ�	0)S.�Lz,�Ž?�]W)2Ed
��
����x*�"	<�/L��Ӳ�H!z/<�"�J��/_�lHw]Ħ���f��!�*	�̾���+k4 l�@�`���9� [s5ES�~��jf��n�z��8ʑM��J�ZT}���c'��ťt0�GQY�b���+&Bs1'�B!{&w��֥��������Kf��6k�'J3��3��'S���Ռ��J~|�;���%�t她J��T���x�	W����%h�ǵ#�@�8� 	�H � C�?)M�`�	�^PO��M�sKs���;wM�"9�O�i��0j��,�t�iu�$�����Sc�Ԅ{�9������S��!�#ʅ ��5��ЄCkUۨO&/l8� � OI9�1��j�:���I6Q��,���,@B%#�����CBʦ�,��V-��~��� ���>Q�QɁq�qq@r:y��ܧ�i}s�8��/�{O���W�k1�A9@/�]���2]��;�[��$���^�:9!_!�$�&�'�e�\��R�f�'i�66a�ĭ��}�[���,�j<T�C���
q�(
�O9R��fz��8�*��R'5$2�:۫yC=��;3�}�7�Yj�Y�Bo[��~���]�^��*F�����|hws�oW��8�53��?�����S�ew�T{�b���#lt���	<\������R
���sPa�'�D��=�M.WA��Gq(v.!�+]b��GOU�}bI�3����)���S��I>�K.��Q<�Y�'��w���g�b�u�r�f��V�'��CM���9ѿ�%Q�X�[�	g������t�/�G��^�}��AD^i����T�ࣲ%��������5�	z�
��K�aD�
M�>�yQ'I�QJ�EH/��@@0Ce|20�r�@s��+>�X@��4'�C����	��!$7+-�Ne/���JL����@2[A����e���m@���o�g�D2���f�の�K<`R�v�:��#z6����V���k��������{�z�$��O`�����!�Z�X2p���)�s���M�[�c�f�b q��x�b��95
�3�!%j~��dF���G�rN�{�T����,��J�[H:Fz ���1���lِ=���	P��(��9��N}�޵D؂���wO�#��60���.��X����bq�b��-8�iv����v�/<�f��
�RcB#�jJ^P���xTL|x���e|H�mҌ�9�J������Q�٭z�Ҷ���ZW^��ƲA,��.���p{������g�87r/�wrQ�DxV�����GiB�g]��?r
�Iø�S+�]d;G��W��VK� d��s�)u��c9���
?��O0���x��cf�t�XqV��jj�@<�ĝ05���Tyq;�������f[��^�j��.-i�?����p��r����R k�F ��pˑ�S�w�Ԏ��F��׾05U�|���uEC�O�9z?I�	�-�R+.�Z�m��j���;����Tp5��1B=�}f��G4�;��BW���Jn9s�"��a���7.sR�m*D�n���7H�g�0���8\v��sQ��D�{��Ϩ��՚4?g?p��OOvZF��"�E�iE�	�V�D(�T��xd�!ͫϨ�R��A1���c\O"�uk���L5+r���f����1~�>π��� zb����!{S���-���Uʰr��ta�0ڻ��<�_|�����5Nr����2��FM"�P;�ٞ�M9fqHL��۸�pôXN=l<ҟ�&Dǃ;x���=D�C�S�)���~��E�HI��ř�7͊s�U��t>���j-Û�}@@C=e����r���7�WqXLKv^�lf��\R��Y�Rz��1�S`��'z	EZo�EEQk(^��&�-� ��v��س}���M�0��-�hNm�dl����AT�♟�Vt�KH��/�{_":I@VY��0��Th�g�a���rYN-x�}vf��^�j}�N�=�"uu��Th���|�� <y(��EU�G��W�J���͍T�TJ;�2�"���|aj�/����O�����fw�~�5ʫoڬVz �o�������U�$l.DU5�8���FJ�R`�!�֡-k��� n��,����t��!dT�,u������#�[����;Ct�ϳ{i;5� ����1;����ne�2�s�>| �n���[|�Zy�΁D����Z:�,憔/����yUI}���U�7s(FW���uQA���"{���q�VIO�" !�U�Xy@ x
�P�j���/I ̓�?�ע�#'������t1.�z��"ϟ��f����k�
�w}tO��vAr����K��d� ΄O���9�7�7� ��P^3PR䦉��`��m�A�؟K@�~c������X
50��� �uN
w�c��S�v]<�b��h7�����k�U��B�V�����}�-���nR��x.��g�n�b���{��}o��*�H�^��`XY�
�|���&���r,Vg���L�O��M�/�6!|�z;Ѕ�\���(Vᕬ�T"���*��Ɏ�3���?a�ݨ�خ-K�H���a��;+�\�2���o��[����'�*O��B������s�Yn9�c��`y��fK8 �>� 7�R ���햘=}&�y��{`����K�P+�����͚ϙup�k-���ɗ�z�A�����ĵv��E3�b*���A !��`!,�8�>Je�!�1��:���TI	�0��T�y޺h��a͡�@y'c�g��a9�g�;m�TEt�����=�ʲ_��XsWH�L�I($�uvn6�a��uh�� �MMU��s��G���;�-"ֺ�6Qo�:���HD��^@޹�Y�Q������%Ɋw�1Φ�LE�Y�Hes�	��1D9*^�"�I�=\rC<P�(��Vk�r�55�P��!&�gW����j�dVՉ���w�anSך=��~ PL<�ٟ�<��q�Io��gH6Ri�	���W��b�(ϣֱ�A�Eyv��}I���F��fm5�?oӁ:��S��,)��-8z���C��Q�Δ:�~�{��c�LSkE��������~$k��IGv�ҥ�-!�V�}-%��0ꭾH��ժ�_s��Pl�iCs��,j�������z?�+J�m�f�zף��B��7��t�;몝9�g��:��oT��t����z}U-�h�3��B�yER��Ԑh�R\ѩ�C�1h��쥹G��FF��P���W�A��3��!h���,�i8y�u�0�y�BZ*��BƖ>����oum�����^E3�έa�d+�D������1N2c���}�{�_n"��ņ����.Z:ʁ��QI�e��P�x�9�'%3��_��\䉆ܰo/=�]�vI ^�S���~�H]�#eCt��N5�1�2��˟�&�k^?Q�b)�E��Q�e����y��n�ZH����s�ǂ��Y(u�Rm{����wQ��
��&'��c�Z$C���Qu�7��	�qw�N��u���~זH�W�汣PJI��|��r��85-�i�7�U5����Q�z���Nʓ�s,%�L������`og32m����pX(�|i�w���hu�����6Ks��R��c�z�уo�i�h�v+�kH>SV�ȃ/�#0�����e:�쿲%r�	�G����퍂�a_6H�g�i�QW�l%|�Ɯms�ܢ*�䉁�#�xM����ࠕՒ%$�u|I����){�Dm��w�Y�(��B>��--2�
u<j��qV�Z����h�Dw|,Bĩ-��������?��ʇ�梭���P-�ZB��)� P�(ϳ`v[2_3�vLzD_�-G�#~��0SL�E8aIĘ�g-M�2�H��ѶJo�z�˪���=:��y���!�`.�mt�
���p�?L͗a*~���l�p��J|�.#hƘt��Fsٱ,� ���������0�{�//I[�9���l-�]6̓�
!� k��F�т����� �
rZH�㌳o� �T�sQ,7 ���Y&�Yk���j�|�1���
5�sb�˵����I�v�GH�����R�ht�3��g�o�����AU"X����i�������q�=��t��p�����,J�����NI��S�_R�R�0�j��;�T̯�J�A��4k��g��R6�w�1���JP"aB%��Փ�u����8-�2��
�v�ad�6��%�n� 1��h���%��s
K�b�y�V��Q��������=���M�{�z�B�-��$z2�s��g�z�ڬ���C��qŗjX,�����ml䪴e]7���8V`�P�CH64�w�a��ðŮ`+r�Js��@�j4#|��A<��V��q3` �����1g�F�>6�խߨ�?��6|�8��&Xm\˘��8~b�ձ�@0���V+>�P�o?�����>�jN��i3bۈI<�F{����b����fo��;j�[�d��YVy%� �=�=ʃ�)��]��M�:-㗮����7�>;+�����[�4��w)z�����S��b��b7��/X�
��1+�"Ck�BDQ�}����G��H�w�Š����0e��&�e�<��AO���K��;]��q�m��#:=��Җ/׀+�,����~4�1Z:�p��$�P�	E�^[*�25�+�I���5е��=�Z�ŗV"�Oo�:G��9ɀ����F.�Wy�r��"-����ƀ��R��x06c�Q<w��ҁG3��ס������`��e������л.zrM�ݍh�mޜ>����/!6haE�5��'*"� �_��}�k�������rR:3d.���(y��l	�a�.�]lShO�n��a�l�c�'Fv��jtA�0���M0U��;�TRe��F:x��;�x�uRn�(G��L	�K��os�3t~JN�7jM���aO�'c�Pyt���iT�`&��ÌQ��K�{T=��;��4�'N��B����0� S�Bh�
�x���q���������⵱��[��p�`s��D�7NՌ�����Ƣa�˯���n	E&�F�6���N/���2_���:uiHq�CʌpĹ����sYJլ�ϳi?r���d���Y��A����X_�V�l�l�꒨���AҨ�镳��W�OϦY1MfE��}��_�l����|����p�n������Ѩ
ܕ Jӭ'�o���bс�If�B�I�eAg'�q���n��'y��aᶐ��LksY���PX>['"Y�3�����=t����:Ά���o�+vO�.Ɖ@�k�=�8O��i�~��Ɇ�>�L��Y�n2Z�;f}�7g����lO^��j[�%T�9x��O�ťPKL1��`�h��,+��Rp�eiJ2w*�Z�c�T��� �֦6�?0aљ�����g�9����ڝ��{�J��$���'+��₎_?���H+C�`o�k�y�h[�Oh�2 ����(��E�*}�'�ks��p��z����P������V�!�k0�X��ҰL�=[y�P�W�PI��Cm�,����#��0��l;�oz��oq${�e�|4�f��	-����$b��\cǆms˩��h>��&h0ZL+K�V����(�0�;�ePϚ�ٲ��+m2����ѡ��$�'��N%MeQ�<�K�/���t��5Ԧ��M�H����w�qץcB�:��K�XJ�%h
[��8fj�v��qS�(�$����S�,D��OH��$���e�I}�H����n�L��e:��ΏuN�A�S�~&D���xm��9w �"�2�8Brv������o�k>����Z,����nj�,b��|��ƪn`x��Ƕr��y� ���?_��M�a�Z�?����&�rÄzT��w��W�2uԻ\���띫P�_6=v ��MZ�.��.1�'�I"*���/�I�;�ħu?Yh�&4��1���p�_s`W���Q�S�vH�ȻR=�B7(h�>.���G�m�Y+�I�u$u}�6/D}l����!��h{gL?3=�}as +�~�|=�'GDJ�K�� �1��G:�M�
c�2�f��\ӽj�I�u&�5�|�F̔�-{���fB�k�%K|��co�"�!�KN0����������k���^)�5��s�ԕ�0�2����=N}Op.�1־l?);��j���l.:P���8���H�EP(x�����I����$f�o2Uٴ9U�cZ��{�
�%5��_�#Gʉ���A��nG��>ӵ�F*-�Nti7�U��.��V�T��?{��
y�Z�;�w�#�����~')#���y�Rs�I�ˀ������I�R^�� ����-<��� ��ܭ0�����֫������c�%�[2aT�M�n���:��s�|=0`�Cwei���&��D���S>	�d�)��m����χn�	�1� *p7c�\���[ $����@��-��Ӿ��h!�q�^B��Kc>d��H��?ъB����X�@rS�Xe/��#�UMm�/��ۃa!A>�͔!�R	>A�H��ܹ��%g��#�&�B���TAgs�A�����<oEUh���n�2� !�Dx�o:�҈UqVch��4(��3�X9��k)�è�è�wG����c�hV���x�xࠬ�ӹ~l�w�o�A�!&/�L�r�㈫{����O�$�sT�/�w8É}@�t�a�����z��(,��'��UDi� Cg9{2�
<M�ܳ����6�Б=�ka�����g	�Cx��:�ϴ.��QĮ�p�����qX�Q��:v�]�}e}�����J���U8S�:*yH��鉅�Z��