��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1���e}ʲ��cg�t�ϙ�a�:�KR�%���ݧw���ȼ"~m���7",���2b�q?IzWf6t,nk�}�|_��6�� �g�a���H�c��[M���,g�6M<��%��u�X�,�A�]���DtZ����p� "a��R���Q�uoia�sR˩LZ�ʻ�g.�iB��X\��fny4�`��9x_���.X`��$�����?�����I��>Z�u��R��:�?�� g@7Xpē���
^��
9�c��'Ӽ�(���ęrn�(��NֶǏ$��xs�S� F'�㡝��6C���ȔTJ��7�H�t�U[��/�i_	L�n��x�(*�#��L�7���x��O��t��;�#'*t��(�XL�z��?��'
:�z޿�.�>He��q�9�Fx���o�`�Տr=�!jX�ns^�4j���T᡿��3�)�<�����w�?���,�u�iͩ�Լ+/�u5}���K�|1D +m�0��̅H�����X�~/]rS��X�s���n��t�Jne��3�{/#f�l���Y�C={)��(�����{Ʉ�&S�a�l>G&0��z��c7�p�i4"m}��3}<����)r]r��-����P��A���?��� ���vuQZg:ya�� 2���!p��8$g�<��+��$2՞E�.��o|���\x�V]Ꮥ*��I�	�Fx���;Pퟱ�����
�h0|jF��r�w/'��u�� x?��ѿ�V��U
M)z��Q�s{y&����лsu0v}Z]���i��[�	��,�T�~�fx��(�%&h���L�!dm^���ʚ����X`�q�ið�M��u�Z�y�
��~�fu�!mE�]�9��+�J�`xE-�O��|��y������z�	�f�gV]q3�?��Лo:�f%�7"_�̽�������1T
.�sD�v7t؇�{$����j�L|����B4](5�mt
'eI���w�D%��|PD�y��Y�N����0��^K%�S�V���gՇ�Az׳�IqEPQ��b��/�����=���?C��-F���!s_�M�ˡʉ�8����"�9�!�sV�|���Cq9@�x76��#��_6�8���	{5��:��¥���N�n�ez�S'���!O�BR�_�	i�"��$������{3��)޶KC?޵�2���;�__����p#ɖT�b�8�~	Ȏ�Շ>��	�h���y�V�|��3���1-}��p�5!#��DT�����$��7!�B,�s�aښ̚��5d�4^з��M��[�}�H=�ד�o��)�I"�֎���A�������F�p�>���Ax�8�����Y�>���b�#���a+�3Y�!'�3Z�k�GJٖ�v1f�VgӘ�v�7�u�y�M�?F�7!�-�V.��U�0�V�ef��TH���h}&�u��WUݗ2*K}��J�Jt�G{edd�"e�#n�/�s��v�a][��[t��bn�� �""=�<���QF��ь�{�d�A�H�Im ����� l-����
'���:�C�r�T��2�b����	���rb( �;Ɋ�}�;R���\����ߕ�̋̉��v�	%n�� c�6����YG���^<}���ͬ��'��(�����v�Ȟ�l�T�e2̿�>�W�5N��w����N���J�Ɍ�y�Z�F�9��;�trID��Z^N�և={x1�4��#���l�'4��d`��L�@����c�+�D 3u�����-/�������[�r��y;DGwY�����=|��y�u��3��۾]�1B-q<��:yψ���A��<���O�k�T7�b;���RA�9Ⱦ�%)� ���!�z�G՚��kG�lΑTz;�4bGn�r��ѢB*w8W�~=(�_��e�BDߡl��a�\��Q�4�3D��A��ˬBM:��d��g�(�2�⻰��W0�����} M��1	'��^�+P���� ��鈑F0�\#<�B}�bn݁��T^<�N�Ѱ;����:��^����bS8wN�[2����\�1�J��o�!�+=��F5s�$^ޏ˼ ��H�=y�ݴ�ZU��s�>}�'��"Ż�r{e��[���Vv{a�ؓ�F�|��,��Y���N�2��.j�p���7y~ 4�4?�s|ৃ�\X]�K�n(Z �4�����X�.oB��0co6ӫD���ր�D�ѩ(��D��%�� �m�z�%_c�](�wx��ٹl(w��c���f����(�rk�1��p	��
����(���=�#F�y!ENBI Z��"����S9�&V���7�V61��Ncm,����2 ��l��\����N�$�'�Oȡ=l"Z���Ç����4��f.=�O(��+����d��o�z#�YE�v�	֌��0UV���-�!��[ �>�M��<�;>%B�{����<_>	�8hx,d�ɏ�6T��m���v���kA�>�?����C�.�F+=J��w�#��;B���&������7��gl�)��(go��5�~6�4Вao����^�
Úh�Yݩ!�̔j�4\�2��a�&uQ0ݦ� 	�����=�
�O��}�"�:�`�٣������	��wo��	l���;��,���
�`��lu��6�S;�X�����nEa�+Cb"�g��=�Zgޡ�@�'l�"Ƕ�Y)�cA��QPi�,m�(pi�ٗ�>��0ۣ),Ec����+sIQz*����r����v5�8�ٜ{��8	:����H0\�1��쎚�OE��z�T��?\2Q��4��Z?�Q�~�E�qP�Hf0r~KBI��ך����8ܞ�$�`�R�.0u�5�s������P*X��Xe�вt-� ��S_@]01����!�GK3�?3�F��A?����E2���M
s��8( ΐ�D��Vh' ��]�vq��|pj����E��pw����*�񠕵���W�\�K�d����7�N�Ѐ�Q���!�o������"�{�p���{�b��1�E�%.���S0�n!��.EэJ�[��X\aeۤ���Z{lᛊ":=5v��.�N>���_��_=�7F����l��*� 4��
�� �WFpm
QU9�p0F,#[Wap��X6�R�4��%�fC�`�\4쑇���m�`a@yڒ���7 �R*-�[�E!գ[⧜�I�i}]��7.z[r�u ��-]?��3>��Z�'���J?����U�G��h�/E�K#I�5�p�E�P ����6$���6d�}{��ږ�)��$11s%s�w���[Z#�����=1 ��2v��ה*��6�\�2�oT&�����G;�ɜ�)w����O$�������%�Oڟ�b�n���au�`���iL��*�E�}OZ��I�XC���s� XE�3JE�֊.��"�	y�Vn���� 	1^s����0��|Va�^hf�LhᰓUYY��rm�!���rŏ��jA�YW����ҽ�@	�|��{FAU��m;�֘����:3Cs�8|-sz�ܡx٠��)�k�u�z��Z��X�	Hp`���1M���ʤ��3K=�/HC���)ðF8Vr����d�a�����9�n�C�o�4���5w�jxӅ�)˸���\�x)�v�ǥ���9�e�
qy.L@w�3ߩ�fbc���|���r��=2Bѳ4e�7���`�Rt�M�ƁËe�g�C>"
�B3I�|�� r�#d����6&lR�K�r<��/�����So7��[�o^�-����r�V�*|8ufǰ@��-��o�j�;��|q�gE(�Ì�[�-�3�ѡr/#�s��v8"���d�SIϝ�L8�����n�[��L��i���>�$�S٭r��5��V����Æ�'%A!M�t��\Cq90消��V��"�;����ǘi���5[���=+��O�a��P��������
�[U���jwuH�D���De,3�ٷ\⷇�n-���8�>�D:j����f������\E���+Sw�Y����9H/��5F���@�ӹ(b��א��ڈ�.��>�����w�u�33������Sr�YƖ���W�7����\��7ìE8ڀd��py����"51�"�XT�Ķ���&�y
;2"�Z9 Mq���P�%���P�Tb�	�Ɠ�5����2��"���'�+����<� |G��bE�5���d\��䡏����>����Z���y�L簺��cy�`ӓ�Mj�U�����(o#�epY������E�&P�K7(ax�I}�O}���>ߏQe��:+�ЩB������K`�m-+WG��Ay��sg��/�����3S�ۜȁ@x3\�I��3��E5�<���ԭ��o���*��*�.�z�I� rڢC� &/#B���3J9,���!�d�<B�H������;=b����OqԮHt?#���*㘤�)ީM�����l��j� �� f Q�,�+�O��#�����1yvz����¦Uc�1x�[h[��( �w���O�2!~Amc$�}2�1R���Δ�K�g!���{0�H(۲�4�(��E�)&w:8��(]~��,��A4�],lk�	ճ�Z�TY+j�Π:Z�H���\��F@��N��C�y�����U��NZc�G1l/�R�"!�iC��`��x�Lt> �3'�4D'���ӧ@W5b|r]�9f�� *f5��5kP��Mˇ�D9�%7��a^n ���>�b��{\�nJx*��,~�I�7Ɔ��[�D�Ia���Ir�|�⦏�'�#\2���mȬ�<A��P��ȍt��Ƈxܴ�s�9�Q9�"��	�K
�K�:4�U���3��u���&WZ�;1>21]y(yZ`��E� ���z=�Q�%�|Y���-�ݝ.����t����������!_f-��� �%����~yM�.L�"�w�r�ZyE�E�&qO�v�l����;~�N�Iޒ�NFv���0�������K�����ѵ=�������,�0��^�(v����e����������['�J誣��t�l��	�
B�zH�
��U���!�> wpD _���x������k�.k�3�9�y/���c|��,�7����\`�$ߚ�;��ڔ�?"�TSw���8�WdsJ,�%�L��
�րkS�4�c��]s��{仄Ƣ��m)���(n����^�|,zr�q1�thOz<4K]�e1<��g�T�$�  �@cڙ���l���6;�P4JD�M��x^��X�E�{�rѼ���O#@�9�H��	n�ȥ�t}��C�殭�>@��D_�-���tZ,�kj"Q
�"z�x�z��x��%��Yو���x��ܮ�̝�o�:�7�E�>-�/�M9��aE�'��`!��I�% ����go�vg��r����&${���'�4�O���f�ӷ������]�:֦zpٿ^�]B�!�`km�|��0��2D9]�f3hu�_R�{�!
��K�$'(���Ț���{��<$Y���8�Rx*<A�R��lz�c��A�CςI�x��n�	��y�B�v�Jr�@�#����%��n@Z�glU�#2Y��j/�]�����	e	�RR�Alp%���Ht�9'`�7mv/ol��F�%���AډyZ8�=/��PA�Mrd�ς��<�����_��k2?�H�����L��� �BY
2L3�	 ���B��/O}��b��Q�ہ�&	[�N.�J����]�\ё"��g� z����]�x�eU��]�8�~a������	�k�K������=g���|�]Íp םU	���4!d�0��d|����H�M�]N���;<�?$�.���{�<|��E�qn��*G�у4#pv�V��D�h��2�V������M���p�*a��}�cR�m�e)����R]�*7��<��cn���VE5Fh��9Z�F�Z�P�5N<��';�DZ�`����<�;~��|�)f;��x�eN"�]���HOb��*��,�M�|��dx���rƔu���#�u���|j����j[-�Qw/���5�[~]Shj���n6� ȭ��O�i���=��{_&jc�����q'Q�P�5���+'�Z�WM�34�m�eo�)�v�.��R�i�N8����ܵ��Nĩ7�x}�@~��� ����Q�)%�8p��[=�0_v�e.P��j]D;��Uƥ�#s�Cu��H;��J ��ȕ��PJ_(l�s�{�]�y�?�RE�[n^��Hٔ�O��r��7zp9�BV5K~8����c�?0�����p��/
���qQ�w�0b�(`)u�* �#s�ȅ��$�D���c{��_�n��5TdP@��D�_L|\H`�HvdA|CΧ��z?7�u�.Vz�i6Z��ŵ���6��B�+_ǐCw�����MnH0X�|ݛ���Η�ثX�|��`^kD9'8��W-��B�Y#j������|�k)E���f�τn�;�+�E�Y?H�	M���,�c�.��|^��{h�P� ���J�(�m�:��8�hw�D!�&m���7~+����_���y��4k�����z�f+qj�����v�:��8���$��9fK\tf65:��v���U*-��2����b����=���8�dy`�3F+0�Λ�'�2����*4"���0^��z�)�'W.⏏2vl&,(b�g^�V?#�Va�{p��)ҡ����� �����y�^��+OO���ý����@6G:�JQ��h����Y�B]�f�C?e<}K�J�F���3O5G!Z��[�?�)�9���I�wR���sH��z��I�p�B���
�a	2��[��S9���.�b"�8O���n�ڃ���?���<fiP*+GB�p�E H�eʘa��.��g��j�����FiFtw�A�I0���Ǌ��m�v���T(BYl����N��\]�=�=lӼ�&͡�l־@2t2�?ٙ��[��wd���8���Dͩ>>B�RP��旾<LɞТ�\Pz�g�Ո��S,j��V9cz0�e�X�jT*��6�>�����v�G���3S8s��ڈ&��xz��xZ,&eN��#uH
�k��rF	b;���,��a��w0Ho�"�A<�q���*7�	��{hm��ø)z�\c|���` �FY��%�}�[1����:�!s�lW��Q�ޭs�M�ctqbT�]�����`�2�2W& �*'�oŦ��nuJ������ j�K
�=
��)���J��E��_�U-a��}"eC���RCYsA�왆�//�R´�.�B#Nv����v��=^�$�����c�����e��L�^�1`��L��A�<Y�L-���6��hVt�tڌw�ͳiZz��Z�K&�2�a�jAH¥��~��+�s8fo�չ�j������cƏT#��ڠ������'��٫8�j����fI�_1B�b{���6g�U��$�������>j�)G�������j�+2q��B�2;X�O��1D�p��챭$�#�
�#1�ëDnT��^�@�\mt�q�/��,>��MPEG��#��i������q+��/]����YFB7zc篌IS@��-���pY�D S)�R��+����4��'����F������Hgn�Õև���2�W(F)#D�#�`v�[���v�\DW���)�`��9q�%�N����3���'�C֑��3�7�3�
B��w��%�[��n���]�t�SH�}�GN%�S�����~�Ѷ�2��7.$��K.t�{�Rx@��Go��� ��}R��7��>*��MA3��A�x��f����u�����LBpX���^��iT��*Ĵ˶`����w����Y�N���WrC�D��H��`\_��:�K�[�?$6���u��g�T�W�W��['��d�Z�(�ɢmT�۪W\��1`�=9L-ͭo����粡���+�Bw+%�f�� ?]ϣ�C����1&�]J�bS��lX�gon��tZ_�a�-}�I����W���ӛO�?y�=�z��f6L[���m�����k{�o?*5lh~ߺ��?"�"
�<�����}�=��X�#R;ߧ��:����J��2^	L<\}*�j�����A�B�	��^�n�S��(Q�X��}j F��]��.�7��_�P�*���
2E+����������a�R8�Z��к�3�����K �L����+r����������%���?�q�!��g�4br��$E���-(#�1q�]Ẉg2ͮ8�@�Y���H��Ӿ>���9*~�C7�	���%�np�o����9�,O���غzp�d�c��h���y��q���هϕ�ք�3�@�5����N�&�7Y �]�S��W�bĤ��B[���/b+ٙ�M��A���iܳ������e��wR��/H �|`3����V�o�`&@u;wqS����Sz<����XB�@R�lv�p�&��?;�#�r�ם�3�caC��`��T�U��em?��aI�m�V� D��qF�E(���N��<:�����{?Q��*UH�s�C/�,׫>��V����:袩�j��T
��Y��r����l��9����h�iڬ��/�9�md��i��`���Ue���λf��=O9�/$��ΑЊ[��ة���n���fE#W�\�F>��� ����G��w����l��t��B�����د7�$�	& ���7E9�ӂ�n��h��m (�D-�E�%�o�#5}g0"�TH���\%����țt!3�N��N���n4�Sv��B�b�������$vk��ť)�W�N��fu���J-Cu$Zu���KvEJ��k{M]��/mh��JO���4�ݦ�V��DD���w���oX37B�Ђ�ʧ�����&랚����\n�M�ߚ���j�a��V_���5�X�7���yH����W%T��!��)��6�p����*��k��g	�ok|]�3-qP
��Dw�y Ri��KO���Iϯ�QoU4���,\�ˉ�RA����X�����{?˛��md_����|٦�^ A(��!�TI�[7�NF�2
\�G��I�c`���U�wuãd�w�ǽ�ќ0��c"�LXN���:.H��h=ɡ�~����+�q�����W� x|!���m,�@�Pñ�uߏ�
N��xa�S��F�?R����̔�{"Z��y��V�����xjЋ�%}"y���m�'�w{�P��Qƌ���x�󑅂&I^��vA�@g��DOq+@��c�^��\ĕ|�3A\�H�;:'�q��I��i���髝����{�ő%����B	} S�Ҩ�	܏:��ݽ	ˋ��Z��H婏��ys吏��Ά'�2��+�ٙX�����]�D�}��T�=R�'�s	�Lp$��Y���Q���~��^�P��t���d|�C�;�"a@5���,2k���pg�.��}"s�'q܇��x��Ou��@���R\2�AF�J5iv��]]XJwȫ���H�-��k�-�'�- ��c=��ltT�A�E�N{�����J��J~����2.�Ё�o��g��/�2��$X+�{-���V��������=j���wR�����x��eXvY�������<�����!�KN����}��H�.���&�D��6����~�0m_0������	�as��xfa�����}k��ނ$Acn^�-��/��ބ<g�xyέ%z'W+eo��i��@�HP��W�X���+)��(8�K��Ʉ��
������O��к����7��i�|�H���&�I[
da�UJ�ʾ�^)�ue�p�X>�'_��$��"���E��k������u�0e�ĶM��c���̬rTX�P5{ٵ�]g�(ߠl�0���D�d"O֗jlQ�Atz���^>�hJ+���5�"x�2$�����5�����3ۃ�z����H˥����s���/]�s�WK���#�~͝��J����W���\ZOP�� [�ak;|�i���;�S�D��S�nZ���x&�%��.�HHV��{pF��AC���>�=[��pd\3�y;��ԉ�棲7`ƚ[)���&��!0�q'][ڇ�VB�a��-�ּ#�|��p�u���&dM��������>�V���|l�W�Ҵ��?ՖN����h�.0�n�g�V�m�hu6?��t��څ<8�q�a���XB���;��=բ]_g�C��ω9��Z�·�E��fΙ\�T��[����<�G�Ӝ�S�|�L-g
�x[�9��%=�lG�A0�5ލR�ˌ�T��([��2�F���}�0�3��[O��E��fhEV�6,#Q��,5X���7)�o���g����r��s��@K���
EK��5T�Dp=]����k�Ҋ�������#ĕ]ſ����
�)-f�AN?~�I����c��g9ђ��m�z�\���C෰�xQ_�!�9nd�ŭ������O�|ߞ*�_��V��������a�~�?]�8fEH�wa���6">|�u�ߪ߄J��a;��|�|��d�<f:�R:Wo)kVUF�����|)|���W:Y{f��=��:D$Ρ#����Ijr~xB�+%8�rW�47�x=	��S�| ���[�ꓖ�� N�⿚\Z�?�=�T�@��J�f9�\�*���t�@�>e�$���H`Q	��P�wa�[$��y�4��)S�ǈ|ˌ�p�<[IH����73��ɔb�o�0��um�R�D��s��}�IG������@�tD]W��3猚mW�Q�⦕O~�s�j_7��͖�`���ͳ^\l���?���yU�Rfe~v*H�gvZ����7Z��:�v���nj��	Oc9:_*�?�]��_�8M�F��r,���ʗn>y<�=R�&-�Ó�4q��ʂ>��-	3�{��~}y[���6O���x��t��P��Ѐ����|?˔��r`1��J�N�C@�pU�ܑK0>�� �3$��������d"��z�Cqa�]���j�֍�w��U���߹�ڷl��]�������f���G2AT�0.6B�ue��������/�%��� �C���Ai��mﾂ�6�ַw�:�������×���۬��^遄�,�L x��޸)4��撧��>衉���L��I�Q���,,L�Gw�������u�^�)�s 0J9�J�m\/>w��&�%��v�\���1�q��-uo"Ź�{s��Jy!T�(3���Z��^5������K��Oz�5�-�u�!�\~�:^�[
X���p����ӨF1��>!�/]zǄH���ӊ {�ʮ�b ��x�5�_p�%2c�`9�P���b�,{�P?�,75EcMs��%�r#��/��ֹ�`�0N��?��Ա4NfVV�VcG&a���)�!?�+ul�0Q��q�`I���>���z�e��ѿV!�Z��C�"m p0}:啪�E�.tJ�Ujwr=C|HgO]���S� �OV�.�ZEs�b�����"o�ϯr,��X}�&d7⤨.{W��o�G��'.sD�&����� �����f�.M��:���jמu�zl*OH]��$q-kH 
	ny�Y��s������Kj����:�X��9e��X�\( %6��R��nR�䙕	實��1@������`!GA�2��{*�BS���C����R�y��$�T���h`o���q|���o��B��B
�5��w�"�;|�eBm �+I�F�O"_�A"�W�8^�.=�"�7�X������Wz�!d��;�S9�p�6�ĥ`���O�b����᰾Pm%������eA��F/#WS��7�]n��wL}�O"E=R�n��w �xXg�z����,�g�@
n���
��N�D�v�m�s�8��X�7��� ��2��/�}d[]��F�Q	���r��?�����(��Cyg����ң��/�l�n^C��*p"��D9�'����
(zh��7N'���o�pb����
z�xgŭ {*W����I.)�N���T�����]�I񁓝��^�[RK��UV���oE�P��soe9X�^ߠ�JJ����搧�蟷�xκ�^���cH�N����`]� �7@k�	�0�_������H��ei���U,���f��F���)(%>7J��Ą�x!��Do�
r��.4X���4�|����s}�:�i8?^�>�V����NRE�P[����k���eF�L�D�_(f��K=:<硢�&o�n���b����Ŕ׻�lh���f�߯�ҭ��#�(|I�1 �"��jć{�6��+�y���f���R��^}�è\�8�|�}���%8��i��Π�`�̧v(gH I������!�eVLV�#4��e9�{�(��-�/�y�8v���ǔc����x8B%����o�H�"�����; �΄3�]�	�]�Aׯ76:��]���X��n)�*b�)�fk�w�.[$�i�W���c��H1���Y��nz�xz��QlԹ�R����9�� �Z��b#���L<��D �@pN8x�䣄̏-5�u8-��q��)�2�����!��C�Ԙ�D5������BJi���a�h��;I���O)(7ȅaS���ōo� �6x��ug��|VnH]dtG/lЇ#�������E�� �? l��݃����(+��?��0 �dM��a�hr{	E���>9-����gt�`���Ҥ�̹�5���5�w	/r��jK5e��=��M1�����P��v�>�� c��/��$Fȯ�r}�J�<���l	� ?����צ}�bW�Aƍ������c'$��]��F^'I��W;�yyY��;�}�jW���*ֳjW;��H�i%W|�aMW6�<}���Ҽ*v:�����*��AC�̐�R`���b�*@��!JN�/�n�y�MY'�IC 3!�!L�AcK[V�Tn����1�-C9��0'�U�J�L���
��'�B�p�0�+��Ȃ`�3�#��?�Fݟ��ǔj�q3c��[4��+���BOJOT�^�p���N�Fnk�� ��O|
�$_+L�&�7���v�0#Pd�.�2�|�2���Qs�\
�Oć��[q��v�#�\??y��-�����=�>��Y��F۲(� �����h�ͳ����T��"Ͻ�"Q��b��u4]ɕw��Oa��?Y&!�"��ָƂ�<-��Y\��i#rEcUC�]Z�L�O���1�b���6w�9��/}K�H]z?C��C3�̳p���7�Ɔ�[hGV�A�P�"^��!4� ���ZH�3���پ�x-��������F?��Q_Ͽ�H��+��o ����L�2���gO5+�9Yd�E��=`�*��JCH�xD�c���΢����D�Ȳ��T�)��(S}�N��J���Q� +���Q�*��a���&��x���
K4*: ]r$�bD�_`�,��5�Ь�q4�����S�'6@��)�#��[��!��"��²��oBz)72GQ�p/my+HËq�$��ȸ�z�L�a7ЫH�[��QlX�����=%�˃���g$f�������q���e%8���
 �-�q�O:�؉�D��j��֑�u�!�W���U%�cnڤ����8���^����e�,KSR��B��2��Px+<���^��K��e���LpR[;V��z\;�bm�a>�p�n����9 ~9i�����������I�w��1]�ܵ�Ew�9��~@5֪LS��&�3�KƎ��S�$�=@�L�g�﷨+�%9�|�B>W_��ɉe
�4��̥C�qK��*lH�4j9Ly6e���)W:|�@}����{�;{j=�BaU�(6�*c/�
wx�T�b\_�[��jÜc����T��+*��ni��T�X�c�h�8t��F|cx����e��{� �i�j��p��a���d���b�|N��"���W�aM���!?�'�P#��
a��-?�0���u�{;./21ʬ��o�W0��b�LSM,��޸���3o5����\t���a0�|��ױ�Q�0�;wȯ�ޘ�Ce���:9_�c�$�͊z��c�Ww��2Րm�$4E·�@ ����H�GbV̭�-�K�T�*yۇ%��3 ��x��q�� Wc�x}��I�f^����߷G����|cm�61�T���$x��O�Jx�3�:k��myR�k�%�l��[}�d�aJ�Q7���V�ݞ�ߥ���3JIaЪ�%�׫u6��Fd�U�Yo0�(ǿ[�|&E��M��3&K���>��*�0��I+�"���'�0�آ��B�:xi2�Fٳ]'b#��f9'�S3'�,wJ]qi�B���w>����b���{��q;k�F�J<�HFPg���7ݧ������ԏ1\��w��t����$��*�� �k�tEe���9!��M� �[0��xz	'�b��e������]��[=T�3���	jb��$�W���$;1yI�	6LV/Ɨfy,���:12Q-ĸ�;���P4��{y�&�gn-��l��Z��Ag���h�qeh�S��?������u��ݾ)�����,�B%����!t��0�Q�ԩ�.��9�7U������gv!̼ �=�m�j���`	S1�)�$�}�����8�]�Cv��9�`	X�X��@]�_�h�E�1��·��'���=�
LP�PY5�.N�ip�~1����J[z7���_�I��daDZ�!�R��,w����0U>h�ɯ�r���S�s���f7[�{�Ē'���R�o�1�l46���XypR`q�\ZW/�p�rq�1���{R�9���A6	g��#���EܩC:7�_w0M���a�z��틡<8(��NY��t��&��'��L��%z-`w��=z��J��R|Q��*�Sf����^�/{�2?��m&43'�hW9
�U�Ħl=IK0ȑO��#2} ��c�c�Z#ۿi�x��b��3��m,5ܘ�"Ag5�y�LH��M�V7��0�4���zx�$ u�s�uI���R���V���,�3�L`���D!�#3��Kl$�ZS��Л| �5�Pdۙ�qHZ��/��%>�k�rP����vW@��r��C�*c���O{
�k�^�0��જ���	=�tr�ܫ~��ng������s�k�rU��7�/$]M]��"6�[v��V�3������J��o�W�����t7�&�#EK԰P0�!�8n�ÜƔ��ӊ�	���F�J����V�<���p��H���*A�'ϝہD	:VH�S�S߉��T'ʹ���啎�@Ju��X>���i��zd�$�X�3���R�Nغ#@�=���b��}���h�)7�t�Z"���(�9J)ѽ���N�;��f�P������_>�6�s5��y�c1w灟O~ ���p@�c�f<f�d�\�iwJ������YLm���r��jpW��߷�o��fzy8�Qi�H��&&hfT��<Y锖g��~�Ł�ڏ[Q�M�_3W�Z��No�%M��LV|�!�l�����i2�v���L���[o�������Ӈ��n������R���C,=���ǩP�>�r?���W1�ϽC�R���r�ǐ�ď�����
\��_s����r�ѵt��܄�>l���𚿬���v�����#�Ч0M~�j�x�h+uȓ�^��u��a�^/�=��|���^�9����uN�D�9�G�mᩜwd�G�_Fr�&�3��R ������V�C�V�j%j��q��|���4�����^ְ��b�y,=��q9åK��U�@�ey��`��ӥeEi��^ћUJtg;N��v]'���G9�h��}���3��GYg�X3��#��ؖZ|��γ���am��i$�����b蟘+�8.�w+mJ�<�Vwa̜$"8�E�wo�:6���4���=������{}};0�]���"jA=n���s�5���q�������
P�TnU��0����.x���R(Y��������^\�T̯V|P�	�n6 �F��X:kc���S
tSfk6m�|� �jas�m�7a�P��̴���|t�����ѕ���hxX�zw+~�QR!��cx�q0�ë2ń�{:��L���)�c�\@$�ɺ�A�:[����������H��A�|.d}����;e���?�'����A�$2��Ȟ�C���"�F�V_&�>��ʠ�a���7�d��=r�ݡ�%A.e��
"1��)�j�v��&�����M':��mFAX�x��KF����vb�mlp��`3��c��v����9p���3A5`~\-��x��p[�$
8h��G�\�e.}�f���|�.��!�Pq��m��vF6Tw�SJ+��@�i���e1�`h요���RLEy?	8�1��!����dT�����E[�l6!�Ku3�w�N0H�8L���O+�:z��8D�p�˟ &�����ސ]�y�%T�� ۸ی�r��y2����d������=z��Q�y���^��x=kp����? kjE�?���R�f�����v)�\#r��Ȃ���z�5 y���B>���w���-���G��m �m���ړ(�V�TmmjDj�]ކ.,]eIa[�D�v�06�v�L۞f��?���,ǅ�l�Z�z��MԚ4%L�N�2d�Y;ش�S�ܚN:볪���$Ċ#�N�: ��_h��󢽆"J���YIn���!�0��Ү�&��}�pAJ�� �URlI�m����4��9�I聍�qё��jJ��4m��Ab�@PM�I�uT���S��ai�C�r���3�&#Sc������:Tn��ۋQ��?�vn�*�f	J뱵B?9�W~�[`��WѲ��,�:{R�t)�mrd�����`�._/�I�ȗP+*��et�i�I��AӞ�h�;�E�0�֎S��o����3R��T���l/���&p�4`QL-���v��4�&��J`��>��װnK�P�}�0�?�v&�kJ�\��^+�z��"�F6k��(�p-��u��ӄZkyj���P��_�	���{!'�_��߇���hy���;�/(�����xLH�U�ɸU��M�Π>����i^C(�냔��-)�ɩN�R.H���Y��9򯸯���o�Q�\C-���Z�>{��r:����.�A֭'����h�A��C5G$ބ�If�$3̰�m}v��z���[�$�_��!�ع�?NR%fH�[1u@6F�A��`]U��:���l��h;��us�0��X�o�2oPŸ�W�i��7"u��S�)��+�R��h�*�Ѭ�~[��[�}dWd���	�B�ǀ�c��P��>X�}���ӳ�ձ�v�33`d�.OF�6�g_���ym�s~�8�#��xN��k�uD�Uw�o,���l�R�(�O��%�9��LsX�:�q�xܫ's4�F!���P�f��]Qb#�Y�>�i���h�>��v���jF���5΅�]����-}^Â&`��0��q�z�+IS��KO��<��$V3��&�3���ĺo�g��oq�yU�}�����y�R"B���;q��U���iy�Y�"��-���h93���g����[˱>�V	jXl{�=���4�V:=��ee���CV�iD�	��$g\��=����*�WoLɶ�ۮ����G����sg��@
3#�2\t��R�*���Y
C|���a�X>`v[Q��(~if��y�o��-�	��p3�d�9s�YtM�;93���q���V�ٵq�<�k�wp ��2�r�3�a1qvG����Oto���������~}��)�AU���a�P�(��h��
xl�n ��-t�V��ɷa3�AWC <�ZY�+Ԑ��0Ix�����+u*��/�����
���3���_��0"j��&�b���2A�gtu�be��v�)�x�/��Ty6Z˹랓�p�~����V$�K���6,����d���ƾ���,��27��['�z��[��:@T����_��]q=\=��5c���
�'�(�<�A.���qS�>Cj��&��+ך�S]�.����$���f��ϫ;�@	m���jv�1���0p*yOL�j��֭��	>�:H��v�;,����c;<B�\�4=�5��QRA�&uf"�׿�[�W\��櫢~���^i���U���E7��Hq�ҟ���=z$�{�3�8��+��5)������XnMʕ9�3���Y��^�@�:��ڊ�#R��!�,���܊�����q����8'7SOԉ���=�8�K���e��vKջ`KX�0EB텻��\x5Ӵ��z�-�p�"�n=�̐�Y��QȮ*��5W��E�>�Y	��Q,�"�vI�t�G#ov�A���ruR����	\L4������(�h�t�b�ww���E�G�<��+F�8uq������w�0������Q�%o�F�H��6~���M����*BS7UA�Vr��g���0�<��`�x4���Mj�z��z��V�X���ua�-j�xG�fp7��\6�SQ~Zqm&�,��tp��.?��zܑ����q�B$�W$dl�B-����M@U�~����%,Oe��i?i�A�G�_>TF��wp�x�o~6����N_9j�ȓt玶�����������OϪb�ϲ{��!�J��H�&��/�'�m\
��2h��Y6X��pS��8O��L�$�P��5*��Q�,�䅫��w>aq0�NC ��QU��C7.�[�:?��PH�osi�E����d
rُ5�Oif���HD]���SLK�W�^�;�N��A� t(""�&��%������g2�ҠT���
�Ry6����K�����q7���H(Lecn� M�x��)�Ӵ �p"; :��e>�s�9��O;��y��3�ӹ!���X�$�q��9�ԁiϰ���z0�K	��"��N�چ�^o�@��ժ�eQ�Y��&D������n�AV�����N	E�	�Iꀕ��#�3�e֋������M@��SH�R*�L;�v�׾����R �5��"Y�@��=�uB