��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\����q�?��e�I8�b�Ǽ$��"����ׯ1�V0���9��";/sE��ƛj�n~��ߩ<Z:񴘈�.�fN�Z�K����N|ǈ���)m������Y[L���a���
o6�ך��Ms7[=�v�j)n���3B-OP�*�B#�3c�kl��i6R�|�xJ��2:e�3��ӯ�#��s���w���'`H؆�ͳ��=^R��9��"��{��l!�/.�Z5�8n>o�>ڟ==�~������D�Vw$��'�g�J���s7�\�xF=�Y�/��|<r��;�NF-F��%�����HB�D�wfrI��7Qp.�����`��q8
�����b0RIX�v"�K��f��8������xJ�Œ�{��a��z�y΃�M������X����av$�k}q�d����Yq�A���\����j�d�Y2�F����E{����&�>��i|�ʬ "IۮG�4 ����$6��e����*���,3y��F�'�Y6;U�T��'�?�]2_<4Y[VP*KK �*��[���ڙ���h��p�Ńn�Q�)Y6�>ƕ�%p�=��?s�=Q�0lnh���N"т�Gtk�/Y[���ېL���0���ҹ���lR}��a��uN��5��5Ɵ�(�z]�Mہ�rs��A߇������~����=t��x,80?8ן:��K��ѧ��J�f������0�>Wf�S=|��I��2�*B�m���GR���K�|���O��\θ�O28v�XP�Hv��Tz�E�a�Յ�|�N jQEd7A_q������ʍ�B�a��&�]G�ii����������h��_İ<{Y{�������%ݜ53�Y�J���=h�(���Y��0���v��p�����(���lΪ�J�ԛ�4��b���m�Ω�䴳�<y�=��4[�C`��!3bٝ���PZ	h� �p3�mp�N��S�I�H�¨�p?L�J����[��d�0�;ԇ��|)��v��L��+z�ݭ����G�C�|i��1Y�[Չ;�&_ނ����vT{J��e�-�?�Q�z�L��d���gq�s*�b�V4��}wM[�Q+�>�X�hu�:�SW9�B�簫�Y*�<T!��Z�ϝ��&//�gܧ�굮�^��zZ�f��t���V�x�'�[-xd��������g]�)\�&�=�&Wuv�R(�����{��n��۸n�)��s ����ro++Ҡ]Wj��=J!�����jÑf6��Ij8,�6У�z8��^�L�OTD�0f�@�����20�Y`���$�"f��$�U�<�P��w�ҪZ��V��@��S/��,���\L{�Eߩ����Ѫ����3��hm�V�Q������_r	q�Z�����)�:w&����
��9�h�b�ulՍJ�pR��T�1W�V���g��k���^�C7����кc���l #�Wq����!���V9!ΰ�-�4�n����.M��>&v4�%U>�5"O��˴�/��,��U{����Ul��!i�5�0EC2�4S��� �S<��b&�W�m�BjR\H�큧7c�ႤI$/�C�f�_{L����>��V�k�e�2 �Z�r@z����6U�Mz���iX	��ooc����4��2�n�� �Ĵ�ڙ�HjT���_��	. �f��#�Φ�������ު2�K�@�Q{T����( E=�~Q33S;އ�JG�mm?w-���<�Ϭ�Ư�7�S�z>P!w58<ɞ�l�;���3��ܧZdc2#��қ��� ڨ@`V�@�C�ɯ�)��ˊ~��� ��٭ޡd<���6c�'�s]SS��A(Twf���u�V�����wT)5��٨<����n�>�5;3����UF&�y�c��3�-y���\6���M��6�K�]їb���r 7���tGJɹz�E�(��C�Q�9�y�����i;��V��2��V��v�_����~���R	�'�Đ{f)7��ˆ�-U|IiKY���5���MVV`��;�l�p�`��z��*�̳�|��l ��H����-��^���;Y+J��r;�Ɏ�7=��`p��.L��������7]nF�s^���³z����w�4G�F�X�0E��On�壧�֫�;-ʾ�{����`��` �RR�!�u� _{`w�y�L�v4Ls���ݭ�������O��eck�Wc�GrJ(1�o	�Q^�v�8�?�[�eÛ�Mj���P-�K���Lh>�0��b#�z���j��eN�"@�Q��0�5@�)��I
/\��`ɻ��,�����+5�|*�k��NPٞ6�%��O׀���+$��V�!�6�A8[~/��YM+�����T�F����Q	S�_c�ѩ�v� �6y/e�L�:�Rg�O���G�D�+�'�?�#� ��ɯ2��ڟ�S�IC�&�e�叏\�������@t�Ag�(b�kn�� �g�R���PE 4Ŭ(G�lA�~��h��k�I����a���&M��;��xsg��S�!���e�3�3~ב����.�u�~��Ix�2�O�\*4�&������i�9��\\�~3ƃ\��χ�A~.��z؁J��R����	c;�����Ṃ�	g�s���4�<��E�Yt.3�t�l��$N����v�ZOʞ��
U�X����N$V,2 Ms��?�k�?!�&\v��ҏT�r-�! cx	���W�&_�}���M��#���H�����#=j����\���$<�\���1�u�
Q��3�t��"&p�g��gk�tWi�G,V��Q���4C�RI��2k�7�gj
��6�����~��(�����+)�I^�*Lde�z4���]��(/0��KX~Z_D*y(������ȥ�̦�m!i	��[{bɦ���\���i��\����_1�.d�gb�Y�h����)0^�/��_/Jv���G�2&�j��y�~@�u�x=@�uY� =���C�Zh}��"%���U~mV,�ʌ@_}�� ._s�|�S[NfH��6;+#��2���<�����,��2.��N�J83U�Wb�iX��8�H7`tM�X�p1�3�iO�-��L�Ě��>��w�dm�֥պ(\/�FQ=������C�$��i�π{π0M[
9�VQ�(���zn�LU�[�Ϟ˖(e��{.��u@Jj	q�O�q$�;�*��ߙJ�C��@+'�j,:q֩���<�N���wc'�[u\��.��wT�JN{� �JcZA�L�PK�c"6�qqC��H�39"|2#8.���"LN�
WlҌ�9Q��7p8t�7��DM�tȀOn]-$���+r�3ԯ �2��Pp���ά�nB��X�����Ș�j7��s�X�S1�Зf�7���	�^����焐�>4�"!EB�����Q�W�J��Px���x����r��¿&BX�qt��X�rpb	h)��[���g���<�i�� r�D�<M'�(��%�o��6�\� �"3n�0�=�����6�����Ҁ�G��l�U�R�XȨ�J~x�pԈ1�K �%�Y9vy��Z>u v������ǥ��}���/�z��nW�i���/��e�6u��᧎Q�Q��Ӥ-0B_�$���~;E�bk�����գã��!Yf�rX}P��zP���(�A3Cz� H54�]��h��b����8)�9 "9N���nK�|#ŲT3�M�7_�F����D+��?o�b	)���CCm���~�����%���|ً<�����qH�9\�0��GT45�b"�L�o�!}�*���"_r�׎�EU<�˰�����([f-9�����:�OΪ�L_�B�k���t6:�����%!ST�~)Y%%·�f!��c�}�3FX5����z>C%�ݿ�ae���A�(���fʈj���g�����g���R9�-���J�$��hQ48�}c�^�zr	wQ��\J�	*n���)edu����4�z�f��ˮ�0
f ��ԗ��J�]w=quł�V��aMu6%t�Nd��b�?��E��><��Ưq�7'�� 3l�+����mr��|��( ~�L��q�]��Q����+o�����O�^��o�k��=��+ѓ}.�"�O>�*sg�nm���W�JJ��	���y��路-��f7^�$�,�ӒU\�#Q+q�yf�NB�2�Q�� �VUg��.>��+��C�AC�q�<>��f���p�PB��R�B5�:�G(\�n�M�+�b����HO��lf�,��u����{w�ZI#��d�}Y��Q�_�a��N.�М���Ǘ�¿<��M��o��T{*��*����]}	12�J�VU��8[G����?:צMt@���g�A�l�ls`�|vY�J.v1�Ni�Q���ivE �$�E�M��)��B=��+���{Wq���-�e��2�e#�n�<=��bD��6���β�4�����h?s]2���&sB%3T���U8�br��!�D�GtM�?A̴��$�������a��7��^��� D�Kfh/X� �_F���=���+C�e��A^��f��p�Sy��w��$�ϯU���א	xf;8�L�IAF�PJ��}e��v �T�zoV�%	�,`���d�B�E��>e����i9fZ�e����E��;"㵰"�s�&{�zǐ�?�1�[�������������m�
�%�цjc�� �N[�,��#�`n�O	��{�  �����F��5�N*&zȮ�X 0tazk�Q���Uw��������8�n�9���H���.U�'�x�k�*t蹪�U�6�|g�N�ϚѵAq)+����6�pS�E����M*[�D=���$^�x�t0�Cނ���6�����T�P����qo���YN1�5 �b' ��������C�m2e�4�| N�^�ޢBT>�|��Zz��c0�B��"b$ٺ�hz����
h`ؠn-���xF~��t/Q���:Ew�>y��3����������������j$,~���a�k�2�g�I�C��w{���m/�A��^�V�����/J��� i���a��S4��L��sw�X�i^q��ea���*��M��p���E���J)Jj6��\#�1��	�`5��o�!_�tz��"Bt��#�.�_��9a:����̬YG'Р@)�=���]�x�aE��2�_�ef+�2�4h�#�	W���0��Jr"F m�	��\C���MB�h9S�'Vv�ܱ4���9�9��2՛E �z�d���l4?��~.����,~���N�Ң�W�-�<��=��G2�����f���DҶذ��5�=t$�O�!&Z��)�{ ;~��Ӵ+��Ĥ���R�M-]�u m��%�;T����i��C��뎵����c�8kwO�C��c��4�05��-�8&Rc���N��c_As�.p�����:$2b۠~�u<��$'��>\��=ǻ��?{;Y�n���+�X%�Hw=�/�$�H=j��5W��9�#}�������&Z�{�-7�0�:��"� ��@$z��Q�����UB��t	O�A���4N����2�|x��b�wj��7SU�f70�C�����*�B}�ov�n��Ж����l��/�*�5DY���'䡒�L�Y��0���h�
'#+��6�[u\ڲ�4h��c�oC~�ΣY��L�ݩ��|���m���&�͆�臢h����Rhw��Z��.�|�>�n�ۮ[R��תG}&�Ӣ�Y��A��-|M�n'�Y{�'����7�n����8�QaDW�ܑ�Z�S7D�=�j}��5+_��#�|�K \��w�3X�MňX/o��8�{p�ʡJh�]����{жH�,P�a�ʚa�i�WF��~n��tc��lv�n�Ӭ�L@�dxe\���Q�\'G�����K�ujBY[� �|��E{
A64��t�3����<2�Y�Ik�8F������;]Ö ��FMx�A]�W�T��?�i4R2:+G%��K�����w�\XIM��w0b�uX�}x�j�Q��0U0�63��f�џ&t�� �4�*]O@�Zo����c�(����'�8��]8iNE�o&�u��ͬ���z��Z^Pr�:*����~el<�1z���@,8��Iװ/As9EÖ� �O�H��*yq�@444U
:�K���t @�D��$�Fف%S��~�h����h���k�wP�X"��YXo)���>�p��a40
����I�UJ��z\H,�^�F�~q�s��U����4=)"l˂� �SZ�B/	S9n�o��<-Ԅ_9!n܀k��п�Ь�Q�KP�X�l*^5��>R��Y����n�q�ȳkf�R�Rh�Kx�G����X�L	(�Y��O	�w�ԅ b��Yȿ��l�x=|G
Zչ1۞�������&Dc�ߔp�{ņ��������s-��g�ïO:3�(������:��<�7��>�]�͘�nR!�yq>��CE��Ұϵ���>��op�7��i⹵92׈pBds.�#�#�u��۹?]E���� ㎀9��r@,B{��y�i7:ߞC�Q�n��M���>�_��~�%���ZoQ�̢���H��ߎ�b����RobLK,
c6����X1���u�.$�|�E	~�6�R�<$ C"e5���Pr@׺�U(��ST�(d�)x���������&3�M�Egi�=�i�Z�z��}��Y��q��e���g��p!Q�@g�F�D;s,�\'/T�̈́eH��
Q^�T}'X�y ���*C�����o��"�;����@X!��Wi�2z�@��,�K����j�;(��аB)6�^2:>���܋%��14�_���m���A�9�Y.���A�>���8��6��-��C>��q����u�g?�b�Q�Z�=@�k4��'f�U� �z)�u߾����=v��]L$�~a�$�a���+��ܢ��I�P�xB��j�-9� D�?�Ƣ�l[��/�����i���",��@̧0_ ��&GĮ�줆}ɀ�~���Y;J<Q+�S���ul�|��rH�"�G��5����r�V�uď���%V�%|ٙ_֒g� b0�����"9�d����'���*�>e�6���YK:���H���Uf&�"LP
Jt���x������wj�h�@[�h��C	V1#P
	%���܏@���D}����	^8ĵ���[p##��m��܀� l�?�u��H���c{f�cN28i�L�p�LL��$}��s�ݎ;B�[��'"������g��d�P�/Z�=�R�K���Sk��EȠ*qc�y�,ȷ�g������H�cPa�~�������
9`��v��9WS�����^|���E��fg�n���R[��Kмk�z�ӊO�n�My��@��ܙ��!+
��p��3�S���[����]\x>����R�}�ɒH��mi;5�U��9v���FV#�{��=IF���&�rd	OF����P��%�]��2:^��@k��suwSPd+��N�ci�bD<��E������X)�r���ffvf6�L���`a��*-�쥀�ҋ�&V�TVS��f"�N��&�~KH7 /�膢�Q`>�IQ��������%���u�n73�L��ꂀ'5�J@�w<�f���h�w=`"檈�h1�������é�����r�&\2���P{Y�wI����t�󦗣���k�?���u:��Կvf��7g�CS�"�wx{Ȁj�BY�VW"�:�"�S��Yg� �k*|G�=[�-�� d|Q��Q}�`¹�L�}�u'�Nd��Xrt۶I��#ޒ�`�f
��X�p6
��b�$^M�&��.��������������@�m��������"�A{P]{�.&^K` ���^N�*i]
e���읐��׳�!��ѝ�&�  
�{U�G˸��
{��9@{�������5��K1fY�cI��蒝�kK���y�K��� ~C�����f[��N�M	Ǆ
��I"��F���Aj
��H��d|��/oe��Q8b9���y���)��W�t����LF���qȵ�=�gz5m�*�}�O	�����BG�v��}
��Z�[ i�2y�L�<����?7�����7��c�u��ּ�c�"YG<��;}�&>��"LE�B��?)G�:鱟Nh�!HN&4����v�ô0�U��<�H��t���r��m(�������e�Y��hؽt�f��D�ǿ����s%F�mu���>P�@�)�D%4��Ղ�MZ���]�pR���C�?X��(�Sť��ܼɥ�`�b��U��fO�. o>|�}8YD�-.ڀ�#Y��d������\��ȷo	H��^	)���#T����w�ꮅ�f�� �K[&3�zq�S��N�>#���4e�e �����B�nJq�uyN�?�(i�Y�\�5ޒYJ�}x
(��u&,�e��N����=3��{�e��j������[G�t��o�N�ޗ��I��A�Uq�N�y$��u������|�\�Yv�R�S��`���ֽt+E�����.yG�Rx]��h�1�X��I����)m;�����@�WFkwZ�m�<��xܞG1��䝇/�F��{�׌����'���ט�ńER���m�n�������z���#$(1���������!�>�|m"�]�NG#�5pm��%@c�XJ*=�Y�?WvÐ�Tr̽B��NmY����7�Ϸlw�gUm2D�M�	��J��� ���X�O�Ƈ�Ϩ�`{Y���Ƭδ&ȩ���985���깑ג�sg�J�>	;]�	*��d��+��x��A�&�J˥ �ȓ�סY�O/3��sˠ$����9�����@j�p����l��zF�VZ-�ת�C3��Oؔ��8���vbgy 	�]����$kȞn=���+�ʒQ�kn�@
]��U[{'��Q�~�ˤ��6���5
��v��~Ku�yQ9搏�g#0��ڦ�f��#�)�꿞��n]��(f mE�ÞX$�`��P�`����63�Qi�)���: P#+��#���l�e��m��i"��)� kqrf���rQ�c3�(���^��.�2�^U�z�R~�$l�0(�Tf�q�Ԓ}�ȕ������u��$��ʿ߅K�%��c��}Ћ$h����#T�j�_�M�z�'��8��rǵז���l�f���.4����,��Qz����B�L�vPLʪ�|I�_�O7�����q��%T�]�S̢�����&�azĽg������s���3�z�R����/����o-���������t�~�!AhE_���qE��`v*��`ʔ��i���:����5�&�{��ͭȿ-��ߧ=�f����h��q�j�U;�2�9M���ɐon}�N��yX'I��|�Ҥ
��.ï]�V��f�<Ş&޸R�kV4��	Sh)
����j�lڬ�����Q�����!�"�凭���d��O��mf^[r�]b��ڪ����e�@�4ҩoWXE�z�(k����y^l�$I3.�=��e'� }�+�8���"=7�+��>���O7#��Er�'��Ѱ�JJr[ |_���_}IF�:D���B��drc>��Rz��c����0��Akނ��9a�|�ztߕ�>�C�zx^�V���"˥�B����fk�j�Za�qe�wː��;YL�}�X�T�Z
Gs��os�"$�'�6��'��(1 ϐ������֒��*ͩ��ŠʹM�k'�"����yv~�Jd�D�i�l�9�y�~��Z3�j��I�'�dk}��r�w!�K{�(2br�w�띟�n
囷���_a.���}M��i�D"$cf}���:F��tY]qm�Y��Dl���*��b����s��?��x������tO?�>Ҟ���}�jX�ƭ�l���)��yo���ּ	h�̫e�.!��H���+����kXV�y.N���I���\�"�B�����@�n���*�V�1ߙ�3�`�=��5��������z��w�-�����Guv5� �a��;�F$W?"%���F���"�S%KRλ��X�k���gw�xbB�K�ss� _4>����"���Ƌ3eg�EZ[ �&���E� ��'B)�aNh��T�r��[�[G�̴���z����o����02>���N�y̆>�1f�����&c��1���mVQA�e6d�C�b��:Y����$kJ�@��js���XQ�_��~�sd��7�ay��P+�^��倶�=�*&�Y ih4�� ��~���2���$WK��N�:��G���ȟHtsLٻ�!��0��bl-�	��]�����ߒ���!�6��'�)I��澅kg��iڥ�7�o��� X\��Oo	��1��X�(�`�d�?_n���(��\!��l�G�5�{�EnEh�B8�t���l�}����SP�5���HG��/�_$!�V�s�ҥe�n/�@�����{3����ڣ̔��!%�q,'Tr��B\���W�T��7��C�`�(�YeR�4T��I蘟:�"Eб��|�7;8"5�s/��O�"�%}�@?Be���͝O#���,l{;��;��MUD2�nT` �fH��Tq��&*��Y�zl��@�v��Z�+?��]������2!}aN�50��i����|�Bqu_�;�C�f6P�f��΍ic�&	�W��܈188�W�
�/�zr�Ū�_�%�(%�lI&�p��d��UE�]�E`,�3�W2fQ�&eQ_��q��L��ѹ�9�ǡn��b��x��L��n#6��{�=���p��^2�\��ѓ��-�������[Vܙ���^k�d0&#�6YC��/�T��y���F�_Q�W��!1��F"[���(���ni1�NU`�����P\��_A�ơr��g�i�Α��{�m�S&���'�0Oj'�t�;h@��7�B�ٻ��e��*�!���v�);EQ>X���"�ݺi��
���
�ѿ20N ��y<��wn��՛�7f�˸m���lw�K��d2"��p��}��o�s ��t"����,y�~_����ȯ]�3+�H#��M�A��%�XW���;��Ms+�	�U�vxQ:��!��3J�Ri�תq��u��A/B��q���3S�VK�J�~�6vpG?*�8�je"��7�<�(�@���3����U��PI�[!g@�V*���gO���Z����g�Ϥ,���}��O/�p���5�(`X.u��w		��ͤ �(>0�� A��d�,��hنCr�n��iH,���v[q4��|7�k~?�R���`n��V���ͶO�G���d6�	��m��"�!��BT0��A�,�P�U���&);Yͽԭ��B���k���Z N���HLW{d����!��S̅�:��?�ݪ�"�	���]E3�M/-��ſ��I;�I ~�h:� ����s����Uy���0����3�˻������)��eiCC���c�f�5�zim�v?�^�l�<�g�J���6\����e��\�y�B�tVnm=	4�_�B�Ho�s�{zN�T�����x�N�����6Q��s�G���W�3� ��K��L����z��C@K����T�}�:��/`�
F�.�Rh~�SA�W*���:R2ߔH����d]�K���Es[k��Y��9(�:V�%�N�3] �O ��Ҟ-O����KJ^��Z���#��rC{q��mUA@E>�چ��^E�1�O�k��9����|ڹ��n��&��@�V��[e��|��1����?�U/�i�/n�\�n6N�2�]-��-���|`��*�����9>E=r�֩����ķ�x��&^K�Ǐ�������~t^ش�Q N5�|��u�z�nr�Wm{���-g�L�kC����ә1s��a�&Q�8�ݿ�>�.��i,��n&]]d�g��FBj/1u��3N�+^�Q�7���ϸ��<��Yt��۩Ŷ����]������r�!��*&��nt�O��~_�����ݙ�d�-��N������f�؄7�9r�8�]��f�� ����k���J�!�
X��B��%�x�x��M!��2��)s{�����z�T�]j	��#rg� ��[y�'`�� v.�d�<�Q�|�
glJ��@�T �3'��N\ ��L�`a�}��h��U��T�n�$��Vͬ�኎�- <�Vd�ڒ� ��09�����A?뎦-i��$eNQ�B�W�?�B�E[�)~Zy8A0��

�o�
�+�|W@������ɾE�/5N���� �b���������޼�?���Ϩވ9�9H}|�)ك�4H��rE�2>�,���Bf����b�^l�=~����+Z�^� �
�����=������}���2�H��cG�o�]�����@(�**�@�s4=ӑX���J3�5���S�4#�`���S�_n�WB��j���a�&f�K\$��:ty��rc.�U��������T�]���DR)��yd��c���{9Y�K�{C��O	��%�7�/��U�'/v��+1�d���u[����<�޷V�ɳ�Oҫ�l����f�yTS��ʅbH�N�J�U��C������_I�2d?��x�[��R���f{�z