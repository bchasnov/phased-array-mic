��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|8���e5�I��d8<���*�kƅ(aBj���K�/YЌ��G�������y�:F���>��fF����I���p+3.�Fj%!�akL^E��4��Yڝ�ͧ�blgK�`�Ep�� �T�ʰI��?�9��*������N�8�F�D�r
�����zo�k�>J��)$� )/�y�*����[ű�=�[��a!�q�H�4.����RHuӂ��-�tȧ=�H��~��Y(C��(�CB۽���se�Q[���S���Ok}#qs>T�K��`;�p�TH�sA)u�"&�s�Ɵڶ�ka�>z�,�u�4�=AkPG���grt��F��K���n	��){�gƆ�4[|,�&�6hCozi�����N�d�H7�הe��+$���hk9���j�b�_ː0�2LX&�]d拎R~�w袶��"��~W����ԇз�!a�Ӱ�F+b3�2CQ�|1�Y؛4�?&^�w�F?Eh�Q�N9��ʵL�-�Rśݸ��gOw;F	U�u���uȈI%c��|׆v���z�����)�6�K|y�_��Ҷ�3�L(q<�",]�I�����躌�`T-�i"V�;�J���l7�e�ͽ�è1�@cjn�x��_@=�_����.����f ����I���ayX�~R��7|m�l���|�d9gv�FF,�ЭI�3\L�6>B�;!h����ݻ��'�^���H�h��H����[H�A<q�Ря��5oϖ1���RF�g�<!����?m�Ʋ�8@��#�QĐ�9%p鰥��_8/����B�y��:�s]!W�\O
�T��SB�do���Vc�B��:V��|�u4*]u̾ENk�s�M�.��7� �Jp�f���:�餮x��Ni�Ty�� w����dG!T.s�*�ɫ�3ɸJĺh��[�M�23�}��:�|u�\Ў֤��6��&���8@�;�����Z.�X�j����N6X���y6/�@�`�F�������}�
�<�eX��ۈ�3�^b�U�ҥn�o1!��J����x�U=r��{no�V���Q�����
���ӏP4`�Oܩ��m���E'����]t_!M��1 ��r�������$���!�/׀���T��m��\d0�(�S��|��a���c��Z�`�f�mD�1V�*�#)o�$"�g>����s��{1oqT�������fzn�j�+:j�~�ޱ�Q&%�����-r����ļ�J`��&&x����/�{�!���N�#8��G�>:, ���9�2l[���'�f��*���*�l�W,�����^+t��,��K�sm�����T +2!�P޸�Cs�uY&=aY_2� ���)��x1��/���o�lu��Qro����~n⒰`�P.�:�f��42|�5�I����	�L�k���*�DUD�~b4����=uGX��>�W����_� @�A{��3���7�G!Acj͵�E�N�E�y�:%��^��޼0덆)�\���� �����		`BI݈)J�/J�)�T,�|E_b�p�	�0�f�V�e��;����w-��-�����;���+�^
�+?<�Q+�6i�'&�:'�!\���2`�e ���ҸĊ�p��$�cs4��Y[��ҵ�K�<�f����:�P�[���FL������T�;Ox�<ta@cg1H+�j1o�r���������'BlU����ŇXK�>#��/��Ed>l}N�tۛW��h�mW�	��޴�#�U���P���Lΰ�_tR!��jv�ɪ��~����A��͊߬���*�d���Ķ���+3H�$��+ �S��/����"�)�+G7�]�O����)��'5aV���!�d>G����x��-T��lu�P��GQ�.*��ę�fݮ$���e�m(~�]c��ё#0㳞P��{ŪM1�#>�C���A���3yh6��9,�oh��B��w�ڳA��`��lK�/Tr��ʊÖQ�'�#�>��ݖ�$H��vZE�.9��=w�.�kGG���?�h����W5� Coa�����%}��\r%���o�;D�~bln$�JR|]q�ȓ!�ĖoB��r�bBJ�޴������C]|w�p7���`������;/�o�ӈ�VS��3T(w�*�qB��S�q:Ekxڶ�=��0",]ֻX��?�Ծ�%,dP�g.�d��Q%�ᤱ^-����1�.�֘xqk�$@�sg ���ē!�p`=g *��_���m���G�m�wg�f��FƝv�0c���zñ��Ւ���ǟ�$,� <�Sj�ٍIx��1B�����3y����6�8�eߍ�g$J`l`8��Q�e�L��q%n�� א�����ѽ!�+K��E��d����O�a����d�!��i`�J�b%+miB�8@����8!^a�t�+n�EOI�nFE������y)�)�9uDO1fx�l�����2���A���3�"׬%�1���f4�+)�֑�l7�;�ry��f���a2��Aޖ��5��1M쬺��i|�q��B�2JQIS�*��������UF�%�Ma��T������ِI�>fcүzQ����6C.	Q�c=]6�yR�C�IX �3��;��R��ߗ�M�>�3��<�����,�j�z��A��U^���.�g}�>˳��9�P�N\��V4p��i���"DqH��D�F%X��Q�:Z�0V[=tb��c�3J�_�.�	~�.YI�����)M?b���UY��ұ$xv�T2�P�}n�W��)��Em��~�{�]�މ>y\�k�Uk�]:Q{R$��pgn��,bs-P�ҳ�v!�hm�YK�A�)��܆�6�]� jd��rv~}�d[P��*�+�y�h�Iͩ�N^U�8a����t��%g�,���������=D�U,�Y��;�	}��������q����>��o'<�<����I�ݐ�N�7k~(a��Ԉ�)�JEZô�W{$����Qp���s;���^��D ��Fq�k��@�p�/!�,ׂ�;9�W�6�'�wA[�Đ�՛)!N�Z)�-~��(	�/&:o��ٞ>]�|/?�@��
���@ԖF[��W�������!$��o/�Ź[9˦���}C��ʀ�n�e������3�\C��̿E�x�TJs��)k���]�����\M�hڜ}%�҆��.`
?Y�b�� ����2F�o1�
H������S0�"��ȯ>�L��X!�����G�V� �ѧ�Z�\�O*%U�5㖺�t(�a~Ϡz�[@��z/k�i��N��GN=�![㋒����Q]*���$�E�kk�����x�,$��U��#emn\b:���8��U�X�$y�v��{eʣ��]=��+��WS�em���H2w�2��,I�<��	�g�(Ue�Ʀ���'e(C����̤�4�?�e<U��-�u�!�#�N��C�8��Fqo��`�(���1xd/Ec���.��#��`C3��Y�[�a@g)c�;����#�hm���~g0���T-Jh�1��Log�檁�;�3��CX�S6!�h���U,��ko���F_`:��kƮ9+�u^@�ryѭb}7�3��PN�T�+ ]G{� Y`�e��_���yK���0�w�q��d��p�~�.���|��l��1�g>N��NGNc����KY��t�_1DZQ��<����W��U3f��F�����gzF�t�
�!�.H];�jfFT�m$D��j)6�x�l������:�n[�����s�*/��# 1|"�G�/���yS�!UGm�l�к�s/�}7�.U%}s��Y|͵���y���^5���t~6ߒs��э�	�V��1�}S�X�����Fk�;��{	m++�s���1���\��?x���p6B4�_�S,V[�>
���3�k	qc��J�M�s��hl��~ׁ�2H�v49h�Q�Lw	mS�*�%N[�vBg��ǡ{IĲ,0�j�����>�=���YX�4,""�D�P����
l�챿IM,ӧ�ƙ�
�D��+�
�Ϭ"��u�	7�����ߐ���gP���r���i�@e��ѻ��	������{W4��yq��Kӣ�_/�#+Y.#E��6���.��DIֆP}�4���o���u�+�d2?��'T���%��0��};�6�>�������ƅJ���ԙ!"a��j�����#����*ң�#v�$��@cZ��.��$���O賭p[|�G`�T��o�W/�cFNT�e]�a���y���^P�muڒr~e�$Ӵϻg&�"���S��%��y�Y^Õ��z�sA�dA*/P�_��b�Z������ ��T˲!A�F�7A��ӭE9����N9�h �j�J)NNc��Cm��e��V��!q,oJ�qݒ�9��.���M?]�+�C/"�=��<���_�9&�﻽�?���j�T���$�P���*�2$�|O��5�eл��Jg�����J����a�1��i�Fj��qGt��Z�k���+ӓ�E� �	���$�����<mk���&�
V��Ľm����s�'?%��<V�a�[(U^��t�2B"I�6��3T
���U��u��DXeo��Y��9���8���ӄN�4�)����0��]~�
���|7/�7�\��S�FR���c���2D����d�-d�m�Φ��
�l�g����eѲ�����&�ǂ�ȭ�7����c�3�{N�A�Ыi�6"������j.�'7sp�re�]d�A��o]\K�Џ:��dB(�������{�B��y$y�~�	=ݭ���r�
�9b�d#�1�8wv/�:���� �a�1
��<�
�a���'p�W����)����O��T՝.�'��R��7?��ꏹ���"�J5I[	ɏU�@%�P��Gw�HYk�T���eH�b�ԹݼE�#;��CD#��
���I#��ΆȦ7�w���wEkL��2�8����հ��M�̧CfӰdb]�������l*ᾬ�5Mo������ 	�K@�:��;��I�^����4����(����Fco7,�WȂ�~)MnuM�z�C���1���Jƴ#�g2'zf�{qX���';2�8u�K����vQW�4�!����B�!��}3H�MY?f}�ҧIm��$��f\d;>�).2��N��/�B?b�P�)<T���e�砡{��pW�aV�_#@1Vm�QE�uB���4� �����s�$8�q�|
irȤ�M�����Jr<�Se�H��yN��%^���'�d!�G5[��x�Z�sj!�SV�>��!E��;a�+�ڧmx�+/�1��F�Y���oh'�n!eC^������ۼ�C��A��岓1�SǶ u큾ӯg���s46o�Љ%�zA��V�����#��׮լ�ȧ@B�qU7��4k�����x�o�j�Y:��t����|�i�}�Z�4&�)6���5(��v�$�I�����2T5�L�W0�ȨM	�Vw�5��4��L�p�i���tI��N�n�l�e���B���E�\���ʻ��<���tX�u�f��.�Ǧ�)����a���xm�"�~UM2��on�+2�V���=�Y����r��+��:9-F��z���Db�����8�P&q7�s���J$�^�8]��2��]�Cu,���t�k�H�g	<�>,Bκ5km��(R���u���5�qi��τMH��dN*.�]������X��U��t����֦����ﳓ�-���7�0q?��3���@����xՊk�Tm�(��� ���}"Rt<���Z5��u0hd�m[{Ņ�kJ�#�Y�2��Q]��=]������H��
[��-:��u`���v;�z=�u>�*�$���Z��<;��r�������	�h�uҝ2�A\z�~Bm����Ρf�M�%�����G����0J�c��;Gu:�hE��'m}*�i��K`�M�Z��M ��B�}�u��RF�&���E�'HwNϰ�o��.+����3�V�=0\D.彛�@1×��&eI���B���O���o(a���@a�╉�a��}������:i�y{)��\џ��eh�kR>� �G2A�B�X��	i�@(��2�T=;
�/>�:*�If�&�o��~�lg(�c�:�%x���v�&.�Z�$��n�����%��8����7,��rE��gu�$���&O}��n���j�o�<`#Ŋz�=�2���3�W�E���q�8^ g #��/Ϟi�y�����3�E��0�(���B�SpM[ ��ݐ���Wy�8`z��IރkN��=K� S d?��B���E�fK�^���i�Ԉ�I�"��"Im�;��(��s�8�F�������7�je�{���֚�8c�𚵼��vڹ�}%�=���2S)l���>k9!^������vp�_
�� n��MHH.��d�&�KA�~>9��s�.��0�FK�:�T�n*��-gГ妬2!zAbQr���9��m]�%�`�����<FytP�r������p&C�_�I8ݹ���k>h����]���_9���O|��ນ�vҚ�z�ai�b�T 7~��u[��,��o�reh��3]����G�{��%͸�f�'ab�7QP��]��q�	-_��o��*1tCKv��Y@_e�{�kw�怒ʮ�4j��"H�,k{?��U�k�l�U�2;��8p�[�٩���J�E��ꡥ��*��K0銐;qp��OH�����0�U�d FT����\9���э�{¿�瞌������n��;�!��VE� [�����[�Lk%�����0��^�M+�>F�݀��+�̳�������UZ��Tc0x.8 �兄}�Xi<\��YLX�FԉK��R�l��o����'�ix"t��*Ky�d;8$P/��V._1[\�)OV)���Q�QQ�<-;��rUK/d��#���,�α�X�V��?W'����)�ѦZoMr���Be���(��0�i��a�1>�B�G���'��EtJ_;����n�le�tL����5�X��T¦XI�6c����d�<7��`�)Yy'�?��1;���+�k�C�m�YnN�X]�`�����_ �
�L!2�2j�V
&6��OZ��[� �7r$��v[���I��q�Q��g9�
sN��r62���s-�`��X��~֦���S����9��5zD��
���|�}�=A��ԠW�i>gPT���p�?e�2W�;g���Z=N��R��&��C���Y��S��-a��0�������r�ZH�v�,P���J���&7#C�T���Q2���=0��?���(�tɫ�10|�\S��ZP��Y�{ ����8_�*���K�-���~yw�����lۧ�׏����w6�?�;��o����h��T�^|�l6��4��e3�k�MH0/R;��)N�a{"]�J��w�^\,�j��mE�w�71�n���%)7x��$)������M�.��$Bf�`����˾���O��$�3�ᄚ�o�Fn�_g�ߕ=2���|"���x��mj -Ή<C�Rr����\IMI6"C~�G�'V�u�q�-2�=G�e�X���s���������Vh��Qm����d����$�����D�����Er?'I6�g�C�]6Z�_�N�#?:jB>��	�;��+M��Y���Z���8���Y��uYe���G�<�� e>~D}���jdǻ"2CY��p�'+jZ�����*]}J�1b��8��WBHg�Kmz�rfj�b��_1��$���OZ�R�U�0_�mx�g�ޝ�<ǡN�tۛ���f@ 1př���oa(�q����ׄ %��/�;�3�U��y����M{w)�j
�_6��_Y*���ƴ�L�f��>�"� ��<O�F��\�ڨ͙�C�L�/�����gvA^���@���	n_�кa����lZY]ykѲů�l���ZZ%(L�M���K�3f~�V��A�}�uq��^mg�?d��Ƅ}Z�����Y���TO�R��[O��2��+q���I2�p|������W1N�xfs��S�6����f�0�w�6�c�w�퍯H��k�Z����m�?B0 @�r��w����v2C'_K=dfݸhȳ�8%s���s�#���
��� �i$�Α���,_ց*
K=r����vմ�b�b��r�N�P�^��oA���]�KA�(�����cW�Aut�[ݛ�4	�����d��[���ѿ�i\���.�M$�8� ���g�����bd	1��#�D0����U��z�D���oTkb�ӓ�@S`pX�y؝���%W�y��\n�[�+
���o��!�fh�*�k��Gj~h������on�5���ͷψ�G�Q�i�*��r\�l[��W��łn3�&�OZ齨�]����h{l�F��3�R������&�eZ�2f����b��k���I��I2�~�Ǩ���a]��8q�� �x�4]�I�� �^�D�lHF~�W+�h%M��
a8�]���)F�b�",N>����SFs��5q
2�z�g�B���8È۞�a���gY[�b���'��P��zL�:��<��5�O)ҝ��P�L|qim�`"'I��׉�:⬯���^1=o(CB[ЍD�᪁"�� vb����풷�������ǔ7+�R9�×��Úf���`X"�&�9��Ob-�ώ�;Dk��&DʯRQ��5𱘄jŹ���&�{t��= �I��u/o}F��q�1n`q2k�;Mt�b:�W�9w���k�j���!�w�����M���Νd�e��9���G�@)��!/d 2�Ž�a'�=<?#��um�%����z�2����������i\���1��MY��j&�q���Qv�E���� @�@�l��Ѩ�IeC��&���N�[�PMg��Z�" �D���#�s�x��N�%+���ټ�,~�Q�O���M�u�tλf����ooڔ�dX����|�PW�C~? =�9��v������t�� ^:�\�m4j D<���.�R9	Zv!.�����`rFL��t2�Q�8�� k��V+Y7y��_;�tI��?ǁ�Y�D�߽X�"��0L`&&껋ѵ�L#�� 	�dc(��9A�Z;��h�g[f?4VOyJat�+`���؛�u����~<������
slr���:��B\�L:����އ��/����t�E���_أ�9�纥@aU��aD��e���Y.��&�ɷl��Ј͒m�����p�E��[�S�)>�U�63 j��W���&�Ecf���A"�4=���|"�>YK�k)1�e��2��ʺ�&I4�>�pZ8�~���7�e���Z�DT\F�{E٨�]F� �R��ۜ8����K�V�?�A�#����[K�^�
3?t�;Ãp�C�BT� 9(e
�p�S�";
��݊������>ml2ث��6)�9�	��+:�g��c7���)`�Ž�o��H����2l^/��1��ӟ:زC�°3��g���[1b������u��J�� �rI1k��/�\�]�HiY��;�<P{��Q�E���6H�HD����q���?�m�`&��y�{bN���r?֜O9	�?�%au��|=�q�*S�0�*y"d5՚�?R���`[����S[+��M*���J���7�!!p=R���6��q���󨯊�	�ǁ8��E���qIT�D�z���H"M'�C�9�HP���>��ni2��o�t3p�{8f�$vF�珳+ˡ�W�U��d�$�h+��-���{��b��e�������g��Ud��<��k_������3�#�>��[�hA�Ä�3���2>�ue������i�;��b$�
p7���@�t�M쏯{����4�>���MЀK{��t�
��|e4H����xBO}��8��_��2rQb����6C5w�4yC����U0kl,�y�U�c=�^;G��ӕF)f�zB�rA\@T�So�/"�#���a ꭆ���C�@�`�7R�^Y���Nf���n��*��ՠ�e(��"8"Ƚ�T�� T�)��ق ����[]�A� X��P�ʔ�/�I�Y�'Du���o�#7�C���铠+��p���!X�H��� a�ȴ��d ~O뵾Oo� ��>�d�n=g:S��pY��-�����h̞I(Z��E��dp=��f}(��t�m��	��f�򢑵���*�Z�i��Ƿ��g4o�c���z��X��]�t��zd���u.\-O�z=����	;�!b�7�����\83
a�jY6�,;���b'�$�7���_ȼ郝���:������$Ti`���c$�����S!�.���/������P���%��a��iyw;�rO��ϔ������R#hLhDz��{ݥ��t��0�((ɵa�����akG�˵
�j������ꦂ���IW�ҝ���T��Yщ�r�x#���~���ƥ�F엞�1�e��� _1���U??�����4��/�l���z�;���8��%�Tؤ���&�q�Z
�x�A%.%�6��
�1A��{��E�Ʈ�o��N���g��ԧ�L�
6i�������;�pn��i�[J�O^�/o�}@�Oa\8;#Ye��^�����J5\�M��ע"��X�1W�Z"�cz��6ʩ��uɂ�e_�5�E�܈�=�־�])��U��b�W��R�[�0�_���x�a�(��T4��+5g6ɉͮ*f�X{z���v�J>��|̒_!��O����zqG<�-,���@��t�}-is��c�}�5���e��s�7k���-X���%5�����n�YnvV�]�ۣ��N���@�X��2�*R�61�o���V�V��2��f�P{9�f�h"��զ�Y FV����.7U{oW��=��p �	#�t�����
��Nб��4Z�֡�܎��?1���!E`A����:� �{�����)����6����S}�z{�� �"rՕ��!��L��C����y���������q�hR�'j�N�['7�[v�畾�{]2�?����l}jK{���2�@�nQ���3TT끐/@�"�A��������Ά��Y����~��$<J������i�#��U7Ԛץ��}:*m�?�"v�yI<;��<��G�f!�J���Н@|�d���9#^'o"��{�o�Ӈ)�+^ￒ?���4:�4� 7}�W���b�KF��,�=����Ɣi��tٴJ�¦��V	"(���e��45���C�R$�� �ϾX�#:�.�aJw���BC��l�
Z� m_�?�ׁ�"�����f�X&�6��1�$�r	�t�Iި�����V�*�d�viqX|�2��� �0y	�������+`��0��9�_?;$�]�F
�u���&Uw��3`��-P�[)��j]r���J�˕��^�r>G.�qz��6(�P����P!�d��L_[�O�!�[0v�C>u]���6���8?J��P~�OsθL���v��Y<�E�A�f�ӛ�a3�W�a��$_�N�.516Ƹ���:�s	�2[�:K���ۄ$��'��Om�jO~�s���3�K�wL8�A�EzQXC�z��ɿ�a���}/wʃƐ����Ô�8��ݹ�w>�-׶�v��h#�;��]K ���p�2C�G��c���������Ǔ�5���k�R�/�K�7O��h������P���, E��B���m�v0vа�s�䄮3�;iKչ�s��ۦj��<6�[2 ���,
~֙]����es�=��0��̖��k	n�+�-���B{�ݦ>������n�6�����ܸP���

L9�	H�r٩�=�aШu[wi�&n9[ߙې�+a2x��Z8+̏��4:�Ȅd��԰��hҨ���`��r�����Wg��UD�x��E��L��>���e��L��*��X�L�Py�ei�Vg��2�gRBJ�I%��?rٺ*(r�a��5�
� �kq�;	9�gp���r/�Q�tYE@���k �q9�L.��m��������x��V�V�Ə_��F͊�7��_��ME)/��nhU[qInF��Dj���".GlJ��4X��z����Y���]�!����}(�G��k坃YC4t�6��D��);6 1��8�;-|�?�����R��$���i�M|�7��d�9m����의�����	��N��^�&4�p��Ҕ���a�JM
��\���mqv7�5���<=ݍ�RhUq_Ó����&�l�-����&���5�B��oó*(Q��D`����g���!��j���Cկ��"�1�%�Ƽ~ |W��T��1���$ w�H�<k5�0%{!�'�EJ�f��a�=��ׇ�B'ë/ �hZ�ؾ���=��ӗ�ٷN�3�t
p�����?��p;�ȊA��D�j��}ew���
<�d	�����h������\��s����G��T�)i��8�
�m�f�~��^�7�5x	���c���=���X�:p���a�Q�1NJOI�6��ҵ8�3h��	�{����8��rӈ8�2@��f7غO�л�ks�`�����j(|�	�nM�E�7���3�����5�BJc�׬�_(�3�[RG�A����p��*��T�Wϥ��� s_���˱�ÍQ�,��v� �'�X��/�$B�$�ݡ���@�_2���p}���._Z�����Art���|]�[�E^I�j��vvl��e�9�65�c�N�R|5n�hn�(n*�S��F���`3JG�h���2O�MZ���c7��ϗ�����-27�r�\L���X�����E���|�tW���D�L'7mz���%�� G�Ӌ�N��eA��yMap蘿�/�KMm��	��'~'�0��k�c�o�k�������D�����e��l~F��p�ɹ*Itf�H�`�8 ���&�[I�<dK�!��͓`�	�0��	�����e�NR�c��ژ��Y��.�|=uL�t5\L ��TA�L��%V�q�,t6����വ�aA����5?�Gת&٤�C����M�y�Y"��
�o��v�$8m4#�ju���7���D}�c�h!ߦ�EY9AZ��(x��@U�(1&%m��+���=�}�b�3�S��)�eCC�}Y�$����۝���Z�w��*_�[*�:�b�1(s��få�%�ќ"Î�F"O�� Xlt�����a�ȘDX�h�+�lN�?j��#[��V(��Ut��`����"�Fz+� &A��ĺ�K��f����T߁(�N��!6<�dG�C�4k,�C�w}��ZR��e@.�w��49��75�F~�����c¯��U�w�����Q����<e���H���/��|U*y���1��#e"�y��{\#;"A������#�]F:���
|G���{��T�YnsК��8H��������U�<�����]�P��ni�	��� ��#��;�V����f%����L��B���L�_���d-��ߗw�uM�<�89M�&@���B2�+����\4t��EV�j�Q�Њ�F����cc��ֳ�����+�X���kSϓG7�h�G�P��-0z	@^�ε�򊦩C�^xY��X�Ҏߘ�L9���e�*��6r9�j
]�j���#���|e�����1�����?�R- R
��`e�_7ć�9�#��S.��M�n��C�E�H�$�Zl!@�A�T�G�����b��w��j��}o�=�/A��~�Mj=���g�/��q2��8?w�Q:H�;}|(��]R���7�ΔyaW23�$��P0x3��I �����k��M�#Z�ڗyQ�x�۸���D��IaTl&/
����g�e1�pD��EZ�z�2�~�up"&AwW���'�8�r��DrUR�%
�{���5�����g��@%K�J=Z�Lh�K�����;��PJ\�M���= ]SB���ßx���2�p�!?0uQ��7jT&���4�wAOP��Q>l�u�������m="f���3�*���I#-�(
y����y�$���W.4
lM��)��ۿ�$�1�T�"��}�����,ʷ=�kd�W�s���"+'�Ԙ#qEЕ�W̩�AXM2W��=�[��	�R�����v�ެƵ��t���1������)��?��u����x�}8�6b^J7��?�#����d@�H�]�IoY)H[�;�r��11t\�P\�C"�
��@�GԏpB�#���iL[���*���5 ���BY`K����0�GG��T���!��@�?bϢy��Zim���dR��������y��/�6UM�$T�|�sQ��z��z̼�gDU��)���Y�����q�ʡ�f��cq�*yc<Z\Z� ��p�Mm�*]7l�>�w�Z�I��#���a_����g������f���U*�)�Ƨ�?���0����®`�3��� Rϵ�b�65s�6J���7%@�1�����_l�z�yu�=
�h|�:�Ι�v��Ya�ʗ�e���Y���Mm#��R�IyoG5���zˣɬ�&6��2�w����U�bɡ>VP���/]&�ԂN�H5��' �%������y���S���ED�-27�wlVA������D�2;�{��]Q����~�'�I+U�)b�sĞ��
✍��C����t��V�W�P9%���<;5]6aHF�ݡN;M�3��i1��[�P?���B�'�Ig%�n�xiֿݽ����=Լ�ᾕQp[��8�E63�������p� J�7���Up���qU$�{+�P�]�\�
�<
������W���Ade�dK� ������.�1m5 �\�O�wh&DZ��� D�h��RkK�8>�&J�hlF�8�8���c̋�e����'"��$P��Yk�I$ጁUZJ�U��N��^3)����O7�����gD�gƐ{������L ���JB�g���Pp}��N����PkOI�sNx'�i��p�������.:F��F_V�3�+EV��Pg���m��O�¸��प�'	�y��Ud ��ĥmh��7漷�����)���ż�+)�C������;L'��Eb��2�:h��TY
�ƂP�>;"�fD�K�,E�l��l��S��k4�ߔ�D�΃�[��W�K [�w
��_�;�M�2����'��C��)�'|+
:8�?�3��<]��R5ԕ�yPݪ���4U2sl����M���s��w�i��b�����{D���n�[�	H�@A>��5t���D�1fC٘�|�huyNaq	�P�h�͍�;e��L���>t.S����6����;o[db�g0!��-�_)=�n՚���A���� �>�xx`����%O��D�0���iw��7��8i��I��4���}M��p�PAYC�Tq�o�,o��Բt�k	�c��=�P�Ķ�� .v��b���T?؞��~�j"-/& ��hJc�C��p|*G|܋H�};���a�,��M+�C��K9�H���:J;Y=�s��>R��h0��� "e�'��%;\Gp�2-?:H}7�h��=f����J�����;����JB�?T�(	�mڎb|�O�ȓU��.m'��JDu��x�~�2�G�����,eg�@鰄*?��C� 5j�i5<i�k5���9!�"6�9�&��ʳD��'�^<��2�6J���"9'8�ȱ�E)5>Uoǘ"���o&$�ziI�7�y�5�0����6����:��s�l���E�jZk���Q�T�
��i��dF��>�Li?��[ߟ�7��&֥���$M�K�i��Hs6�Sc�y�����N��r��6��9���bgj���X%�+^sL����=[4����Ղ���f؊9A%�cK$zۆ)q��ci�2�S�]6A�52�X���5e��j���}8�e���B����M�U�YǛ��!
(45�߿P4(�QU�����)�Hc(��AĿɴ\]�Aa�P�,-!<��Ԡ;�V��� �r,��*�XX��"���x�~�� ���޻V2�s��
6ґ�������.֗��6J��5�u�U�<PZ��A$ ���-�F������G60Juc�vY
��`a��M����:u��,�l�o�&���D��_��W��՗�j�������;�H��B�isr���h`+�>��:*%�$X���:"PE�ۼ�2ɰ���~����#/zc�/w(�Ho����LӖ3܇�XԠ؟�7}�-�/�?1sJc`���PP`���[�ǔ󤻦�^J��>%���Ǝ:��e��Vex(�?S]���OA�H�I<�X���Z&�7�D�oTn#�����K9�L�t��?V��G�Tk�I#�:��*.¤X^���"z��7������x��e6~���_=���0&�1�P5%�����!�Ak�/@���M3����f�پS�Q�~����{�8\iX,2&=�%���L��������pX��rn4p.�Y�:C��8���	�Pe�<OI9�Y*tH0�Ⱦ?3Mkm�[e����Ӆ�|����y���':������*�pu/�\� A3�f�ɩX-w#&d�{�� "���r��`��/�Ѫ��ȴVL�4��lZJaJ�W!h�|*�����$Q�Mx���#�����;����Z���1��<^O?��5;3;WQL�8a�<`�0ZD���]�.Π d�
�l)���6|2R����!���3��o#�[i�h�����z'�Ƽ{2�c��M ���B�̝�v_�7�"_�Ov��F�B�t>JQ��m��:�}�#z����)Q7@�uj�!�k0�a���mW��E��`�o�<nǬ
:�z�ۿ�ubݖ-�l�GdA��"Ȳ2n�%��`ą���6-O��k@7^g�%�Wᣪ�H`��?m�eCǃ� �) 6�0�:�p�6�8M�H�����l��&�ºnJhu.Ynm〳B�g�mpݒ4�`p�W �d��G��?rZ���?�Z�!��_�����y�.t�Z�Y/�j���8�f��O?������wP"�z�(�y�f���<�13^	B


Pj�odJ��Չ�
J�"v:�&t%
�B:�5e�v'ｨUB�ʸ�e�؁P�h��ť!�"9!?;$�Ȣp��]��?�fӻ�3�1�ҷ���B�dn~Y�n�s�WG:�hNVP���]��Y�U��]'�a�3�A��*��lŵ��=u��/�s�;�r�����	3�0HP�Ӧ@ d�8��;�x��7�m�XQ^���x�QRǛ�gE�b�~�ջ�d�s:5s����L8��8��[�
��P�5L������vTL����/�ذ?��{yU�}�ԸT\w�\-:�@cX,$t�����t�X����b���uY1��"�,�tw��8n��)��f�>�ރ���oM6O��s'7�!N�5��,�1�.� @�������s3a�{��K+��[y4���ZZ+��ǵ8�P�x�vڿ�tx��i���$�OHӈ=R��c!`�K�,g�S	���DaM��0���&��s�n�������8�3��y���qq%�Q�8=R�������Y�/�"!�%i��p����O[^}���P�@m|,�=+��o�3��9�� ��=
.MRN8.!͌����oAtؑၐ�N����Ё�E_;1�Dwr�V����(]�fI~�9�Kv�Toi���ЋZ��7)�%����y0� (���iE��{e�yE|&�LN���A|�'.f�a�,KH�C�أ�nZ�)�����QN�F���D��Q�����y����l�@�'���흶�|wSX�o�刊�Γ��
]�ⷂQ��֮~�d�Mڒ����Ò4����S�O��]i����7nϗ��������P��輍U��i?iSn�LV�QS��s/�U}�\Wl|����3���CV{N���(�(�����44�Nݮ��I3��G��e�.Z /���L6����$�v%����Hʇ?�m5�9g�=�
P)�p/+!B�d��l�*j���[Z�� ���V5.��-M%�-2C%4��t�Ow�7�"�C�e&���*�᝟
i��j�||����H��	��EM&`�0�ޠbϻv�����?��ϸ����j�U���.f�[�\��D��<�qy���+�	�=��I����&�i���8�^�I4�5ˆ�\�݃���a��U�˼��P�=C�T=��*n��qM/c��Ig։lE.��3��"��������[+l�i�Q�QQ�?�7���~�3��"ɘۣ �M�fHǢfEwյ�$+�h�w�'pB��Ұ{4����瞨������3pB�-뮌q��Q?���fa�ga��k�h;�IE��l�g��S~V���� ��ĞCmO!�f"�R�	�n����a�٪��,y�0v�l���
�q8���Cj��ә��f�h�RF�I�� ��i.�V�����/R�n�l L�i1	�H���9��B?��z������w>h)o���ۍ>�)��ʇT x��0�u�����^q�1������Zf�@Z��C��R�a-U֦�҈)�Z��V��'�#=z;���}���x4M�U
63(�~��+ <,�t����N��i�v)<��_j؇���?���&-�����ƃG��lG���I}{$/���!�]�;	8�<ܠ�]3~=�(M��{[���F�/���U[�j�Y�
���=C��x��}��T���~�P������$�L@v5 Z/�FPl�?L,U/�z���K�Q{%�]�C�Z@R�{�?�iZ����`�$zn$r��k��&wv�j5���oŝ�h�Ⱨ�zG���ܠbc��X����f�V�f��ױ��������f�Q��ɥvl+xW�iT;y!]jp�\�P�Q�	q+F�y���V?��Z����\ @�M�6]�(X��d�jpeZ�c�������8��^k�1�������S��ܛ��$`��B@���y
_�F�ȋ���f ܵۚ�*�vt�R$R��5�b�N@&��C�e���K�@��Qb����O1��|�cT�y}<�/+D\ґ(+�aw_ �B'��Q)k��wW�?��7
^
���f�n��)��P��.Xp[���� �%ԝ�{'����D46�b����i�o	�d��9��4����.u��h2'�cV�5
��UY���8�Z�>Q��yӽ�z�y����CiK<�mJBF��lrL��p�-�"�Tb�,��F�m0`�6��uɝ]��c�H�"�Ȭ�1���	�8����C���Z@<f�X���!�P�9��ZE=����5��K�1�[�k�����6����{^�݅7�V��}r<��=y�wx���VH�KB�j� uxӊ-�*��"q��N�ߕ
{i��cF#�1:���Wr%e���{�Ds��R��W��L�� �������on~���� �`qߎ�� �b��9�"�c���n�+Cy�L��oE����W�YVg_�*��=ޖ^��+�|󣢋x����($k'{�����H�0����.)zkFw���w��V5��b����?��.��c��Bk�.�^�xCf	�$X��y����6]�\fy�|�i��8����B#�.�G�,{q��]����ܦ������oȕrK؂X�+.�2�D���GyPTX�k��YIJ����.�g�+-�4��+�R��h$���ni'N�YJ��4�G�����oqVL[�=&䇰l�.��X``k��Fv�7��n�QQc ŕH?����|L�I�dbm8���z�}zn�Ǎr���CPn��4�7|��Wm�Y07
s-�K�>�_�+XnՀ������o�t�UG�dhW�ۺ�&�Y�d�W��!��p*gmx'�A�!�7� T���kboD�	��4���NA��i��&\�~����.+�/�j�
�,AD�Y�ͽ�Y�a��1� q�S���� �N�5�q�	!�����TC�G��a�������%UMe�BnP;�;`�d��-�Ų�bdSQ�zl�H���}�f�ɥ��8[nF�B)���h/�;H~�[��J` &� +O��ʔ�?KܺaP���j��5�0���=ҍvx��JH*�tM���5����?Ȟ�j��JQ�X'���1�s�E���Ї��[Tx���s'��bO��Kf@�j:���M+�����aa8Ӿ����_gD���f��mmޚs��w��g���K�ù-��PŻ�/���YF���hʛ�l�:�?E���n�>�4�T�O���H�d�C���Vp�:�4V2��/ԙ�k�������GB�F��_2�:b��9'�v�x���fE������}t��vĢ��������t~�?څ�p����r;�֗Ke�����e{2�W;�؞�݊� �֕���q���գxx�P�䈀���E���{��C���b�K�:�U���&$��T���|y��c��T���|���a�j;����%�͐���啅���*5WZh�;��[mRa�IW����{ќ(]}������կl�c��[�ָ�y<?!�H� J��Mo�˴�-<�#�lמ�;�I<��GvB�n�7h�����trAoFy�ZH/ }��@h�l�]�A����	}�!�{  ^~,�3��U�k�C��6*p�5��}L�UP�%��F���W����u_>D{L_�����h��v{������������~��/�FR�,�T����a[�*��@��C�Y�h]��	�یM*?���f�^ę�=�K����w��_�us������O�R�6��-X��]	���g%TK�̩�Q����(Җ��O:zvM0����)���]t�if�W���$�8p7F�.;H���3�P'[|/�+л�Q���Qj��z��rfC=�W��-�[��"�(��.��:.��֣M1�"@c��9;
r�b������n���M�ʑV%��pl^_)pL)�P�bpA�G��݌a%������e٠jA�k�n�#�bzA��(���/#�����B�2)�e݊��A 蔗�nd�l.]��*XE�?�_ش'T�^����Uɢ�V�!�G�"�N�ozQ.o�&���[��Fp\7X�0��@⚳�'L����t����x��t,���z|0�w��6(��v���3m�"��z���#���W���6�i��>E�ZW�5wq&�rE���e��yDW�GH�(N���I� ����i;�%�����e���?�4��$�kYq���gE�,Un8�ږ�U*? �ߩbD>
�Q �ţ>u��T�����i�bV\Z�ې���C=���r�_Ɍ�݄<U:�	�Z"��}2SfarM�l�Imܪ߽�|�_��u+o�Qȼ��pS]�K�S�zB��	��Z���٨���e����-0a�@r ���F-��_bDKlu�k�t���������l����#��G�B}l�p �ɷ�]���1�؅������Q2o�-�\"��j���d- ���RMՌDz��@��K��Lm����|�ӓ6������H��a��p�k�0�`;�������7��4�v�����1��M[�#ѤV��MB}��[�uY5'�����ծ�{�"�/o4��`�d1�g�����n-@K֤\�䲗�Ì��f�Ѻ퀡=�p+;z Hs���-х��{/l���>�a�yo���H$S'�ϟIt���/11�����辑�
��	>�	��bݳ���H�������WgB�JD}�䪦h$�����}��[�.fH�M,�ܲ(��^�E7�k^�.��Sm����G}o����m�����(Y�~��bY¯�Gnfn���Pe�g����� ��U-��jg_�8�O�`6��l	B	�F9��@,� �H�w�]X��QxĠuNL!bN�S6-�S�h��O�yRl�i֣�6ڰ���R��?�g��I*$��{N�s?��bߖ�3a�mJ+����B�+Ox(F�O3��ilϵ��I����Ie����^�c��"�l
��ݷ�^nj")jź�.�.��%�mϥʡ�j���\نqD�ؿ�Zͭ�?$��4�0�8$n��'��p�r:4�We��|.C�`.�7��=��t]�O	��JHU�ꮥ�4h�4�]��{ P�
�+��2����x.TbӱQW���U�h�Q��@%X�+H�]�`Cl��.Z?㣑������s�(:�ϙ�;rٟr׋�?s�w�����qP���Y�����~N��wK��wW*|���/L��30�?��*��LL�@��½��|usT̾^��+���\����|��>ĺ�R����K1��c#�t��
��9p��}5���J��*l�=+���hM��3��7!�)��iuI�"]��/l�f"�z����i��+��8,3������hV�Y��f�%KpG ��*�:���!^��wE.,��e�i?��N�j�E҃n�h�����G�q_;<��s�!�S�VG�=ѵ[@|�#�Q�p�)���A�g�W(�j��<�f�p�0]E���G�sA'���QM�_��v���xU�l��,�$<��%-�z��*횴8L���}vdZS�r�X�*AX���w��aL�e�.��ߴ��}.J��p����M^�Ә�j=�!��l�j�(u:�~n)�<�T�#"�xq�$0��} s�AΊ�>�}�>( ���5�]�2 Kǉ'�z��.����A�1�/"D�4/��Mܑ@<T=��;a�l��L���1�̴�x�&v�B�'Z��kw� �`����I��M���_T�ODk"v���ّ��9�7��}�`��P��O	�W�%���kG����9���LD͉C�Ü��7|PBc��Gh��E!F;�lIf����5��V�k���Δn���F+�������鯃	TG�����; �<cW�H�l�囵��JAk'�(vp�!Q�?D>��W�kG;;	w)l*{"O�f���>@�ˎJҝ��B���2�3N8�w�
��D��&F�S������R�>X:����,�ˢ�|�k8�����w�i^Y��7�w��fyM��0.�:j-"��?}��nz��
e��1��ZI2p�����M%�1IBL����Y����Ǐ�a\��dP�!����0+���$�D��'`>U���C2t=�7��߮|��C, � {m�5$����=�q>�vS��K��`�d<�x��U�������G�+�8��sϫ���o?�y��z7H�-|>����Ш�����$0bw㲅�x8��-�M�
$*���^��۬T��i�	F��Y53+�T)�j������1�$a� ��v���I+�"�C�z����d����TH�Ub���m�D��$a�k2�)al�}nv�h��>��šˍ����)`�e��d��}�G�]�]�G��(3�0��T�z:�����u�}�L1}�AG�<Pt �[|���
�ׯ�yx- xT���f�{ȫ�)4e��:+��������5ZhA�[�&�>��G}>�q�Tg	�sPt��-���^�9�����ԏ����M��_rCUWe��[̋Ӗ����u����+�@��N�s�J�<DY�_f��f��6#�]�m�?��~9��:�׳���"��_޸M�듔����,;�M���i�-2��I�ۢ�á�9!������|�c<�$���{�����C�mB�6��6��C(w([�Q	���ɋ�7�1,)���x��S��x�?ĕ+��H�O;��w������_��R�<�q>y�s��ϦB����Ԡ'}�t����A�M��c�ٽ��l��2�/*�N��1�@+���4}�0y��q�,��@Y�{���3x��� ����bȎ��]3�O�/z#(2����+S�H0b<�|@Pq$7�S'|Wh�D���m��>�7���1<�M2��y؄
1�Ү7��"�l�ѥ�U�")��=�wa]����	ˊ���ʀf�
���8-����hD����S7���0ͤcގ-� n�8"5Q�ϿY��n�1IZ2����.�Q,e��
1fmp��A�ᶧ	f&7H%Bz(���C]���(߭�Hi(�eHbC2;D��K'���W,�PM��Fv7�hZ���.wp��`��YmxES|j���$H�t��'��_b�@J�DP�w(�X{i�0Qjh#�� �_W0	��Q?d�<���ơ'[K�{�*%��q�ff֣�
�~�^� ֮)�U�u�M�����t��+�#Bu�<oU�:�(Ɯ�g���e�]{QH��`^ɱ�d�JL����1�B�h�$ j����kf��B�hl��B>��{�P@Q�2�[ۛ�p
���V�O玐��^4�ɢ�����.U��G��qmd�X"�nBZ*W��>�T�Rd$q]Mϒ��]�k�]Ĭ�Ј�c��b�]�H����A9�r���w��+_`-l��$F�A��z[��`����2�VB�bt���."�HZ�7��!q��Y#���Cf�{2
V���Cb����5E�@���(!��A���k=u�$�|��z��w��8�T��X"�z�3�LW�
j�yF��Qq��WTVk��$�/�VNַ1�FQ�`�V�?��	@1�HH,�z'(Ca�W��	O\�� B�]b�Y8H��j���z)o�-��g���p~�Np���Ǵ���-��}��kN[�|W8����q���������#��*Vut<�qdYUk'C��e=N����c��4w����e\��L���g��%t6 ��N�!���j�i�]�Eȋ%�W��b�e�V�ěp)�B>?�<��C���H%΁��H�}�W�u�3~����wlА[G�A1����q�ȅ�Qr�i��B#��.*���u��u����aV1�j�-�HWc��oeʧT��Y7	���N%��>~Vu�\Wo�g�̆�j����"��
D�D�S�x�0��
���ŭ%�`��wj;���$���;\�< �E�)k-�'�s��秱�
�G嘪����U0���#��ۃ�Mc���+�0{]{��r�oP���_��Y�<��������<E��S����?e��n�)B}4j��u)M��J�P�eq�a��!�ɀ��QF�
!}ovŗj~TDS�/^�F��Ԗ�^�16!����h'�A��>�)�l+�.��.��h�+ӶU�e�O�<H�7��,N����1�p�@a�����_Z�����/2�uoV��F��>�p�yy�h�-�R��^s�F�|�|>��;�������]5�c4��5���V2�f` �ۥ��y~���kE��݁���}�Ye��_��Q,l���r��ym��ęM2~z���S��?�*��ĉ5����(8���oA?��?���3��;�B���U<DgEdI׭�p!p�W�u���bN����P���t>�����cm�A���g������&��L��0�ѶA0��xu$N��_غ'PO��"}��)r��|a��Pt~l`B�ĭ&�ҧ�tw��	PR/5�O������>�=Q�qf��㝶):�k8H��x�I���s�YJ"�R�L���,ޭ˛0O���	ien'a}r�e�s��$���(j�_�"���ً,�&qGP��..Yuq*�K%�$:'\��I2=4����堰��JP�d�|^�L2�'X����$r�Y�a�EC�g�i��p~統��׮�=�tK��c�4<�z�C��C�i��O}W�l������ ���k7��I��`��h��%���U'��4#�£~-���G
{*���I�aր�/Y�ǌ͉v�/�u�q�L��9�ߛ��t�̬�ّ�);���!\��Q�!y9Ц����/ϓ���+���.:PpE�;�po�,�p�-��DR��ƕ#fՙ��ƈ�J�Ʒ���V��_����B1?�'վ�$�wj� pOՂ������!F�sJ}r�*��(�[p����^��'��݊S>͗���6o[�& \B�O+�9��ɉU_����#���M��>�0�q��
,�5�a��YuI��/v��E��^dgG z���֤"��e��u��q\�)�Zs6�z��2����5g���`RoY5��<W`k�ڢ_��b��;�%^w�� �*��E;1}S���)��f�Z�U)!��~#���Ѳm���~�v/�oG|.��a��]�>�b����KW��fa��{E�WʞpC�����T�;�Ksŏ9,i��Rfh����o���4����x��n���#��_���?�6�1V���XYeƑ��H�y5USoܑ���i�\660^����yI��R8<����}�a�k�'�H_830)Ȇ>���F�?˹^6���Zd��jG���Iޥ%���=�g�hj{?�`o���M��ڧ}����_P��S�OF9�g<����G�*���M'�i]���m�8���V��Џ��~c)��-L@_j�]a�fS��T���C��}����d*.�M�2���ݍ�/�/