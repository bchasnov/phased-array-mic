��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\����q�?��e�I8�b�Ǽ$��"����ׯ1�V0���9��";/sE��ƛj����Q+f�
_U7y�5�YJi�]|L+�ۀ�N�3��Y61/Md4���w|"2�)�3��>u.�s����5L9�a4t)8סw/D{�
�a�]�+-d�hD9��B.#T|T{��Zؓ��@q�k�H6ԅ�.U�h�ɜ9��,���C��~G%��뒽�8b�v��Z�.��6��p�~F_Gz~�'[�E�T�R K�P���!��2VkM����.[���몊?�PD�>*O��񓢭&�H_��6��4��<=+�|p��������h����Ԅ�ų�Q��������rf�*��}�q �_�nUP����yA�=K�-�S�o
��vP��5�-��vEq��'{�2�N\�0,��=���>�z�9ٶ((��ٻ�@��T�s�8����F��զ��8�W���-49wh�����8�ʹ\P�<��o�Q��J�ЛR>�R��^���p���j*J�0`v�\�09�ʴ=�as��-tx��IFr�j�Kb�@�_uv����,ai�D��;>��)�m���/.b38�x"k^���"����TL֐$���<D��M����^�K����v�0G$��xGE��S��&+\V���{�4N"��SYK�*] �y�~
�Xz{k��`�̂�͛IRɹ�=�=
R�^<8�jЮ�Q�E�"���T��2ϛ�����G�ٶ���X��$�c��
�ck����L�l�G�(�~�����>�N�bH�'�0���.\i����מJ���bS����
}5�6H4m��c�lM>@K�ǈ���4Mt�k�akhRt:3�Ac/�\n4�I��?C^��{������lL|ә7u������!�?�cg ��%�������}�_�H�r#Y�r�1m�܉5�B�#8��K��$�WI*C�R4�yGɫ��[L�
��z%�B�
4~�<�����=+�%�:�l�����-6N�e���6�]�L��U�jZ���+*��h����Z)��@$�@�({x�f�W�FtA�l2?�O�ye����-Hy�%˸���1h�'��zx"��
q<6���s����njYn-���X���gk��?P������
3�.%#�d�`W"GGX�����t6U������F� EZU�v�(��XF�n��4���P�W�u��b<�Ѻ;ً�8�CV=�}�{"�Wh�q���ۙ���ճ^`|9Qe%	2oo��dzu�@Q-c�f/�����[�l7��*1��e���X;b�,k�D]D���~f�
LLAVH{�7���988�)���b�ȣm}V�]����h�kϥ$��l����zb����>��A0hHDr�Luz��¯G�g�)6ԗ`g�0ց�F�Uz5bz�����y�0�)k�w�^�#<��n�	�����~��#�:��$�1"j��� T|ŵ{{�S�Wg3���/�r
R�q�J��r��1����႓� ��p�N5SD�`���f��'�B� �Z� >%��.p���/̢��$�]d&)�+�����Qu�j���sb礽vH�Ak_]�tH��'Y(�f��<�A��>���\K��L��JQ+7�ዜ�͑}G[>�sy�&��Q��h#Düǅ�:�5��B�F�s���xF
+Q,�����4�c>�}
�<�4"{*!��C.�`�(�t�@WM>h�d�?����p�r1�'^_XkB*�s����+k����Ěo�%c7I�����anR�/yNS2�&_8.����j�
�Մ�Ê���O��k��.��9<�<!��v������>��<C��r�7���
h� b��횞�����5��l�
O�����OK_��%b��IA �O���;b�GK�V]����I~I���D��d�L��I�P��T��*�1�/x+����9j-)�!ib�\n��{�do��lp��"��O�_�|�\��t�<�)ַf�'{�3_�F}�@�Ꙋ
���	�I����6l��&>f���|C䔺�q��d[�sߦ�ӆ߱P��X.���ě;� ��m�zMW�e&�kwI⺔(��*kW߿��\��%8�_�I�y�ܝ6��S�}���_h��0����DW<̫'��Qw����S�ӄ��7�op;����_G�zm��<�F��p�^���9#I�(C,,���e����q�a�QqN�a��Dޫ|6}ћw�	є��j��v��ix��{��A2�_���/�O���g�ܜ�X' _�S���
�w�3طh;H%��*v��v�\��:���4Z�o��4���y؞A��*Ŭ'�`>.j��(� �@���۠��j��,�z��w��m�Sm��G�lU�_W�450�]; T��W�@t2NXw�{�c����L98HCp�m/0 VV�O�o�k%� ��V��7��8��+��E*[L����{&� �m�P-�=�6wo2�V��u��=!���T
|6�;���D$G�42����'fq$��|#�Y��ۆ)���t<wO8z��Tb'hf���GgὺL�p�J��L����|	<:@X�3��0tV�1U�!�&>�s&d�od��?��腰v�ߊ�^籀��uHG�>���6L�����|��
ی��1o�<��'v�g�rCN������<���ƃ�P@�%-��]���9o��<B��`z���E�4P��#�AO��#��	���l�
��;�D�v�Fe��W���� x;Z8�����h����M�m��?��9T�'U}>q��T���P#�niW������*L["�X����NƔ!�:)���8%��2B o��(��#yz;���/$fOX3P9u�����u�0[^$��C!����:���.��yz��6�O��0���X�Q�P�	.7�Z5�q釨��ɪ�]��S�LP���ȣS�bl 	6@|;^��c�U�wՍ�O��p��.�3�/i�$��a��"w\� ��ET�К��w9z���
)=*Z�C8�z�����"y�;#���v95'$L�����Fяo��>F@���x�P��0���.2��j�r}*}@��d�����ɫ*�(.:�),ݕ5b��4֗��\��nk5���s�>^cq�76�"���ka!���m�0�/E�Mk�q`��������Š�צ���y��4�a��c=4��+t/�p��`xǏ$G�q����z��r����)7U|uHn�ybn���X��(��=����s����T�	a�|��!��<3���E4CV|���J����Jb��*�Ɋl��AF�Z;�CNa�W�~����Sm�cXc6����f�@�=P�ǢEE���`w�o:J�=Q�e�����'9�3�"�V�7�����p�b�3k�*�[}T9)4�� 3�g>���u�h���&^F��ҽW���ѯ>����W�|a�0F����M�*P9� KX�f"��P�,6���[�5mX
ѷ���hp�_��E�>�(X�������A��G�o��2��
�����5wm`�|��c'IS�Dϔ@s��R'�%N��Ɓ��������:1���B��wa�-� "E��23�o�[�qH�1H)�d�������$��<���V��\�����1ŕhJ�W2]�/V)eڣ�k��O�q�u���fMZ"ft+��y�h�8M�hҳ��>�6��к��b�#@p^��H:�J�i�5��R08�т�-�-�������[KR���x"�y�5N��,&��[9m� �=�f���L����I�)p�� ����0�U��p�?JG3�չ�E�����X���B 4a�g�3l4`e�/��Q�������ϋ�|���o0$-"�����m�k9	������O7�j��CN��yAK���F��V��{�S	���hlÁ��S_������9f�钌�g��8"�����*?���xR[�{C����  н[YJ'��=VAetE�ޅ�d(�$��+<&�q���c�@T9:�m5�`��͂��ɁZ>	�/Df��2�>c�|}�%I�rGl)� .�������v SV��RI��ǥ��?P�NռT�H��I���z����.3�{턩�R�)�V��J���1�1�A���s�-D�l������5Ұ��U��0���:@%�04���}�UD�l�j�k��&�-E�����8�^�l��$����F��!'�v�"�Rh�ⵧc���k��]��6V��r㎼W7w���](+�ڈQ���?�pp��A�������g�i���u�8zgy�<;xt&�z���f�6e,���+�J�t��>��E�yY
g�̫��р�s�j��YE��&���@zdʞ�N�Kn���	/��$�w��PW����\91��HjS�^>jLk~�h��FH�#��� �>��g}�������v�LQ��s�E�4�GÈ��}�u����rq�վ��HlQ���Կ�M�'�����	���6����b�!���
N�l.c����g�4o=~�� Ɍ"T ��Ó��\��4�����%y�`+ ����]C~'��Ԭ��W�ɺl��Z�9%W���W	�F9�uÝW��<���3���-����9*yLy�f�L�p+dɍ�d(��THXv7pΑ�� ��I����v��I8A�\Fך�A��xD�@۽���$9@ >��·@�����y��)����owAŨmϢ�c�	�w�����NI�:u �gcA�%����Y����[(Y�s��b���糋o�+i7��E�^l��>�<k��˗>��a`�h��2���?�=kb��b�� �����N�	��f^m���w}`"VAIJܝ�1�q�p���vw�,q_�=���YIV�,�1ٽp�����<�����A���� g����́�g�׹b�5�H���@X�=�Hؒ�a���� �"���-�܊32�|ݾ�ԗ�O�e�ت/�Xl>���6,�"���I@���
�~\b� �N�E^�h]�������Ƙj��*_j�v�N�7��4� �~����B�����N.-n�*���W�";��Q�>"�b��t�$mCh��3ك�aaG��;F�z������\�A��A�F��;�YԮ���߫�T���>�%%���:ky��8�PD-DM��j�M#\1��l����=������/f~$r��WGG�aBʉQ��"��g��L�O+ޥte��vm��.;׾*`��Rţ���G���!u�D��ޒN
��pA�aT����1��	�"rC�D �V������O����i��+�ֹTB�k�V��!�kd��a�xN�9�<�n2�Y���8ƀ����Hְ��9�P�[Z�7v��;���Wx��熴,�:J�b|{�]���=����*��Z�?�W�k��e������N�Zj�b#v8J�*Eʀݦj�OT�i�[`� w���	/Q�:��ᚎP�M/pKN-Z���9k�D��C�A��9]k��@�r\�!7P���wݎyA��9�46���Bgţw��!2h$}-����΄�Zn�i�<Cp8���4��g���I>!��!-+��i��ڍ;ɖ�֕]���F8� ��@���E�F�������N�l#[B�#�E~�-0���9Q ����+�����W�bq�,����?�Ϡ��tm�����.��C���{�7ɭ�/��t�Z���pe�6~-��u^v�g�i�ΰ����A�CA�r9ߔM�Ϡ��4d�C�q�z*FF}F^���{wf��n: � &_��l��q�Ώ�5 Ԫ�8���SV������
�5��6��]���e�>�L����ߨ��¼h\=<����Yl��5�!��e#����Ҏ�`z�xutџ�gMiO�$�蹍��^?�HV�����/����2?�̪8���f6�À�b�Ni&�iщ��/*�[�w��![�
����u��|i5�W�u_�j���Ņ���O���R�.*��>{�G�_D��У{o��0�@��$/�8�U�������9��U�(p�_[k�ڪ1��,�E,�=&���̞B�;��=�L���4Oa#�l�=G!2�{��?,��4��Jy�������g���	�Q�Y�{1��0����;
��}����V	ޒ�Ф�.@�������#��w��쑴.xk��([c�k٭Eo�C�eV�.މ�w��<?��Fh�����|%�t��ֺO����".�W3���&��)��W���>�M/:Q�W@��t݌����C�c�B�A)��%�?�Q���%9�GCUK����kh��`�>�b�P������1֥�h--�k�c�%ay��G��~�3�6tx�u���@�n�N�wL�/���G��H ��D��@�	F��X�"߅h�BRx�i"$�F�l5w$��H62�r���Ÿ�K{X�dՁ�I�g,>�|��=d(=��
�C
�ͯ>�Q;���,��F���� F�h;���B}�.�.���%5��i���T\Tj��%��y(jЪ��Tb��k�c�`�*����w�!��.�A4�z!J��.G����������3}6h��� ��ܞ-H1�!��{#���7:�,t9n
`�g/���/�ÄT=o<h8��2�v {��� ��U�S��