��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��/��Q�w���a5P��B�~�/�'̙���S{���^�qѝz��'�hřD~dVr�F�!5�=��[�\�bYzy��d�(5���*������j M����J����Cw&�u����Dg��>_�,��o��3�9=]�sn��5���A<�-��Y�,���AU�G���̻N�	�Ϩ�g�ϵ�w�Ω�k���R�9HO�o�u�(v�W�T�yVL �q^�Q�0/�����)1�cڵ�E
�W�D�t/�Ș���~x��R�X7�]0|��?ͭ�m׭��e��%\rN���H�i��8A(_�P��0];�ű
�0X�����&�Մ�"<I�L`���`�����:�������>�g)%�N���g%ȟ�p�tQ��[���@��f�+�p�!�]}R���Zy �V��(|�E��ӎ3�zx��|�^��ws�E�.ao��~P��i���0���J�4��:��������#0��9"6�ѵt��L��80`�ڡH� }�l�p�2�<�|J��Y����e ���B��!NB�,�P�!�o�n�;�*D�J�@y��!A�-
8�oUEU���(<r��1l'b�=F^~�~3������#�8��f}�!B'g��C'^����W��V��u��𪢕�/(|��������R�P�q���t��y�1��>U��x,�*|��U�x��@��K�c���i����Q������m������9��޵�f�<�AC����e|�$��+�z�%nD�m��$S�h!|��e^�~����2P!l_��Vܷ�n��.>w^�eﵼ`�k�����Q��4<^m�4��@����~ͽIZ�{l��(��%4��d3ژ]����7%�;��	�8�G3=LC�-S�p���k˟0��U�T��F����8B��������K@�4���U��/���� �����nL�]X�wY��U�Ȥ_�߾j�:,�ݲ�6��}췗 #{&�V���$�,���R�$�L8N׻�	��v���ctLf�'*"���>g+�l��{�q4;=;������p	��<����
:a��	Ԇ#�#�\�:���z��QK��a��Ӵ�OU�b��xpH��#�y�oZ��#z}�R��Rq$z�xeRf�Y�|��Z9Aĥ�0֝>X��:�! �O�����,B,!��u�wgc�㯎H��V?-a�u����6��/3ŧY����z1P���VN����ԝT@�g�p&��c�iF�Q�+v���^n��?&	
�h��ѣ��FoZ�	�`��n�v!��>�y�G���\F!����d�ݻO�@��I	=�������E�L��&y�]���Z�y����Ŵ��M^�{E��a��д��45��R@�.2�[��+�Wun���N�=��ANh=Q�%֟���=[kك{ǵx�'�P��Z5����J�y,���HE��z�\ؼ���FX�{z�2�m����KE���4.��M�;�f�ސ��*�&3�U#���۝�ΫƦ�8E)Xw��$���G �`��qՓiF�9��r}�[��[x8�B����}�D��J��F�_a�h�{=.��-A��˧�JK�NO��8�[�����kd��u=������t6Xg��̞�&����P�d�t�J �����ȧ�p˔�to����vw�����9Z��V�?[��H��7��%�B��U/Lǁ�-pP��,J�������oJ�!��TLS@�Q� ��V�dg��}�ҡ%*�G6�)*
�w�?	��� ��)�[f�h�f���WD1���GH����U� �&��f 7���P<ڀ��~{i��]��|��Q�����`�E��ʒ�	fWα��Lg^e^H�+��}g�hy��G��Y�.�Ґ�&$�D(��tw���hIӼ*4�2��r��G�j��1Q0�9Ē��X<�	����1s6���	q�W�{����Zj��c�o�,�9�g,��� ���q褕
7]��Z���	Cy9�J����'5ŷ|ˬ��2c���Y��E"� S$�H�c�q.��}���Գ��SW.�5�e��s�vF��I�#5�j+�׼,�2��o��t�#��"��n�)E��Ƶ>]G]~,�a�P�p7�E4}0�j�[1�Q��T�;ٰ���o�3E���Ǩ���	(R�3)�4�~��~�@;
?v� r9"�*G�n/*z���
�$��#6g"F-�,�Z-H/��D�M��㋞�k̬R:�M��;��ak�v����g�r1j%���T���u׶�h+��i3�*��
G[������Q��g2��-��~�_'���2W�?z.�<���������D�U��Q٧� oJ�*	�aTO���l���ЋE���8�_qlgԦ�뽛+@�2l��F�џ\WvS�����qo�m*!��������Q9��f�c���7qF�	�,M��*}p\!�dlɣ�� \����R�:e��q}��V0n��!��7�/����X@t�O+���Xa��?I�����݉�`�z���pg�3%f�2˵��C��$;�/���?��2I�Pނ%�d��h�֋ʊ)�h�HI��({V9�6Eevs��{Wu*Z��;@p����S�~g��O�i�N�;���dJ�
�3@���@��AP����D��|�,��w� &��QZ:D��p�P \;���YO�x�K#�`4��3D�+��@��P�Clp�{���p4X����WM�K3�+h�-@3�:@?�;ke�a�&��;��Y��p#�PG��ĚC ��c=bC��v�Y*�l�+b>�t��?	xGP@ӊM$S�Ja�=Z\�R�� L�U0iMv}^5�yR���c.��H>AB������$l��:X��h{ 2N���l>`d-�$�/��	�{Zu)�;x�I,�X �����D�/D���h�Y3m�z)�uG��V8fc:vО�>���!dp�����O�r����Au��7"u�<O��DƔ���v��5v�`��F���g��g�e����S%���Wa�y��fFg�B�� �ݼ�N�����`��@�R�2�~��Rf�sy����k��������|��b��@mF���*B=^����ϱ������)!0�ovy�HtB\�C5�̯�7[λ��@=������#4
W�BL�!ƛ��4���|�E�*F�ҁ"�{���9�(��ce�݁Q7�s�4\yβ*��0�~Ն˕����sn���PP�,e,elY9��0��	;�^`3M"{�pNh2d�o�&Y縏��E����=����z	�ظ3���e������.Z��t���D`gE��X�>e�F@��I����A�`�Dv�ʲxw5����s�X�;����(�{)� 0]�U�B�,�G�u�>$gلH0��*���fc��*�<�T��(W5��v����y(7,R�ZޭKѨ���H��N)�@\�0E7��h������\X$��0�Z}>0�x�Sx�����=�Fw��طAm��vY���	��`ĩ�����Z/�C��!S�8+������)��xF�Շj\}>���Ň~�3��L�-Ҟ)F�ݗ�����J�b�Ǧ�%�zٻɤ�9P�_�|�ipc��x֪J���#�:)�\�c
pe%��tƱ�^W�=�A��P*�?���
}mqA7��k2�8Oe}�}�.8�0�Z;p&����b�+�!�ETW��ݹB]����p�������I:��N�����C�ij�+�{u��X��^w����������o���m���q��HTꅷ�A-�DǠfO�>�CO���"Pg��qb%�)�=Vdy�7C���������h�J�Rv.�A`���t�^8JB�a��n�V�x��IP5.�# �x%�""Z�&[8�3��x�Ա&8L8%Y���Fc������%/���]mQ��ͻx�>�ϩ��B�b�Q*3�	-
n��w���C!�#���@W�ΛC�YO��IFt߁D�wv,��(���n!>����Y�Mȥ��	��`�ھ�Ԅ����[��o�����/+�*k��0�lE�Q�.�ZJt�^� �Ż��cs�;��r�����c��%	�6}����Ĺ�wJґ��2 È?+����s��.H[\��ܘ�y����G3f�k�{n���̔XЄ&��&�%T~}"����F�`�sF<c��̇��0��E��)��8�����X��:d�hW��>��9�$R����������$šz$���g�5� �Ó!�4���)�g�'���3S�/Ē�.DЈnQX�|�q�Uo��>}I��?m��+�\O���z�@?��6b���W
z��8Q��PిF)����qUJIVП�;ce� -F*؀�n�.���5��w�#$<��2��X����x�BZ\���8+�4t�t&-������65=ߟ#�H�Zh����$OXm�;*�u�z��[���Dֵt($Ҵp�ޠ�T�\�ؿ�F��X��e�g/���2T��jU���id�i\jC�[�XADZ(�)\����V���-֤�k�{8�`�ױݐ8q�yN�	�y6o���b(r�t�K�\�������`����A��Wy��|�;��/��8iZ�j��� �N�9]��W�����s����)�k�;	�q����22�B9uyx��g有K~k�j�>G��V� ��p����|�l��hB�/��8XD��<��#Ҭ��HWTd;�&d�%xhQª�F{�:�V�}{�/?&q]���L�z�齔���8Yi支�e$�B�t�� �m�lx��4�d9x���0+mQ*-�l&s��ֳS-�f?E��4i�0��,���XI��P��'���b���`\2�8�:��͕D��{��`�X�D�y3rH��D���< ���xY7�<�گf'0K�LpSG޼��KT�Jt���\T�0/�ۄz�L�����a�z��8�aiBe�d"�]���:���1�9B[�MuA`�W� Z;�V�Ǡ���"���2~���˔%��?�R&�	� v�`C(�LZ�\lB�h�v��3���_��i��mS4��G�X}_��M+s6��6bk3�i���������~���ЛBR��W�m�����%�9��|H�#��u�����*� %�20�[]η~J�?�Ӧ�L[a�p���,�˜=��yc�t_<8C��=�i792�֦rio�}n�)Y�Q1ނ�/ �]Y�� ��lӛ�s�@&��\}I}�?�LIWvc�}Ry���j��!����fL�C��Zigg�p7�S��'�T�s�&r�f6���ʵ+k����_�� !�� �E���	�k=/Is��e�-�tݳ��d���z�N�ؒ�7%��:��^ �B�E߷��P�.�k����΅�Ik��USb˗F �H�AJc���ӗ���{��=�N[=��Y�Yr�"�XNP�)�~�GH�21j!=� 2�./+����5-!���o�
m͊�tC�V2\��9���)͵�-\�ِ�[�̧,�ǋ�oy �a*��
�7�/+�I��]��;D:��H�~��,�KC�99~/y��� ��ᬆ�Y�ʡ���W�� l�4����e�9��MC풏4�I
�"_���X�����ӏ�� ��e�d=�D�j����2��El����~�����CW(�H0�`����˄(l��NS&�%����l�6P\<�AU�� ]h����2��\:�`U(��ء	�D�NI��D� �ώ�n� 1 �驋�zB"{�M��T;(~F86���Y�����/q�T��aὕ��0EGB�e���y��J��:1d~�'�G�_Ѣ���~к��	W�e#/.�vM�Ϡ����e�a),U|cX��:M��Qas��毃�B���k� �h�7`��R����������#��c��܎>WGw7 31y���_+#|$�N�tO�o�T��V_EYI1��pX?�w��$剏�H\�-�
��.KX�L�����q0w�JUX�yt�T�V5�_~��dz�܇����c96��~���Z���CD���:��H.)���MF��{h�'��.b��mXw�M��d�f z<��"A��|3jmf� $=���n��Xy����Q��&��,1��3b�)�[��:��ʨ�s�&��M�]����h��r�)��*](�j�i��w2�"b$^\.��8�%������T�p{hH� [{���Q9Ŵ�>�r������N�H�H�?q,5Q�*�� t�{������� ٨�y�-O��w��zS���lLH���֠l{���� �������~c�{���U�Py��<�*����`������/cZ�T�U��������N��*�8�[��u�W�g���=� ���7��V���!.LBI�.(��2R�p�W�Ƒ����}�KPt!bK3�U�~�XOp�xv*K`:�~u# ��Z��>��2���*>X�t���-[}��%_:�{��F�D�/{z'��5���-�g����p�h;x��(���{�i�q8�:�?L�m���,*�튤����}:�A=�Y93`�pW���g$�rn���X�e�U�=f5h��<�ڏ�mb��C���k\��R*�������7�_����JM�0�DA�1�r��w�%͔Y�D����5vlN�Q��P�����Hɕ���Z�f��y�%��7��c���/d�.�x��H���7�ܩ[�*��A>�G�Ӑ �=���E˼ؘ�F��uma;VPp��L���Z��L�����m.��_��8���$k:KP�pr8�_?�,�qE=��� zC�
��D�a���4VVE��=*%���#])�9�~�ބ@>��^ll��/h��>�]�E!6<
���h�8����}�弿�r�՝��6'��ɠ�x�pQ� ��3��}���JҽG�	���0����R�1\�����e)�^���� /��0#҅a��x§��7_�,x�č�w��T��?2?���р�9�(BUPn��>e`��j���MA�8��W�8]�����"Ӆ_��Q�c02�'��A�3O��Q�UD�4)}�✔*Β���Q" :y^>�I�����J�YS��h���M���.x�U�ڜ8��T�f`�Z��ۢl��X�z0�gt�)��\�D��a�d��t�Y�6����d���(es���%��
�e�K�o5�̨i]ϵ3g�rn����� �a�GϿ}��'� ��]����3�
8�(���ɥrK7�J'U�Urgzp7��++@��r}��+�j����?W�#"����;c�KE�������PE��I���+�*Mq�6�LGy/�Q�^EH��?kR�xS��/��Z�#%)`@:�r)h�/zwK�X]�#+��c���&�3���g�I��1f�V�c�_�?���5�S�oF%e��B�/�8�Q�<&Bi��J>*.B�TrV�E�����K�P	I�:�E��I��H��07��D:��=_[L���a����A*�L5�}���X��+$���¥D�Rr�l @�w�7�R���jcnP"�[�hy�i����唖 �h��#�g�~�yXRm���!��%����K��-0�r���:�M�5Q�����E�T�n �I��3�Aϟ��1��G���I�	�"&�u�\1��`7�=�@(�a��c��U��1���1�a�:�КB�"�Y
��TaAn ���/z}H1?�����^^�ٗXe�|��V�6�_�{�?��U�����Jn��\"�J�{\�N!��E���@�@"�p�Tsm1�8�Ģ�5�8`l�q6�z����b;mn��I�rEeI�DǱ�?�̣�����Jh�0��F���O���л#���!Q)b�̓�{hA�/���.�U��)��,HgS 5 �
�ߞ�"��u��%�]�|	J����V��I���.#g����x� �a!�0���"b�(����v���1@�p*��La����1V|N�~�