��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\����q�?��e�I8�b�Ǽ$��"����ׯ1�V0����1���=ηE�˟KƋ�6��em�`d� ��h��Xk�esh����!n�*�>{Ɔb��@�x=\��L�c ��� ;+ ^� ��e{�؉ #it�����ZiH���
� e��<W�"{�#Va��v�J�ڏ�f�������
o�\�H�n��mY��?�Ȥ�v^	��x
��ۓ���j�h�a)'F���5�xqg�����o7݅r���Y����X,55�qr���p�uߥ�<YM`x!Ft�RDSs�&E�t|�@8�i�e�mP&����$�^�|c�;ك�4lp)p�y��M ��O�C@^ڭ9���A��A4��Ā�e-�Ld��%�aQQB���!���2��ف�h�f]7���:�Z�jZ=�� 9��6x��4~�Rs�A�F,Р�ٹ����|:6��}v#����d�O�vV��y�P�ͬ�� </*R�䓟N��W��������k)I�@>�]��v�\���O����{8+�`=�F<�/T����+/U�WO�e�R	��Ϳ
=fz�e�i�5�	+������� �7F�AN(��N�{��u����U2\�%�A	�C=����ǀ�PS3)w�#]gp�u�3�R��-"=�u^��o�5���$��o*ؐ%im����p����b��s9���e���������#b7����^^o�oU�܍W�>?*��
�IZf3��#	�S#*��TK�S�g���tO
�{�^u[	!�9z�:4��e*8_���V�@��.�p���nh����ܧ��&1Z&>r�=����yd��G�Q`���bb4���`�0p�@��j��Q��X�����I��Y�w'�[k}�R���ū:#Q�4S}�Vw�l�Kc4O�[[�� Blo. ������`�!C��O�c�b�;�&C�TAk6�AQ\��d//QM8'�'/�͜�|�h�x��t������uU�h�h�5V�Sr��F5��}e|RK�̿\��p��;=f�����;+�v�2��+Rn�����\ϹӇ���F�QP������ug����e1�3*O{_֑F�[[ғ���[�/'2�u﹩�s��\��h�	����[6�;���ݡ����F�5Ȅ������!�`"�A�:k����a���֯��ɩR��F���+����{��V/� �&$�m�3/�8c��I]{b�����X����N�L{c:Pt���-EfN]?p��bw#��S5�:<��%��E�)�:v���%��+Mw�ۙ�~�Z
�J�u���N��	���"r��b}�Zq$��|��&�+����~h�ʳ>��]M �?��f�{��6_������|,�1]�����?�J=iӾr��Js5'���$9�9����hKj�<�Z��Q���5�S����V����Ň���ڦ�_�~�r�+;�]^�4�	@�d�d~���i���� kr&�3\��@�-�囔K��;�'�C�(�2�S��V��n�%oX��J�"��a%2�s�6�%�]'�T�>;��T�|X-�5��]Vs����I��ei
� y��Ik�.8PRs�^7�����4��1���WQ}PrՆ���p�$�#U����@h^��MH�3!�g�#��g�ʗ���G�&M����ˍ������9�Z�;K@h`/��Ʊ �,����R00�D�L�����G�t �z�΀ߌ깩OR`�k��&Z�^���w��G���j��ZZ��KL�v!w�l��!��~1:��<4����vb�ob�$��'���j��E5���BSC�=EK������߮PB����l�,�H����8���@�>;-3)>ԩ!�j���cd �|ǷD�C@�t.{˷#���ޔ�]y��n��l��+��t`{d�y�����{�)�|�@�� �R�<����\�>�k����Y��X�%�?CNe�9�^��ɏ�_E�2G�gԀSj�7���Qa�	W?�03aR��d�>�_Bpg��5��}�dߪ/���s.�>�Ta]$�p�:'�u�+������h��ym��#����1�����O��\l4=ӥ� ]*�+(�X�͘=	�{p5Z�A��y��ID��Ȕ�&P7�$+ y�,X��SȶYm�����B3���{��/��"I ��u�%���VǷm.U6i�%�P~gH:����|M1 �*##x��8������m�y�\��M�?-\7�8�1H;�|��)R�#6Q�/o�`��ɽ�z�b��UӴ��-%�I�Ep�!�QH쾪`�=͎9�mW�Gb�\��ȷ�{��15@�}M�#����x��v��^���ɞ�O�;�N��Kx�8���ҟB�M��g�����n#�4�՘�eR͓���%>���!���' �����0j�h�'T�B&C�b�\���uw a��ԋ�V����闝�C�T����n��t���I�������4�i���]���q%m�{n�<���0��b|� %o�E�f�sU����*sտpZ��'٪ƽ���x���?#(nny���]h�`6�Φ~��t�x��*Svs/X��˖e��<Jrlw�o����fOa!(�<�Q+�l-~x�[������z�aBc%��q��w���"��
�`�.���l�~� �����Bð�����2t93�߱R�931l���K-HL���P�R������S`�����#,�C�y|�-�&S^w����dy9dN>#X�7�W���S�~*��CL�DL�.5��3����%Q���_�~�)B^��\P�Z�S�j��`6ٷ2Q	��;F��R�om�s!�h�|��
�B1����q���5�����q���$���=���Z�{����ݚb2��I�)S�H���va�L��G��tnD�4��OSqJ4|���b�� ��j<���n���>H��ͪ�5��&�*Vs���<�n�Q��9*V�{WUfJW3���q�ma|����q*4��0�XN��N&��R,=�>��.����9�-�mp��5�?��VB�%abu~l�`�Y��\�S�ZTYމ���H?|�%1�}�W���hB��f�[My��.��d�7d<���C	.��ؗ7f���FT��RER���L�ߵ4c ��j�� q|�G�;�F�&�Y�Ԟ�W�^��Q��S�����-^�M
��:o�?!�4E��� 流cކR5
��D��ߊ��<KE�������]r�^y)�f)�#��aݷ�L��� ��������ũ��;-�+��w�u�z��wT�{��2QH�`�Z�)� λW�oZ	�N�y~���*�w�I��+�}:���+P?��0kI3TH�.%x���䅤b�nq�:sRS^������ڙWX�G$�m̄u�jyK9/���~��â�q��̇'����ѯ�u��c�I<�����ʬ,cGjV��/� �������zt�Bl�(��e�;�jS2���k-(� v4���ΜPt��\�R6q�{�O��orľ#<�O����K�AE��[8ֺ��_q��ǥ���Ɂ�م�	�,�Idv9���I���/7E�@y)�H�����.��5�`�����h&����0pT,�v���We�Ƣ2��=�|�PpfV
L b�j�u$��g�rm)U��k�Ô�2������#�w�����Vr o�W>ic����c8~�0�˱��'�)�@XM�#Z�\Հ{��w�\o�4~̸l`�>��$�r�m��`̔M,K(��W�����b��2�ѻ��G�ʩ=t�(���~�^��D�+�s�u�w�>�	��<6���kU9O(�н�C��M�[Z=�F��̊﹠�r�C�F�/��n��'Tv�"�����������&���A�R���`L�.��[0#��q#� �~�m4o��G㏱ZL^m�0�t�@��g���j�s�"���!���HO����V���Aْ�j0aL1��O�j���R�y�Zӟӊ"�m3`jӈG���2�ޤM(�p����>vv��&�R��"g���Ә rˌ뻪丐
����n	���ԃ
s��%l���kT B���WJ���01^	,�?xLs�����d��!��B|�A�U�d5�<�R��݇��1��=q���Z�[H�g<]u��wx���΃���'�ì$�x>� ����B�I�⣵)1���d�]��X�G�!������Tk�[��U�H��U_3Ql&�Ǧ�2R1����_�^cJ;����=�DeI4���fu�L��A�^+̮����~s�iUm�AQj����(:��d��p���p#R#~����,!�� ּ���V�&0�m_s���/+MR�ߴ�ֲ2�8G	e���	f�Z�XMЮ��v �h	T��q��z�M����05X�"�m#�iT��2��Ň�_��P�.��y��n��T��?	"?�(܏{m�q�ޟ#�/�:Ͷ�&�n�����1+�ae--��
�M��[\�l%ۤ���=ߞ��3��*��ߣ�dVO�Rh�MG8�G;rSD���ފ��=�a�V�yﺨ�95z!�T�`�{��{ߣ,3�Y$�,��kߦ**�s҆.l_a�h�!�<���U���t7?�u|��x�X��G��q�&6���EX�	{'a�����	]M1LÅ��j� j*.|T|�_���p��c�[K�p����C��NO�݌JM5`nK���j:�z�y�/�;5��a|�P}2cV�� �i�ɛb��]6�)�E֜�u��Q0Ĉ�n��`>��O�����'���ͽ�8{cC�mj	�H��x�Ƀо}�p���R�4Ǡ��9�Da��/DbLܺ%*Z���XCU��(Է��^�����w0Y7bﶘ*�̣몶g�Eٽ�CSUM�J��F� ��j��iM$*%y؇� �e��0��;)U@^ A�ca��H7Qٷ�5ls��?�/R�e!�	q��4A�A���q�5I�����ژ7����Ѱ���x��n?Ŷ�$���Dg"u�%��(v쾸Cy����%��E�������~��d�����_QȦ�Ԫ���DK�~_�U>,�m��I�z�9Z�]��X����k�u��f}��0�l�:W_��!���&������>�"G�@�)��-D�8��Xa�=e�B,�u)��.F������!����>o]�;b����ϔ&���ǭ1�+ d��g�=I�+�
��'��Y��|n�M����DS�~�c��/�їS+e�^����wK�e�]@� �`�+>�~_}����r�<X>c@V�)���5����_�v�f��@/�i.1�Ti+}d�,�Rr �'�Y��n>�$QT`�x>�=�y�2ݶ�~�V��7Ն�)bU6ԻqţJS�1jI���aC:���Qe�A%�.	o/�8�]pQ�6�Y�˘��-U�(�auΞ礒��X)���,V���?�A�㛎Bj���7�)Z���|k�D�K|�B�Tl�ITe�zh���u�~V�%|�8vZ��*��y�u��PIr�Ux�ٯ�K٢|R�
z	C��ڭ�,7O�'����n^fNB�Y���v)Z��_��u/?��']��fC{�eʥq&�����[B�4�W#_E�6��
J��<���;@���6����?�;�LP��9*}S�gpڧ''9�k7�^�SF�i��C�K$3_��&�ܤ�N��#է�f4F��T����A�K��gL&�O8�X�����m4���t�n�n��ȘڂVQ���� RN�����L���>�S;A�J��_�i���*�s�;ґU���dF�N[K`S��QWcy��^����g����~���-$߽�m�D����3\GЉt��s�K\W�쏔�I��4\�	� �Ă �&|����TGyp�O�>���W9�����;>;p�	fᲰup�! ������8�K���5's��]�-���@
��?���F#�d����9��I,�����w��ta�.�!ky:�[��o}y��p�H�q>[eu�|�d(Bi���fe��b��A�� �h�@3ڑ���W>E�� �ͶH-+)�'ɇX��O���<p4��@�4�hc�W'CW��B�Y�Л��b+ ���^����0Ք�ԯ�Gj	d5ۖ�:(�vn/Q;��Ԕ�|ὕkp����k���X��K	��zWs�.�K��&�t�6rU	�yz�O��Ez�d��u \�g��璜r�q02u��4Z�[�S6�"4;C�l�3���Bpm�_��pi�����W���_��`��,s��Qz�y���,����.mV�pmR:�3�h��]��_s�V���}��Zg�}�F�)䏋�CH�=EJ�B٧�(�2�4���mvn�M�85�'{7���BJu�Iy�6З����Ӏ�o��#�h�LU2 (�jΘ�2��29���%��L��ṏ�b-) f3�f���D~Sr��n_P�|W�#}��㰼�Q�E҈x2� T����̭+.��"��#h ��=��W�rM�\<Ůh*�k��#N�V��1*��]�QT`�iԊm�<�����d+�qAd:3���9:�ދ�N���Fȃq`̹k4�"�ނ�}D��$[���n;�I�uW9^���q��9~����F���1s����IO
�f����G;-T���]H�\�K�h���1�}foj�Bu�d��c�xg[�N~�+�H����r���6'��zT7�%v�'��bл&��y1��v��GI��,+�v�˥�5��w��ZL��3�w��n�V�\\�jA_���H�}�,��)>�;��4M�ˠ�U�%�i�U�v��&�Q=M��R��'(:���ǂ�Q�x���1���bv���_<;�Ld���Y.��eY)���,JE]dix��;������9%ӳ����C�$p���[$If���C��?E��w���ds�I;A��_���E�J~��av�E�P�T@�Z���s�*+�	i���2T��i��U���rs`���y\2���/o-�4ż,����qj��#	��s�
4�vS���3������I�V��$ʍ�����`uɫ��C~��s�Z�ĘF{ll�����eC���$@��"?�.�ӻ�$�AWE�)�Y1{<$�=]g����H�P$�4�'Gz�kJ�,a�Ǹy҂���T��{P�F$�M\�B����G������q|���+jk��X?�{6�t{���r#���40�x�z;��$�(v�U�J� ��U�Ua�J��d9j����q�+��0M[��@�z[;�j���V������vK�N�1Q��/�0���f,�`#�0��%��T���:^��� =:�D��W���G,/��g��*WvFs�Y����lr�Rd��3m �7��*�>^�XoaTښ�%E�s��_����W�Y�|g�1ڍ[ۄZ���Y�x��$�;MQtO<�r]I�����������3g�Q�� �S^Nn����v=���Z����c����xW���Ata�Xq���J��n�[h���dv���u�Y���8Ƒ&ޜ����j��c�C�e�hg�=!fZ��_�K��L�p-c���DL������=����4�`?@��)	6P�w/N�9S�N���|H:���q|Öw8w�ۍ#����$��| ��fO@�ߞ�hx+풶-�~ן�&'@Mh8l<|1wpv_�b��䱢}���uT U<J��9�+�P�;HT5�m�_R�<�[�m��^�C>@>� �h���0E���ث��.�Q-��;^��኏����q���1M|M�f���3����2�b2:�ȿc��u���!:���t5<&&�*�����4����V�GˇC���5)���CX)�О�f������vf�ʚ�l�_�I�ǎZ��w��A����o�v9���č9��C?���`o�|�s7_[!2L�2���=à?�t��^�� 1>U**���1 ��&s��.�v����S�N��>��^��0:��%+��S��,��</*|�	�����XD��t6VƆ%�N���8��ᘿ��zTg����^ 'E��5�	�/�H6������f�B��v�F6|V5��nLZY�Q��f�? V��q���7$�^����T��ni��@���6���f?�QD&`����_<�*�K�3q�֍�$�'I�
W��Dζ<�\@�R���"
ч@�u���L�;)�+�I%���:D\y5:���M7"G�H��nCa����e4��k��A5
�U�`՘/e07v�T����O������zl���jf��9t��۾�
���?�[�~$����)OX�k�Bw^l|������� ��&�",�λ�����-"\dj�1{]~bI�+{:�0�>k��{�,ä꨼�>^�A��3:�#6i-���XtC7�Ve�fsZAB�N������v����Ԧ�w=������StR�5j�oF��t�fȆT��9��*�
Z�.b3C"��u����|dl&�'v��_�ї`�_V'����AUp�3�9�{�&,?T����,94���!�&G�株g~��$^Ҵ�F���1ϭ���c�=Uv�錨�{����b����3�e��6E+���6�����l�wT|I|��JGHԅX���ںo��#�����yO�~$n�HT�R�Gk,��Z�SP�4��Þ4�v����9/��F�}��
6������H�1��_��o7�����|�[��ㅙ�+7��vD�$�ͱ�:�;���%�C>1,�9v��3�J�;*L&Tɬ�`!ޅ��8\�5&�׀���V�cF
�HPW���n�耋�W�$>�lI��{� �i�Jч]��@e�!פ׈"#=���) ���*�"L��	�&<����di2���mJq���a�=���|�$D��������Yܠ����Z����TT��j����C^�ٚ�y�N��( &��{q=�3�3F�-��L��d'$��v9�K�\�5r�Y?L�X�u�{W����	����%�T`��e�s%(}�Z̐	��a�푋F�fN���Q�4{�Mr_Dm��Q��5�@FS�d'.V�� ���B���������˴��=aq�:3�g3�v~.�Q�����!+?	���,����JX�7�<�(ˀv���6���O����\�����zbT(|g����F��M���IK�_?8.}���*��[�&6%���};�����v��q���@�	��hW�oM��,��~��e�	����9��V+��	��`�8�n:ă;Lљ�5���`�E-�����/�R8��LZ)y�l�.K؄w-AP�#1�t��l�>����E�0lj�f"$ow	�[���U���U�ɬ!�?��*�Y��Q�3���:��:pd Ȥ����ݝC���	 ]pτ���>�7D��X@rU�Ї��ڼ -vۀ��xM�04�K��X��	�l�u�oB��[�g�6��-pO�ۺg 7`�4b��1�2<�ɗ�n�)���j���r��;T� �Ƕ^��&�=���k�Ѵ�h��E4��ͱ�Z^:y�R5��;9���
�7����r��m��՛4V��"�6��x9Jj߹(5�6����)�X8W����ܥ�	ۘ�R�y���Pض;wF��D����U1G�vn:�dt��w2���h_g/1��&E��ec^Q�h��7�+%rH7 5k�#i6P{��Kk�M��4�E���.փ�g�~�Q�Z<�ۿ�L��/+l�s֙5/��	l�0��[���r,×�4���bm�J-�̚���6h�����!�5�[T�a� ���5��p�J��c$�i>|��#�x���$���i��@�l��VtX<E��S7VQ�,�#3{��̋�Ƣ�w�su��g�J������Fv���e���4�@��<e�����X�'�����+=7�K��O[���o�_���T�n������z;��,��l7��s�Y��KL�x�ZN������#�jh�ȿ}d�{>����lIgX�Ӱj�l������>$qZJ��$�7�V
����;%��.�ݱM���Z��`�T�������~����l���93�i�`�ꉈX�E�S��9a��q3�� ��G��u������p��� s4�C �&�\]��p�&��E�/�k�R˸�:�j�%f��~a���-�	" -��\l�N��l��Z6��y3��ܒ�*�b�?��%^?_^I����#�a���4|�FE�k^��4�����3�ݣ�y��T1��M]S�d�P&/<d�v^�]��f�N�<�s�����V�_MmG<y:s�����(�<�����(��L0VS�D���^$���~O��Ќ1/o�������e�M�o䅽 `ԥ]��)́{M\0�R@fh�`�D�=חg���bγ>T�����뱽{L�źgf��;S�zA.bFaK6� A�ɖ���h�k�x���jz�9�(�^?����YCʈ�1Ce�=��q-q�B��f8� k4��,Rm��9�qñ�##���~$H�wH��}���P��0�M ���nwC����n�y��W+�0�d�q,}	�z�R��W 7ݹ?��O��m=����з=~5�!�V�~O�6��zn�Ǻz�_�kc��:ߊkM�ڠ��y�8Q��s?rk�Yl�&?(H�?x"Y��x82�'�9�ؼۿbc�al��5-�Q_�t��v�j�=p"��9�=ޭZ���f�v+,VѺZ�6�Qkb7ic-#'�}�����ke7(�3���cM��ѳbX^�A:|��'L�x^$KcM��=�K���z��%̚�%�8��_]CYԬ��c�.��O��ḍ�MaՔ�F���>��(&�gX$ L�^�U�=ņ���; jMi#BZV��pC�G �+��s�0��������lu˸�J�-!�W�� �7�YXR��[�" �44y6�"�� E@��z�f倕�(ߘ;�ɸ�uo�3�C�~�R[��;�(�kM����}���ÐT�mCib������>�/��;����Q�cm�����ì�{��fia�V�bk��
�E$i��՛w'�],�Q��Va [Ѿ�ZtD��C0��"��;��Y�B8���8 ���%J���\_EeNCOS߆êa�����("���x�@v9�6�|�@u�����?�D�~`U�heEZ��a����RFDshZ�_�[3�c�q�������謸7�?�uYIT�܌��Z"BR�R�����|�v���=�L����� |��e�m_L���/9��U�Η�8�:!sjN�-_�$��"E�<�H<��ov��E�XkI�uN|�@�j�dE_�KqW=�PAi,A�<��Ѯ�Pep�Z(������)��������Ӎ����{.o��\M�D�����8���3z������t���.�ؓ
����5
�"]C�C��_m�FMK������e�'s�Z�Kz^�\ݣS��R�gK
q�J������T�6X��f��Ԑ
Ȅ��!����$h��|����Ll{O=:��x5����ϔ��Z�1��#��d�n-O�o�4Av`@�o�`�
nР���YU�Y��sB,�R�B*mﵓ^*���<�%t��N�"WF�Q���k$� ����U䲚��&��#Gh'`��t���A=[°�dԴ��N"�Q,���T����>����t�{c��w���R�H�|����z��������j���I��g���i�'�2O����rx.��%�$����K�Ć�tDF �3H� ��5O~����A����/��,�?A�s���葳�bޏ'��N���?g�̯�*��·��X��@��T?Dg��qq�NkRyr2��6����ǅ��={�U��"^�vQ��Gߦ���y/g���_���з��{��h�)����!#�RZbo��(�Q�����	1��Ê<�u�S��D���g>D�4s�M:w���㦘�v����<z���2#����Bc�������{Y�"]�������x⥮ 7�(�2��b�KR{^$!��a���έ��������<j`�,��B��yD�p$�v=�*�o1��YX�|�h�C�7T�!!^9 �]e3��}~#E�n,�*�a$u8ξ)�J#s���o��2Eo>.k�?E�8U�L�-�k0��[��K�+>�]к�`�x�늏k���n`r�&��DL�������Y$���_n�t����pke�(T���t�;4^a�RI�g?9`���5 (���;֑ �n��+�g��'ҮcK��G5�Bd+^���������Sc��\b�����`4o�װ\��g��V\A�QҞV|�� F�-W6D�[�֩�a�ϧI���%v�Gy���UIY��%n�����<����@���Z�G_ޚDd��l��˟#_q�u�̬o��R������������U>��VE�i��1�e��2(��D\������O��,�l1�{��A��
U�PF^a�L��xKs�|ܚw�8e�����t��ZMͰ��`,o���|UV�&�T�N`�pt��nr��{�קeO�[��4ڧx�l�Y���l�Ѽ���iXy��2�d�V�[D�;[�sO�����ɚ�����A��|:��tACb���X�B��։W����r]�l?����{B+?	���u�k C�T׳��s�69X77k��pa��;h ��v�?eřܾ�1�A��s0V'C���@3j��"��o�zGal�M��b��G۲����J_�kk�mV{7�����#�+����sI�\	�u�����@��,dQ���_�%͆�@��#�j�L�z����j� ��.���9�ǋ�Vͫ��NGi$Uh�tݪ�ڛ�0�>7�uB��Z�N�5�eT��PU�=_�z��˾��8B��y�_}ra��դ@z��H4�K'���TG��Y,�%7�l�[|�e�6�_+���,��CΜlU�`���GE���z�^�z�SX���L���p@űŀ�Y5������W�h�S���g���}}�\�)Mrύ��a%B~��V����ۡ�'qφ�] ObP�m�5`��ko}dv~h�����^��:�J����ha�L���B�>o�<"`z8����,�p�b��c��w��b�f��ܿkw<�u��Fd�����W�߆�9��F�-M�]z�5�Ml����3��U(�O&㱓��s�[Nۑ��S�W+٢��*Ƣ�F��y��sw� 0]�J��+<Nǿ�F0���L��u!�LE�SZ9;g����6���-����[� c���X{���b���?�J~�g�o6�CQ����{��y��+_��
���N��hIv�Lr.+��H�C�����l������ϯ^�x`[�ֹ�$I�4�K��1���|H����J,�q`-��$]WBT桷��k|t��V��[���|�}����1�)B
b~���@��37�m�������uA���#��:�	1���lѹ�x���Y��Af�ǍCK R+=��n��\s�xI��rG��N6�O=>�{ן�!<\b�}�������}v������A���+�������m��Cc������{�o(�� �
4�iL�D'<����>�ku�&T�}��~_M���W�1�n�Ñ����絁�\���-'�Ә������:K�������4\eE��{���[N[���2��I��6���ޒ?���� ��V�e=��Z�]�s`�`&<�da9���������rz�Y [�����W�`��3�O�����H�I`�M-��-����O�EL�3��/�v��Ֆ�ؚUZ�Ɋӆ�X�8��s@�� �U�z�3��'�ӎUE���ɽ�n��9�/�N88�R�Y�	P���c䞐��,M�TD[���'��N��1�G�Ѹ��kݣC���-r�?�6�AZF{�$-�^�Y5<V6����_��ƿ�FbS��<C��X�0�:G����;��G��8��O�a��]��ն�Өr7z[�/L�MXR"
�SἵF�������!���7��]-ɢL[�3�wp�:�3�>�q*����$a�d�Z��	�bX��(����_�7�������8J�9�κ/cO���=�B(h�4�$	�Ş8�q��ue׾�gμ��t\�{0�>RH9�7`�{�)�`��M���H��r������b�`c�h=�[<���]aۻ���Q�Oe]��U,+�鿙:���կ맺`����b��JH�=��`��s�Ę��K�Ƀ��:\���?V�/����ً̿"���j�J�숮t#�w��$�E����ݕ���Hz�D��D��M�Ah���wmё� ŕ�n��-��9�7�� jӌ�/�P��PE��ʬk};�k�w�IjB_�9~�b5l��s6�
�`�i���sy5qr.�Tj���f��'Ԭ��sH@n�+��q砫3B��Ј�Y��k���z���g��bPZURϕ/�KJL.��V�'�pi�~H�ȄW�\~�bf�%�N�F[�r��ߜ3FL��-��>���w*i�t�Jv�J��s�b�N5�?��?����ak⚋�����,�7ADz�6j�R9LJ�ՔЗ�(�������r�/�"��^���F�	��b[p��IB9ܤʦk�ɬ�\��8��%��H�8����oX����&<I	.ii�m��!�f����3�f���\Vu�O�z,QN�5C�[���$���&;��h.�g#2x�I���`�����s��^�#�	�;˝�32���9 ��jT�C���0!�4�HЎ��7�.�S�(P\B��lvP�}5���o���m�X��0~��e�m����w�\p�	������oPs�l�C��*�2N�;�
�4������e��s_��Z]dr�I��i�E��3�ȡ��s��E3�T�<V�"��dAe��v{�����/��Q���r����o���8sH��KQ��~Y�rE�^4E�
69$x���w�8��Av�C��L(EF|�ƴ^P���=��\��&p �/�T�Ѻ�KE"�C",Y�)*Z����,���vfkDQ�e&�Oy�m�Os��QQ���������r�֚�	�q�i��伿�3�%�Y��k5�/38�
�>&���O�,<ǆ�>:���a��щ���-�R�*�Y=:2E�c�?m�32+HO3��Y�ј*��\��G�B2?�ȜB�J�u�fO�,�hĸW���X�`q�ֹ���ԅ&����K ��8q^#��4�౅#^ӿ�;���P��B�?]kS��ZWf�ړb,�K���mxJ��f~K��&s�B�9��ɲ�s�Շ��F��V�ޖD!��e��@p	���$�r��syΰ���NH�k�=/C\�9q��X��3G4������z��?3q=L���x[<xHDE�S����N�BU�3�(�  wv��������4�q� p�+N���h�	����)������Zv/�yk��ڠ�?F���D2=}/��nÇ�5�[��?V�C yFpk�6��Q���x;�i!�����<�Qٍs�5$�𐇥4���Q��
�<P��}8\�������������о!C6���#����a��Jkj��K��heK4_�+Ņ��'f=���Cĥ��x5���=Н�X>�K7v��L������g���$PB���gDM������hK�,���Ns(؈�[�1�=G�P��ȵ���������ˮq,����u�/��|{�&�2g���: O̠�pQ����d��Կ��9�L(y������:a�B��t�̪(
��#:UD0R��� ��I?Y���;���"��7����шW--�����NRa�v���E�����y�!�7׿�eh6<Eq"9�c=���W2�+���%hCa&�b�Bë1�6C�P)RIf ��Z.Q���"؂�'ǯ6:�	r�2!X�fY&A�H����.#��$ ��P�@�ϰ$C�SEB�S�%�u�!�&����^�?��&������5�Ln�/�-^����c����g�o Rݚh#�=�/��QSDKo�ڂ;����i!�bY�]kM�@y0)f��H\�]����H�LӾYmR�pPM|�������۩��Ds��h�Y���O3�	R+��'X�D@y�bV�:p���`[gAj��K
�gۜ6�z�n�� G����ܓ9�'I�_D���,|��G.>���}��B���$	+��r<�[S釸����t������XE?G��~�� �3�%�}���`㧞���� |���y����π�RJ <�M�{ښ������V;լ��������{$j�:,g��cn&����2�K2c}�X<W��"Zz@� ��^깭�;�s˺��XX�m�z�z�F[ v��Ĭ�f_�������K�qjݶ��k��U:���z�)��<�t�	aL��T�'�]�w�����U�}�懶����I��ܤ��wEh3���.������S ���_��.8Э�����E5��31�ƀjhqȲ%:"�Y��|��8�0$�%UB*b{aP�)S@}��H�T����O�����gO�FK����Ƚ�L$��+�6pT�$ᴥt�'B��k���^��a�as�T�J��(N���i�{�w(�i���a��T�4H���J9�P�q�N��8��h�ƽ����_�j��1�Z�; �e�B�${Sby�S�B��U���B��6k�xd�w�=hB{díbm-�W�0/���?D��.�8��Bb���H1+}V�������
�ݽSѯ=z�Iְ���G���i�X^����*2��N�ʨ���F
4�M��Y`�sDA=O���z����k��B���y���|l;Ў���l���R}��2R2m��W�� ���,D���cM
�]�y��*C�
%i�4I�!,�3���=*R���wA���!d+�w�zx/N�?p��۰�H�4�����S'OdH62�I}��
 DWx��U,�S1��4��my���j8�d�w�s�I_HoI$��d��.�sV�Z5b?���W��������mj�am�'Y�Q-�.��Q.�#�ؖlP��y�*�ܥX��)�¦��2Y7��U�E/��'�ʕ�@ۭa�m�<�C�j�h~�<�T@ʼ�Gk{��U�-�eS�����Q6���,�^=��7n/�_\�K�?H����V��C� b��]�מ����]�,j O�q�K P(������,�U�\�=>=yv��$�׻�ٿ4�������#�����=b3Vͅ��Zs.�}ڠ����9��J0OۺCe|Z�ŗ����=G�k�n�4k����N�� k��%�Bx�[�Q�� ` @�@�����8b�����,���Á�8p�{k�)��F`���C8>m��|hbt����Ki��������li���NdV�� ��I����
�r�R&��3�|y2u:1�`��'�~o�x�6A�ɖ��{m���?K�>B�? x� r5����O�c/�TE!i���]�����^�"�2ppy������F���-�VR�!���rE���؎���k�]�黉��L�|.jC��$��H�:{�����i(,�Zܚ���:.���g�@���.I�E��Yt�N�H���_jv`2�}Q1'�.#�1�����Z�%� Q��)OM)�E��,��j����y� p=���O,1�~a>cxΪ��̪.�hC����H.?�E���v��8М���\���`n�`,[#�b(�w8<���&�¦泮,Vex�'5�ھon�\Y2D˧�2��y��.}�U#j5z���9�|�&��Ɍ@8#� ����I�N�o�}h_�|��O���
E���eQ�=�i�ِD�A�����'�����z���;x/0Цc�a������jK�p���3n����3Y�LY�J,�d�Z���|�X��b���I�!ܰ������h�f���Z'�!�C�	�POO1=J�e�kZO�P$ʻ>�26n�޵��Uzh��m����0�	��������g���AX��a-�)ڙ��?hͣ��o'�����e�^?!�W�7����OV�/�{1K��A�rh���T*#))��U²H�ߒ�$\����7l|�D�2�~�C�H&�ȉ��)�Y%�f����
�>1�~�&�tZy��-n_Wح�
�J0t����o�ZVv��~����F�!��C��.�6�v��s43��Q���~�Ʌ,i���'�T�kM"���s��?�sE
_Nz�+T��#�٘E;�
���hV��p���+ Y�.����J6���J��u����]"=m\݆�R�Ά���h�VA��ܢ�&Gay�@��ό�4	�{D8���Ʌ��A��d����@�lKz����1��4���������^W��j����LP�R�u�[N>3��hz�jW˫=��G�C��P��RָB{2�
���%8����z�.e����	�bʕ�y�f��#�̇��ˎ�����o�`H�b h�&���kg��o���2{��3?�EQ���:�������,v߱�m�S!��&������Ǽ���m�N\$:Rv"�g����(�t����{U����k	�&�x�v���-֧Vk=�%����m�WΡ��5K(U�S���Xz�
���sq��vn��n?]�@�4��O)��ϱ
b�K��-P�*�$�VKF�?����?�A&���hu׻zAk�B�q��(2SQ�X�C$�-��#"s���h�
WRI׶i�6�`��P�TM�����, ��I`��Q�5م!D	�(�^;d������s��6f�)1jd�v� k�Ů�~(��ό��YP^���X[��$�1�,�z�Q���"�xa������>C�I/d�z�"E8Ȱ(��X�ηEH���84i�h;���V�}�m�Q=�B7?��FVyj��L��yؾ��\N4`n����L:^�sB�����4�d���w�_\�\�yA�cc��r��(?���}�S:�YYܜ~#���µ�`m��|Q��mF��~Q�f\d��>�L	O ���I�L"��@5�"���>ߡ��x��hO�U�[uv�)���n�2���½�Ɔr�Tn�e��m2ژ��r�C�kU5�JΉS�?b,E,�nG�S�l����WUѱK�i0�t)t����w)��c8�6>h�q��d
 ���I�x.c��&&(�gY�>��M��o�Ǎ�f�y,�6oQ-Hԏ�O +|{�b�c�}$��w�
�u9{�Y��P��M�&�97�^�}��hU�j��=Wkf�l��m ĉ�%�������"ĝQE�Ob�H����Ehw3ċ��后���vj��v�|���|i��^���Hs4�����R�J��"�D
.�G!�z���� ��a��MVUX���N?0��όl�aQ��T�/�[}��Y��SoT�"O`�r�E򺚛�y���t���<Z��<�#]7��J��3?"oԬ��\�n�Ρ��q����T�W&	�"6+�~��^#5�YO�ac�э�����S�Ta�A]��2ڨ�1t}��l��� ���?��>������ ]�9}�p��[�F/��bL��������ʂ)D�Q`F��nB@����~XjwL�t��E�°ߚGg�?�$�1��:*dx D�VK}xz��W��y"�Bug�W��bA�����3WC���#�!�rM�����E4�WI�u��w-��,��Uɨ�O<*m����B�Y�i���E&���Y2u�S�l�@�^Q��k��l�oGVO�x��gIr]Wڙ��K��R��M/�Ϫ`%�>�Ͷ��ѯ��)���]���њ��El9��b���T3P�"M�����"�q�;��T6��*�C�e���`��<�C�F�QؓBvJ/���m� �x���T��±Te�e�[�_�wV�`�-��Q&dFX��_����� cSt3�B�e�=R�K�IS9��7zC�)�@���K6��DF�Y�t߬�k�<c�=7�:t�š9?���\}ʐ�� �((e�wZVN��Ľ:��9��Km:4Y;�&fE �TSel�Af{1�b�N_���Bs��Z�L�_��D����;����BE����s(Nn��<��;��=&���C3�G��f]k4�B�����c�&J�ۀ�6��̝k��l�kv|�?�(�����E'f��(h�(�Lf�����nN�Q�<q�f8;C�_ֿ��<q����"§5�Ev�P��e+gO9�~�ٝ�@ � �k�(m��1�����?n/��9`t$�t#�	�;^�mG���%��Em}?Vˀ᳗J*��`dB8��!��H���+�"�cG�DC����IgBb�U���HІ5YHL�p��t���B9�=@���\P��������\��5E�����+����X�	���f4���j�S�Vn9p�,�]e;��|lJ{
�~��±K��(lP�i{�[�~w.+"q9J_�}��^�~>t��$*آ�_q�D��lcY��m��y4ڊ}�q./Be��iJ/W�@����?{��H$�IO�M���H��1���j���¼�:����E)��
L's>3	����;��s'���Y���]1GAb��f8�2��2Nn�+ʆM��VC0�a���[���P��HB��>�*��+����$�!��?;�~�D~��֌��Rh5@������a�{�$�E���¢�	ˋ�',+	���:(����=��&�_)\x�S�m2��c��T�����ys�/� �l�
��rL�J\w7@�x�4����U��˃��$���R�ǌs
_	f!`�Y<���oȫ�<:���;t{��X����fR�z�L�%zͽ�����(�{��Y]
Y�}�-
L�� ~DtsMWZ:��Gn��߬�e��6����P>��I��l�j��*1��?d�9�e)�1�L782p��m?����̈[u��l/\�#���T��B�Ž�����
f����c'�ڿ����Y2��0u�.�
4��A��ϩ{J ں:�be{���]�{3兴Z8N�?�A'RX)�&(�ƹ�B@��}���jKz��G��3����0E"����A���&QI�=r��p�Ju�S�w�`)��'��C"\�F��v�$J}k���1N5�Im͠� ���SA��M�Z�I�������(Q���5����NN�ؒh	!ƩTy�jj��r�Y�L�Xɚ-%�5SV����`l� �zezMMB�ַ�QS ��+g�M�O�P(aa�1Q�n>)�\:���]:+R�!�i*C���'_��*�;A��$�ثo�����H��Z�p�Omcǩ�(
�L.�)P���Y� �������B������༟�[�{q[�}T�F6�KۚP����m�x
U��]M�����ͼ�ߌč{_�XH2X
k�N��]����++f"p�ԁ�nn��P�H�xq]F�4�w�j�ފ]ۯ�Y_��A��q�m2�(I���ؔ�^��������8�W����}�R�A�)-z';e�I����:dK��^`��[h ��`��<�b5F�!�"X\�I�޿� �"S�N�����>����#��}&up�*U\Fe�>�JS��^hگTࣙ{���lu�� ��U����ʇH�I��5U�"SÌ�p)L�-��'���I�IB����3��]X�S�W����w��.�6��1Z�<˰�G�ψ�f�Cf��H�D��>@�J�N�Q��xi]����L@RInN��8#�~�}թ���㭡����)Є���f��GXԷס� �`����jq/�n���,�hb�ke��`jd�囋B�m�H��9��~K�	5��=��a������-*�	��� �����b �Li{�醘��uB�~0���hn�b2�#Ӗ8��;�qXi�qCw��-�)!I��z��n@MP@����8��E�����*���iZ�N�w�+��]S�!�-V�%9gC*�r���zY
]�-k��w��-�J��(�R�����)ҤYY�($�{��b�������%_�r0ɏ_�4���3	 �K�4��2�7�x�Wm�vC-��W��o��J�����"@��10���G�@,��O:`�X�+fwn���������\X�6n`[O��(�T�P`X�^6l�d��L���_�}Ӝ�b���f'�g�p��U��g���:��D�E�Im�[�/�˚�J�@�P�.�xX��Gs� �@�	�E�K�Ѥ+*�%�c�+E��?y���C��)T��c��W�,�\����ąe5�3�>(G�U��S�`u�|t u�X\�����'H��;��?�N��0�#-����"���p܀L�ょ�
|�0��A>u?HOKʁ��1�8u��3����;�]* �f�+{���K�7��|�LYPd��F�<��Fn�X:Bm�3�ރ�������x�
+iҭ6���;c��f�A7$qs0�t1~�5|�f�wu�W�
�ȼ�fTbY�i�(w:�w��A�@�L�����p�C�F�1���%q8��8���P�7A��*�-i��Q��:<��<�\��9������Sp�IϠˀ�_�א��߿Ap/��S���.����X^SA�tR^_���H8�</񥶚����W lSR>�
~�r�ӄj%�*��4����p�#&�=�	,F m61lg��;�<��(ݷ�Q�P�� �$i����N��䚐sz��"�r�HC��J�4�K�<i������= #�Y����h�E�E�=�H,ʻ�E�^}g�D.*��KEL�����4m��=MN�r(�c} �b/G���'����_��H�G��بȧ��{0�ZQ����ټ�GD�)�
�*V1Q���k��=<=������-rc>\�7�f�*���[J�0�y��0[�j�� ��Ofa'��b.����%�ե�>�
�;t`�>�ރ��So{Udׅ
f�C�� ���IS��p���M�.8������{��g����t���u\lv�wI��q��v�h��:�[׀��]]���d �����%ч�-Ƒ��?O���K��g��aÍ=������w����.��-�U��7�7���\~�Go�_m�_��E`V:P3�=�%n��8gjJ=��c��'�˺<S	�i���a��j1ohc��M�E*�M'��>i�VU^"ik\�:,P�����*p�zI
�E�#�8�2��у�Ɋ_���q*��ߦr�����N*z1�5���ճ������GɎ`�{�i����u�٣��z�w�QƘ#��l|���"��(M��!O+�f�v웮{�l�΍��l����=6|�����-?�"��|��d�	�>��s�]�p���0U&	X���]b���z���k��ฯ���lg������1�%3	��N�	���-��cJ�����Ǵمs6}1�A*U�.�,U�e�`�IV�)f套H[߯�6�T��S}�O�3�[}%]6ܥ���4���#�$����� ���ƹ��_"���G�'��X�_���6�|��6�KvM�IȮ�������%7���"��ql���U�׍�1�~{�����a��wi_s�B�Y<����;����%��q>� ���(L�@�t�1�©�p���t��mU纒$_��6��K7=�]�|�H�kv�u8�]�ς�� ҈����n�C�)R`�2R�!V&�b�A�äW�CMjh�F�����bmK�#�ҿ�kF&'d�ߣY���{v��~�P� ��9��'�K�����5uIK�$�(�9�B�G�&��j��JlF�ck��,1br�Ƹ'��Q'�j�K.��"�Cו��׮m��uG��" ���"�*���ɻ��[��$`
��ҧBY�,=U��ٿ\�=�ީZ!9$��_�g�~�+��.kSN�ߐi�F֫��H61!P�O�f�e���aƩ����JZ@���7R�z>�������0>q�H-��ϨY��4�;^»�B皢Q�N%8�*I����U�Z��R���k�S�C߼kT\q��(�|q���ў�.`���H�꧛��D��a4��/�O�D>Z�\�v;��'O��}o�Ye��<�X��0�VfU�ւ�ѐ�]�dB��p��n�EN�Ǳ��H�$�0�4�Lx��¢�_�,R#�0	��Ҋ{��Pz���\cӁhַ+�7Nf���A;��rJ�K��ĉė���6�e�q|/����Pe����@,��0v�ϩe��rJp����y��c��B�z;3�l&��hb���j��|A���@*v}�뤴��Kr�7[�M4`�	p��ğ�u�G.B"(��TM�Ѝ��,0�lo��-�$�O;O���e8@�vg�f{[��f`Wl8�(�Ui��^��j���
8S�M8����/y�a6�k�7M� ��5�����;�F*&�����t�lpj�R*#.r��<���5`�|�ETY{u��G/���sbd��w_E�/it^W��u��D��i .�{�ġnv��Y��p�����G�|l��Mjɣn�(�&�i�����:Re0�#��܄�~*��֑�g�;��<ԟLh����tb������݊���`�9kZom�����D)���&�1��+�ʝ��^��e����uQ�l:��MY��cr��\����1���7�{�m1L�����!���k0E���rq��Gp�.v]�m0k8t5e��ptub�r����ZmG�����SWVǙ�4���1.��<�A�d���i&�I(p�?}10iXj6L6?��q������Ëo#f�2��6�f�C�E�V���)wt\J2��'�N�´�`iN��2:,k�����]��	�� �&���ͻK5�>X:WA<����Z���F�:��$�oŝ�����x�R��}�m�P��5U4���>�C�M#-ٻ�d�p�^0m$�E�r.�����iJ��_��_8=E<�%ń�Gd�\N6��ʫ<w*M��Û���.1�)P4�1�|ܡ)+{�N+��t(�8X��u�d�xfv+b�����|��l�Ul䚛�C*�U,CX�>��n�Z��3d�qBǜi2��X����9����q���OK'8��5ec�Y�s���M��G�Mh�BD
�3�|1�bE��F��ޡ���J�n�\�'T�٫�:�zbB�eǌ��$��	�X�c�j-.�r(j��f
�P��ED2/��/��a구r9�p�e�ҵ�P�̡��KBi#�'E0(%�?\�u���'0[��Z��4��e�&���.�ͱvM�6Cܩ*uGe�36&YX�x4��d��ǯ�����s�L�L_r���dn��7h���F"]�{��5�s�$ #���ĭs�q���FV�Ժ�3տK��%�XQ�6��:�Tزa��Ņ�o��ݺ���"�c�JI 1�/���>� I܍ �o�6�A��YWAװIC��;�	|�o3)��+���b�f��w���F�Dr'��t��M�JѲ��SQ� Nl+,F
������&��짖\X��+20-Ss���fJ�pR�]��i÷=�{2�׊Y��!I�wjڰ�v���Ԣ�_^S��X%oB�;�uW'P�ݰc׆I�tu�N>s�|֡�g�4��C��L��g�N0TS*A�tRs��-��7�J#�N�+��k>F��O�K��ȏ�#�^-zA˷q*�El����d�����ٲ��H4���]������nU�[��SY�&~�V��C��XG���t�����o��YC�����Gc��H�p�D͙v���{���/]TKI]R� {��hx�(�DШd�sb+����L�L�z�%$��׎��c:{W`fm0��#X&5��)��a�F.�-_���F��z��L�Z�PO�Έ����A.�O�6&{���Z�#epg�d0��}]h]���h���bEa�%�\�>)����pR�KE록�����Y�pG���G8 .!�MoN~��nn*9�|۬�f�N���U�݊�to�\�w*��@k�HC"%ي��<�0X��r[���!3y��n���Ѝ9%'���2��)��6�������z.����	�c��"�้�����8����gYdqg�*�4���;���8r�����e���>�K�3>WD6��#|�Y��31�q�A�Y4��\�3�hhK؈Ѻ'~����<"��g
M�2���:]�R�g�B�ĝ�{��?�עd�u������!KV#�����s��n�f�bv𢬊aڇ�	S�к��s��9`�m�X�gv�З"5phL;c��<1NJ�uG�w=,)r��Xf��C��Kt.S�=�֤�{O��5�&����[����*6��u�Mm]� ���ʵ�:y�����yV���}��JAjc]�>t����(��@2��� /��#��a�0x� C~�6J��!,>�MZ�(�e��,A���])��o/NP����ɨ�b��ߏ��AB9�����gt�n���	G�o�9��]z�M���c�Rr����@#�"�y�5`�
��=T�+͛�$ux R�[��)Yڙ|[E��<�l�x�5�#�`��y�
ť*g	�l_u�c�fІ6����*�3�g��@���M]ޚ�f��\�y���j�l��o��-n0�0�
�d�Q�28Hx��B����@��Sx��DF$�F>qH�ͮwǷF����|I$A���7*������2�K��[ݑ�����m@�\����1Ⱥ�n� ط\#��ס*1����7�}���_ʔ�[����
<�zs�e�� ����^�{���^�.����c�G�����"�lzuH�EW�)Ƶ�2������.��e	���2�R��A���8k�&y��L�k�����N��l��y�'Oh�V�מ��	�>�$Fݲ�JQ̮��XJ>�?�Hi,7���k՚$0JW�D�=#�8��̢��v��j��1��뿓�-�R=��^쯇�$����2SI���U��q��"���.�xȱf���T���<T��W����ȥX4gm1w�x}J�Q�.����5��R��/YyT�0����N5��%�NM�%�ގ5y�r��9f�E`��Eaa��;�'�e>R�n=W
QZ2��m������On�d���e��Ln�wg�Pj�y�I�J���f�:���� Ò�q��5<�n�u�79�EM�CZp����~��f�D�W:�5�^ 8�;T{����"��� ��d5@�����*�s����+w�ڧ�g��X@��t![_H_���Gj���o�陴ִ������
4����e���x9�qƹ�RGa����:L��<E�d���F�#�35=��!�:���s:�9�p�Ϣ��H�_1V5y{<!���,���\�9��aA�J\��
���?s@�L�u��;�;n:]�Em���s�ڗZ,����\��������Y�3d!� �򙷡z�j����>�Pz�!���C��v��R`obޒۘ��Sǒ�*�P�D2PX�t�]�>8	�뮳�ǵp�_&[�2�]I���R'�x�IA.�m*&i�Ӡ�.�
��2�"�r��1�Z �fZ��I�y풭F����^}q��#���+
��D{[.�O9�<�d���̒��� :`[KAU�O=(��I�Mz���l��K���wS��@F"�����櫓+ ֣���]��v�w����i)��A���7����n\Q�Ա�B��Hǫ� ���t'8���zWV�C��-Z�L;�h��A�0��\Е�h=.�Ù�ptZ,!�-48d-�@����=葒��h��1*]P���
���
4#�2%�&輣q3�h�R؊��WS��A���y�2F0�d�j� �g�\� H�P�)s'��Yϸ!յ�����}bHo|=�����?��0���G�j�����ς���H\���Q*}�n�Tk� ����n�O��?ٷ�6�����n�]�' e��ȟ�|�2�Y6f�X��"ɓ������1>�p�,�L�������L���i3����EV`愂ൺ�6|� Ϗ��l� ��% �փ��e�n��99��:���"F�$��U�	/z���s���:��{U_>�?]u@:�݈�e��2jנ��˕l�Aߚ�Ȍ�����n��5T�'?���%��RPx���֜��%E���r��'�H$��DX�g��
��c�b�e��ixR�
z�Ԗ���+��|�Cv~{����Ȋ��N�>��שJ�lu���bq������0�Wa��A���;�|$��Z�_�K�Rz.������D����ʿ�.�	���;�$��j2�a��.��|�"or���	+BW�w5rJ�¼6LDJg�Ж�|�.��`q:�%������u�L�p]=��@�����BB�$L�ޟjx�Y��1��B�/�S��n�I�C�8�?��h������}+�V�x�6��T�t�H���?�Q, T��o.�7��ս&`��g��E%[�"j̖�����eL���~�K��-�9�zQ����4H'����?^(=NϥaI�cb�x_L����W�>�kv�i���È��4]_蛙�.ю��́�,�8�������x̼��}t�]A�� �P<G������'��!���ߓY�uq�Q�s�-^�~\ր)d�� l4Ù��ޟd����9 :�tq�؞���| �{�!J]���9��}ݨǝ4��_�!�q]r��D3�*��}���/���:ώ�?%���)��gٞ������_b�(�W��ۋ��s�Ҥ�P����m:��+!��D��!�����DP/�@>���#IÁ�b�f�X/�G�|����h|�T����?��p�,�Մ3��u�3�J��vi0�'�r�	\,�&�:��".��1c�7Z������ݽ���HxD1��4 ��좦$�}v����	�拼4��Gp��wn�4�~Q�ͥ�L��6�8}�Ãӊ}c�I���_�[�9a��yBV;Վ	s��,Z��km�����T�6�)�v��&�hx��U����u|�����>�U�*y��V��ց��M���,�x�'+����}�y�"ٹO��{��a��7�h��Βˤvf��bDRPyYF����l�9�2�a��e۵�q����Ym�������tȬ��� �9:��~W'(>�KD�sd%e0s����h DJ�Qʛ�{;B��H��~Gb�QנC�O2Smа('؋*�u��������8�w�#A�j��C���+��㈫Ա1m)i�����<	r����4��.
^r�A�a
�z��V�|��3�Un���p�fh=f�7�o��O!t0�+�Y
a;1t]3C�U&X�&�LS��-*%G�[vJ��X*�4��s��b7	c�U~.���O�m�B6z��A��P�4"��jq�:�'|��9��7h�?D<�S���	ۄ��ZC=R �qZ��f�J{V�xhV��=�H �Q��~���g�_,���a=F�iSJ�=�6u�|$A,Vn�c�M��֣rg��%�����x�&S�^W�Ƅ?\�~&���>!��I��T��ld�dtX8$���b�fI� Š
�dȊ�Um�$�!��i����=���26�3?�	���]ڶ�?����D����i�+�l�K_Fw�2ͪ/я^k
�9obR�4��+�	�Ш	�(G�˫�]���.�[W�o u4Щ�Y� ���&{�n��!��z��ɑ�"�Z!��}l���������n�c��ֆ��9�V@~��C�N����ާ�$c���Җ�|_��R��
x�D�����#�ʸ�z^N�)JO��m���t�?�D4�7����7��$c�,���bc�ӂ��������ի���<�.z^�ȗG'�����,p�M(m<gZ�cDn���۔��8�N:��q�c�c�W��3��y���c,�����S�<���J}2���M�f��%�40��͢���m�� �F���&l�y�� �g{�; �T^�E�F+H�H(����g�t��G>�����@���s�e�8E�B�!6,]���/c����w�H�':[�����_�����A���Yp��^G`���ROޔ������wg��K�bFDx��\x���h�3b�M��{*Z�b��O�2�3��,K&=��1ԮL�t���w���5�,��-:A���3B9D��v�<̊�C[����������s
����r[�+
�bE���þNŎ���e*�xY��6ud���,�eMz�­��B�h�<ΎG�<wU"m�+ۊ���?���\���HTv�n�$�2��~W%�J/��l$
&Ul��bҮŽ��%��݁�΍s�����g\�դ�Ou:w@nd�&��6��]��b�����BF�$G����R@�n�ؐ�8����{�	|��)^��Sn��苣�~�Y�4g�ţ*�����q��p�L���>�<�}ٸU����2��4����~/;��\��v�|�,���uB�X�;�:���-���岳nT�vԗ�4ވ��¾�����������(?������[K�����Z�J�[=�\Š�?�����*s�O+L�`E$��B�6�C{�$�,��]��V���l$�Ngi�������Q�d����N�Ъ���;n��8�)��ّ�j~��@���inϟW���V���M��0�\ٷ�ot�A'f
��7�I�i؆e���QZئ�؋�6�q������]v�,s�_%]������7����$��!}��K�c+��<�=��Þ��6ꊠ��5p��h"�8�G�.9�����R�Z*7q��0��� RE�6����n5�"BVis����4�ܵ����L�c\na�_�m�H��p#O}GI�o׬��6��g��m����u��&,�)_X L���L�5;����9�P>�ĭĕlN�(:�M�W���j�N�5��X$�)��^�¹b@�o����*p}(���t��:Y�I�$���2V����@�S����z��8�����',"R�IW�R�.V� e�E���?ܢ-�]��,H��X�rY�
T`����ѹ����!Wu��v����r�73,�\�ߗ�����c��(��׻/�ڹp��,[F��Hf����0����J~7p�伩��*�\\����;0t���vRʸ���Y|����N��O��Ѩ<)e�|�A�h�s���Ğ��'���c�l�)M*�?�� ka[�B	=����[������ 9@?%�p�����R�#��:�`�֡e�p�d�IO�m�j�K�N���N����~}�݌��M���'0�^��0���FΏ~W,{]�z��[�J������;m�@w�s��J)u+G���r��GC9�ā����X�/%Cڂ.��ra� �ϣ�K���"�׉k�0e��G[��ڽ�)�N`�a`�j�tVQxF{��ھ�RH����F�
�}�	i���v�Z־+? �J�t��V�K��Ӡ|��~��k�����2�j���|	��LRZ᧕�ˋ�ʡ+�]�2�Z����&����N��������;�c���Uӻ���!k��L��R#��z	�(�~�#�l��Vk��ly�nH�V�E��M��Jm�1i�CҪ���6�P����mZ]F��p[��aH�����v�m��r�J�K ����*F�g�}�H�x� �3��s��j\�\Z���l	M4ۇ�}:�4�K�u)c+Z�n���X�FU��kS��-f�Wb�v^�c��j��j4=wyg�\�#ц*�^��W����׉a��̧(��%A��\��i�榕ҍ*�w)��
�?x�`�@����M��������X���b�V��#Xz���_�cR\��R������+�iv."O�������G���b
Y*k"fd�֝J1=a�{X<�G
6�pX"0����:�%�n���o�#A�تa�3�Ľ�5+�~�����x'L����q |M�]��䰖�/�����9��	�5(�rqD!�r�4Q|��a���@���L�li:lH��m�������F:�-���;�3)yҪ�R�2CD����^�a�����6S*��� 1�$t�� ���Q�o
ޠ!I��$�$y�JHP�1�U�gDz��t�--~��	o�1:\IĆ6a��1Zbf�琜j�2�*,:��ھ��} Sb�#3���x*_�]���ngh �Q�	�=�İ�s���"�+��K�M���a��z�(�jǑV���E��c�IP����@�6��x,ɭ��I�Z��ȵ��e`�N����!��i*�G��Q"�j>�`KF;��TR�Gs�O�^U�g��NDS"���LC!W�=7דn��E���u����j����
�+��3.�I)b4[S6GA��#q��,τ��T��2Q��7��i]�8���9�2<��jq�'�o�Pٰ sMb�S�F��@��k�]���{t����l����PL��7ɛ��0^Fc,-#���Ԛ�,���m���{�Oh�� ������B^pX�x1 ��$<��!N�5�tǦ T�C�H��D|/�$s?\�Q������_�;_fn�8crCY:�5�@|�O���!����0��1Ҏ=��~e#;�\eܖ	���B����޸�%��2U��\����C�=k4��'!E�?QO���h�'���J.t�)xX�g��h�7'��d���������/�	�a�$��۪�=f/r?��mdv�? ��	
� ��C��L�����#�9���G�yeW���-�E'��� ���6�������~���˽QE}�ݷc	�,4��a����I5l��U�:S�۠%J��
.�'�\��j�ǭ�$:ǅ��α0��e<w�5��o�f�ɗ���}=�����m|�[r^���6
�|�BT����Xs�C�ɷY�=������v|pd�
 �䃮]n�+",�3k�AU<�{�0p�wSI �8�<��~X@R �`��<Z�� ]����Qu����
�ַ3�V�w*ʤi�fP!x���|rN$�.`$e�V���=t0c��1-��{�k��DB4�,0o�je�� ��⇋dG��	U���|A�0��*P�7.���+�]T^4_U�~@�~g)"%����J]}8]�RL�j�)�U�+�Ѕ��L����fc�r�S]C�,z1t��+�`S��3�_şr�)��S�qj Z���'�16no�j�u��3%�3�.s ֧-�F�{ݽFb���цG �Ts*@N�`*m���X�&:1�R���Ɓ�*��Ҳ�|1���@%����/�`�A���`��Pȏ]k�a���D4��t�	qT~C�6�����0�h��¨���+�V�]��Q:׷9�\.�w���IԚp>�׀D9J����4s�{lLj#��s;,��ؔE�GV���I2��!��Ԝ�H1�fn�>�Ŵ�E�p�B��1
/�4N� ��uN�K��,K����-��*U�L�f�
bi��q����ŉTg o�����ŕ5�B�=vHB��A�/���I������QE��8��9��Qb�6
~��A��1a�&�$`�AI��*�Ľ'�׻�1\A��u��#��>��K��D��8�~!\���c*��)9-[?�+mH|8�|u�C�f.m�~p��pj����ZpN�9ꣻr]��3�!�I�5[4!��R�m�X�u�����(_�,9yORz��y����]���z���$��;��e����r�1FP�����t��F��m��}�<qsP�;��@]��AB�+^r���/��;���xo�6�T���5 ���6e�xl�Yd@װI��g����2}�b�����-���G��'|i�/=��7�I�x�cl� y ��N��P5�ɉq������;ep��?�����{�1�~#�qZmK05dX�W�����I"��s�q��+�c���x�!g�7�+<S{�/�@Nʹ˵Ku�H�\�=2� �7ͺը
7 ����dQf2۰�P�j��/u(�W��C��T�Iˁ(�� vm㈴LM������u`DP�Nrբu���q`�����W:S����U]�U�́O�O	xoH�BV������Q�o�^�k��o-O.��.���φ�9f�Hx=gs���j�N��N}��]Z�ҩ�w�s�����������y%mv-E}.ܼ$XL�m�=�)B���c�gTÇb��׊(�S�O�1�[�wcK�-S� �`�c�(m@a�Z�)�^e�꩙EyQ�吧	��5�R���p3��R�����'C2]�D���?GY�ͱ�kC殽���&���w�<�9��6��Ej���5��u�[V+%ktA�u�`P��9�ǵ���2ˌ�p_�ۋ:�`�O`�큈g��{�E�E�k:�-�3G�*B�:�f���.���rk:Ղ��8�?LϾ��K3q��L(�>�i��m�ET��5a�#4�����\�'��Wʵbu��?�p`B����~�zKS��m��A�#���"��~�b^����J�Z�Uc��=��ۃ��c#�S��1D�G�%|N�!�;i@���B+�C ��&#�j�0���
�T��/�CJ�JZ:P�L�ݣ?��FtzlH�m���t��3����։�P�pȞ�Jm�+'�WJ�h�����3��������vp���`��(>m\D������!��]P 4Bn/8��#[�i���}�;�"�Q>��a��Q�A�/�ҭDM��NЅ$��q�-��>\ߴ��Wїr��i�j ��������oDI�^��8�	�/�MJ0Q������G
�4���<�@��xO���������;(����7ۭu�2y!��,�p���	UP�C�]{�e&'�%�^�Ф��@(����C�����c�S豜D���6u\���+;'�d�r
�l�$s=�t���1,�����O�%���d�9Cz�M���Gk�j3r����]�Bxm���ْX�/�]ֵs mx���97����2�iλ�Î:��&iTQ��u�cT�\�N�����1,�i��k�y��?�	</Y9�Ϫnv/}�\���i_D�P�bN�����5�u���78�S#�M������H�����Y	�k(L��[���s��q�x��!72��	B�f���x��ܞq_D�k0?�ο�����\�S6t.J��*�6ȯ��$�9����p�">��s�cN�Oy�<o���S��zP�Һ�����L21v^*x��7]7�h�ۙ}��s�˖���?.,ܔ�Y�X����~��i)o-Tc05R���?�^O(����6[G���)!(�]�w�q�Piǰ@[�ѧN�.+��"�r9%� ��sC��^)�Ļ�V�>-q?��0I�	n���e���lp�M�g���VP��j莟Q-�Sv4�+���n�E~�˄Q�%8��w��֔�s�T�����q�_�m�v�;Q���$}W}�Uu真�i*��'�,X33_bd�?(Rn4u1P#C1m���F��1���mN5A�?�zn!블�l���5%4+ݽ���LE��).� ��B6Yj`Rl���Ov>�,�2L@���>��4����� �-n"ɳ��L����;��M^�x�lz���1��B�y����L��ڹz]��T�N���6�sr�ڴ׍��\J����ٽ��jLSb1��s.dm# ,�&Q8|L^�6DT�����f����� @P蔎�	�d���)j2��J�4�D̹�Uc�kl=��NJ��K`/���]��q!��΅�;���ltq�0MWpr��-7;���jeA���z蔌�f0�~��&K���	W\��]xȡE�>z��c
������FS
#��!2�fiV!w��@�s���&�zp3g�~���p�B ����ȉ�!�C��?@��dw�ݛm�TS��5���9��X�&N��Q���x�>���;1N^�����y��C�a�{Kd]�=U)ZG����k�u�Yn�yJ?CĨ�U�w<46؅]�𫭱�$�hۑ?�$���ƎQ��)�b\��!|���I�U�a|]�XU8ʌ!^9yi?�jл
jX"Ul_!�U�=������?�)N(�]�I�̆�j�J��5�\uZ�R6j��0U�=]�#f�3�Z«�����L�:!��W*����u���H�%%5�\,�1$���`��/�� � ;�(��v�n�dL�����,�ؒ�
2�w�Uؠ#�}u<��gҋt��p��Gv�(�������$1/Z�$5H�(�1ă���UjZ>�:jjc`�-�h��؛��?���r���>���ƙ����Ew�0D;��.�$Bg�o^:F�=Q�F���{cf�L�ߎ�Lă�FcIa2պ1�N���dQ4��A�N�dԪj��C]�N�+]"��J�<1C>Ŕө<cAJi�7�+J�n�SF��¿nÖ�f�q�'.l�(��J�#����W��R;��� �zl�]U��}����^>���J&��*ŤD��y=Z<����C__Xh�0 wkB��+�/:ǰ��O��1��G�����t�щ��So��̍��΢W�:7�q�H��:s?�'2� .�N�wD�s_N�3g��^׉��0Q"P͖�P/��atK� <����
8>�q�ž6�a�d$5+�_�]�?��̯&��J�$?;��_�m�b[�AA�K8����D[IV��:��:��a�KY�G�"�p9x�V����2�9"�(w���f��P��ֿ��\��Tg&�� �]kh;r��8��S���d�B�"L{8�gB������j��}M�~S�C46-a$�3���i,��|R�4��؄�7��#V|�C��u8�Ʌ�}�҂,4�P%G�Ac"6L�́������`&�#�¼`�h�bn��)�Xb�Gd��٫��*Ne1A~1�ӼVC<�âle��g���H}�����Զ!Βb��k(�TYv�����ڦՅ~5��,���v�IK�]���L�?�W�(���$�XN�z����k�R��S�BB��;\ϧ�m!4�`�u+p����h�\�Zo�)�����.��B��~=�n��ȼ=�7���g��eU����&�U\AB�x����8�poc�!�G�;sC�K��s��Hƫ�ɉz����v�M��p>��^(b��bʭ�M�&� �/e�|�o��HqPZ1�ܪr^
�.�Am�W-,�S�pM(��/�=~/d��LY��Z���>�ǢS]~O���wCe���Qȗ]N��0`_�	����fo!� 3�%�_n��f�o���)Voh��3���V��ag��F-�\�<ܼ����:��ʰC!�&��CH&�#0-� �*֦!����&<c�}���2��yP%h�0�ӕS!�	�2U�����Җ%^I�@\�cgIE9&/KotSm:bL�����b�R��Z^s�D��
��W�D؆�"�����>*愗]��3 ���N�AS�f���_�њ�]� �-��_L)�g�g�X��a팄z�ԏ�:��"��"�Eu)��*%��Q��zy}CL�X̪s��h9���te�|Y��%�q}���2~�˦N������_�i��,�V�N��N�b��
�ŭs�%����$ʜ�T�ۥ�l�`����x�t�$�H%�S�yh��˙�^�q+�o�4qV��L��4�2�tC#��Z�̩�9�Q�H����8��Ft8����K��v���j1����r��w���$�"qwLZa&�3��aAdD�T%~)��qqxs�x���¼rVYR��c���߅�zs����|����H��Z\�&h��Z9��4�r )��^���\p4�{��v7�Po��,���"����Ѷ�>��:�D+��Όq�Q�մG^?6�u%FW��ʟCw4X�*�����39NF�-� ��Y�㘍��z=�@��3��m˄��'x�`�V|f{y�.��Sˤ���;�v��ٖ�\�_Ϣ�ީ��O����7���#syl_�V��I&uc~M�ۆ�0�+�N@��g͇V|VA�M0�	%�C*/S�߁x��l�]x=;��ޠ�u��9D��,�W�fj� 4K�1�%�K�c���aOT!A��H�;K�i���_a״��{8a����.��f�����?�����m�뮍Tk�찆Uă�zx��xVǳк��;H�Ǉ���_lB_?�ԑ��:uL�,�~�.(���Sbk0b &:d���=!�cWc�6�l<q�Yb٭I���7y�e+sH�f��jl�����F_5O#gz	��E=��j�$H��n�m�Q��B�YG������[�C�2|;�;P�'�ǭ�o�%��T�O+�g����4�a���:�s"k
�8�{<@*�.��u�(J�=Y:�X��8��T;|S�Qz��GO�n��E�A�U?u43H�Ҹ�W�$@!�a�uMbP�KԈq�"|.=?��W��D�ޔgoJf�q�����rH�s���2+l�(	�C�Z^��6#:�ev�᪟S������o���zЌ��NF��l���, ֠I8���	
z/��64�	��T�,�-�}p���>y����xI�_܊H��yh��;�}1{2��Jc�ܦ�� �����yf�a{x�QR�X(M��]�u��Ln�~�-�/��/Q��ۻt�h��9T�f#�W������+A_�Bj��A4��|D�b��)&��w��&@�&�HD�;[, �!�V���4�q���VX�9�32T��k���m�B�u���M4���ھ�;�@9��~�����+��VF��SP�56����c�ǋfl�w���of�>��!��S��T�!�w\A�Q`����5��L���H+EPx�4��SA���G�����ME�~oZ��ytu�2e'�[BD��	��k�&���N�:��UD��[�=W�0>&=� $SO%:?Wq>]ǣ,�[�߃Ɲ��o��?�i#� 4�9�l.�y��9T�Һ���ש�j�å5Y�\h���4���ݜe\�G���		nOmj��SQ9s6O��3dr��ڴٻ������G�5��nv�2c&h�?3���>�F ��W�|��;�a�	jT�IwE~�� ����+׉�Q=�̙��0b.�O�*Xu�;��uΖ0�3�i�O��U#���.�E�;�p��9��C]�Մ��$L �����GWj%QnL/p2���o6���L�r7h!�
�:q�KؒZ	�a&��\{�^�D�'N�u���K�9�Gk�7�yr]\|�G09]���U��C#�I.����	�j�*H{}�y@�:��{���^wy�t�Ծ�u�Zl!��L�C�i�Z�:yKH�E\r�1��힌�#�����������&�i+�^�J�W,7˓��YԜ�ͅKw%R9Z,�k�����c���"����hR�:�@G��Mi��ݎV
�?v��E�-!�4�"��?���8�.Np��Z	Oj�/�'�y�ƨ�Lh2�莽�@���{��`F1�n%�\n��sI
��ok��2D�K]Ț��[���a-n���9ax���7N���;o��;��u��0��9��!�T�O�@(V	LP^��T�K�R0�7�c��[zv��3"}��Y�#��Q̻�"��T��]��x+te�֭ .ҕ4"����������zCMW
A���V�찟J5³n����"��J]W����}ݲ�`�;P��7T�'���=�+��QЁ��5篃Y�u��) ����f+�|�|8O����w�y���oޖ�1����ö����J<q�|=R��������Hf�Le<�=�t�Yu覺�w�'����ŪO���qTl|����t��V�������?p�z�y6��ރa�GC\D�����ʓ?��F���PFj�}ӻ�k_ ��"����V�������#���9�Ƌ�.쎡���l٥�9����S|�֝G�R�ܨo�֗秎�e�U�����|<�F|��@*2\��j��ZR�
Ţ�'�CZ�^�V{�0�!�Iz���\�Ջ�N�}��%��ޤ�*ֈKwfH[�r9A!� bБ�
���0</멼�p��U��2u��E2����4�ώ�&�`�u��i�^i��X���A	#�4e�+x� g�3\3��z