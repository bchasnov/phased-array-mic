��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf\�|Vv �[h��U+6�6}����b�N����e���`�V���΄r&�Lw�+o m��肱��m<�w?(v��h6��Rz����8M�VX��ЪQ�Jcs��9�p3_��ݣV'XӘ'ٜ#'6�gr���^..�5��9�33��8��~kn�쀩��Tȁ/;�,��T����d���)��*��8��L�|?���m�<�A�o�4X��?�02�6�!�HϨ��F��l�;vHe�񼷆��(V�f�ڌ�W�!"���L�`'{IF���h_[sF<����đ��w�5�Y�U�[�`�o�r�O"�r*����IB$�H��©y.I�����N@j��a��m��?�-�"��r��p�?�~/Xg:�Bq�1�ӓ�n��{^i��q[��Q�+z�b�VY´����Z.L|Z�9>i�3'�<_�{�mhS�-K���a���.#��鉨O�7�Z3�l�iq�+�:/Nx�>�1;���&��6,�n�u3G:F�	c�@�%=�(�}����I\,�9,����m�m�xŞ����1�M_���:r�EG���ë�K��x*����D���.%��N΀���8��	�p���`#$*��u���+��:\QO����_�#Ы��tÖ��nDmJ� ��8TK	�ӎu1�5I�k���R�j��D������԰[e��QU�:t�?��Gx��r�k�e�|���WZ�J����_y=�F�Nc1�u��xg�+���r��	Gn�de9�5wTDKqh�C+Z���"����3����Sn+=��nG݇�E~����O��ݩmcs�&�z��A���U҄���e�a�D�Mү�� �����KNjƣM���S�x5=�N�9��f#���؎u���0.H*6��
u����L��� %	�쨅G���R�r<
��B�G��ڜ|F](u���;!5���0�x����c0w}9檐a��d��n���R��-_��1(�`�G�p�<F��*��˼Ԓ�39�¨v%=+�y�.�$�2���0�}��+iF� 榈L0��D��5XX9SpX���ة@S\z������h����{=�*y"=�xn���+ϳT2Ũ��\���?�M��zO����!۪�͘ed�~2lD�ڃX����!�A���f�
�rpz�4<=�X�W���\)!n�%�RX��V~�F���odn�\b·�i�u�����%x���@�>1�O�L�j6��`��f�Xj�;vM�=}~ 0�i�Qn(	=�M%wx,�; k�n��^u�*Hs�
)u�Q]ʗ�����uMf��C�w`m!�YC)3��-�F��Q�P�� ��Cu�X��Փ.�(~����k(\�۴ u�C� ��%�&쌔��:�:V�:;o�Z�mO�Z�E]�<�Z�\�{JAV�n<{i��>@�j��eo�-;I8��[>�h�ʺ}����|k;�=O9/��%}����pg<�A��vKm(`��PL�IN*^@�����2]��j��Ъ_;h�����ol����LHh�UY�&��Tr���5&�J��bɻ�G���*}O�yD˔]�ƪ(�qCs�qܛ#_�� ?�.�j���ʶ�V'd��_��b.�^l�o���v��G���EؓH�|����88޳�lV3��¿�o�޷Zxq5�P�)�[�V�.���0�b�nOAqL���xms��� �=꩎[��ڎ��0�֗V�}���"u|}�'%�f\T����a��17�2���AUE�Y}*�H~Ȁ9t���_Mt�L��̫,���nQY�Kڋ5�0��/�0_�㿵'��µ:��c�m�l��	D��=�l鋇���ҳ)�`}8��'.�FILc�7UZ�̊X�/:g�ja7��aT�!�5��|�]�־\��"LeХ}�N�^�ˤ�aS�a
1��Yh~�{3="����˅�o��&�Θ�� _bX��	�'��փܸ[{����[���*3�<&���"w���z��B
�8v����o#Ɍ# d�ƭ���e�gTt�*b�<w�����}*ҥ� ��%�Y�ƽ��$z̈����ڎ�1,�!�օ�fIzj�w�m$4�Y`G{a�*��4V�Ӭ�V�m<��|���b��q�ԱX�4^
ݝ�ݨɍ�,��Y�;k#�$�zC�k���)�,�N��� z�ȧ�dنJζ��L��E�@��؛���\�+3�k{;�>ܪ�D�����U������=Xh�!� �2��e�I^����Z�Ru�e3҂ϚR�eu|�?�͚Q�{L��瀐4�?���E�ߠjĐ���^?��~�_F;44H���(:wOʰ����Ñ�v���G�-l�M��[���1�;�ngMAL9�ңC?ܑ(V��zx����^�2�c�b߾�E����k�d��+x1�ǫ��#A��~2�����V�_��c@s-	���ifɔ'��� �����ʐ��ʰ\���2lb�h��g�k>M�0,��p�	�|����|�~c2�c��zg��5C���QNo~~���@������	��!��h *���'����k�i����
����OnT�:�ǅ�I��m�h��Z@Ye}����|<���``\@���ډ"I�t�Ć�:�BA�����Y�أ�LcX,�KX��$�6�
7���.������_~�b�����u��e6��7�7Oˬ������	E��L瞥X`Q y\�q�0��T�G�?ް��}�H��B��Q�������:�W�N�R�w��Z�B�A���e/F{R��B�����}�d�J�4D�Wdh�-�Uj;?ӭɛ|�L�g�ܘ�A�J�vˇx��Y٢�\d�Uf!��~K,9|�՗i�eܘ����m Ŀ�p��a���=�5���ų(ENx}��i�?�D�E��Sͫ�u�G��l˩=�2�8�˿�5iw�p�t��&#��	��7��{e�\@��K�o���ޔX���9�_x����FG��?�~i��41����O�'
U�x�M��yas�x�!�Kߥ�2�`P�TV��

��p��J-�Lk(�e��d��K	��+Snz��5okZ��Z�:$�^�)��w��q��v���a\)M��L݇����A��/���(*@F�I
�$�)���<}��X��>3uh��jp�]T���0��zq�J��na� rʢ;���!J�o�P42vn򳏢9eHt��������_��>�����S��o��6=_U��O��<�j$�(�Q��Z�~����lV?kT3Q<��8A� m��G� Q��D�O������>���SiT��2Jp�,_�m=v�m��S��z�	�TE�]�f {0�n���A��m�f͝x6�QAwvV���ͅyz�I� ��se�@<�c��P�*J=���Tt펡���}f[�~,�'���V�N͚U(�'��V��瑠1�Vڙ�BӍ���Ǿ�Ԫ�(�Y�,�;L�Bf~�8h�вڴ.Yu�Xr��9$�D$��� �#Qa�jyfGX0���ea@��b��#6�I(C;x�
�b����[0:����w�c�~O�E>]��t��9�t��Bb +K-��3SPQ�ٶ}���)�X��� "�D�	��=E�mc �r	L��/u�q��Tv +�_q��|�Q���"����W��Xs�?�1|	u�8��Ӄ=lh�����M	n���K���� ��2�͝L�	�T�7��!�I(�HG���ޗ�	{$�G5]�ح���zZ�����@M�ʔ��)5j��4��r�v�h�G��+�ܝ��1~��,+�FY}_}������P8|�1��p]OW%��f�x��C$k�{��]�΀Ҧ�u�r ��0��;[�HZ<�D!��^nגA�Ɍ љ�������n[2�M�uCz�=�R�?]��
��k�B�������=5Z.��u+i�KҦ%�[�I���A~9��~yJDJ͙7�U7~�o(x~��y����s�(8�$_�ׄ�������_m�+�@��l6_Q\B�҆���d��j��G!�	 v4q�a�yS-c�=P�0矬2/��#?/���������LO�-gtϽ���:�a�@>�����l���D&^j�T�́�rc���@�!w��1ᶓ�-8c�%��B0q�	���$�+{8UMZ��cW��M���Ă�~�s[C�3sF�Z����)>�sw0s�DD��~�%0�����B S_o]?�Y�j+1����)�a���O7
v"l4	��u����my�g��H�}�ۂ'�K9\��-�-�Ƴss�o��_G��0�4@Vք;�ͺ�u||@+/{?2�������*!�\��z�v5�z�.�C�f��{������(cR�K8ot�Ж�Q��tbC�мs�h�&�?��p�3WZqOr�bߛ,�ʴ=�!������A@���f�L4e���uT����Yn���XC:��̭EC��q�\�MU�?�y_�$�=�����z)נl�y��Bp�|�XI$�_���
�$�4���(n=h�<b�?�ʴ��R��C�/;<�]c��r��)���(�o��M�G�=��A�����/�#9��Î�[���&���}X6��D������Y�:�2�O\5�?���)-����A4��3���)QM�Me����G��'�A�#�d���-?�D�����o�����9�X�vD��ǃ��] �Qf�}�bLņ�TzZv����#9�\R��<�Y{�)�9ƘB�ڢ(��7�S��s�A�\%�l}yT2���W�$���Vy<�_�Ўa����F����z�+��c�_�m�GA�w����֩������Ӹ1�5���8#'�v9��{
qB
�"SC��}�t��3g��b�6y�a9�xu���|,J�*���z��8��OKz�p�6���|ڸe�A���H�|Wqn+�?�0�֢$3�Xx<\�t�'�y3La��P�9ɵ/S��M���aG���q�C���{e~�C�S6`��S&�Aш����?S����+`J�����s��	�{��z���������3��fa�5j�8��/yTd���������k ˀ@>
���J�Z�N"��
�9͜AU ��(���(���R��p����YY|`u撄N�m�`� :��ߌp��>f�+�JPT�p{& �8��������F���E�29O�A��P�Էm� z�����1h�j�<��
�5-:�
0*�����L�@ȁ���&Sɇ4{=.��tͺw��88�y��By�%3Jg%'�z�n�gt���f�^����8��?�2�>���]���q_�B� ��-eH�f�<�����QI����p��~4K ����N���p�+ϊ/J+��*�|�7n�K������T�fT�x��*
f�����{	��W�̦�2 ����9[uI��:ĭH��)�K2�Ff/���������NR��#%���\�Q�}���ed��Qn42�&n���Lḍ�G6�����Z-���_��4e�����'-9
y�(��E�]��L��ma$���s�w�Rn�먿#t�}H\u+TtI� N���E��D�9H�b��:^;� ����,Ǎ��;��S��~���Tj[ǖ]C|%1p��5���YN&��.�f��@gq�8�o.^� N�}a� �|o��kj�[����jF�.�ҚO���	@H��7�|�H���~i;`����{�#�})�\ݾ4�1��7s���l\C�qj�,�;sV���_l�3�V$�t��j̣��}/vpΉn��(�ʴ=Z�)z0�rm�V�F�H˽̯Õ�����Pͮ>�nm�8v���
mZ���~z$���e9F��ve�pKR�*�n��A&�1}8݂}|C:J�j1��=-�k�Q��C�� ��K��-5w|�+������{"�J��@��V�C0�s[~*y�B9�6u:���Pߡ�dҏ3LXԳ��t�`^�*L���ͳ�|�X;�Ug0\J���1WX�b�����b�x��R�߇���[yw�r�S���=�"~�!�B���'ݎv`�@B��
<l^����T%:����h���D�}��֎?�v(M>A�HF�C���u���++Ƅt06�G<T�^^/d�x�f�6��߄ԙۍ�����P�J��-���U���X�����<0�K�՟�Unf�g���ˍ��8��;=����쬔���{<���^�o@ѧ@r���}`@�j�'13Ѝە�[HK��`}:��bǟ�]]
e1���5���)7�MH��q^6X�o1����Q?ɍ~.�GxG$m�o�d}��o4&����#]�aJ�Zi��;��F�O4����$�7�$��tA���l��^^�5P��$r�L^�{R���=�y(�.��;��rC�CJ�;Ə8	֤�|�n��t3u3K��?�@i8^,�f��q���LTFT�b;�-�l�NY]]�Y��}ß�i��,vf4�C�~.�Z�:뛶�7�g��.7��ǋ=�=�����W4�h��'c��՛��@��)��V"�#�/�L�6�Ż���I�w�v~no��5[qXu�<J����Ӌit�g4mR�>hk����J��@�S�(7�0�{����u���zy6阮7J�^o�G���#��7G0�|{��Y�y%���+YB �wr���k���6G�&)��E�}�?}<�՚�w�Ь��_��g���:wj���Q=X�~?s�c�@nMX�ä�R�l�ׯ��p�:q^��M��*�{����i1>c��_ C1lVH5� �|) �'�j�=�ʫChM�5�pa
c*���ůn7���Ձ��{�k��V�
r���>�&�����ܴ�}�K�7h�CY~����?6���(����R�8z2N�(4�P"d_���R���P^�F���O�����G�C�YW*1�����5��۩�ӭ�jmOv֊�;I�z ۏὉ��M�#ً��-D���[S��P������7?��XUEH}��� Cz�. �\(!�4��GM���&��O6�	�X?j��d����d�R��}��ϱ*�>���s]v���KN�����)�5�}��,�N����F�+�Ջ6���dW�Idߣ\��ꍑ�ܵ�Ay��Ez
���:���Z;B�f|�7�.�����&��e('��E�Y�e^l�2��y�w	�	�L��j_�Dc��ߚ����O3P*օ�;���$�j������EU�\�i���:�3��(Vc�-�B$�y�@���z�ع)S�?���*}�/mЁ�WPf��õ4!��)*L���S�pZ���;�Y3���R����P@h���7�~�#��C<#B}T�a	�)@(屺���gB����X�����������@��[��=� h��4ؚ�o���sV�?�wV�(XS���_�-�[s�7xv�0��:��O��B;`P��k�K'�Ǘ�:1�ǜ��I��7�Ү�&���V�@��gZ}dz�O���)}�.$���0�Ӣ����&�C�t��H ���}mL��A!�7�%vh��c�$�T��sjx�ɢFn6\��㐔��n�A�^�q�q����үF���O�0��9w_�@�G�Дk.��&cM�f�n�c7L��E5�:ϲkҋ���J��H���g͑b��J�2�bU��<~OqRg����1�D�V�Le�
�=ī
��.�.ua��"p�)2O Bq>�BwY��y��n4��
�Z�xH˥n�ׯ�կ_���F�]-ˢ���(�S!Ԁ}Np����Q~ߙ�K=V�G�6=�q��M{oξ��7h}`�7V�oP��u�ڧ�,�*�T$҈�*��7�RH�Z�M�*�Gl5��+��,�i����^�h�
�XW[�֑�L�㔣h7'�k�xDҧP�1G	a/C�����}k �{]QEx	���r���X�>KE�)�Oq��#0haz��;�0���h71�z��){�Y?�7�~�<-��B���u햽z�y��� H����*���9%$�嫮*р�~�Z��"��1U���Ż��ۛ�:@����̟us9^��$�:� ��Q�Ć��:ɨ�a�B��;�����P��%I�e]-���ݖ�����+���AN;���f{���tr�zS��R$?x���d�+��6'�D�Hsd�����;�H��C^ȳ|U���q�.^[�Lw�=��eua�l��6�^�
���w��2���6M3��WY94�'jT1qٯ�(@���2~�����X�,i��]$��T��>آQ]	�><���ܴ��7ݩ)��_�hYU������vN���r��'w6�E�ε���J�*�Sj 	0��o�#�ǫ���Zh�ֻøN
	����O�4#�f#�3�L�N�Ɏ?��'�,P?0J"�����u��'���PN1�l	�-,t��X���ݞ濮�?����P��Nk?Ь�d�rQZ�3'�p,v��fy������T�nw���k)u�y����@�7�}e��/����'��|5=ٴ �+&���[���{�^�A��S#�9�j�1�\��(�1;�s(Ɨ0�_yY3.6�>c����x�"�:]�N�oZZ�C�O��Z��ꁼ�����Y�]�+��u�7}�{���{��@�	���°��J2}C�pF�/���O�TL�~�j+D���MO!p�A��A�>������,>�\i�9���V��s��`</K�;<�=�����N'��(�<iEM�E��*��je�&��k�֍�\r�f�W�=;s-b������
��e �l��Q��i�*t����h���L%��+u�"�:��z�"u��:�\O�q��-���cez2ȮED8vzM�I�3`���ΜV���Z����{
�k���~��"���&���?|��CµE���hFW[$�;�64�b�3�0~$�w�ʭ<b��@D/:���� Osx!���زuw"lx�08;`�}b�X����.���s7yo�L��]§4m�4�L���U�c�z���M�+��B����)���_�ݔe{�d��I��}^�S����Yc��Ɲ�W<�^g��ct^�Q~��r�H��E�(Y3�j��[v���:�a�C��ˑ�o�}�<l�<�>*��]v�g�APyg/MP�13V/�8���=�j���9�Y����<ʋb@�W�@{"�nU]1�S��]g+	*I�Q̛�#\��39��L#J#�?�E{$>uI���D!�AĮ�U�Ph�`��@�q�0A2�-b$m��^�4&�{�hmwD;��ooq �4i�}�i��aеF�,��bu��p�Г&�㲊`�*��9����ᄓ�����c5�k�oFz"��(4��z��/{b$�-�!��X}^���U�9�湜^��sb�>���^'�zW���;��L"e��{���d]��3���yEg#F6\�Vs`�}H�Ž����;�h�"'��Aj@�c�&Lu��)�O�񹣶�|���)B>u����L
)��[��5�<���wS�
ŒB�Nղ���Q�b`z<d��G���2O��{�]V��'����D3�K�}���ܤ��u�+���gA�G�F���oiJ�'���I*YŮX�j}�3@�-?�/���	�@|�ŧ<�~�"a*��f#��+S9��������.	EM����qW�����Rņe�mֵ`}��M��x� �~�d�	��}y/>	�b�]�
Z	+�˚�{��+lu���i��z�������U��j���ç�I\��(�H4�� z���{&2W2	�4���'�#Kt��1Z������l�e�M�#���#Q�6�G�d��e>?wu�S)�D{2�����-8̨��`�[ƺklX��y�id�Re� iU�ՠ*a�)�?":c�M����ˋ���iA�9�6��_k���!�:�����;�������ń�^�޼c�����n��GOe��ͥ���W����4�V%��F[�g����mH�Z��J��r������Ύ��o ��X���ѭ�g(=�[���mQ�tk��W������x:B��^r��U@r���|�:��F�$N��r��^o�1���v��A7\@\��t���XV�%��=���rE]���F-4������U�9��8���)d>�EH�x)��UA����{΃X�#!�Kaw9ߋi�S@��Ra�d�t����~c�L���0`��I;Jx��D�7TW���T<�8*p){�h�
��y&Z����@���\(H�L)�����m�	Z3]>��8��c�ب�� ��2�o㧇��T���gY� �k~��u�fX�2��߶���e�= �����p�h؉VQ,����,wx���U���W��!+���ox�z;{�h��Ѳy���]U9i������?Cdd��uZu�X\�EԷin�=��S�ٰ�����'��(��l*���ÌG�����l�TAf����wa�D�3��뛳�9���M���]�;����X(uZ�gDd��c�і�b�ߖ�k7I5(8�|Ip�q�.��B_��t%e�����Ku�:=?��:٬���k�u�10�F��(���u"v	|�W$��N3\�Ͼ�sA��A,dS8�%�T���1ʧ_�B�]Ѫ4L��%=�$��@E�o0���,=jJ'�4�N4��/�X���&�C����Q�Х���;3[HU*i�P �[�����A��O��k��N�8G���c�k����Z[R�n֓�������FP� M�z��{�-�����ŲX-�Gl@x�k�i��j+����ݦ��	�kԢu�OrTٱEX:�O
C$���h#�U������5�cQ���}���,|{1���1Ŕ�t���jG9�WL<�U��X5u=����Io|G����[� ��2���qߺ���H���
�vX�O>�����#�x7x��,4Xjx������#'B�p'ze��-m���s綸�����m��@]��MJ8�c����5epG%?��\�w?ED0�$�N!��B�[�8��ә���w�s
bl�g�Um���G�4�)��Eބg���+����r6�Д��d��D��C��v_F(������WG]���?�;q�̆x��Ϛx0(?�D��ц��X,+a8q(IF<���%oH~�.L�U,�pPAݔ�Ţ��Fۚ�&C$�fl�Ń��Jt=�2@?h�Ol���ۊ�hwn�D�D�X��Ȕ�L�R#�'M�E���ǜYN�&*����8�@T��o*;��Qj��l��m�	&d|��"�J����~r�����~äD��z �����O�TI�]�F���Y�Z������qyd����U��qf8�Qj~0��e�[o��y��G\��zqA6{W����\X~�(�`�r�i}�hzU���;�MxT�b��Z-��;u�Ю�@�{h���
��~�Rx;���>�Їl�EA�O+(gOF�wY$�Â�u�e���]�m'!�jz�Eɡ)�²������=���nz�t�W�;ڐ��}aWu
݈�7�ub��T�g�F�|j�
^f�R�ͦ��JP�M��ٯrv4��`�
�-E_���K~�9k�s��I��K5!O�������zOn�Z6���[�
1�ˉIF^���e�7l�����Q�P܀��֗1S���겼I�;AQ��ޚΚ�L�\�d�wǽ;x7�,�.�$�h���,V�%A�#�`_�1Y'z����ޕ$����k���>�HSI|�ڬ�ɟ� 5��Q՗�jލ�:̾U���͆�������%����:��n��4�<����[fv\��S	�R��-$s+R�<���9��r�SD� �����R������ǒ��0�����ǖ��������`�ȳ���v�, �m�'�̄C�-�z�p򣲲��c#OT�!�$�������(n��쒍����sm�47M�~�����a@�s��T��p�p���W��.�>ԙ�
HN��M[��5�d�&A
�!���Roj��N娛��+�!�|�XE|�NG<�F��Bp`x��*��;���{8�,Z�~�-�=���{�xnÀ��nf���T��#��Z�{�m��Sl�j+�<�Λ�����}̩��W"%�ɇ��Ma�Z4/�E�$�I@Q��a����#�D�����\V��ܨSN��^�;f�&V�|\](����$5�˔˜^�I��KfhG$Ǫ�d��
�X�p^�u~�m�<Xy/�PP-�|J/��PkˢW�s��]��e1'�x=1Zk>�ݺ�]�xy����
m�STb[��_8�Y�i[cG6���f�1�-�P��X���PZ�Y�Q{���Q�7�T��{AX �*M�	<�� ��S��v��_wA���
���os�ns/r�<x�6�Znsp���/�H5k@��}{^h2�����US�
-Es8��}*�Gjɠ��Q)�b��!� �]�SI� ��z�.	�X
I������C�tb�����g&$��X�I���&>ml�1�P��0��g�]M�p D�8�#;�E�`f$&�wI��t��Ԩ�CC�u%��C��4�H7�Ph�>�#yJ��1�G�]�<���w̮ h��Rm.Mj�|>�(�B�+�N/���2��CO�S!:YN!�e�R���,�i��9(�U��_.x�}rXmJ�������	E�߅����K:�v#��z�!�=i��Vx��aT=}I��f����l��q�7(���q�w��f3���,����	E�wڱx��
�ȁ	He Φ�!(4�2�D�>�ױ4]8Z�Od�z>ϖ�i�
Z�74ɪ*�g��cՓ��tKq��j�e�8q�gHΉ�?"��m�v"�����6�r�Ex���"S���pd8?jg�4�����)ПoK=lxoX�-�$<3�CM?�(�4*Q�|e�"�zR�qƙye]�/��yw|�����������L���`��UD!k���K.��{�-J2������{2�x�u�|H�e]�w8`I:���	[���6�ҍp�;t�Z)i�چ��gDS4ܗ��B�UoeH�_p�`U����ﷃcIg�Ϟ����'P�g :����yL�l9-B��&1׬�N��j�)E�Okx���j`�����l �(@�?cP���9��'3"_�j����d��H��2z�L��_�_]���
$��x_J�S��BO�CT�[N^$�����R�i�����������x=1��n$��dg�����[��ʍ��Ş���
)Ց���k-������-��,�BѪ�B����j�_"%�@�a���۠0FؕJ��(F�x�J�bNlG�yf!�ʽ�rP�!!f��؁�>�1ڪp:��"J��kU"�~�n쫏EN%9ԏ~�SR)�2��^����Fb��v���W'�æ�4Dg�, _1}]@X���v�T���{2 p��Fg��s�(tkġ�$>���
�~�v�T=��y�nCVk�<�޶���G��#	��.P%F�JG?B:I>\�yj��<��oT��Ef�Ev�� -a���Ib�R�9��RO�԰T��H呏��.�tܬ����ccnt
,ɓ0��W�:�U�M� �^�̥��"i�w	F8t��A�R��W�`�Vd4SLFa(K�;��"l��3�~|��ߨ�rZ����%l��Y5k���fk���?[`��!�|����09������*�b��V�|�?�]ߞ����=>~�)����D���I�
y���=m� ީ���z)���������\�pF��=�����K밭�(K��݌��F�SL�/�$�Yn���JSO_������֢hf\��O��K�aB��7�X���&.j�.�N�Y������)��0n���Q�����L���x|������3>n��7su�g�
mNk��;z���og�p5~����^��I����J�¼���kS��B��U�e�X�I����u�GUn�=F�N�I�\�����x���G�~�$��f�պZ�0'��~���ũ��XA�^&��w]�f���'w]��b�W��Mnk�JA&�]�1�	F-
���E40£Ծ6��[�:B�����=H�}xY��\P.2o��o��^���dg+���D�+�$۫�d�>�<Wy~X"vB�PO��.T�͍{3e�t���������1��$H�Xv��d۲ѧ���'�OB�1[6��K�t�{{Ta'����Vv�a%�b�(�8��5����x��8ʥ���m�R�ؘ�Gt���rK��U.zd����|`0�#%St��;�G�$�XGUi���^8v�AȻ �1�:t������1�����}�`}b�x��k�����M�ڄp��1ʮh2)� D�ô6j?�U,����������rI (��5��}�[�>�Qe�uG�O⎱F�S�%��V˜{��ߜ�qR��!M�*֮t�De�j��cw;fQ�E:�,�W"B�7+���5sW��kwW�����f.H���3?��Bz������WPھ:�[�cW�#�e6��e���_�6{��,yF���}t$�ݦ�A!4���2k�.�=E��7��#���c�#�40�*NlhN�+��G����sK���2��9�WA��sDgP����3zO���35�������@�{щ������"���bS���TWG� C��F�펫'ꓲ�Z�I6i��B_[��Յ����יߦ�-k�U~��s&��:�14�oK�d�GsЛq�����a}��V؊�~�H��xdL���BbD�+��(jx��}����l���������#�w|=�������_������&:��*��ʫ�u<�1��m5�,��q#�#;�skR0�ѐS�	V+�:���o?[��������Y��|�M�̼�TU���n��L2��V}r�;��IZr�\PG�CYqA��QQ0U��e�"خ�L#��"7"$�H�N�;����7�+B�#�y#���\��߭P|>�<v,��W��ln6u�IueWĐz�ebg�R�
�+�}"/�No��gI�M����i)Y��Z<�nT�Tw�ς0��q���%�y�H�T됱+�dFH�a�Kم�������/� -��C;k�_{'oa����>��Lq㦺vk�{Ӧ�٣�O��K�*�_�C昁���39�$/�lg����,*yd)H�m�/%�.�ᘢ�H�� c���d��ҷ Z�yJ�w�L�axܡl�a�4�7�4������8t�JF�s��U��C���Jv�bR]�1��ܝM$J����[�v�q�A隐�:k9B#}Sz@Z�!����uj�?�AZa[�'%ZDÖ~��jv��Y�,)��Mv�bj��������0b\6`��T�1��/3fT�ar�A�H���?*<v}I��
�G�<ַ�����.�m��,*�ߓKG[��'�� ��a�� ��.�BC#M���o�n,���Hm����'�'������>�4�/�m$\%��� Xk���:�OKܻp��}4	K6�9�Yz���+YQ J}����4���i^�e����l=�s� �<��Ro޶P��zI&�7'�)��01%?y�U�O\\�X���󆈒�*�F��.�leK�s�D���D��BB��%���/�z-�-ע$%,�Yb�mn�z��Um;���&&	�<ZU�;�^gIU�6�"{�:a��'���x2��\̿B��G�O���6%�G�*J�2-@T!*K��Ll�S�v�r�?�F���Ե�	2p+"�yV.s.�*o?��/�`�H[Tn�;x����z��8A�Ͻ<g����>�#�l�3x�!ꯍ�B�")��)2�L��p�ȭ�j-��Ś!|
�H�-�;������K�On�7�col��xBb��=..�f�@闣z��
��ʦ���'�_%��:?�r�՚8THQdsm�X���d��H����{�����)I��u���S��\��c9Ȅ~�?w�i2Ӗ	oO�t֋�;�� s�4P�5�Z:n9m�qjP��vL�3��vez2�.g��ec�)h��>g�Vu>%�XH�U�[�~���Ĝ�&���?�� .}6��߻ZӉ@�$K}���XQY��Q�B�x�7DJ
g�
����ޙ5PŰ�)g�1�ƌ p%�ro�8n����k�L���{�a�z&���/����pp/^�etƅ��$jnN���
�(<U���UI����˽�L��L �Y�*J�;�u�u�
։RM%,r__'�]{o"���F��-C#��Bf�\�m�Ƃ�&q7��ʉ��� ��	{��k�5'�VF�P�bI��L�_5Q	�O=i�J����>YB	�<�4�N�1���<Ψϗ���Z�1%�#p��}�ň����?�9�4�ӎ��}����3�oRC�IDx[z�ɞ��&{%�~�$&6�q�\i��9߄S
�/ #����M��;�0C��g� �lڭ��ta���s�۶"g�U���;u+fq�4[\�8:���O��3S�H�D��uj�&W�ݏC��G�>�&��J.q�i�%�E�*�S�� �5��r"��9L�
�]k��~\L�Zc'��B����>B���!F1G"d6�����׫�x^7�n㍂�"�W	n�lں�B�AK�v��,�c�i�������9wLá��9�9Q�%����|�P�N����pչ��
U�l�/�׼b5�X�b�B����E/Qs�!��X�5��ra	�4#�o���{O��Kԧs��9x }�=襷���������W*g����	�3G��ٲ}����Qe(�T���>/�w��yk8:k�wH���}Z� <���N���;��6d�h;H�-c<�����B�h�NFǚU}�
U)����W�+ʋ����h��fA/�Z��)Nc5;C�����@Xb�}��oB�62�W鹱Zޟq>&cW�Ŵ�rJ��(��peL����gG0!%ևl�R,�[�D�S��C�b���!��G*�R����!�(�H"(p'.���9�Ʌ�6әݣ�N�rp��J���[�e�F�B��ԖH���n�u�zy�I��X#:��dY�6T��\�������:�.��?5uRX�?�d���?��!ǅ`;�d~��C�Ȯ�t��O�ӄ�msNX����r�`��_��9��i"YR����Z�,����p!�L̄x�ƋmT<����z�c"�b�#�Ba75喔+�ɪ��n@�w
�j�/�߄�F�����(6� `���eq@��gc�B4��t�R��*�5>�Q��H�48���E��ڥ�c0$�.�Q'��G�}8>��R20/�*��ʦᘷ��Y��Y�H���hF "R��
�w�-ôN�;�y������"�c�H�j��K8 �59Y�Jil�q��D~oi�J#���1��}8T31�����4v�g?[]$gon�#�Kۅ�w��-��8�aͭx��K�:<��/
��w�O&#6�ӻep��k@x��E���Cg��Ժ\�3JB�����g~�{6sc80AJ�sxs}����e����v�,��������2���Fz��R�EajH�Q�&��5�le�>��{8�y�{�P�C��>�p���:`����Bj
kK��]aX�N�o�Na��O1����#7,�]�Q�t�]��HA`�9��{�� -�=kƄ��M���}$����w�2Q��;܉t� ��h����WD�Hi���T�u���7j�S+��~6�A�A)�&�"ua���Gl$:o���-����Q��>>���̸�0 ��o�7�if�6W猖����:x��5~��
�j��F�4���_yѿv�O�ΕE��9����)rXNx	31	�y=��Lu ��ll-�p�Q��÷�<�؍TVܵ�4�Ԡ�K�={�|����B[�~�ӌ�|w��H̽�4���'�R�+�E����1]��V#�](��qn��㐳�U#w#���`��dT?V��������\���i��� ���^P7���o2�J�ف^1_�P0��S��?c�M��T.$t��-��T�D������m�h���Su_��|����"�q�1Hu���D�`KJ�aw]b	�8�	��&Jv;k+�c� ���Ū{rz�a�oK��W[��dJm��Y�;�PEs�W܉�|��
M'�x�Z<�0@��t&��@u���K�-�T,��T��Ԟ9j^��&uՐ>��s�~��rj`k�"��-] ��G�Y��(��[)��"t%f;�+*�됭���	�f��)�����O%w�Kd���i>ux�P��x|�`�5[Wlp�� �tݫ	t�f_�}7[v���<$��'��6��G�ڂ��]�f�� p�$W])᪼ ��K랚%Q��0�q��b�����	Qx5.�|�R��8�E^:(�ņ�ވ�����}I�4^��͒���{Rb&b
���V��8N3p���RKn�?��f\���t烻�/Q.4���H�Q�Rs�go������h@;��^�9��:��fl$"\�6~p}=�
R���L�����I���cq'Ô������è��)7��i�6�� ��ޟ���s������\�c���>�Ă}`�"���o3�aB�DQ`��h���f�?eǾ_�BKWa�S
a'�Rry�8^&$Ze èy��ud"?�Ն#�Z�#-��p_>�}��
�O��ǡjn�k��8k.8��k�Ӹ]�MD1����^����\��ar�(,�ؚ#�m<�X_�����B�N_�K�Y�Hx5�@m}t���h��#Z���XLiG�I��T�({6�b'�I
4�vM\L�Y7r�<5~����w���\��6n���Q�(mL`��1!�nm���M��0��ԕg�pB&�/Xd�"�r��-��5S���� o(n�x���2�o��0�M�s�~ߑIxf� x��kة�I��7�X�����$�Z�`=�<�"V�g��� g��C�Bi�	$�����d���vD�>�f��aSVE"��&���z���RIesT���E�k�O�D~L������6�T*��W�/2g�$E�Y��N2z'�e-�!���@ߡ������2���!�Y�9�k�֘;yv>qh�%���S9?���40"cY��x>�⌥W�Q��,I��z�R��2^���u�x�^��)�S[+l�ZL�B��[2b��I�ֶr��fqo�7����c-MD	m�>�ǿHKm�b����&��KO���̺8-�4k~��sM0۹[@�U���8��8� �k���S�r����\;2���&���t�QS��8l���/� ���|ɢ�[�in�,N.��{>y��j�s����{�bpXj��h����EIc�"��F09&[��-��`qPޑn(/�ƁM
P`��!_A� v�����}���� �r�`mRhm����3�u*���wU�?dI�\�s��V��� !�M�f�_�0Jb�YA���@��%i���2�Ax%ӫbt�Y=���~���3�ި&���mM��Zs� $Dޮ�28b@��9j����]�n���3�?��b ^?Z�t`b�Y�7��j�� j?aF�;k؝!���[��(��ޖ��Z�]QՌ,�`;c��2hԔ�	�k��-�	|��9P��8�+@b>�)�'έʋ,K��4��kq�%��1��svx�d/R�K�ٜ>65s�u;P>^a3��|\?��и�۝]4���j�C�a���#M��_63���\4�.rMY<�^��̖�i۔���n^@���,KB�Z���Ƃ���Ԭm���<�Y��Q'�à#����<�J�&�����;kL&��Q���ހ�3A�˱_�%�'����I�a����ߕ�Qg�3���W�O�k�e��͡ojx�K"����.H��]��F�@s�l�u���ɩ1e��.�(�<ݲǑ�9���J�k}�[@���>���W�H=��}�]w�� �%Ƨ��o���?X��A��/U���|h�d�?y {�*��h�@_I�O��! ���hY�����zw��/%8�%Ɩ+��63�[��e	?�e�'o��8��N� �Z�y����[~;������vh�0�/�g�tU	!-|�KL�	����q+�oƾa��ۣ,�U��y����L��O}%�&�<��!t�e���ϹA˞g�
?˟�!�� �C��=�F9~��#�;�W���X��0k\���������]ih;q��33��{�x�_��u�X)�q�7�oεq7��eoeƙ[��D�7�2�a�Y��4Lo�Q��K��FTd"�Eߥ���[�7��}��ݠK�6I�P������k�iLe���{$t��(���&����8����]��.�ݔ=�I~A�\��9�P�
|�������~|?dي޸�(�On�"h	�@��H����R� ���O�E�S��#︹���h'��5y���wT��%W"i��c�^Ʉ�%`������*�{i�m�v��%�|O����{]bVs^����WHgX����C�����a�ǯ	M=��JB+z�0�:��_w�d��k��rl�GF �봭�����K���%W]?��h/�AH_S�p�Uɮ���P�%���Ȑc�n�����L �����)�:�2�������Bcl�W�?�A��1�_��&�T�ǰh�f��C�X���L�9���U�<y���h����/��Y,:K����'�ٴ5���ŋַ��i�nVr��O��h�+���lbc'���g���g��gY��Vs�:��W)%[����O�~ΘNRxc��!%i�^�w^�!�:��P���fh�B�V���^X�Ҁo.�R�ʵx�{�� ����I�a�ş����.U+��[��Z����U_4�	�#���@ar#�5Q������n�O:�E���A�"l*�~���2����<㋢���{o?�����L�#XU�jH���랮�*�#qq��F�l��a��S�"�>�����l��U�x��Z,'���S�+X��BG�T*���t �����-UeT�B��YS�;5k�!ٺ��Ɵ%����i�����ы�R\e��NI�ʾ�ߔ�q /�5< �����Z3X��uP#P�8[����ʛ��W�e�^ ��df��#�}�l'�uћ�l�_/��FF�>�9�#q�F[���C�����w����L��oT�]{\����U�!4j��{��#�4@�:����N��ݛ���a/hrr�L�}Ї�z�s�6��Qk���t�W�O����W���;D�F�CR�x�أ���.�~���=q��~�8ހL��-�cc)�\�E7��ږCM8�pE<��k96�e�j[�oD'��\��|��x���F�3GF�\eWѺ�},�C���N�׈�(�g��>��4x��	G�F!��\�S�� ��_��$|�-��Q��C"!��� ���#�(��3~��S�ߒ9���2��F9���\��x��g�{��״�A�&��T�*'��+虹��W �q0����Ψ'
i�����;�sS09��U�<�`a�4+C.83���y�O2'�`;j5^�Qd����l�����9e�p����I0�vņ)L��m��h�����������	2��{4� ;-dsV����2�F�ݩ� ���"��j-n�h	&�=��thV�m}�M�xG�aw������jQX�#Sor��Ѧ�ԧ��]K ��7�9�U���"5�N�����[�R���|D�4a]���W�`�$��1����5G��p����v�'q7�б������S����Ž����&�^�Khŋ���p���/�\�6�U|�l���	�n�Pb��T�����z�L�SU��m;Eo5��T	���n�Y`ũ�AQ���Ex}�!�Ƚ���pb7�@f�Է���<�3�VL<��{�T�0-V(���l��e����v���顿�R�.P�ng+�/Q@��ڢf�V s���z��/:�ޖe�S�8Ky8���i�r�R?� �� �lW���X).���S�y����>~l���t\���ˏ�L�O'(_Z%��'
xv.]gΖ�B����u��ȫNjI�~�+Ԣ�5$n���nv3�9W�^�:�4�?<���Ћ�*L�*\y��%#�����~�,0�?�x�3](�D&�EP�2ƴl|F��q�{y7�Ql]��&bT�ĝ�����V��>R%�V�lh����ș����S�D�eH��E�D<_�Y������>i=\�E��z>�k�_�QT��n��֙oE�