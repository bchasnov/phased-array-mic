��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\����q�?��e�I8�b�Ǽ$��"����ׯ1�V0�����A0���ߖ��z��M,�[Tyu��9k���y����xV9�Dy���2s~�^��N�9��ph2i��*�մ��~�p[p1w$���n3��������=�?H}����a̽�I�!�de�#�F�o�D�ɓ�\d�S��~*�[zE�����}��{G-=	j���S���� c:�����OS�mUj.���y�?'��*vf:�p����������[��C~��!	���&���K��������L�� �u&o�\�.��^|�3�T�/4�!����iQ6+P�3g����<Jj���Z<�r�̲�.� �T��3]en��=����y����P���$bwȾ�{�tү�]@~\F���w�
 �f9R��<���%���f1��8<�ʋ %�UsW�&����+6��{&R�����#��ؚ�zH��qV�Y�*�R�����=6i���˃��(ZaS9#čy���� #��EPkB&{�r��hyO��d6X��NtC�g_�c�
d���Nc���)E�\9O@l�L���j�r�A;�+T
0��{F3�r�*��,ˍ�.ew�[��CE��O E�BD�S|�͵<5e����D)��%U��%��+(x��~����,��:5��Dm��Y�9��뼰�C�����^	�%Ｒl�7ip�8ӗU��4�g}^�{ �c@�Bu�ς���Ug�{��a��v@v���g���=���7ݑ )r\39%x��u����^
B�Sl�\<a�$���OF���R2���*�f�
�H�����_����S�ѡ�����8'z	��N�V���	.ӖVE!I��xne���M�vƹ-q2s�oq��� #��y����<� ��mq�:;���cw2��-_@VN�So1�ß��5����
jE*O�헥\Q���]�)+t�f�����(C�Ƈg#hC��B{������:,	���aܣ�~��Lˊ��a��������&���9�/�{������q�����L�n'*.�I��������`&�3b�+�x"�Ik:!r�� ���
NY۝^Ozf��g��� +�
f����=*��q�-��;��uϨ��L�J9���1·�����a�q����9���ڍ8s��L��5�M%��/	'�<j���$(��	��mbq�1ɺr��,�X>��~ TȈ9�����tde$��k�+��s��%G~]۹R�ڊ�U�MCW�" k&��=QX�ᔳ��#<Շ%KJ��P���'�/9Y�!��2
�9���1�;�b�6��sO�Jbr%�^+6W,e=��Kf��N�攈<_��q��o%�?��b�0���p��C- ��۱����F5P�@ߪ�K�����Q�w� zS�5-W�0���$���d�r��B)�����o�7��S��ƌ"o�D�*^�V	 �� �p�=2�D4��5BeP)�eĦ�XJg��6WU�ed�1��!�h��tK� ��V�Y��u�Yx�UN+�؎}�;��W���)h�pD*�Ը�9FM�6�X�h͟��R�|b�u�8�"6D��