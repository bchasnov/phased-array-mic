��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\����q�?��e�I8�b�Ǽ$��"����ׯ1�V0����t	����Ve<��`�4�l)�X
�9W7n����t�1���O�,�� ���e�TFj�"Q5�ڡ���$�R�vV�h�����.P!���ə�{�0�e+��I�c!s�=tX+h7$lA'����-E��x�;����yQ�U�U�cޅ�<?�������r�^���Z��J�� ErL��T��N%�A�F�u,��]�NQ}��4m����V�!c�1~l>)�S�h�oQK��_>�Q���"iT�x����g��	��hS��j�$��.��T���U�`��.L�9Bl~��H��^.i��p,H�,�|���T��tz7��ٙ�T쬪��m����!U�����ʲ�/E;��x���6#��0$�>�����ح����رH��w\��e�6�uIѧ������D�����R��:`D��ۧ�v�e�M!����{ʎ\��|u����P�ᧈ��u\���"���׎�	$F+.H�6��'b����3:�-A~x�ֹ�v䎲�$�������Ԅ���W��A �*�)����	/\'�t�55>�α���și��	�2���_��^��!�yl���G����se`l����}�0mٲ:��΃��7T��<.��4�"8�z}���"I��h%�pݘ���h
��k��̟�!%~�
˕�چ���k�Zk���"���Y��׹���1y�|TB&��n� ʾjN�5��wh�5cĺr���%~�����"y��۔���i�-���1n=m|Ea������EX!�X7_�=L۹Q ��[~ ��K6�tB��S{f]p�3����;�s�5��r��3/x�^�`І�ɳ�M��m�ˏ����!t�����P�+�k:��~ b�/��#�\G>���g��V����]�#k�#DK��yx%��{�����{���r9�������y�N��K�pHr��v�i���� �h�P�R�eUmR�j��x;3Q6�ҍNl6qU`RxWMr^���wv�n�}[�L�l�c »1=�Ð���}mxnTa�J;2�`�`c�V�؇>�����_،��Fo���*6EЅ�-��y[�_!�H<i[���]Q�J�.�װ����?!$���:X�q��=.�%CЁ�D;��OFE�����Ԟ[+@����yv�����LN�v1�u,�
a	NB��0p�-/�?�u^1���㈌��Ǡٷ��j�{�_��a*��걀�+�p6Cå?i>H����*�6[�褏g�b��=*����V����Oʻ���_�F������6E)��R�>%ñ�q�/V�p�	�w���a��>�"~I�u�4�z0.Z�0�$(x[�Qu����m�(�/�,RF)iJ�M|��ie����_,T.�ўK����Fˀ��e�yHGTk����kBa�`Ȧ); �M��I2cvE�#�mp��2c��o�tY	4�D�2�tH�=�I5�B��D�����)u�/Q�:��!�8������]|Y.�WƑ��[�a�&����e��s�Y��ߐV�c���j�{ ���\C�凥�R/j׍�[	�4/�]⺻qs��z*LJ����|x�py�.�^,!�.˦ť����pB�jkZ���v!��4���L��Bu���ҁy�:�>��@���1�\/Ȅm8�w"��l�^7awr��.`��׃�˴�q׷>�H�1��{{�z��ur����Ь�ӧ]-����c�,���716�F�E�������m|_�\s�Ŵ�vF���|���t���Q��m�+ĕ�~`�c���J����
�s�J��[��A�����T0,oW�M��f~��V��d������7
2���O��GUҴ��YZ%Nk�d��f�7����	�yF����-��lkZ܀C��^�J�\][��U���:[��{m��p�T����<�I�U]F8"�jb��hx�k�MĔ���<��U)utT^h���%7�\�}������J3X(��d'�軾�����[��1��,�*q�ŠN1�v����^W��?8U}�������P��	(^�?��C��k+�l�V�}��@�1�H��!�c2�_I8�V��%�͉C�k�vS�!�c�����Y�{�
�#2�R�3�g�`��BO��/�����1�-+ ���'?��'�n[E,`�0j�rg�p:g�\��I;i^05f��*��+���e�"g�Q��yb6;��u .D�k�I�ڧXQs���o������p��D���Y��
���7EZh��4#�vܶ����5��*�|���Aq7;����H`zdϢ��=�h.��mq���� ;�ql��iFv\s��]jz�7�}
��YNBʑF$W9.[��]�\CL�҄٧�m��/�n"��p��8��m��NUu�� 0��`���, f�`x��iҫ}J�7� ��w��.U�nX,��ag�v�q��hz���gv�<����㾏UV����7�?�{�p�}�>�f9��KE����<1���X0�΅���n�/L'�w�i��)�G�����S�@n�ӵ�`�a��7�}4E�Z$/�q��4��f���}���46Cd��FL�����^�3�zK2ͣ�ŭg��W|��lQSn��P���D׋Um�������8"^�b�a[��d�J�=�Ez'?6��,�<ؐ6#Ci"j��#�A��򪴇/�@z�D��j.�2�w
o5�"-	��UW9���@�Vo��e�v�'h���k��<�QĿ�nEW(:��<�����DW���c��kF�4�t��j���_�����q�9�������ue�y_�:�f�j1���p���k�9ChQ==�[�2 5H�ᑃl��w����9J�=H�rboנV�i����_�H��値�@}���Y܇ǹf���|L�Ђ����"ͬo���������+��^�S�յdx�\FT0��oUN�#�	NQ5.u�73sBI�V$�����p��6��{��"���I0�*y��O^]PD��<�� �ʏ��D_���I�t�9z��"���6m/Ԗ=�T[����K�dڦOS�-1��#�s�8Q)�1���2�V�VJ�"hź�U�ar���η1zV�y�:t�z�X ����8{���rP��܄uXh���k���"0٪��!����mIK�wZ��9G�2w�PB�x�-��<zp��߁�9Q���Z=��pu�?�{����	��<Cl��-���9�U�n�z������]y�V�Kxv����;��mG7�Q����V��׏�ZV!�uL:Lr��2�1��cP #��]�js+B����^�ei��h��l��c��ؐ�� b��s��݁er5�CS��-E1]q(��U��6���m�*�qq��oN�8�2*�T�M	�>�zt�p�5�8-��9�"�G�y>�Y�ݭC&��R�MX���Փ�n��^s�S@�SJ��r��º�GP�!D�)��E�	�nĔ4|ڄ{����'E��|$�ӐT�Hfi�Q�w�d%�6V�ɧ��G��S�[�D��67�J�F�v����/gb�=��ʳ���7����
.�q�Z��0�W��ˢ���L��ϥr�h��pv{KO��9z	�}_x":�ԋ���j�,NIJ�捫�Q�����*��^�(�,���ı��$`��;�,ү߷o4_�����T��]>�J�O,�ۿ3�o]�0%,2$��?�|Q�lu�Lv�#��!/l"�����nV�^8���ŋZ*��1�d���įq�H�-��8c��\���򲉺�1���z;��' �HT�� �\�>d�����WW���T�F]865� �4�DQEÔvU��`:Z��3�k�ڊf�DBU���6������q�A�[�P�=KLO1U����$I$����h�_�Ӱ,M\��ʢ��Z�`Y� {�3��BRA�Y�־�O��otJ��V�u��*JiRfw`��x�~(ٛ�LjJ0�1�=�=�Ko��[����P���:����Y��`'�T�8L� ��x��q#��W4M�+D���0��MÚÕ�֢O�O��v|ޯ�1�yы ��� ����)U;�T.�n%�7!�.���{�`@F�L^,XC`ˏ��kU���b䡼=c ��;hPj2�]��p�7�N�w�PW���⠳�J����w��k\M{���'����Mj;[*�/z1�9�gĚ����'3�ӡ��0�,��������w'���-Pӓ��<5�ꌠ^f����ۿR��{�t�{�eh�l�,�,'��2�&��d��y�d�Զ�]�Ku(����Xr\ܟ�e�*�~~�&D��=Q��������H�
����^_�tVӐ��r��&<���By%=k� FG���s����H�B�|{�	��\yM���wh��rt�mN�L3l��G�ٍ���jq�YX�4^+J�DP�g��6����3��0�������)�c�X����c>
�Ǚ226id��_�K�7���_qk���Q$���a�Cc�Wψ�b�Q���u�Dc�(�?�S��'�o�ٚ'B��G���EJԴuO�#xRc���C"��a�'�yr�%��(���S��k��r�:Q��a�V�;�P�Pb*�_>paL�m�Xx�,1�b
F�6�O�c��V� 4�_�+�Kјm��J��r4��3�rS�� v"���߸��	�i;8����&:���4p$��W����^G��Æ�K����#����Ө�!x�!�u�[����n�}�7��'_q�Fp 	%���l� Y	kb|��qT9q��$������箸���ͫ&�ɪmIG�8Ӗ��T��vC2�n艤	:��w��_M~]t3������,j�Ah�R��2!�"�u�
D�(}���`bT'�� ��>d���
i�t*��
�J���P��E�A�~3L�H�Ho�5�=��%���G�m1n��sq��g��V�Eh�w�@P#F&+ӵ��E��aJ)t�%��U��R���3�-�U�����( ��$nQw�o���"ۀUe�g��"��NÈ��h�: �"�UHEZ5@�I�R"{�v�3�B���]��>1j����~T��]��C��v18w�;X��<��eg�E$�Ə�����m!;C���0(���W���]�`�1#N`�w�AHAFd_�lL��W=�p�[��O�;]��5q�-��� �&K�N��+}�P�}ְKL�D<�[�")i�|���?]\�ێ�mX�O��(u;W4�}�O�R���QZ��l$t��i*6J��	lz8,�v�=PU�d����c'8�a��1�3O�,��)�c]��f�ق�f��|��[�l�qT��J�d�H������=HgEؒT�B�@^�X�}���t'���?��������Q�X_+���5�mJ���Ё�~�V� ����$�5�����V�m%��܄��{�1zZ��F����!�!�
Đ�U<�<
�
,���u�;��l�Wq!�8��?��q$�k�@ܜ��a���7��"����SŜj��m�тxt�[��ͦc�l�@��6�$�� �䂎�(�K;�X���%���mF�8����&�7,�m;����q��tf�i�v_㓍�^!��h!��}s�aB�uk�z%���o(��%�bܩ���$ے�Z?��ߍJtgy&����m��7��e�,jD�0����6A�1��L������WgDL�!��} ��+Wz~4S/����d��m�+�)(�z�.�)j��|U�$%��V�@�&�0F�]�T܂�uRMν�C��F^��8�KO�~�׀�,V�3N���p���.
� �3���11�ya��t@oѺ�m��E��Ik�8ݣ}W7$e��S��ES�v