��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\����q�?��e�I8�b�Ǽ$��"����ׯ1�V0���R�q�#zf���l%J��l�����&qaݏ( )7� ~��ė�*����}�E��-GD����f>B�";�.�z��|�)����s!��a��ǒ8���W�	�br�_�t׮�ǔ�8�3�ޢ�1����Ģ}r���@����G��DC�6Mmi�*|��Ͻ�_�Pl�50T���c��ż�m�`��M[����:��I%�k����P��_��Ы��B�"�<�#���_6��{DN��T%���=��P�e<��=�$u��:Q�$%b�<3^�����gW-�����U���_�����)���ec�E��b��cT$���a�Z[������t'xn��i��/",81�\�q�)W�h2���=rf��E�t�I�w���x���D0�E({�xvf��J=e���1�qnk�p<M5�1a���g"V]�=quW��=B;��0�v�ٹ��,���X�708!�Cl[
#U��C�n��Yn�d�<˒�������t�媒��>N���D�>�fr_9C?ͨT�E2�0w�Ui@�U4{?���g��!<߮L�� �Z�|
o�_���BY; Z������:�*���M-�#r.�I��Ĕr>�6(�� ��J%�:��N~|��6]�J�)�4��p����%j��g1��G��p&_�p�`��!�*ss� �*"~��i��٦)���/iM��O-nrkg�Â����	�5�wt2;S�l�j�o8�[�d�:�$y݊p$�7i�ո�D��Uz�
� �x�h�������ٙȋ%&,��^BYH�rN�J���	1�IW����� �O���~,(��:��r;���ES�)|G��YH�L�a�����+sE�Ue��0xp���(�$��)�����q��*�jnn���\�z��B�V���������
�@�>�7I�-�#�?ף��u@ҹ��"�m��|p�FC�a���9�p9��͎x �R��(��4;K��H���2?؝���f����*�F��敥T��bQ�eF��M���|�b˿�O�ȿ ��3��'w�E�-�E��� z���3�2ZF�]�����x3�6$T�W� ��G���)}zǦ�7�i}K��N!�_d��d��E����9Φ���פ�O�͉�b99Xa�lIɇ���0Ĕi��ܝ��7�T|V��kg��!�\�!i
�=J��
��0p��,��n��2H�����$mӓC�AZ&�A�L�%�C���0�Y�o�?��D?Z���<N��ǝ�o��@�f�b��Ȳ�!rǮc�tm��,d�Y����=%	a��*��47��!�O00��Pl.m}�5��v�?�rG"S�`ú��L:$8�B���aOo��٭c]hi����?�>�.�\R��tw��[d�i�,M��z��&�2��Kdû��>B�DWb�_�eU����n^��Y0�N,!�Ju���vg��( ;Ś)h�$�Y�R��F�V�mK �К�[B��+�CV�����8�Nޫ�S�z;�ɲ�M�(Ÿ<�ʿ���'�^��9 ���[=����sg�}x�pA$C_!Jnj	���?#��l�i�1�h;�|r9�(<��z�ײ��h�Oÿ!G�V�>�ݻ`��[����M~VAڋ�㽘�qyL!/�}�ݫ��l��I��\��z��ƥ�s�s��ӌ;�Y�w����Oԋ#݊�|Xg�O!��r���u��YkY�rCq'y! �d�4~��Q��?�S��_�C��	1O 6��~
�U[�~&��.lY�xA�r<.q��1�<AT)}
�_�Qd*�q[�q��� �n��ls�=u�2]�4w�@F0��ͺ�����s2�/��h8Ta�����B�*��o����VR ��� �Z:�0�K� �I��ksKo�䊆��,�|��f_6��gs�Ƅ�mg��ɵq�w܃�����S����K�ns$��QsB�� \�����R�SpK�ؒV������g/��0 �+>``R,{� ��#N:���>��ԗ}���ZN8����P��{�K#!-�פܟE������b*���Ζ�Vܖ�~Nxw���1�]��;�uo�L
���1���l T�T�*��K>(���~Ѽض����ե �mv���h�V1"��x�)<o�x`%i(}�� ���Xش��
,|Alm�=��߆�P�ɣ�x�� n#����P�({Ë����S���-�jZ��}"4f����I�B�����i�\��e���t��y�(�qxo�?�y`{"��`h�g���0�n[y�yi���HΓ]�ß�놌ӟ��A�(��m�e��Hr�a�P�V��W4ߨQTt^|�Z���}7��A�sJG���[v������?i���r�+Qʂ�O���j�JQ��OQ�-O�B��J�d+��vh�d6-��+�=*H;�[���i�3���B����侃F/����|� ǭ.n#��|1�t���_{3���Go����}K9ȓ2��K+�D�γK7�Q� (K�>Uƙ�2�:�A&!�`�iO�g���fk��d���Q��J���=�E���\X����n�êì1���c��Һ�u��~�/���
XOQƄMg��?)G�:���I��CS|�ɶ-���������D�/�Eu]��+Xk�Zh���0 �d�Ӓ)���D���tI�V{��n�<)�}C�我��-��D����zQ�eI����Dl� `�K����mל�w
^��KBg0{�\������#-���Z�%����X_�+�:_>�&�4oj��X*�Y�HW�(�̳�N����W�4C�S�}v��\�[XWۥ����o#fQ,�?<"F��V��L����m���~x>�����
?����	�=?�-.j\i-��I�^��{��":����W�?gR����A[`�-��Ayd�m��1Jݞre�yT�6��?̛��= �ӥ���k��T�S��@��M��)9�*�>�p^�W����Q�{ְ����ۿ�3��T5*��W2�<���� ����ғ���c䉤��gp���=�ޗ�0�!M�ͼ�H����r�d�,�n�s�e�!G��=�ۛ�����Y�u%��&���R �.���-L9�6"�2�"��o��4��7���3F��;��cؘ�~5�#����*O2B���'��!b>34�i����#�#r�iٝ
2م��M�@�` �����0Ӱr\�C������Ѿ��2�Y���X�����\ߦ�qj��l�K��h�-V����h��U�����F�{�T����Io�����M�ķ��%P%�C|*�WPL�*�L�='R+f!��д�ClqΌqwD��<�&�@��<�@�t��)��$��'D�ݬE���a���|�y�Gz	�`>���n�	$��#��$<P��n����{�����KJ��M�xO����G��"��m4�n���X��2M��D������{�%���U5�&�Y�� $!�A�u����g���Ugdq��HB*�e1 [��.���W�K9����j,m�ik}]b�>PH�(��}�1���ϐ%��k��W��d�@�qU���`�?G�,���Ya~=�pL�3����'&z[
�<���� ��O��A?̠�^p�g�_ ���*����U��c^��K�ayp3��ŋh�
D�u��K��)�����ĵ��M�f�ү�^�qO.&����T1�;q6���l6RAt�C���㮬�
��f�44V�b�!:���AB���T�J�f �8*il@~O�Uu�6l�;�W�g/�k��Փ{�&M�!L(t�%�.j߶���	�D�dm�������z�:�H��?���~�1aC��a�E�[X���˔SW��ܹ7���[�K3!;����dQ��!gC���R5D����OR�0dt��T�fڂ)?g5x����9�$��xVJ�b4�����E�����J�R�0���Yr�),cu=���6��9�5b+ø����1�5p��9\9�xcơe����`DS�悆a��v�:k½���N��Ej�h��<�v�]��A'�{/uq�F�J�\��M?Ĭi�i�����Sjs�q��������M�b|��Y8@�eg�A0#%���w}�x7� �AL��͒Ԇ�,���I���{z�ƙ���X�Ok�Upto�:�����Q�2QC=�%�ӼV 0�aB�?9-i�A�ػ���X�Z��r��4�"�t��� "�y��ܩ��J��r��iL��j�5hN^`̱��m�7 -l�qx� �7֓��>�����P{��WNz6s��=`V(�K�	aҦg�ޞ��[����~�K�jԢM�'^M;9���"�Ͼ}g���Ͼ��3��z�P���lbP�����軇y�Ɩ�֚K�ф��D����^p�YlQdf�����5u@R��k�5dd���G�W��È�DufW��\�h6�4�5^���B�?h��\���s�;�P1�Z���X�5�_%����)��?��c	�׸N���_xpb���
�u��H��'=;�y��a�[\emn&<���وxҽ߁Ȯ]��Gp�h�������"Y�^93l.�|96] 6
m�CL��Cf���˸�s���T�WK�\���d�����k���;er�C�ѯh3����r�a�ŀ2��W�U��*F?@�F!�r�~m�_
�1�.�	i�-��Q�O�.B���\5��_m�{~�R�g��r��� �՛�g�����8ͤLj�āf����Y�,HW<��w1�)w��r���4m��XO�����!� ��k~���lO'���Sݭ�����yۡ4���e�4Ȱ�+��v��Rҳd�b}v�'���]��#k��>r�F�N�B����*v��GD;��P:�l�?>Bo�y�.��P�}ka;Q����Oy,�jv�\�3���eZ�7R���^z��<�l�?	O:�\\�"?�br��Gq;Y��q0���9���^֐~�^�=	�Ē`�6oJ�t�����|�Ėl�	b=�	�[A�PT�������h�Y�����s�'4�w�Ŝ��?�����:����M���B�f��V-�g�ǅ��M�������ٹj�A�	�$-�;��p�_=��F�8nQ��ݷ�����E[�D��miy�|�}fmA��}'-K���i�%E}'.5<#���7�޹�^�Ug��K��"+�۳�#����G���37i�O��W��rg���Q�os���%�,���p��B�*g��:(����Y���#B{A�tw=�(rTS�5嶵�'_ 2����*��=�r�v������X�m4X��-~L/}uآlsP�X̧�XP�[����T���U��p烛�O"��P+�[���W�=����C ���D�N:��Ř�A~�&������yM)��c�^�����{'����wU�����4%�`�ņr=�OͲ=��h�{���J�u�B�[��QB�.�\�g_��<8��׭���U4�PUrQ/"��
�^	��S��h�܆ŸȠ\��1��\��4SE��(����]r\�"�0��s?:|<�7�ʐl9$�G��f�sFE���]��n8�r�����6<Ŝ�t�G��' �\Xke��d �M����sp����	�Ö> ��O�D�>1'���g�i�ֵ�� h�g��^%+a{��h?h��a.�vG7�X~�\Ц��}�atK��oP��,5���X��-�Pd#P/z	D׭h�t����MD�.,j�7���Ŧ�l��C���,��o]�Ŋ�2�?btxQ���(��������̐=Rub5)�/�k���N�ߣ��!&��s����7����Y{P�������&��]�t����=��s:�
1���c<�J�u�����"��_�i|�$����I>�8,V ڔ ?����/�*��*rBK�X���Yp���,!������l|t�[Ӊ��{��Fe�=����/j�
�BZm��4��`�6���g�m���ە�X�>Z^ˈ)��; j��ӟ�_������e�$D}�(��^H�#s���d��!�������4#���ͷ�$+{e*��,~����3���?�=����/�����
�0O��X��bD��p��VC���';ܘ�b���Q#<<lU�����b6[���M�T̩�	��+�3U���D��[��`4s(Q:1� ��kI�$���&%5� �0�a�Ķ�F�#0zGS�����>g�c���rm]D�N� [2랸חL���璪|(��������I���1��
f����{�SؠU����k�W�=+��s�h���1�J�z����4lF��l�h����|�(����H�z����j̲��"G��ÚiH����M�2 �{IPt������ɤ���!#F��p����w�4	���6j+M~�q�������<�}5���ă���N��6D@K0��f��g�W �^N4^Z�M�R��
�e�X��g�= Zq޾U&�Xx4vvbxk�e�B�]G<�]�j��
�M�m��8�/�'@Ǐ�]��� ���T�.���n��r[��[1An��t��Ig	<�n��j"�0`Ym��W�_�����ƕ��o5�`�NC{R��jӓ�,�2�3����e�ϗN@%�a7�N���Ob��f^gֳ�,ŷyv~����"�P�u�Ϩ�Ӵ�y�y����Dg�q�������c��?���u	q2�l_,+Zg1E��o4�����ة����b'�����F/����5G ���Ȱ��q��d~��; ��z��$��+�5ToCݒ]�Y�ra�����❀��;0;,�N<0@�R&�Tc`7���\���477� ٻ
Kîĉ~@�J�-~qǶ�qi�����5�2����J1����A����P���{�����w1�b�(+
�-�+�ь�&�-�%!� F!� ^f>��F����l!��V<L�3�###��_��N�:j̣��}߲Au7��u༇)�
�`rͼ&���_h_���T�W������BA��H���9C6,Q�YE��H�M��,
�L2�����'r��?��p��������lm�����{iB��&L2���;�U�W��=j�g�����7�KȢ���\�	9�����,���c�Q�,] |؂�5�q���@��*M�;,��*�D�~���bf��IH'8(�������LL���0̣�?Q0�͒�_	m�ו��
(��rh���K�nf�����j$8��v�y")Ӱ���T[ԾEJ����[�i��$�w��_��TH���W�\m��;�����I���U�a�2��T�E�����E�!~�6`�az�ڇ���`p�y�6����~Ŵ���߃�҉�ros��.��G)#ͬ%[��}	��,���/�u�t[�z�9�T�("�l�ڜ���f���*��[��j�C-G������gP���ٓ��m�����]EJQ��{F4����Z��J"#8v� r���ar�8�S8�>��'Sp�m��}��6�,(׀Tq5-`�&��B��D�����o�[뚻p㦯��]S��W��[�O��]���3y��Wou�yGqe2e>�6�.^0ǖ��m6Hi���N�c�K����p���p�.�G?��c�Ǆ��b��^�+��ۅ4���#B5�p�ʲL�A �����9[jZ� 9M��^�	��ݾx���cGR6Յs.����$!�B�}�ǘ(�1>]��Bǋ�;�`�(�[��JĊ��^�4Ⱥ�o&~�]M��I�
�i��."sx[�1�$^l.N�E��h:yZژ�2�Ň�����uf��KḤ_�gm͟|*뷯(B�I[��?O��n�Y�:H>_���K�d���J�zd�[������?W;�ܙ8:e��d~#���^I��{c����&@t��8��gI�HrJW�6pK[�(�z�2�!�
��p"/�Uz�R�e�FFE&�웲=iyFk���@MB/#�R���P�~��8��G�����0��~�����XL ��DR�m�(!r��d-��8`׶wZ��;�ocen$��B(-"���R���{���X�Y��Ğ؃i����P�O��-��ߋc!���ζ���U�<9􏉾�hK��O�=-3�lj�phV�[�GWt��o$`|�a��V�ͨ��?���G���6(@�4��#?Ư:�Xj��0Ӫ���;�8����oN�V9r���ah&���HiH�=�b� �8������PR�۹�ֹ[�<?.�)��J���,�?sС���6|U��j����er�D��q��{+�#�>�kmO	����$�|��@E���s�\Ӏu�Y$�^p�}��Ե<��s<H���v�U�2�]m��S�M���n�m��0ӰZx{�9��G";�^i�!6�Sz���}%��#�ˤ��^[�Si�lTaH�y2-��*���w�^��c�mO�<�����k1����>!��E_�H{Tׂ�g��
F,�[Vg�(툞�$:�X��J��撍��ӈج��g���0p�W`�DC�}��Й�F[&�;ȉ`f�r��ꭓ~�� �Bn�K2�*W��4kt{0��?�ݱ������ũB��J�˩�K�5�3�I�y�{4�MR�9
��W��/�Wi_�c�b��cC��
%�X^O(�n>H�50&��� .Pm��P$d��C"���j#�����$���a^{V~�n"5�I�`T�P;���Xߗɀ=P�&CY�D16W�R��iی�ȭ�eH⿈R���zn(����:�Ń��|	�8���DX�ß�E8�F��� .b�7I	�N����t��k���6�1��&'�	
��[a�M�^}s w_��l���S����]�`V�9\�z�bJD���{�J/I��5��f=�ٽQ�[�)o���z���|��)��-���y�}�!Ԕlf��ٻf�G�