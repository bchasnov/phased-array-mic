��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�k�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������H�W޵α���N-�`��6����ݾ�FF��eF4��_}<�ےA�[,�|{�?r+-��]n?���A��#��Hb�а~�g����o�+5FL�cu�ȗ$��ƃdY=�7X�aH"��;�������cJ�������w3�ҟwTʡO1�Ur�C0����d�X�8z��rJ��w2����L��Ä���>9Ħ)��)b`�Em�(�q5�
�j�.eþ6?��x>qQ�g7�g����F��f������:����4��F �AN�<��K+�'>�m��%��B�rd��`��c�5=�4�D��!��B/Z��c�x9�D!M�o���"�&�/� ȫ���W�\�EU�fM͟1J�Au��Y����?���F����j�n�!�(�ԡa�I2�ڍ��{G�>"d%�賊�K&�2��M�5���S��/O��9����̦D��w��&��3��>��K%����\���(�'L'�m��l���q%��0��Sj/�?P�t��҉W�&Y.4):z�i�ب6��Π�l����JH}`��0������G�o�d�<�@�;���]Uͧ0��8-)�F��dTD�����j�p����Hg��|�yńh��� w�\U�ͻ�z��t���"�@���ԑy)�^<X��g���QOBKZ\���T3�ϫ���➲ ��=��!r�{s����"LF�$7�R�D����?B5����t�w"3�^�\u3/ߑ�@���E��X��kd�Pϑ���<*��dO�g�c$+9��څ��I��d,?z�Bw�¥���Fj�(5�v�ka�U쇦��i�lbrx�j�0�7����.�PMS�Ҫ�ȴvn��4V�������l�At�B۷׊5�Nr+cï��������T��=Lh�F&l�j��[�Za�-1*���ǣt��{���3�  ƬY�����jm��Kߜ�׊J�ae��c�(����q# �2����	��&�h0��b���^�1Gm�&Ub,�p�V���v�$�VF?�� �2R��\���eO�5�cP��U�:c�8о����9�4��C~�cH9�!�Bg�se�k�o-z�&ݰ�6�$8M��%"�v�h�.��1j2�<$��T���-xY�?(���U	�i�eվ4���6�/E��ATZ@�:�T�Wm�����	�8s�#pp��1K/P5[�!J�M�}D?D�F��|B�}OF�F5WӃZv���w���8*�2���=�&%G��gJ_7�f�<\������ί���ޥzmGz^�V��\�Z5�}���L�V�kV��0.�E�NA�Qʁ��լq��߇�:htM���O��(Vw��+aE��-���sd��G���^hf-d�[�S��I I#<���j��>��JE(�d6���~x����u@I�U�p�pT��`@#��k�/c����U.M�������������S������ϰ�Jz7�鱕�������`���É�$�5�+a��Ag=YD�q�v�|1�̬
�4s�Y��Ԋ��Ոl##���p��( 5�BZ�q\rp.��As�(]ˏ_)w3L"�({��t𣑅=��P�U� v�7��е;��߬ �^�Y�FH��!���'�����T��TM�y�q<�+����_�2:N���v�'�3
5����`�Ż�~��e��Ȼ���P�����y�rh����\� ��:^���en�,�zL�oX�uOo�H��E�f ����~�2l#�3��v��32!�d��h��W7@CQ �K,�^�>7rJ���?@h#3#N�� �d���&��`c���w �ܓ�I��Vd�e�ꋥ�&#S���Dn*pR���4�N��2�V��/4%��G�S��D�H3�:�Mƴ���/�ÿ��H&�̶뀹�q�g��f�/�K40\2��CM�VCN�]�:�|4>ڡf�!��bY1^�6J5NJ�c��U[�Zk@t�o��c�P�(5Gp@:#y�7�"ۖ��6��ig��|��PZt�7
�WB�N}iޥ�>_Dh��H��G9��;�]�k�u�y̜��[�J�e����k��!�g�I� �����E��h�ĸ�<߮b�1��@�#���tK���Nq�y�����)��@�G}�<��<U��&�%�����h[�n����i�������=m�eQ��l*�c\��YT�D�r9i}��l��_EF���t�'���=R� j"37��9O��ϪL���;|!����r������3c~� ��+�C�Mb�	?Y�D�Y1O�E,Kko�S`�._��(��e���w͌K�b��yF�G�y��m|�� �L#y'�`��t+���|��re�p�[?s�^5�D��g��`&���G]�YD�9��O	�/L(-���n[���Z`�8h�N��v*�-�� �o��<o��c��JM���Nz^:(Ug� ����ɡ,����b@;s����G��%���nG�D䊐���NZJo�����®(�������K��@�3�puh�&K7����9�5| =�NvES��gM��V��-�K��O��2B��T)/�|5-�m�-G�w��PB�K��4��/�J�_js���(����3H봐����8I�6M-��R���h��^X*����[V�g*ڹ�l?^+a�ܖf}����282.`�u�(
ˠd1���wU�5�� �G
v{V�up�	31�ŁQ�_S�f��h	,3���17��������@Iv����?`�"����!J%"�<C�Ԫ�loO�
��D?�=�����m��0��|�(t��|� �dy;b�,����*��#�~��s��L���;���� �q*����'�����e�.)��?�J�jhc#��r��_�ï��ު��,]�/�K�w��B��>��y43^h=avQ�H��ۭ�k ��M-q���mk�S�<��lg�ʎ�ԭ�v���m�k��ٷb��Y{�nz�-�	��"K��gƻ�i|����ݼҥ�@�"0�}1a x�:\��s��)����iy��l2�������x����v�"��Ǭ_n���9����s�=��u��b1��u����= 	�\����!⑽|ύ!�@��@)v�g�0[8X�K����~I?Y��q��c�����j�zuܞ*N�1� ̢˞Co�,*��ׯ�S@��Y��m���|��ֶ̀i-g0I"t����A��K@����e'�P�Zc�
[Ҍ�4���Կ��� �)��n�z�!ᶽ�P���;��"bG�d��зkY�+{�B��c!T��� �X�i���A�� A����K?K���B6d���-飵�U�0Ik�bi����p[��oe�|��p��[*8AnGc;�Z퉡J�4�fU'x^%����o�
���������㯎�Y����bO�G9�����	Sv��p��]p��W��[L�ڢ+�So����"��3`W��NB�J��E��j~�Ac�}P�L�����c�!t���<�rd�QY���a�l����V������h�4��"Z3:���|\�Ʉڳ��������u},�n��-��@{����U��o-{�Ɛl��'�5� �V�;�Zh�j���>�	�D�*�2,ꛎ�Ԍ؟e ��eOK�S�Y��s.�'���^��[1�&����8貦0��>�.��p=���^�Jd�c	�;������U���#��ri �<�hļ����p�q["E�)T%��5�gQ�ί 0[U;"������m[��y�<�{�@Ao����頲��t�F��	��_1��X9}���ɡ�x)�x7�c�ԣ�B#�����#L/k�@=qHFg�Cm�Hz���?h��
��:��Ƨ�n���£;@�<���o�iKg9l�WLJ�9'��#�:$�Hd�e`]����I-�ˑ0z�_w	Zk�ҭX�~�Zu�4n��<��T$ _�6�?�P����h5ы֏��V�J�3w���5h"�������e�I�jف��aK��ymO�7�d�3�;�u����'�ljH�����KD�-����2���1� Aq�@{��)gŲ5z���b����� 
�h÷�_�S*=K�U�4\�,s�=�p{9^���,���/���.O�b�5m�G:,�Z�K��w�� �a�ф6�C�:D���
6<r��w���|R�#G�'͓��ȧn`�`O���2&���-��s�/�[��C"0��ϡ�t En4+O�T�H�lj����#	�����PY�E`iS�~g��^0bj��r:��e/t+q���|2�&�;��`C��h�D��f(qL�'(�W¹>PA�Ūߒԕ���2����ݫ��ѕU[�F����O{ߩ�cYd���\��[.�_�\6$���c�ޝm1Shy#��f �=�O�ʫs��@���6�����cS��]	����4)�^�=��9.&.��M�͚|J2�۷rƵ�6	�?�$yM����8��J������u/�Jp~hW�}�e5~<�	+�O )�j��cN���(t�G���2���Z���X�ٸ�^����1��a"��%�aK�#*FvL��=��hZ(��OVY���z&�	�ʷ�y�ݴ��%Q�����dMX��d�V{Jt\AI��5�u6����̼0&4�2�/S�~E��z]SYKC��!/�����S���'UQ~��t�X��N�G�L�Di���5L$IE�\���S|��