��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\����q�?��e�I8�b�Ǽ$��"����ׯ1�V0�����#��+e�d����.��]>� ��\�7!*��W�^�~�w�1҈F���0����1KAu��lh��3�u�����t�(=��0+8�gfv�i���]&ǋ�������x���}값�b�eU�b&��S�sኼ;�l�D��Vc²�IԈR�!x��D�Ǡ�!����Tn�Ko�/��jfu��$��2tnɳ��H�\l�)(�(���x� ^峨�W}�F�s>�⮔��<pV_��?e����H��Meؽ̬[�ʷ�Cpo��cL�.�+�^1�7*���mL�fRl�C�\�T��߄��u>��|�DލR�;U�<oJQ��:�2z8e�����Ek�s�*�����A�ѯ�S���x��T�X�d[gE��;�a���tװ!j�����+�|II%�c[����-���|I"����/�2��qMg-O:g���"�ד�@�p0���s7[��I�W"\�]�ޢK�5;n�*"ug�i�?!٣m��^Q!�79��qc��ݜD괡����`^摙x��"�!��Pwxה��3SH�`�]��6m�m�]���zp�u��wI  >߬1�G�[gzX<��(��>����%��1y���c�R^ш����[�y��@�)�N�K��]�Bf��[��nH���2%K��h'�Z�*�
�����801�3�C�AZV�����9��?�3��%��"[�@�h��k���V}��)� 5�����<xH�I����Q���i�_N4�PN�\�W����r��BHw��ޞ毭%X)7[ Ah�n*l������/��if}�h>�he~�\�gU�=�Q��to�����)lP�`j�J�ȃ�t�QX���2o�QesA����61�lb��%�=̻)�>*��uwj��jrrn��1��w�$"=���LL{�����J\O�ܸ����ze���9	]��l�lQ���*9��������ڰD�����j4W<�0#��z�.�{��M�~�,�l�ܗNY�[-GM#��%lTF��s�����_ ����V��q��h��W��(������f=
���$�-��Ui]r �b��ؑR1K�4R�Ե�l��;0�O6�Ɗ���ȱM� ;�U��jÜ�9�jMt���	� Q����4���w�nݺ��ߖ�0�滆�{���������d3@�h=$���n}��<e��t%yP��Vݲ�ԁ��g?�rUL���?94���V�Sj�hn>}nӊ���ڵ��@}�!]2���W���%�Rب-��Y{�QK��e[E2c^��B�rSʵ����V6���N"��<�W�� ���v�|�$�
��nJ* &�q�=�4��<5H����p5�jT]�^ۙ�h �ҝ�6f*�F�)���=염�P��u��%|�: ���q��xf��+��ܶ��pҊ��(f�>����/q_��R�T'��G���]�4Y�W��'�Hm<s%-���'����9Ն��q;8~%dAXe�q���`\��Y�?��ʏ�l;� A;v��	�3����*��3��.��
+�"��/��DP.\?�@�_|KD�[#1hK�
���Ҹ��GX�����JB'��-O��D����[4f�J$L�����5�I��.4�
&��@��֯���.@H����f����2�q��q�Ma���Z[�XyƄ�|y[�Kf:�B	�&�z�r���t�s���5�A$��O�������H^ΔJb���n$ܚ>c[ ���}�񡋱n�s9}�);2����Ч^b��#z�2v5���)�V�{�߉�o�rOſ�[9�)�.��97�Y髚o�.��b7>j&U�lJv�-\j�?���5�<�z��m-�g6I�޲�\�!��O��N��p�v3[G�`]}+d�/�K�t<R!^�~�)/�/pk��ʗ�)l��
M\���[r��k�){Z�~)v��ɜ�A���E�ߊ��4*f�_M�'�k�~��v[�At	�]�!x��e�����D|#%B�W:��&$�2R��P	�����όm���߾Q�m�/!`���J�`�R��Sfr�x=th?���؝�D�}��,�	:�u��-��h�ݘts�_��;�iؙK�/�R�ɴ�;>ǖW�� joŃ(�9����.'H�(S�؉���O��ċ�*�ڄ�"���`�i����.��qfE��������a|"t�U��z�,�|��ʔYhl���`��f3�b���i%�5_�\m�wꐹG� ��'�e%p�s:�(X1��]��u`!�e,8�_k��)��� cM\�â��Ղl���'?�O}Y2@�@��$={ҭP����ί�W9D��\�F����J-��|V��ԍ- '��4MQ��b+Gkԃ�_��������?�`�����l���
Y�����	ɼ�̦˘��SÏ`gj)Ջ��C���J�1X� ��p�5t��1��4P���^'Ht1�u���楤`n��R��J��*�����N7�}�:]pg����t�칔z���T�g?����2�:��%�FI��@���4�`Ӻ�~�w����_�U	�8 �����y��K��p����ߟ[����@�IY�8A3v�{x/�r�P�ќ���m� r^P�q�Q��Z�	 �5��#�d��_8��� 'yݬ�z��\j�n�.��; �{��������?ܠOŭ�B��U8@b� A�b���ir}z�ŕ)N�[�u.6����N�d�SL06�p��5j�N0�޴�S��S���q��*mk"6�KZf�;����G0���IQyA��呤�����h9�^r=ࡂ�wA���
Ow��2�R�"��l��y�N��I:RF��8		���"��K]�r�_ڶ���foP���S��tt�-�Teq�:ݪep@b�B��+^���Ή�Zmt\��?#���y�'v�5�1��k��^N@m%��w�7P�p\#XOt���$�=����JڏY����7Epb c���>�Ή��tI"$̑F-��j�SxmH�z�n�����9D�U��&���^�"��5���$���c�S�ɚ�%E3Rot�?d�/Y2�U�C/�у��a��׾���g�}�>2��սd[ ����ss%��t�&���u��g���dz����M�Db��T<ŧ�I��2`��/��$����I��~�/�40��RP^vhl�����������ԧ2X�*+����d�z����4�;.�nAwx �y�b��A�>o��4)���ɯ���n��-��w��6q��g�<ǃK4�ڛ횣Ti��,'�Kw(��/Z�؜q�sV���C�%���#@�����Kb��OA�2HŴ�o7�.9���&�KYJ����w���ggg��wbn߻�����0����Bƥ�J�2p%�O*�t��@oy��Q{5�5�״D3���!c̑['����e2��}=��ܑE�	8�H�3)��t��[����6d�0�IK�:��z�K���+�p����ӑk�H��@~�G�h{�[XUMhߥ(�{(Ŏ#t!�<@��u[���P�K�0g<r!ߠ�Y��[�\xū[G�
��vz3���F������d��ko!3����}!�Fv�O"O�#�mj�����q��g�[\½D*򤡙?GZn��:wD�yނ���2�,�Nt+:�� I��g��]�TJ�Uv������JmX'CV���KD���4�(	�t��m�|c��ɰ�����G��dAe9&U�߫j5��emC}hr���zH/ÇY�B<^��y�ٲ��t�@Q���'u8>C�d@��ZZ��e�Ŷ3<�N^ 9���xI	��1�+[^�Lf~�>�*q�l�',ua
x�?�n1~I@���FK	(�[�5yh����hu�@4��=Xg����zؑ���� s<IP���,�q	��d�߆wN���By���̢j�qN�^Y��n�Wu�+�K�8k��j���sՉ�w-�uT$����Ӑ$�Q�n���,ee�\����]�ok�#��A���[�i��E����f�]��<�V���ER�ѓ]]O��}�}��������1�7�l�m��k�,xa�XRGWx�愺Ln�?���������(���m�B,q�U�ZZx?Izه�TQ�A<�ܫ�sL� ��J԰�w�	V$�Ǳ?��& ��-��h-���8��'�#�~Y �Q�#����M��&���%E6c�ՙL��m)�~�͠���i�s��W:�Sk�н���3j�:�w7�l�?�wZfeQ9$m)�1Oq�z4E������{� ���Tw�֝~}d���ey*��@<$%�{H�ݖ�ѯ̞,7)���nIx��X�drK��VMwl:7����L��5��壸�v��*\�����Y��$�82�^�Οc֙���WFÝ�u�^	�܆rֵS��A��ե;z�'K�k�����D_Q�ڵ�eLRN}O/t< ���{-R��]�����5_߷�Tc��p�EMR�����RW���%�״R5�KN�ҁ�ǥax�i;�L�̽<o�R�xG����`w8<6h�2W������5sO���{O���4���
���u)V�[����C*Z4۶�2����o�ܛ�W�����0}^E@�IU�Ss�|�}�Ql��)�1q�a�*���᏷ҙ�[�x��Y��X�e ���T��K8�Ek��2�� *鏫n�. ;��ҋ/,*�ѩ}��v��Ѡ#n�s�N�!�����{��i%�| 5�|� �R�>�����<�:m��\kMخφ I:�2,2S�{��7Y5���z}���B��V�'����nΘ�Al��{�t�s�M�o�$	�H<��F����Ѩ9��;����(��N���jWFN���DU`60�����͹�<6��'Ig�~�Q/|��8`݊~Tn�c��_A��D�&��/4�(�?	��B����#��<���R�A���ȗ�֠SN������T�k�9w:d��꼔U'��=Y�_d�X!��4G�4��I��֘���ؾ�і�G:စ3�O���Q�9� N�4��}	�>s_��2���ZR�箠���I���L�w�̏ŉ~dc�Z��J0���d�%۸��,X���j�N���Bt�:F���x���p,���������Y����\�H汤]�&i2W�|����ԁ���.���\V�c�[V�eM��c'�!-6�oiN�(w�U��M9
�t.v���2`�@ГM��Z�/Zǵ�?vh8���v�k�6Wd���4��hO��j�Gp���*0A&���_���9��t�Ōs�}M�y�J��7��kNUJm��^6�}|��{�����>��!��@���s�6 S|U�~�w{�E}�g����ػ�7t���] ,��P�'��zGUkE�������neN����1p�F�ۗhN��ܨj�Ǎ@(�2ε��\���:^t���Agg\4�'Q��?� ��M�1y��K<�8�y���;���V	��FH3_�U�>���mڃ�<���ϔ�<.�Y�qNEO!���(`qk8����ދYh��%{�sm�7�BS����Z:�O�L{x.Pn�M�q����-��V�j�o׷2��
�99	�B�V��gA��6��z,�r� ����Zn<D��)x�X5a�0O:��twu�ӇPQ�Y�5�q`��{]kx��	=�.�Yh�βr^����qE6��z�;.��<���J��f;��v�I�V��{�Gk2x3�YkH��&�'c�S�G6���9�sj]��p�D���9q%yZ���<*�������V��Z��|n�my��*�*��jm!�-5�B�4��>>�/���-�+; fp�_5��280d�W��׵0�ֻO��P�~��K����e�?:���QdE��ִ��;(���=�f�)l3D'!c�y���S�����*�����l� ��D�u��в�rSYJ7A��Y�܆�=,#��>���o���D��Bʱ�\��y^�C	�F����Ǫ���ߺzqꄟX@�P�0cOC��g�OUdd$�U����uIS���:��Nw(�d�C�O���&��DD�c;���&6�����>��U"Z :�����X�8�y6Y�iz0���s�|�q��
�j\I.��Ĩ5	��]#����p���<Ҵ)�'7N�yqE�c�b<K;y�1����!�����)��~�8�(�s_z��Z��e���h���R)� ���
���fTآh�Q��jIw޶P�3u�A/��1���6����i�8Z=t0ԍ��������{D��F����i����Y�_�	ȷ���j�W(��ٻ�d��v��^=�:���Z�j�s4;a���$�Nq�q"��yE�z [H�Å�}��3U-8���"E6��"N�j�?�@���7F���<�)��KdYj��lK|��R{��b|O�'GL��������:�D���i���C�� �ª`��bS�0�:VV�?,z��o���+��;��9J�t{��]�(Ą�v8��bk�k��}�I�t3�u��ǔ���;$c�<
�&����u�Sw����Ss��W*�jẤCg^zrmeY�]��+c���@hG���ϫ1���`r(��D�jo���Z ��{������Q�m�6I����<�'���I�1�I�m��������4�I�i�;���Ga��CY;g��� z�P�ϋ��9�Kˆ��Ժ��d���ς���W�Чo�֫�j6ů�n+5`�}��Ů�ɫ��R����E}f6� �lHW�aF��[k2�K~ǖ�)��r�C�{K�\F�T°�5���J����4^ɼ�����Yg�UNQ���E/H�$oԥ̹D�@Z�[�=wT�LW9���J�^��}D�d����Z��7?�~�VߦH��#�x
�F�_��R�����9�ؔ����X@�<u�ʟ��/���Н��(�'��(p��	����O��Zp���nWTK>	��5��MV�]t�*�� ��d䱍@�4"��]��:��H��0&N�B��Qm�r�;�v1ⴞ�N�GZ���O��K�D��G`� �N?�6�[�r���ť��L'T[���h*%&����XP����$
�������ALI�����{�I,*U0}�, \_>�|`���VSE0�N�U�lU?��L�zg45��g���̡�6�H�j��_��������09ya������ȡ[*:O"qfq�c,��F�6��
I��X�/�鬻�v��K��b��Cv�	�}F�y���1�&^l&~�g骭B�o{w��:�2�'�[�~�!+BN ���;���}䨨+'3�j�d-��\�F~�5K���3n�Zg d}C�{������@JA��9dl���_��Cش
+��x��� �`I�n@���\��q5�������?�ák�Ir��^i֒ �X4���ޟ�d��[h���="i搲��嫨�[�x�u��I���h�3f=0Ճ��-���fI}-K��#�d��ӕd/��؅�x�y�t��a9�s��0T�BW��xna�VZW���]X�V�R��!0�R~����j30�X_\��)i�">FX�R��wU����Y ��G�FZM���qw��Q�O���Յ�����h���V�ԏ��gځ\�d�9\!�O̻�(bX>�<�'���Q@�k��w����K�x`t}�?�r���P�:>�Tu���Li;��#�
�`���M ��|��ID�P֝�p�|��'vv�;�!���C�
��p�B��։xu�䲖���<��^�i�u��"ey�m�zzn���pˑ[\,y@�0����?��8�#�����J2'��'2��$�ZN&��e�8Ԍ*<�]�x���0���t���*�BQS3rz�;�>��e//��;���^>�`����\�x^�@�w�ݶ���}~O��*��w�m����(M��[_EM>j�=����������d�c�R��Zn\" ��]VF�եA�W�v��<t~��8^�ԉ@�d�d�1R0�K��օO��2�P[���!���BP�?AD��9�QeJ�{��}\a����-���~F�Ko
�0�s�<��5K�vH!o��(k��%1Y0Y�����b]��|Y�['#Z��^I�ˆ)�}0�J���&{r?�3��_����
OZ&"DF5[X)��I�"*b�|� G'�A]�j` Z��)X�3�'��3J�@~���������h�y�i�D��f�
R*MN����}|K< ��S����7�!fd"���)��M��0�����u`Vm���u��!�r�����"�37�:'dJ�A�d�+��T�a���a�.�ǰ��>�L�g�a���]j����[Ð���m*�Ѡ�l�,���M���?�zh�R�~%�7����5EI�+z'QA��U<���Y�X�+�Ć�4��*�s�Z�z�5
���dVTz	 �	�zl��A���z�ъ�m��N,�c���g��A��P�2x.������ц�d�� �e��VkH����?���3�oً��Q|[�ƪ�S͏c�7p?D��Vօk�{Ѧ��"�4p:ƛI~I7.%�v_��H&�a���ϱ�*�H���� ���5ĕ��}=�G	d~�C�y�Rh��;��Zk���ej���x�k�ҳC����4��09]n������C���8=���(� �(���@�.=�������a�հ7c��æ??9�͐�L$M� ظ����[}ʧ����j(-2S-5��'�P��2 /K�I}�����~L����e�܏�6c*{��:˳A�-��n�	k�Ƚ�5ŀ�VUx�U����Z٦?�$Md&�nG�.�=G��$��-���>]�r^`���p�F]˶<���)�4�u�7b�h���+�y5�4���%%r��G4Jד��3~�6��^���\^�,���������� � ��e�Z�b4�Q�����U|�v�h?�z�6`����"��@�4F,y����"԰-�7�k ��4�_�L�-Ư��,���2���`����L�������:Rj���D��7N�\L�BrFI5;|���)�qo5�����}{�V����'��CK\4�B�&�h��K`�[pW��=s�fC��#��{o�$d���`��/�5�B�NJ	k��Z*Mv��՟D�Ō�nf�UtXX�0�=e8�,��ǝv�|bA������D	�+�A^UL���_�����z���I�U��q�Ay�ҺÇ���������|NkZ������\�OJ�3��I��,0��՛+�bE3��Z:^5���(�-N����N�]�#�Hh��0�$�5�"[����.�	Ot`�f����o��s�nӾ�] �wZT�|�no�����k��\��F�.��9"�4e!o48����#Zi�d��p����B�,q��DzH�m�L.h`G7��������P��n��q�����lM�yPn��(cfe��܏�����N\��ߟ�D[����Q�,|!R��ϠxT".{�#�6� �]���c��L�m!�xy���揑�z�7���Y$�xðd���vtG)�����<ոW\*lh����E�Py�)SWZ3��H`b!R�h��,�O5:) �E+�p�y�Ů�m��4P�����7�$�w)�D�v|�j���,�A���@�9��m!@����e��<����+'�;���F��.8�����T�!Ǡ���-�LUQ;��|�	���������9}��&'ηS��[|fw���=r<C��_WH��@����m�d"R���%N�e�HM�?@A6�t!�&�g6D����|�%�z�q���(�����o���[�X�MI�)�����|"AA�-;?��o�-Ա�;�����'�B��LR��F4į*�%gA��4��N-���d
wYu��͒�V2k�֔��:s�i�����z�R�|�f��e�J�ȔE6����6���(�K�UR�yZ�M���l�_K�(4`AdR\��hR{��"��7#	=�U�n�p�eC$���ơ �G$l)�]]hӛ�^���H�l��O���',s)JE��C:T�8e��:{芘>�P0���=��������k���'��WZ�?��B�]���6)f���ơ��) k�`!	�!<����~��U�C4��x��ފ^E�a�jJ|�,̜�g��^��n�E��ݽ-s�h"��#=�M=ut�Z��'7y����B�YǙ=&�;7	�j�.3y���N;�?$���ՀTd��q�)�To�l�Jj��	$R$�d�?���=���"���f���A�����(���90�}�K��RYާ挈� )B�rn(K�������;�����+AJ����3��YK�S�`��$�1�^��������ދ�]�D�}�����E8��{�zPk��QK�q�D����h����i/�b�s�o�f;J&�D���	��0���@-٩��
S�o;EM��U߰Ap��4�屍X4ΦKOE4	�@�/��'Ј��#j���ZO����|ӠAR��BSz�/'�ĪA���+��4r����ĝ��(
�eA��#���{�ةr����w�D�Y=��}_�=˰��� ���@
�uR�{L��"^�,:�?*�|_� �_>}r� �pQ#�ᢵ�C�`W�@Y��`��!t�H-iFs0r%RW�Ű��uX��g��ρ��~��>�ҿ̡�(~+��2z,N\�s��0�.$��3��@+�r�K�7�B�K�w?�"H�}�
��h�򒱅�]d�ik���Sq�nV\��3�_��A��)�Z��2�=���`c@n��4����xc��I�.�4���aO<*�c;-Z�=7H��]�u��� �$!�B�NF���rZ5׹2J���r1@ASHmx2ϙ��l��@�2+,5M*�Pi(9���I�!�6�����%��1i�yC ��Ki����7��" a�/J��UDh�3���T2�r��'F�8Y�����vf����a5�?z�)cO"���E���d�=�V���%�Tu��M�/zk���0
Y���yW|���K��?��V���0�<��{Z;�gk����,�v�r"`B���	9\ǜXesuV4����"���a�a�����Zʸ���pi7� ;qm��_HKcn�s<���3g1w�퇜Y�Wc1hH�U��i���#@�� R�`��'@s�w�+�r��@�x��+�q�FNā{���"�x��@NV���{q���6��zl��gοwq��(�I̥���z��%�\�A7�F�T�1ߏ��N�	P�����z�Ǫ
��k��n!-34x��Q���Q���r�dD���pq��+���B�fc9�td��<�OlL�w�FghR#Z�K:��km�k����;�Ӫ� ��ܤ);��ْQuI��$���\��}<�d3r)����ҡ�I��[�����x];�ҟ7}��0�����Ja�Í��/��#ߗ�������DuE�l�D�4���0/��w:�s��R�@�c�LUh�C�JL���&\!�؞M�B�#-�W;�.�ւ���JT��T�\I�}L���ӣ���2ݵ��1#�#���5��˛�Nǵ�Ƙ�b��H	.W��R�b���$��:���lY��������d|�כ����`0&�C��I�#)B��|oy'��Q���;S뭓���L�׭�,�T��񤡼c"EOﺗRPH(��1��ܽjE{�b��f� �e��ӹ �l4��lz�r�r�G_�hkrKa�R��<BMQ��z���L��&w�F��=R����o�=I2��5r�y?i�?���ں�R���گ7i��̳m�7xu��6C������䬦��%����hm�G@F�$�E�X�Pj6&q<3�6+���mc��O�r*�I9\#�D�:O�Ç�P�95p��aRT����L��-��B��B�<��~�(^S���a���f'A��n,�a�a��I�@�8y���/3�"�2R�M�4{���)��R{��p�.�DF��m�4��/�ro�']�Ь���NU�]y���*��f�5>��.8O��I��w�,�
��t@u�	v�j��X���/|
���������wƵ��ƒY�Ȁ�D�I!�R4�����|��Gv�$���\�N�Wp�65���o���o���ʀ{�r�@E��>_|����e��%[R:
�`�u���`�� �䭉�6��?�T�,�~߈�u��лJ�ǻ��"����[��ħ��C��O����)�
�8��k�ȜA^���"o���𧎽�j��)\"���D���j�?!��2�>�^�6y�gM��1x7����'5�������a������S>hI`'~`$�L�tv%)�0�,S�Y�@,4#Dl���G������7�	��Oy]|'�M;)��=	H s�(��`C4��VK��{�W��d0e�}B1PM�u�zU�D��e��w\`�{��D�����]�֬/
.o�Ac��,jn&�S��ݮyc��I�~��Lk�T"�ۆ�Վ�Y��٤�B��Hay�ɜ!f�l��_�fg��T����QR�v�U�m�\>ѷ���y�R0B�����6��o.}�/��;lC
�{��u;(��w��;��j�z_�����м�Yo�^)`�M�jf�۹G|��m/�gb��P��R��������n�_?��T;*	�`��LkN�{L=h y �{$ASO<�^3M",�'Ø㰮�ml]�L���<��j}?�9i}Ճ\rΝ�0�@��!m��k��I��F���྾*�>F�	41��[��^)uh�M���;�����/�g��t�KD�R޹�h0�U*��PYl��?�=CH�^�lD���E����g*�ᆞT�ך�:�O�Dp���I@��FS����D�b_T�h�� ��@��a��'�O\�d�j�lϧ(��uwrJ���p���eұ�wb�J�u��(���������3�s���p�)"�Tp2X��uڪ1�b����F���\���,J�\�y����O�u��d�'�8� ���;rOR��[��.C�eX����ф��.fS�,�3pa�E��wK��񿿁Ð����"%�;r�J�Z˅9�~g���[2ҷM��?�B�&�{�����9v*WG�k�R��a�Ɵ���S�W6V��=��#	OH&�ot��c!;c�}��[��V۴v��` �NP�}$2�T6q���P%$�ؼ,c�|��遲R¾s��{|�	:f���8��(4�db]L,�����vB����P�v7��t䭒��9�U���쓝[�ߙ���R!jOr�:��^��p��͇O@���Ǌ��>����&����k��� -j���(��䤷fX1��"PF� ���zeG�������B��s���j�p���������f�!D�e�m�ETǺr�0j��_�'��1=d�=ۮT�]��tXD��Y�+��0v��D�e7�����-ݪ���E���K=LwR��FjM��e��Bh-���̓��)������C�N��w�s�B8}?U�ob�ϭ�Z�q^	����8��f�zk%q���$��T���|����zZ���cz��B�����qb4�;�tT�`n��o��#���sZ��ݹ�XFI�G2���S�'�|��90��YN��$jtr[W��"��M$��^Ҙ�aUL���w��܁���F� ���l�S�WA{UXv�P��U2O>f��Zv*u 5F���)7�0a�5��j�$V^ؑН�� �����&�=6�c�,�^�� ��`M�p���f:c�o�I��	�,�h��=��{jI��;��P��/C��EP�~��>�5b}��%R�$u���7UNA�տ�=d�M$\Ss�i)U�7aK����ތ�{�u���1��Q3����!���4����YS���D(������*̙��q٘k���3� 4,�L��p5���??����7(�&A<����e��2:rְ6���2T�,k��T��,ǥ�m�+uz4۰�U,�_ޒ��G���h=�3����P��u����C8P�!_�xO��־� p?���Y����HaN2R�9�C.I,�H����� �5��\�q���X�"!�h�@`��7�,l���˵�O�_��1����G���pp
�
	�ᰄ�>���o��f�U�H���6}�EZq�l��z�&ߙ�r��
n�<�'H����k�{�Y�@rydOZ_��O���_�2��&�uیf-]'I��(�nH1y&`�4��z&����w��)ߺ���:d��Nc
T�|D��qal"ҕ����+y+���S�cx����r:�P¹N`{���$�
S&����)����b�Le3�Q.Y덡\��a�Ab�A�����-��pq[��џ7؂t98����)(�Ί�tNK�f8�=��jB�yZ:�^����JC���Z:�FXۂ�3{lk�g+$&�]�l�pY9�����ş��<s�-�o�OǺ�b�5	�9洯/"o���piW�dI,�Si����Yi�;�Ɠo;p���ef�eϓ������T��06M�e������`.u�ג�J��ٍS��E�l��|7W�	�yw��h�WVm��w%{>X�,���٢K��2�r��)*%{�jUs�������!S�~�)5(Ir�gxw3Ɵc��(��a:��:O'W����i�ZS����F�B����~��PX�W��.T��?P�]��^��l$>O�e
�
q���͠D��*"uzW�Z�?�UP��0�,Ѩ/�6jGD3(aNpSƊj�x,@���y�7���ճ�䋎H"���픉����˳t�t����J�@����t�J����c����e%�g�:"�F�����C���¸O�����ܿWå�����kg�-;i2�3��C�v�e�#��K���b�]��&�8�v���j���j�d�+��'�P�dGK�����	��+N����Ol�a��a�тŌ�4\Nʎ��.]t%9N���L��!(���c��WXMҸ^m��N�#e"���tgN>� ���J�e^D�T�ݝ�<m�����+�*��sb�� ���e��g�6$?wd�V#0u�nr�˥�����П0���-�#_�	%��i�|��i��.+��7b�ݱ�e?(vHt��2��4�CZ-F�<�"�'�T�7Z���>OO�)���vy��g�;��Ec4�D-�KT�3�c��̤�!�.iܭӰ�.Y���',/@`��b/�E�@�j����\�0�`C0�І1�.��(_b�L	6x�z|�!Y[���<E�6�!QQ���@r@�t���m�wNNkl�!��p�J�5���|E���F<�LVaViε�I��(e�ц@�$ �?YlR��X��ךw����������}�a������nq�ގ�h��v��d���l�(��/��[���Z"�z�bX�����Du#L� vx��%�<F^_�O���{P��2�����1��EjWM�o���[���K������e�M�W6Q���
�ܱcxր����,��\��[?	�$\�%l]���K����;�O�@�,w���@A1��ry5|_"b/̫F���}*��M��Bs~��!�%%L��Q��b���6�x�	�%�B۴�e�t��_�����|����L�ܑ�i��v��}�]U�ܯ����;�燡b}�ZzA��������n�G�I���� �_Lϻ��:��(�~CXN��CP�@�A94���J���$�^��`�����-n@\�/��	�
��#4��S�e��7�\�J�����ƞ�b>{�7bE��O�P}�e`84�-���د:ce]�o͙�-�s�P�c��I�i�$�+�34%)�=��+"a�Rj���y��%�9k�&/,'�P=@J���!5}H8�_}W��[����HZ�ŷ�	l��B���U \�*"+�e��0���+�n��k�n��C�U��U
H'}!4�;b�75��Bч�Th�p��=%��_�`q���5�䅌	D:.��s?c��Krܗ���꒼��K��Nr�(����>RAn��fS�F��	e��y��� �>��o�~�J^���]˓��<�(���(�X1��ER�o��ϊK��r�!]���X��2Ps�W��PHB�����,R���qq��ʳ'x�~��B��:�LI��B�p�PL�n3�{e�?�+p���rv�ńs�~���E�����y��p�Wn)2ݔr��B��j�{9[H_����i�9�ʘ�D&������r/�y�H΄��R�]�1#�O�Ur}u?\�T���M��^��iX4��#�/Y�$G8�u���
e��Ө1� ���Գ��s"���B��H�%�|,ݍ�v��c'Y�u�Zy㝾��'��Z�hU٩>i��6��0��q��]�}�Q���P�鄋"|����Yl�:��~�:㶸iR
�=n)�IRPaà[f%�G2�ʼ��!�
����h���?�D��������u;�+T��3$�0��h���S X(��9ZA]JP	M��VL�\�I4Fzk��0�O3�y��]ˇ�0TTu�s�?�j� &`��x��	��w߁.i >�K?Ұ9�m�����o6?�|��~B���e	)WJTd��Fga�f����Q�9z�>�L�S՘����c�n�@)�*on��r�v��զq�֭��Z�)ߋ;�MDE9���We�|	�q�pa�x;��(��hC�ޚ�[N�=�k17b#)�.����B��4M7I�YG!�(_$aHč��P�4��N0�������ִ��$;^�&�38}����6�[��d�|"�+�������u�y�`&|.�o�|�<JKq�]�U����L~WM��({!�D���a]�4�}f�Wѵ���ȝ��|�i�����`{8N�A)c1:�.Ga�x��Jt��:��JA�Fh�$��ѱ�V"2D�� vB��D�~��;�`�r�g?��X�z���vJ�Q[��9a���TU}��
�@�����3�Y�/G��x�����2�l*���c�Y�ť	�
O��8.8��-(���� 5�6��+'��[�>���w?S@" �#.��E�\3 �J��z3e���2�yU��%&Ɠ�~��Qd�����3ݦ-��t=&y3���
p�]oе�kJ�jB�J-�"���eNr�:zJ��u)�"�̟���\�Ż�����_*����� ��;�i��`IY<����P��[���=�Zڎ���(����0�����2H�`�����>3���Y���6D��wI&�r���#�W`��/����*���[�8�;���|^�š�Z���*�Gcw�Tܥ��h�i��f�D���qb/�F���gpq_�����[?��f�|���B�wE�������M
�mBw���`�!�.�æɘH�IӶ5xg�&_K$�������m�BI��F�����x���sϕ������>���Ma�v	[ЗW��9��kS�ڂ�έϾ�Pr��2W�]lo���)N��h��7��N�x���ޅ�\�6��=�Ř�[�#��չp%~���� �`K.��6v�I�&	g����	�>oAjw����J@/�z\ Ӹ��v���ީ�0^��^d�8 k���h<���:��GW�/J�/&9vH���nkb�+���ԅrFۭ6M4.g����q,Z�`aX�/�*��˜�[���Z��
����[��&D�7�%[� eU�:ŗq}�)S���@k�}�i��M}W�D�fDO���aV��,2ݜ�A0�ع�)l�6�����<�|�k�ص�T�ʨ�[2�.�u�vl�ŀGE�#y��q#���`�����t�w��a�]�e
w�H3�YT�4�`E�Yto��4kZ� }P�6�m��ˍ(J�â,�a�H�>�����݃ 
#�IF��'W嚣u��8�S��v~HH`wyQZ4 7[hP��h:U=��B����VF�����7d{��:ҡ�z��KG�$���d�����vE�� i,�+�egx�ɼ��8�i"�oF�����EM�N%Wzt@H�(-�H%��(��qZ��Zd�Wo�Sk��Ȣ�e o�,���"˛�_�n܊m*�{���t[�a�7�� �
�S�q)��Ȼ&�>5&�n����&��#�SÓ`�"��,�I�j�0��2�䂥=��[�]A�q�PTn	����f�,RU5k�V�|t\61Cܰ��)���'@?���B4�"[�ŅH��D��wB4!�B�"n�0$���o�=@�7�̜��顢�Ӎd&������Rj���v����%��jP
^{��U-3�&�a�zE�:4�S;-C�=��$↾P���ދ�NȀ��Q�w1r</��x?͍q��)Z(2�b��o<�Z30���QR��\O8b�rk�:ɩ�̫s�o��N�{(�ߝQ��M�5;��{/ OM~��u��	q|g<` GeUA��1�!�#����r_��Ă���(#4���;,h��\.q�p-�����.�>5�Xu31rـ{n"�z���=���ڐz�1�t��F?m/=|I�����m"#���ѬTð�5=���d��c�t�0�(a=����p�w�uO]�K�	���%�7�o�|1�ҡ�˪!��X�uW�y^�W�NYspH�Y�� �tv�9ċ�q���N��Axbw�����Mr�6�m�l����|�}= ����/}E|o��G�$�BU�@�����O5F	�?`������)D����@�P���;	��i�@g�ˬ�}��;QB ��u�Z7��	��!��:�K�x�����˝�P�R���Ք�a슈�q�,���v5����~7���O�.UB]n��*�*���x��������/p���
 �3�h�vxɣS(�� 9n�����2 �Ǉc&l(2��>	�{�`m8���]1o��|*�Lؤ�����ӅhM\�i^�����ޕZ��e;K������v�[��=�#6��W2עM�t0�r��8�'-A��=����k�e:l���x��D�u|s���#nY�D-��5�iS7%�߭4��Y��҆�/�X_E5�}j��l�����p2
�s�]�on���K�e ��rĿ*�v�bkS�{6�j�"��x	�,�β��
:Ʋب���1c��5nnbi���s��7�G��%�&�]��HmwGj8}��R]iT�e��C�����J1�ϝQ���5�G`&���,��Q��i��	�z��ObM�`��K�盤��[h���yk��%�2�}�̎%�������M<��v�d4m�}.�ꥇA�::G��ΐ�_����.T�����o�W���K"D� ��hC�G����o�SM,�U���w
W��b��� *����$ ���
'r��z=]�� 8��-�I����A�??"_h?,�񀽷�n��p
Z�� ��s�~�*�讠D��č�G
z�z~ �@��a�5��3��|�P	�!*��g5rZ�J�!������$��k%��('ܩ1H� 繩�oP����4П�I�c�w_��X�2;9��!���~�����W�~^�?��͊׊��c �a DA��3���Pӑ;8~��W���܅<��
�@Lӱ�\����={~-����ŉ4��N�����Wn�~1	k���*WL���3u�R��<�b���ҙx�����(_�huy�9,gnz�@�Y<9��(�A�tg�5��i��"Oͯ��t�3s	�-��C>+1�u��[ ��?R_����A�׮�KK7�G'p�pg�򶝅-3/�K��fcO���U��A�!k��./��//��>���i�=��Z)x����OU�v؈�:L� �3������\�S3f�(�;n���M�:Xd�*��7��S!�&u,��t'3`@.�2c)�HL��dG|��]�=��+x!3f�'��>���-T�
��F
D%�9�	+2d�����~χ�H��{w\��`�'xzT4RT�;��Q]�O���I^I�v�~�v��R���:#�H8��l	��V�����ыn4�,��H8u�}����[�q5�Y��N_�!p�1���U���D�<���tf��'���1֪$��g�� z|?[tX)䙭&	r�-Aѿ�RF���x�R<�QM�FlR���f-?f#Y���J�x��3;��u�,@�\�i	�ZaQ�[M{�J �!�8�у&m�ͷ��a	�Y��МV/�i2�MM��!]��mL�8���2��
� 6a������i+�f�ZD.�3�;�G�T���7@�V8�>�B/��ӱfD�������q�>ݍr$Z�b�O�#�֟2����5F<���~Y5v����@e���R:��� �j�z����2��Y7�8�t����03�i{�)�Gw��I? ����i}G@�+�d`�nf-ZYY{�Ҁ�;��A��XX�o=>���]�+��х�e�M������]͜��
D<�ȍ_xC�[lX��I;�#��C�����׼�>t��#��c�hs�[� �o:��_�l�nK��-����9I��p؉r����c?An�f�s�mg���^�7~-a<C9���U�!N���,P7�k�D`ג\4��Ԋ^���	dk% D�(����D������K8|2W�1
��]#�H:7���S�׼��w��w��z����YSqIM]�B�\�2�I�����spf���Xm!����Suf�#�2��6���>mK�B���c�#<.�"9�{
��,q����z�
b��$�0Y�?g4w5�F�]����?��#u<J/��U��F�28H���������L�m��^�t����N��C�JZ,���9`һ̯��~�8��'�}	�U𨍌K���'�Ti����Sg�Q�Fԧxn�44�j���"���+�.J����I�m���0�
�e�?����k*f~�E�о!�{��{p��9rjGh�mJCL*��&��J5-T��`�e0�a^�[�����.�獎�6G�]f�\��)�nnL��we+/B��G5��dÛ]��`���pWr�mP֯G����b��k��'z��1���{��9_�#�l�6]xV\��c-�#U ����m�u@|@֍z� ��e�c�Y�_e�RϿ�x�#�]u��DZ,'����i�L�������h/'��wBE��#����[�P9���h5�<052f.��λ�LSc�T>Yu;OϤ�i�ޞ���!��#��8̂@n��v�1��_�>E�lX^��מݩQ����, �{\���eW]�8Tg6�yݙ6P;B6�W��l�P��~K}t��yOz .A��k�$��R��� *�-u��O����b�l��U���60�m�"��KM�48e�+��"���lء��x�&�Z��=F���D��:p1��dY/.x�U���q�S��Y�S��1"P�-G|a��+PQ>�<5�_0���I�7�'NYXhƸ�v�ڊ��.��T/=�	- �s���t,���Z�s`!���RB��"��J:Q=hO�����1�������5>!H<̹o�H]JMCmHЋcw6�K��]����:�+"�z���PI��8��.&��H"�u����qR�E���� U5� �]brÇ�P��
c��E�g�X�Z��G��yk�F϶����� ����iN�x�ρ�}���1��X�lx��n)#�Z��L�)��E��[�j�=��W�G P���e�[��&�����]�.d��F�5k��_�W��7͏�|�1�n\<Z�c~��M���O�װ5�(U�%-����c1H�şj �'��-�܆I��)1�3N �./2$R��fSJ��Ex���|$`�SQ��4�ix��D=�*&n��@&�f�-N�
�GB|��D����q�&r{i<G8��+�
���������w�ܘ�M�5�l_�Af9���'������N��\Y[��nb�= $Y?��4r��F���=E�c�+Y�D+��������N���%�Cm�'
��r���6���][P�Gq�\��X�(��B�\��"NYЛ�>	���)Ǳ:������~�MJ̬.�މ��tK�i��qƎPl]���Y��k?� � �N �2�	��	J\-?PԘ
�Bq8[Q�Ӕ}��_��D��0`����4#�e�}fZX���N-��_rgO��'3/l�`��u�|�f�X~�By��i�`W���/@l�}�ȧP̮n�F�9�{�
\����cE�ˮ��m&��� ĉ^Icm�-��J8�[a��`�[%pf��twa���V=��e~������^�f�5��q!���Ń��'�s�G�SC�̀I�����EFyŬ�ؼ���b�J�q�
X9�xtG��N��p9�ǡ������ľg��lt�68����qn�[��7�d@�A���\͛��� ��I7L1�-��&癨µ%���"�R��`�GzM���'�,�c��e��ن"/u͍3�w��;Q2k�R�	/���O�c<r�(}�j��1s�ãϸ��|Tx�����$����t���D��bMN]k6k���	AĖGvhW�~�����ʤ�����c�j�tWd�p0���9�ݓ��o&L���tE��U���s�L��\�����ї�����Pߏri�~�,~�P��\��4-H���; �Ѱ���ڎX/j؃�M��#Az�d���ǽn�(��[&K���c�L����WЭcG�١5��$��W�iS� ;��o���j
y�G���vc�
r�wf�B������q��z$h�h�͝ JgbQ7\4rk��R�@=X��S}'���03�L�6��o�	�!;
�{ֈQTJn7{j�;�����VW��DzG���j��."T�8�Tx��ƙ�$�\@���j��[b�U�q�]F�bk��	�B�<��w� �Io1Q/�����o��z���J��{nQ��d�X@�F�+΢�dH�g(M�������^^DX�����/�6�v���I`&���RWyD���E�*e����Ƅ���W5�XyORk����:�'�%|���������+kה���A���߯�ਝ���A�e�8G�V~���"W���w�.��c������-����M���0݆l��d�x�	�1{�Y
��j[�]�uV�o��Gc_��q�
i��הR�]ƌ�.��t�#D_����aP��)�'2���H��+�d��H>���Ș��4[���%����6�pMx�yU����zH��*�ud��:6@-����*��S�{��`eR���R�*�U����\x�Ⲛd�`y0,�IA�o�Z�K��Hu8��K��0Ɏ��^�,M3Q�����8i��d޺ۥ'A�u��虐�ΦS�ZY:q0�I��4裄�� ؂$��]�B�cu\	I����Ǜ�	dw�T����9�X|���ln͹�1�����������Ŗ{z���%��-x�o5�}��].���.?��x���J�I�}1oy�r�eY��GH�?�T��������:S��˾E�ԍ�Ѡ�1b�Q{ |��]����M#�tl�!/��@oʣ�!0*]lכZ�x�����1k�$TJq�>d�ʈ���>��<w^KJ����#�9m0�6u��?GD����qC���׵\���L�j����f�e@'-"XR�Zai���*�dCVR���F�?�_M
�-�.ac�|�	w�(9��}��x7��H�ǒ�yM�Mg�v��tV�h
�S���є_-����F�k���(���f��'���1��钑���;h���!����_}U!;��6�,_����
� #X�|[�J���7*��i�ܪ�R�;-���vP�d�yΊ�#�/Э��:��S!��w��@æ�������f��V\�2��Z�2$��b�ڂ���l'mz�	M�<��|W$[�*j?�O��t�"~�7m�����1X�p�E�z�m� �C��%�Zϒ�H7����E��=8
Z�#�e\����f6��6Ѭg������@�o#�%�j�d��T=�o���q\xjD3�2ۈ�;}�ȱ ��d�5�Y�@To5Ӗ��� �+�ȡ����	�?����(,�%J+���x�/�v�rXHX|V�ۈDgAo���Gؗ�)���̙�v���A����TG��[}"t�H^�W[x�~��H'+x&����X�=
k4-���*�ɵ>5ʧ�r7ᐟ\���W��q\��@�I�F�c��6DahH8_��J~�ѺI?��x�6���[@�+R?%��97'q�b`�]R���3��e�)r����:rU|�Q5@=>.�j��7�_��)��8�F�zi��Cj�й֜��,#�FUi�i(�ч#�3�4�,���r�B���>�=����ϢCH:�ݗf� v�i�R,�%���/�+Q�^��i�����,%5|Jm
*vIM�ێ�i�޵V_T%���(�"SX���[����J�beS11��Ai��5j!���ꡘѿ��k�G��H����^7��x�\�����B�Xl�8�{����k|�FR�}�u���c"��lC��H �� �Y��(�K�$︘ &8B�E�f�lI��K;�f�͛N|9��4V7��<�f|T�	��\E�TҎ	rYk��RP�G ����Z���{1 u�!��@V7�2i��yr?��;�^r�s���� �ؚ��<�T]h�����z�dP�����<>1�Pc��@FYͧKu��B�F��^�u�71���B�!�'��d�/lr�j�98i��^�����9+ܗ+��P#ސ�E�/k�G�3��H�^'IK�����D�{���<��,�V��tr��(?\H���K� ?%>U'��e� sA��M�c�0`'A��8
�"�Hj�H\Ң���^S�{A��|�0�V��o,�����#����Ħ�xE��Qf��1k"G��vG���8[S��Z���"B	�V�e?I�VJY<�=m�N��(x���C~�c���?���X�]x��8]y�GA^#�KϛŸ��yoS��S��g��
?I�����܇�h~�
�/�Ձ��j�,���UY%��@�71��%u�l�̬ 4`�@wi��E,!��%g�b��]�Nă�O͐�.��`�y��
ڊd�.��WE:"�R>S�Q�QͶ��P�Tgo|!�#�4�0�����c�l=��x�d�Sv���w��|��I�0�]��h��=yr�r���3Y�'���]�.X*��_���D����X��B���)�7f��e�f��k���:Ηzٞ)�!�gu���n�!n�¿L*n�94���u )�p��������c���p@�����q�v$������C7w�Ŀ+���e.1Rd{\��cCp�7���!�bZ�:�3_�"�Ϙ�~����_��M��ڀ��%z B��G7��Η2'�;� MԊ��~%ŗU���!�R�.�<��+Bk�,k�l���~�ϾH�@�*?�a4���w.�x��sd;��?�M�6�[���X遑�����C:77)���V������eUͧ��m��Ԟis�{j�aڻⴽ�F�Vc�x^�e�U6Y���ѭRg6�W'�����P�zh��[v��7Nn+T]��O}�-�b����ɑߪ��}��`�1r�b��"�6:IBnسk˄�u���F�@�yjY��	���FD��eP�V���nR�u��Q4~ᩮ�8�#��ٷ�`��\|S8��g?��U��ϟ&L�;�ϫ߉\��E�fp.��Q�\&�ã���m�pO2��1NX�B�������ݾ���:���uH��#4�ư�k�K`��O!�4V<�O�B��R���x޶*��1�J"ʙ�/�d[{x��&��1���Aog�$��{��:����ʆ�o@:�9Jb��" "�?_��o7,
�����9����eh��`���H�g~�˕�鯗=x5�W��آ�xM&��~d� �6�?|�&���kL��������;�a5��Ao��f��޸�#�TX���3޽&�n8�����Y8^~n��j�P�nRF�6��Ts�{��ԷaI�����k[t(���M�����z�>�+Y�E=��	�+�Ů�i��P����^cz.5�ތ�[�~NG���!������c�é ����~:?�3�.*6M�K���aS{�	��#K��R��;"ް�<����!~%�_t��ɚV������ڐ�z\��
����ލ�Q�˚���o��ݏ܋?�-�!j�H��'���W�
������I��R�A�x���������[QLѢ`w0 �f�,f�#��P�]���k���虐o\4���L`6O�=�	����5�&y|��j����� ���v�c��il���U�0�q�d|yt]������H��R��ر_t��x��Q8����}���?q�w���Љ�²q�'�OFj�..$n�N,��³{���O	Y����Η���rw�=}d� �pP.�/��۲��"v�N&�CpÌ�+�:���l#l�df�yc;�C�>�H�L�	��'ڢ��#����V���ex � ���b�ϕ�"9)�C�ض�N�:�=Om�x�þ(,d�Df��<��ݶ�'�H�e�;2G�����aSS��븫sbї��YhA<�U�#d#ζ��Q��/{��y�Je�W�X�h�/>;��Z����)����A��݂UK$%@Q�\��JZ�?ȗA}K�h��K4Z=����A�9û�;����,wm�b���fp�K��~<�9厓�@�ʾ8����.�.j���D5���b�Z��r�0���8��)����I=�*�l���@Ԃ���n�r���!���bPr�b�j�nϿ2�V]aW����(?$b8��T���fw[Nz,SM��˟��,����ڳ+o�4����R?�Þ"�3�eX˥뜀�����V{�����H2"܏�6`���(JW�w!Q��8���]�WE	�i�_?`��7g�,fY&$
ow|^����)0�&���yD�\��'w@��dgR�HU�(�~�^�ۗs� � %�?�M��Ou���33��aN�
�2sT-HOC���"v�]���p�/A�d��K2+7 �Q^�]�|�Bp�7ѕ�@ɵ����>-N��#���Ru�xI��y��O��qj�<�Gl��T�B�g����Q