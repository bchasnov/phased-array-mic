��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1���e}ʲ��cg�t�ϙ�a�:�KR�%���ݧw���ȼ�D���9�g�l�@i~�].�(j_�������g�y��5�1_@����ٟ-����1}u������T�$�H6�Ȃ�h���X�ϙ������?��:F�F)�rY3,� ??X�{�E����Vy��R�7z�z�=&��4@��]���R��T��s~bb�J\	��_q���=���1�P��NfOH���m/�z���n]�,��6��d�s�4����j�� ��R��isZΜ�I����rw;�"�@$'�4h��ϽZ�MQ|C��t���w������`wO�a�NRv	�^�W^
���p�P/,�Njn7'wRGx�]W�Q�&������eN)%d#���d��6L/i�kX�g�Y�rW����sg��:95����x����J.�f�ǚ�����X�� ��ok�X!��r_p�7��ƕ _J�WXSƫ��7�B�Iж�J�J�_�Hl�W�$]v�th�gˠ	�i��

�L�8ck�T��ͦ�X}�}�tg�����g��9���"ϞN�������m����"�CksG!�O!����;b>�c͍�M��|��}���}!���[&���n�Wa,�2P���¶ ���J���3�q
���L��"��KN\�1&�6�Вui3\t�*�ǑNձo�F�]�&�x��?�5M�!�wP&�1u�w�]B�3	������NI�1
+� Lĩ���w9R�0+gu��=s��>�6�d�?��{v��|�E���f��+f�S/* oj�[i�4�R�D�S�E�Rw��-���Y-D̎\��m�(v����*�v3���B&���J1a�,��&�xa��lH�F�r��s&?��0rR)�i�����v�آ��&�@"PM����@�w�y��M&�� s�u�g�x'�I iM�>�}�o��P�-���EԤm�U6�ޫ����H�Df�Cx��̂�����ySIE�bR�4�����4D�X���G5ǞK�0��&��(��*5]y��Fdej�T�/a`V˱_�|���5H�aB����O���V���o��ٟb��F֮L�WOwGy3xf4>0rT�&���`![I@��Cf�9��1�No�.�$CP7�1.N5��5ǲv*M%���j�!��b�4�(�,Y��Z�Fa�w�ss-�	��|��ٻ	�{�Z���ε���f�9��M��`[���%(�z��8�{�K��̢�H����g�5�	&�=K[���:�1T*Y�*-<2�!txߌԯNRS�n`uD�g��+~�x���Q�Q��a���E��,��Jf
˳3�*�	�m�F�r�֯��N���d,
���+K@q�I��X�Q�R��o����kZ��l�$��ȷB�9���[��Չ\%c���l�CM?��+%��ro����LrP���Çr��f>��`�z�o��-2NB����,<�H����ۦ��`=I�;�X8!�_���$�X~@�f�H�ֵ��__�г8��P� u���X\~TP�İ����D"��{�KK�I�<�R%�\�q���hukP����(��4P >�ә�C��*�/�I�q��+^�u6��C�p°{��Mٵ�J6d�[��-�*T�ޢx/�6x3Ԧ?�C�t���Z2+c�Q�k�C�U��[��M��澬���D��k��D�����wy��o��f4���I=(ÞQ�pi�s���N�{/�$G�x/)ܦ.��$S��]�Ӱ���+��(&��@|�.B��X�APx�EÝ���x.�"]��v�j3Q3;ڇ�n���z."�=�e�H�VW�,�V�&#���dH�P��?�Ew�O�8��xaj�B%�/��6,2�I!��AJ�0�U��-?LDdm �]�>.daɕc-�����,�ly�Lr�O���O�ɛ;�p���Tc?̨=p�����e���A)���]� �L�'0��י����t$�Yi���h���Wp�ݲ�Mt+�4Zx����+kH�%*���i;ay�'���U�D���|���M�K�7�(��(	�b���D��+BW���̆�V��u���:�F٠L�Z��@�\ɡ��z�H�иW?e-#�W�霙�B!��Ǩ��p����8\m����k�����+R�WURwqB熪x!E���f��ŉ��UO��/�Ju��j]Q�"F�p��wڱZ�r��
X����I��pHs�Q�|���Q���즽���ڔ�8��BK���rh�5+�)g�յ�Q9e�FV�+�xS^4���{��a �)�Lc��
��^2���ފ^��X�;��k32Ӏ��P��/�(�/1N��M��OعN�8�0 �U�d������ȼ.�Q=�28��6�X��>3��kZ6�Sr�,"3��,Y��6;���D �\ˬ�C�E@����:�-�"����*/�\�.��h+�Q��ܤ�|�U��nr�Χ"�-F#	C� 1剸w�A7H��H��R�z�6Z~��kn���&䈟x��7�<~d'�=�_��޿m I��|�ڪ�`Vymʱ���]Y>!�x�9��gQt##|�����v!rp`�������eO6���IsD��~��5�K�Ϩg�n�n��qc޴n�c���c}�q�j��KE2���H���X�-C�ƴB&��Ơ�X/�2�2{���X�:	�?�j�W���業���N��3���6�r��%p�Lċ��[�g|���C9���\A\�����]�"��vk3����a-�>9�1{�;گ�I틫��l��uI��Ì��s���ş�A�j!�~�CI��vH��g���1�D[���*��ZPvJVx�JgU��xݧ�����<��ܞ�k�U��>l����|�ڍ+�,�]�	LE�K��=B�kOmd8��W#;ֻ<��h��gG�E(lk3,�Ъ% �ϋ2���.�=��z�dW�	���Ķ^�к�D`���@�4�p�N��i�ґ�:�$��D
s����z(���r�{�!6��S8��;�*%��s_���G�p̫̓��=�z�(��Hn����#���,�оg��e�c� q
*1L[�w͙�׈��N��n�0I�|E�^ze·��[a��@B�U�T� ��~'���N�m��G����Xl��܎5c�D椪��B�X��NV��҃䅜=i�#�M�"d�x�#���D��a~08r_����L13��;i������%9L���7�9����Y*�Ĩ�A����9����[Ę�]�K��' e��w���C|������d�P.WU֩Q��=�y1s��[�YoA/dj�&��E�bJ��&g���)s&��uk�N�S
:Dy�S�~ǆ��b�����n%*�u�R���g�$�aچ�f<9=�=&{�pLY�� ��)j^E��R���M�#�b����\�s�q�-��n�a,�6וh��k8�r{�9�X٪��Nb1���ɨFq���}e6E�!�s��)޵S'S�n���� ���m7E���~E�@w �K �E%� *��Ȫ5����L�H@�ٖq�ʛ/5���h��_h���S�B��� �f�2���f �h.dwo��,�ǓB�|a|�\��z1sgE_�{�uN""#f�%�5�U+�@���<X�G^r4�/D���HN�5M�mA�p�O��ʬ���h�K���(b%�L�2���"�{����j�!���{� �>����f��a�/���/�m
M���~�mRo'�r��'h����eR}��I)c&ZD���{�}U���`��P�����<-4� ;vb.�J��������{?%��R'�%��}�$�6S��Z�WX��w��r��_��j��J��8�	��ש�� @�D�؄�U�~��%�� ,N-��n:�����5��.c9{��
Láq�Î��(�/���H��9��E�y�/[=�3�RKfAY�_0��NGG��,$̥m5"%��\li�s���E�J��g�����y���? �P�D�{�jJ�ٝ>�ohۂ�e��>���RF�"~���`��JO��N=6�8�oq�\?��~���6PĒ2�;�����Fk���d���e8ep���n�,�UG��F�)���<�e�NLɊ�����ߌ^'�MzgX w��H��X����̜/�)�:��lspk����`+N�S��po��HϨ;�]��O�����Qˆ -�_�K �ʊ=� ��XL�3���@I/h&�@KJ�	J� �ŏ��(jO��ct��2O&oW۵clB�n^��q�C5;�bA����cA[?9�'n��\2$��0�8��!'���N �PoY[��x�����-���*��u��w*��WE�+� ��QJ&p.Q���v�	zM���U%KQkS��Ŝg_�Yj��
X��&vc�t�Q|���JL��ɫ̱��K�.��\�B�P�A�}�,�`�߈R4�-A���:����c�շ��'��͍OKo��9�&�!ɻ�1#�~kk�X�D��"�&9А��������\Xym8Y@���<{�uy�SK�Ɠ�qE�R��\�<�"Mq����Ѐđ��w� qz�����O�� ﶛ���]eVd�a������:b@�k�UM���}͇A�[xF^���-��;0��`X��7�5s ���g���6�V�D�԰�ҸhO1L61N��a�Q�M���+Z���P�C�⾝�g�!~o(�	z�֟���z���V^�U6����J�]����jmF�L�cP�U]���%�za�fm;�1Ӷ�p�������-f�^id�Ԓ�Xah�"��B�▻J>��Xەպ�2ⰩЯl)�L���V��$�lW� Ns#��� O,�h�]�l��vʝ�v7�ц��?\n���Ӟ�i��N�JN��>�T�;�) 8=�>�����Uv��gd�z��d 	
qSUx,���z؅���i��y��Il�Gs����{��*�j/ˮ�g�qngJ2�Ӂ��٬��F�s����I"u��\��_s��%��=�B�*��W�T�q��m�x�N�i�<�kC�. ����e�f�-�Y�=
s��������f���^@��Ub4�.ļ����V�#B}*R����(5��]0�ہX���*X��~'���E(�E�L���}��([��*.#�"!�͆�h��Xq�ɹ$^���4�%<f}p|��iA�cN���MϠ뻒�:S]Y6륑��+T+3�Ejg���"ѽ	Z��U�g ~%�2D�7���T�\;|����j|��ol�F>�[�����璷J7ݥ�[ng�mn8�{�����D*�_*sy�8m�c�Ɣ���=�=��O�7�f�0�E�O3���� ��ް��죗���c@��{޶_sg�6[�<.aI� p����*I�'%d04En�%�&���~ɛ�̕3B�S��h�F�'��6�ۄ�VX "��ݭ��j�2�3����<1Bb�)d	�n�`=��J!��0�Ӏ*ިjV
ã���7u7���nFrt<-�Y4���I��a���hS���$� �bt������E~^]d0��6�8cL�3N�L�i��;lbAy���%�'�Q��BEI���6o��d�Mv�~�	�}��6����Mk/ K�?�K�&�¢o�,f�ZL���EbL��NI''�_X�6௟�5����oV'��֛ҧ�
9��e��T S@��UT`�|���6�m��\N�ߒ��\&͎,r�tC���K�A�D$��{ o���eV ��	⨜L�a�B4f���.���d��W�E�g6���߶CEe6��ۏ��1 �׹֍[nXQ|@E��H�������%�8IN�*
�P��ތ.�R=�J��@��U��g�����)�9�i
$�-ڑ�G�y�O2ɫ;(.���\V��Z{��T�w��� <�e��<��;�}>�� ��(;;�z�C�~�����~>�jA���`��g�2~y���1�����~�+T�'H�����['W���׌�`�^�:�.���9� ,#�K�s4�W\��'�����;Lϩ d����i�_�C�|)�1���b�3���;5����s�xh�|X^�8�x��������& +9�i�I�2��Vtuy��Gŏ�t9���o[��*�$�/L�S\D���(��s4���=����+�m����0Zzʠ����d�Kq��	�}����V���ԡ��K=��F�!�̴����Y=�r֦ ��F�L��Of��z��9õX�<�n�g�2�E8ȱ�	�2�����F��Y�ꖭ��]F��y��q�Ô����&�q�2�ނ�ZS 	��l�Yst�E=
�j5�B���nx�5�Q=t$���z�gh�*�m+��ԃ��;-�WB �5�$�L*�����#>��&�-�`�jb�_�R�/�Naȇ��s�|���)x�0`���$�F��>�"̢p��_HMy�~��O�j��%��/zv�:��R���z�*�)��W/�i�v� ��}6.�U_x�+��3ODK���ʤZ4<��>=�	�< يj�g�	ʩ}4ٯY?�$� q(��G�8�4�b/f���\��U��2����{���0�f`��Ps�+JO垳L����u�r�D*�a���R3���{9��Z�C� �F:*H���D����������Q�1߄n�C�����?�^NO��ď�����b��l�)#\e�v�L){ƚte*�!�<sY�\����C�~�����kGȤ��Śe�G����e[v���Ҥ!cD�C;�nL���+�[W��mj\/ʘ/;�iF����WZ�׽��}e^�_�)��?�?)�jc*��
�cͼ14�� ��t�5�^D�.
�D~6Ya�`���ݸ��`��Zɻ��D�Ls��������<���za�w��f��(4E�Zt=\�ܩ\��QO�|���s�w�G"$�b�C�)Fk�t�؁��CƆ�1آ��3j̪��ۇ4�l�雟�]sHRAK����Opp 'j.f* ��V��	�?86���E��[�p�{L�&�d� �+�do�`D����8i����jY>j��<2@iQGj����Ch���}W?�WUB���S�
��� ��
�J���Ά 3�;�%�vt�˩�$�5TjW*p���	�v%x1�tt\|��H���6{�Yy�#v78m.������ZA���Q���^�C9�Bݷn����I���o���9v�W��h^Fvb@7�����zb��\z�P�����	�<����K��G�u�Ǎ�����)�A�������D�hJy˂����*��"63͏��`�'Ω4�zg�9曜�����U�>#�P����0N��Pxm
[���m
j�b9:>Y5�]�x9��[d��6��櫒���%��9R7�&�vA�(����2,r$�\L����������ͅ���Ж�s����4��l5�m�T.�e�w�$�ܓW;�|E9ܜ<��e��ܺ�����l���|g�"�D��B���J_�2���V"����Y_|$����*���*�۵X�~��ŝ��g�	g:���,T\|�k���?5��!�FnV즳��\eqS����i��5[U�m��&u���D�[q�)Q]�ɔ_3hU��IOvK�DA!""��6��$������}u�ܓNh�
u�[3�zU��n�k���+��z}�=CF��s������W���0)�qv�����-�xq�z ,\��:��y��㬾��g�ޘud�7kx���5':�8���K�x������j���$Rx�^V3�&��&s}���k��C	�w�WԫE:gK��w����LW��@T�L�OXd30ӈ����೮����Iʤ�ሬ��F&���uÍ-�)(wa&�[�!�{ͤ���e/=��>������ܹ�S�� 	M.��U�z%�*u�kP�A{4٥��N��?����p�a�[=�� (��M��Z'�틼T���ǚ��?N��><cÒEpL�J�Js�9��C��zt#�9:d�����hc ToP�7�̻��F� �t��o�+Q���P@0ֳ���� .\-��
�󯔉���v	��:O�yur�*�n)7NSr��-V�mH����,���\)�S^���mmu:�3F��D3k���Bu$��m<�TQ���t�>F��j�H;�I¸���#���DP�h|����m��S�nh��Q�u�$v��օ�71��u]%��Wo��(�Gy�R!r�C�-^/#��n!$�}��^x@�m帨�2��5�{K�$f�3�^���T�&���ل�]����S1�D���Lk�֨�_ ���kO��&V�5�fa{��sظ�"۶V��/f���LQ��#��b�	���kh��Ma.�y�U����h*���	1�Xqf�~��خ��+�B�6����	FlD���I�<�{�\-��nL�ӏ�g�� s�Ͼ{R��<�U�	i�JYAGɚ�"����3Ӊ�F�չ�����5���1��_�NŐuz��AL,X�"�mx��6y��M�BZj8�2krl�ϛtb�\Rq���1w����2
�x^����U�\�����<\��}@K�&0���b�4}��0l�fUB;��/>�9�w�8`aB���2�)�Ҭ@ao�JȒ7�Ě��D���W%r{*���s�x�(��ju������'�Բ��3��hs�;9��C"�&xN�����z�ǹ�ɪVF��6�ELԼʥ��t�:`�ǗZ�Iu�؛� Iz��d�߾V���Y��t�C���yWN%�MWT�~K��=������Y���D�Ml�β>r@yW��#��E�����d~mpM���j�Z����e�W�2�2�<ak��_/g��|�ĺ9�2����R����|������4�H!��u����[Q�E)�D�bZndf}���d��B�'�/X��s��T�f'��SC�7�L��11�;��i�9��zۦ3BI}�ex6�$,���ߋA�R�,�v(xr))<�l��~�*9�Y dI���C��x\M��8<:]�{�d>S�۫Sx��HQkXh����9��(7�>���zH�,EE 
�Ȇ �$���Te�*B�D��@����f�{7��2���T^�,܍`��9:`߭pkӗE��^e5n�U?˼?-3����}�2��W�A%]�x����	�1�N����[�ڈP̤t��r��;=�Xۦ2����ڔ��>���<��G
)	!ܸʅ�t>[�0#B��vN��k�
b���5 ��gd?TA��x�?�o�{�H,�,B.�"�٥w���
5Ʊ#���G����W˩���o{�o�}�����l�~�g��鉑�-����5I��\�#6��N2�gF +��&# �^�}�'�5ck��׮͉B5Z�E��g�&�u�	W�=�Cl��L�rkToݝmf9�M<��RG�����������j���e ��0N{O7+p�(��C{��i���$�^veɉ�v��a�BоVF\ps��e�G֤��i��P�i0T.Ǥ.
]��%�����T5��G��O�O�����q���کE�k�!��	<>�0����UUxw� 	ӑ��%����[�@��?c�p�C���� �_6�GR��j(Ӭb�*F�@�#?���h�"�0)�,�u�n�U;�}>��犡�嗔���ŵ�c�K�S�Sw�yTJr�\#�!�QXZ=q�KC�ñ�7�.EE"U���!͸�ȴ)�PZ����s3�����q��a!�,�jB�0����ZAE��m	�f"r�\�	��v��ϴ�:�&y��P�^�KJ�x�?�)� Z?x�Z��˛�ܭ!�X�q�^���{� �Ӄ$�M���9݆����_L�./us�!�b�u��"cT^C�{"��:,�Hv ���j��fr4w��@��5�Ґ������1����(	=���C=w�p�t��[1�;���%h�s��U�EL|P;4d(r&���3�$D���%m�x�tec�LG�5��tKT��]�ȷ2�lBiv|�%�`�n��.���kz�T|�{�hN� ;e�8y�gK�(�����:z�߂Zw��qX�B|=��b�M����~J0�ޖ]0���q$&1P��ך��+��>�9��e��9��Q���`�Z� �Տ�0Z��k��|s�����6j��<��l�l� �R�� �@���I�j�a���%�V9��ff��>���e:�Uƈ  ��3d��C���Q�b�f����W����M��?א�Գ�^�����*����=���KB�.A��Q��B?�����Ų:!4����+�:k����kTʈ9���&�*P=�㇕ۍ���ɚK�h,xW:X����g·[qurܪ��>�6����kޓ�ԟ3확��|��ͨ���������e�F	�7�9� $���|��4����$�|~�Fn�x�,����d���W�l�'5@{�c�ǰ	�%���Z�_ћ����J4���V�����=F���O )��ʩu����W?�6�����Ct}�����iϽ�ʡ�Mԍpg�T�d;�_Sz�a);ڶ��˹���q���0��p<��+�8w�F��-�fE��q.��CݎPY�1I�r���u<�$�ـ���5*��{���r�W8W�mb�\.ޒ�[wH�c��;��YEt�̔Ա����
ˀd�8sv~��%2���ʭ�ɣX�O��t�+j0A����rr��v�WZ@�Q���]���)]Q:��Î��I�\IݘG��v�r�����w9R9���M�>��z�q��N�*ȟ	X�}C�,�uW��K?[ˎ����nT"T�&u� ��詣��f�V��mJ��L�ش���	�S.���*:B�o���|¸�3�po`VG >���Y;�@���{a��"�M�O~���C����.�K �vCF�0F��j"�) ����#}zJ-��rǻ�!!,9x)��q?��u�k�7C�N�D���[����ŋ�V�u��C&;y�0���Qs��"���B��aw�P�
@��u�v�0Z*Ӻ�3SU�@;~����B҃�lv["qʟ�^�fon=0����?ZO\mTW�X��η�%������;���"�kǣ?���ƫn�%�T�_��5]�KQ�����D�m����sN��(3��]�`���x��m�ˋ�i��p�Ix��I�O
�M�*�^p��Q�%۷O��p� Lq�~�u��16�Hk(1�f�D���J�u�� x
]S?�=�H�\���������m��J�t
2�Cm�Ǭ�[v�X)���(��U��(���P�Qjۙ�3���J�M�)����/K�-0�Y>'q��N@J|��fF[L0�u�h�f�z=.��9L�$NL���q;��D�ʐ����8��N�����W!�:֎���N�vԋ<+�U��N�n�D�/���u_a�&Vq�X�)P�jQԋ�����8Y~o��D�f~!���<10���g��(�6�սB�[�;_Z�j����֦n��T��>�d}�vtP�%D�O��&PJ�g�|���~�8	ޑ��-��o~���0�$z+ޔ�����̭cSk������u�j�_�u�Z��;#Us��2#&�{��\l��*U�ߎ�n.��A��N�}��oU�)��=)ac����9C����(��6ׂ��|���)��e������b$z"��{���v�dc����<8s��,���#���uޅ�Ⱦ�j�F�<!Ca�2C��0(���P�:��dm�1٭��v��
I)����v�� 
�iKʭR��0Z�� 퀞xD�.�*���uE���ѩ�S��!��i��+(�}�!oE'v�aJ�>�z�'dH�N&7 6Y��>"�6k��w�k$U?.{˨$��Γ[�f���Jz�
�gͧ�K�/A�<泱l"܁����H�z9/������x�I)}n��"�m=@�q�,,�"�X�� ,���?�_�'���~����t�����i�O�)08^:Ih��V��(͢!��1�X@���5|*C�����\㮟{G�t�AU���-��,όٳV��)�Y`��y�j`z�ܷ����X��B3�H��+W�MIJș�B�j��8^3��WH���i6����R\�k��.�)�L���7xYm�_��j���Bb�/\~�"�)��P�N�x.�v�����z��?M�B��YN�S��c�EyFN�*[56�6tyx��y�z!�ΰ�����('�e&�S9��&b"~�M(�sA��{��f`��le��ґ�o`hwÎ[�,<6i�V�[��՘����Ό���}�x����δW�`7�9���p[�(��H���K��hqo�<����Շ�;���p��A�⮏��i���{2~�&)���|s�ͨ_4ŝ-C��S�~)7�Zb�5uXW�>���v|��~�������㘭�dd���E�F|�N(�{��~eUn��#�����2�k��rSU�3�_*��V��\B.��826�o�8ّ)��7��U��ɕ��81s����s��yņA��%��'��#/�Yeq�n�=��t`�i��#�<�)kٴ\z�]��/�k��qN��ʻ����6j"���X�(LI����%yR� �I,қ�Ј��,~���33O;�0�$E�0�\iв{lҺj�zMQ��i�����P����?!jm��=<X �ʉQ?�k��F?&�Ib��b�Jw ��xF������/����{��KJ�p�r�,mi$}ԩ�{~�b�guQm�,��/O���S��]����!�������׈`J�aW�'Vj��4����ͬ�U�@�_�
'Wj�]���I�������=�7��U��W�
s�jo�މΊ�û1�o�Bs�b��)5	�2�,��Ez��E ^Bl渌�q�����(�-�rq)���e���B��m��p�M i(���Ȳ�7z����C��,�YȪ���¦^���7�ڍn�}t>E0?-7�B��Mϭ��M\�;/L��ǔ��g���>S�PG��ב1f8h{��kG��(Λt[��x����/��s>x�>�i���	��Xl䱶P��w�T+a�K</p	�y��!�ֹ �Jn|LŅ��H��;�Q��|�6�6B�5�*ł-VnSkԚ�M��f�;g6ՎQ���4t�F�`�w��6S��+Rn!V	��fZ���;������D��	Y��^�3/8<�m�Aand5���w "	q�	�=!�y�4w^^�w4/$S��;�8t�*vF.�
�R����[��G�3C��"Tc��^����9n�B�؇��JR_��K����2~�����P\��Y3�J˫h�����G��aІw�MF�����Mk��չ!�b��Z�N�fğ刽ʰ���fn�/ް@�j�X�m��g��� �G`AR0kd֭qԑ˖���ݝ�%�R���K�>�)'h"�!�%���6�9��"���Tj/������6&Ʌ�)C݆�$?��Ӣ����2��KVH1�8Ya����+G�Ջ�S�Rv�o7�0�6b:ő��A��J�	�OW�OT����'�hv�NS~)����Me�ũ��q:��y8Ҷp1M�>��އ�Fҧ��>K�
%)["@�U��- �>cbs����x�߾Ԝ�����F�>7���u^R�6��7:֔��?�'j\9>�S*��I:�H�:)gQۂ|��a�2�6o�zF�.n��/�/ 8F>E�l��f8+YBܜ���z+�2�b6�}/�io
=s�Z�h�J���9�p�8L7���O�~�1>��kp���̇��ֈ2�%-�i`�Pg��g��`>mX�˪,c�1)ཹ;`���ۘ�Dw�"7�X�ͅo��*hv��K��|B��	�B�	 �`�O��m�FuV)#��Xd�7�6��$%��W [2�Ƴ)��!+������$�/
����2{�&F�:J	4yO23K�i8^p��s�n�@k|3�~�H1�Zjԡ��z����vK���SS�c��8�v59�vOF<{��y9����H�����L�o$���h�h�
��[И��bp��ԥ��n�]@�V��r�(��;�֞x?~�ݹNM.����m�މ���_m��)r�Py	7��4�tH��e���0:β�ț�_+�qv�yyg#������h��|
������L[H(�(���;��S�h+۷��p�?��*`,x�$x�&�?��M�v��jʊe���Q��%_�9�X>-trbD�ZW]5��a+���p�"0L{@$�ˆ@����� 9
Z��Y����mcٹU�h%y%qjz˿Sx6NG<<�.�	�T�b��.T��Kl;A"�L��;�E���U�&��>X&�x��@8 B����&�E�v��;H���p¸n�O�ӻ.�.fgkV��f���V�d�TP�NL���i$ڥ,�����EȊ��Ss|�ڠX�2�Xc��Tӈ��o���R��@P��WN���9�ru��wi)��r�	U߃�"�$0=��\)>���$i�X��25�ϭB�#8���$��*Y3�*�l���օ�1�K?UO��Z)@�[u�d�<|V�c�%:WO��c%d����:`��E���ܣ���5�
we]�@������U٨����W ����\�h��UR7q��E1I&���|�$&�Mvm��q�	��m�f/�I�ݣj߮g;"<�5_��Sh��ᯇ���z��3�S���B��^�������1)�?w�57�>�|�@�R��h�4E8>H2qC�����K���ɞ��j�/�wG��b�]h�<#Lc�����1�MG�����'V�;�ԅ�+���-�U��V�N���\��k���`7n($ĭg��E�G����E.!8ɧ:ٸ�>���ġta="�V@]+m��8���.Sa`
�̏ �$���X��4��W� �@<�N�cΧ���L����|6�}:�ݼ�z��$פk���,m�D����b�8%���fB��/��`]�t�h|�/<bd�.�� �	���1�e7 suC���*\,1`R.�����Hɔ�~7��-2#��� 	zL^��O����q'�@��5�O��N~F(O>l���� Iδ(_w{�ڞ};�D�#�V���~6� ��6RYo#��$�V�%3ZV'z������y�,���$��[ހ׎S�]S&�B�Ty�v����(��OB@�)��|�N�Ϝ��e.�{ʟ~Ӈ�~|b*��D�}�ۗ��O�?g.�G��u�d}�G��K��r/���;�������)YN.�\���M�Rw���-���g��ճi޿ ?�R|s���q��"+�*���XZ
I*�U4='.�7E=9��I�7a�h-�X^�R<��Eq�s��v۵(��a@Z�Q�tM*:�ऎ�m��s���0^8�Z���yw����I`	6~ل�@�s�ӕ���^?�h��~2}N,�I�E���ǚʉ9[:�u "��^
�~�2:��M(8t��â\	"P���򄔙zN&n��0��bQl�9���i����u���1W��]�!>�5۟� ���S"ü�a$}3c�M}�����"ѻ���L���7�Õ���T�K>�+P��w��!�X��^�,F*��\"Թ@�m
���w����(k�$���#��a�Pa�ܳ���������`�@R�r�rNa��ŗ�Ф��J�`YXjh�k�i�n�-�� ���~��q�ʡ�\��K4�txdח���kHV�F�I L�8p٧zŉhj�uO�z�g�i�1�=+�*�;9�<	��P��9t��>,���h�h ������bƇ-��h$K�A���yOI�� sR%s�ZXx�cmx�{@�  ����ĩ�Y������ٺcB�̍>Y|�/]�	h'��<��k�R(��Iڔ\#��_X��n����C �ɘh2O$Պ��]��µRW��y�̥�+Ϫ����z'�K�)Ǆ�
e�,�@`�T�^d��#d�� 
��~B��`�Eb��`��i�%C�Ң�"�eIgl�5��eօ�|<c�B�^j2��dE,�4'P@q���>�Ε6b|B���/.JǦYJ��m�ׅ勴hʼ��	Nb�����_Ֆ�4M�����-�g?����L������#)Î��\1�z���~����z/DF=�A�\u�.��ۖ%�H��ƺ�D���(�������^Fih�XP�'��\BNhY@"!/�m�\�a�\�8u%�ءR� j	(�ӱ�g:O�۪oZg���*��!mY7���b�V�d����W����Ao�,C8v��:�X(
n�e�w��Ȏqk�zC���bɠ1�^�eƹC��t�w���xob7wm�k��������7��� X~�>3*�E0��&��5��?��n���&Ɇ4��p�}f_(�'�K&�*h��Gb�q��C���� �����?�<�/�C�(�dȒ�+R�őO�I��?� ZD@�2��1ܦP�f�bS}�wӻ�ې���U����n� e�] �hw���츪r6�UB�d��Zp�6�� c��S�qJ����W�y()ҵ��`[��h��p��Y���hT$L���_��aF+�$����m��qK�Ǟ?�'��Gl?��59�~��}d:�K]Wj"e���ۉ����G�͹~�R�3^=�F�t|/u�}�rP'�$}���#;�)ׁ��"��SH,�{M-;�����2�.�ͭׯ�@�9����R	��'��wl�>R+� �sz��#9����.�d�KM'��J�(�\�L��W}��W��V,���!�=�~@��'v[,��
cY�3��lȍǅa���U"G��d�����g�(�����t��M��!�?�ft�(}t���<3	0uCv��}�����[�T5��������`��ǆ�Yj
���G�EI�Bz!��*�a�-�n.�p�[胢%R�П_~�0�k�xHp4a�p��~.^\�d+?�*^�=v�zݷ�d|t��z���'$��>���Tz������|�����A��G���@*�4&8!�d��*�i�=���F�ܷ ���6���k�6�߬<���ו2w�̦�K`y�fo4�q��#U-�w�W/�5_�G*g�(�|:.JJu�"[�u��xR���֣� 	�q�TU�.[R_x5�Fr����H����A��7lIӎ�2SV]@	��f���|]	�f���
|��.��NU��p����u�XVo�B図�'Z@ZSj� �����L���_�6�u����$`�����3}M7��¨M�m�{�V[�@�`���U���������k�.�X���������+թC�׵w#ӴD�u}yz��DN��R��EYv9|����~uP��3t�0|���/���:$���,:�Hkح�������H���E�����4pu�^��q�vtj���b��'6��-1��P����q6ҁ|\��s�|��.�b톌�7_(��h�~إa}g_=���;.�G=m�:�v<̦�E�^��Ę)� t�J��g�h�r�`KkoǢ	� oJ8f�p�=y�G��[3n���}�^s�>���?j�>tč�%gs�'�х g%�+vkt��|R��Zi{�`���GJ��
jgǳ�f���ZoBq��� HMɞ�cq�	QeG��(����8�ޑ��k�>eF��d��F!�<�ÿ>����ff?��������_���+���l����Ʈ��K`L�
\���n�9��9�f��9&��X6^|{�i4�WP��� Ӱtl3��U9u�z<���?���0�`��n�����ou��L�g����@T���+�F{�M ��#Yw���f��(�Tx��j;W�A�ާ>>��h)_�1=�#�'����K,ɷ��dԸ���F���>��9,���p�l�j&=
8CA�{����$�/'���jx�� 3�_�����LhS�8t�:��V���9<��d��(lܴ�K��Uo��:y���T�{���:��̔P��TA*�`x�Pך��QSb
�-1>h����\�K��XL����[�{aN话1|�ۙ.���� prO��]qS�v��C��?d���5$.;�ַ�3X��-��#�Br�M-(d	y<Ƥ>���G�U+��$���m���F��.�h\к��7�Y-
ֆ���(�o;�7e2��9�`�٭��z�oJ�l��.r����[���WI6�yj[��9�u�qdס+�H�[D�Kw{(�儁}Ǌ�����05T9a1�>t�2\z�:	���C5������i�Bջ<�!K��w�Cf������y��}5���i�Xc�a�*�^�;o|J?�W�X	�z�!����{�(�w]"=�>�w�X$`@�o/���L<JG�{�J�O����7��w0�|�����_f���ր!��:zݿ�w�4��ū�����^���jx[���y~��H�	:��@l���%)a��Vwu]�3w�$�9������,������aD�K�X(͎��D\F�[h$��*��f��q�Y8��/�A�fp��=���=-���mu���ƼS�T/p5a�	�mDb�#E�<�w��,�0�*%-ݚ���ף��p�@�8|���*ũ�#�%U��F�q�p_���
l�Y>_� l��9tT	yTp�mg���It�JppeW�o��u�R�X��4�u�H`h�����O����	;(��X
�=�Br�,c�Ѝ��ur��gz��F�46c�'(K�D�Qc�I��%�FQ���V;wܬW:�^+���un^�j�� ˥ԋ�\U��т�b�$|�:�e�7OĳU��Lш��i�D�����8���0�<����y�n�~�����!��4g2��S�]JUd�`��ż�G����h#�v"�ْ���H�@���w�]-r��)���w�b���*�C� �̣�h!�!��Q2����A���-��M(5�,�/s^!Tv����E��x����%lZYwb�����~.]N�F�y��[�[�=�	-F��M��.�ʖ�TD3�K]���C�ZX�E�7D_���z��0$�$�1�Ml���N���i#߉�ף {�hj����;O�2�n=>��a�E�+����M�,Z�u��'���;����G�o��c	t��ُv��cV��"�y"~Ь��<���OL��j��f�$�7�~��_��}������U�;-�O��bJ��Мm����:��b|�kc�9�>�˅��Kf��S'+�=�� �ݠ��Z��n]|��;"5i=�%:���W'��GQ�s�a{nrxpɚ
��(��tj-��@ ��!�Yf:����>�ձ���7S�.S�|��ܼ�,�s ��ܜ
<����N-��dA�V�G�<�#Л8sR,���W���Ut̐9^%bPh.���
�xݯ�����*�z<k:�\�iz#��M���7����jC���W���*,;�}��B��m�Z��)��;֊ʤ/��?�t�:�7� �l|�P��;D��}���O��BA1J��>L�M*=!P�KK
���8��@�3��@�CBԓ�.��$�?ע�Wcw��\ �Z���� ��NvL6��cigъ�A��������!�&Ui���=�j�w�T䂢P�R����T���嗾Kk�5���V1�a�G'��/��1,Of\�+Ł�=x���dW��n-ۅ'�A��7�Z��ƽ��,����kx�US 5P�}��9R�����~�[���$�T��Yܪ��ąy��61_[������C:N"���E�կ/C�=w�O�uH��6D��^�|T�5���°$Ϸg�]���c�}��1���!ڀk5FV�4}m��\4"oV��]�e��{��﵇��UѴ�@�8��5OA���op��!�����qK�Ȓ��d�����Q�`�.J���j��c����g�R��[��ց��Q�{K��Y���Y'J���>hc��d�~D���1�Cv���ݬ�_W��q���/���J��dx^%��`�A�6��d�w[���E�i8�����'�kH�e�1��2�ݗe��AHЍ9�1��~�d,�5oJ�gv55|�g�����0��Ū�I��Hpa5�[i�� X�6a_s���(3#�Ҽ���S��Ȳ�:��J�E֖�uV?J�j�j�Ӓ�&u)�6�W��B�-6��D��;�je���� �-ߩ�K�����
y5A���~k���<���~&8��g~6P˦�->r&����p?�b�&6M*�&��u�pV��n�'A���(�O�%��O��}B܊��ʜ�")w$V����;�����;�a��豉�"�y�$�&cc�͊��ŕR�v�z4, �!����t��� '�yRo������`��N�j��
�k�ǭӴ��zGm����JklH�t�v?�����֔ ù
fG3��\�����zĳ��
_�0{2��\�#a���ls�E�tFR�}�j�@[-T����=l([�}�͔}}���p`�7��^\�زeȼ�L�/{�}=�����٘p|��6>��=4��'ۤrǏ���yDS��z# ��'C�����ȥ�X�j��>�yQG̺���i��$d�r@���R`7�	WE�:w��[o.*�aW �(���V�;H���.�a;�ҮKF8S��T�X��@�MH�<G�y�&��K.8����*p����4� '��wu���fCI`\�o�~+�A�*߆�uz�$k�/�������N�z����qH�|��z�`G.5��2�,H#��e��iW��u�����A�J")��X�kR�@���$4� IO���u���eN1,es4<s��C 5.�ς$�'5d��a�੅�64�=�S�\\x/R�4��L�q��~C���l����=�q������j!%�F%J���Ov׻��\���њ+v�,����T����x�y+@�"ѽ�Cah�Q!�Q�?�C�s����=�g9`-+��p�f������h��R�UY^i�fB�H&fR�8&�@��Vl��:i{o{+�e��{�m�]���O��fl����Ϡ�ᐃE��T�Z��.���E���U�x� ���ߞ���D��{����N�%���ah�f܊@�����+�����n
X}��{�#���έꄵ�ҷb��d���Ԍ��R���
��-� ��r�a�{2,�!���-�8�)4����ۃ�fj�~g����o	!�������V�%�
t�W/c8�� �A��ޡ��}z-^�{�F���P�}��Zx�I#��$.���lo|�u�_���Zk<�&��ΐ3�1����o(������1n�n�� E�{~S~x㲈��
)�dV�e4�w �,�X��5�C�Aȹ-ݝ�@=ra��3�V}���Ķ�X�M�=���s=d�K��%�-��z�HY�ݭh�)��3h��^����hIN���j�O�0U(�m; 6��FQ�"�]pũ~�ͷj-�|��, �����9k�a!�V��p�@�ef
�؀�0ִ��A�#��$ #�vb��ʔ�c^$���7�+se7�����=D�����	(Sƍ�0��FZ}���ܙ\�˛d�o�C	�w%��h�WEy���,!�D�ѐ��I'�iώH��M,D
h2�`~��O���]p����3��贸�>��r�������v���m
�&}����U�Ҥ�hD!��وv�S�f�{Ԑ��/^����qMcz�#��H�5l�u�u�1F��x��#�/#p�҄O���)��*Q]�>��v:M��ݏ@`N�A�}��ɜg��4N�}(���� ��c�u5��ў�\TB���.��·�\�F��"bjy<���D��nX�����?������@H��ru�<!���5��r�1��!�+4�),Y*`��!��a&Bڔ�G�\(�줮��z>(1mR��-d�-Yv{B���߆�fƀ^�A_7���E��ox'���D�20����f��t�JF8]D��"U��P���[��?hHf�友�=�2��]�F�>c�:k��Q���\��g�_^;���vf�zv��!�ȭG���{w��)�qx�H�$������!��s���(,[hk�¡C� 0?Q�w�`�=��7����=f���K����6V�$Z��%.���[�kҜ��=$��$���c�}繪թ8Hq���2��n�B]�������>�����c9�|H�ͬ����g���*g����kq�e��P���z�Y�ނ�n�E��� �kQ*��8�����6��x����ğ��G5b9!b��8�K��[m ���R�-q!�g�NGv.e��q���2Kk�5��H�!�FA�|�2�R<��DPl���#��Z� �x�Jm�{r�h6�Y�t�SC�Z�>�F�v�f#��&tЗHWJc��ذ+A��֋h�ߗ_��
Tys9�n8�\�Z�'�D�#�/�ƣ��0��E+�����[�w�+��ڱ�u���Dć��Do��C0Z�V��a��~�%�0������mv���A"��9�Dn��ɢm��z���/�AC�ڑkV�����������znH�z�腢XY!8uHr{"i"5��~��a�\0.���8�gj�0<Ϡw�����tODe�Y"�"Ӳ�X��&Ef����+	��=˘٧Eҧ���4�X�g�r���<B=S���԰��#�L!���p�x�c7[B���gL�vC��뭴��'�*p����(:h��f�c-r���j2�`���^I�F��%�ɮ�\���� b����׵8_i@0�ٵ}=M�9������a���X�0��T��^ �5�]��]ٜę��^��zp�c!~G_ѴWp��ソi���i&�။�;6eY��&p��Rb�����5�dYc�+$O���)�m�@��n�����J��g�e}�f�%�a�mvo`�Ȓ�����	�
�=�t�q�H��ט2!�՘�D����B&��O��<�Ĉť��(��}�Tf�"xXf� ��@6#Y�x�p�}=�¬wI�!j,ka�w��5���t�5��7��z��B�8<��gɀk[#6t��<k�rb|*ȍ��^�[�c��}����K�?:�΍��R�ϒ��L�Q
ߵ��)��(:$ʍIJaf��l�ܱ>��٥j:cn@�)���)R޸�|�q;<�C4�ܚ�+���w�V^{���I^�͇M��d��[�`Ns���um\��T��7Z �L�ŮYԂ~D�c�e�b>
�8IA6�Op�z���5M�����/�-[�o��{�1V����?�K�â�+5Ч$���iN�cy�&���k����~s�ѕ��s��r��w;c��g�_f����cp;���E�UL&_aX���j�3G`V�ac�֋�����
l���ҘneUӨ�,�Z�����xx];�3B�ֽ�&���Q��J�������v�7�A��]MB!崱���sY�y��d`aƼ���!����:��Y�S���{'����\F���f�GS���֓Ir�c��]*�HxS��7�?�xn�|#���BҘ
7��Xf��k���=��p�IK�јq�����<�t[��5��g��V��5�����Z�����W٤~�l�JM ��LGʒ3�l��K�4T�d��8�o
U�,�f�I��������?
؏h�։�o�c(�1��`��"R˴<�f���ef2���gأ��.r�6�i��0�Z��=� ��za�=�!$��V\bH�w���`>l��K�pW�4{��MiH,XY������O\�z��0��|�cV�>����Lt����n:�|2�#�K����]���i/G�a�
9<�ҷ��U�����lW`e�2u�K*I�8x�4*�����=P�]��Q���&R��Ja����-n���<�V�w>(䊌=�S���W6�@@K��Զ����m�"��掖�'G�Z���Y}o�X2ޗ�D,M+���+3�w��cW�8��"�V���6	�D�0R���A ��MCffj��xDt�"\F��/�ހ��.u���7y%Z�\��k��}�9Ǆ���F��.lVZ�`ױQ0�b��~4����&�{
��".��װ�˾0�/ꈉ�3��U��G�����Xd��:��$Ǹ��;�e��>g�௯�����`�y��ͅ�m�A��ɳ!G[��T�SQ&a�J��ǲ��<�e#+`��?����ġk�mF.z����Z����W<��ǽ�	�W8p�ѓF�9��պ}ZO��6��@PE�����b�RmqZ�ն��x0�hp���7y ���^v����j��mCI��0�}�j�b�����Q��6��#	K�	��N�����@vA��p�Q�7�w�0:W~zj�;��4uR榑o�P�r+��4�����>�ϥ�[�&0P;P��ޙv�
�Qwů��Ξ��Կ����Ga��D8p��$q g~3v	�)�wc��-Ld��{N�1�#�\�R�������������"��ӻ`��*���c������Z�n
�������>�Ó��W,��M�BO��+�_���ʏ�8ZM_|�lt��,H�*�N���'ꦩ��������C��O.]�����e�8��j�I?N��5S�1�r�-u9�Gc��.ѧ�)�uZf��.��_�$���J"��&6֊Wn�7�3/�	[�4Y��ĆLe=��ÎH;�������k_�&��h�w�9@�Z�
�����<[�VI���}.U���o%ã
�<����7�r��m�Y��	�H�6F{�}��IN����J��� ��(r.�G���gVza�f0V�eܹ��}j�
��Y ���,��VM�)�>��'b��eA�*&��L���Ԋ�$Y2}Ȱ�4��;!L�|/�ʯj�GU�y���=���6F۲z^���6xf��:��Ga�E��Z�%���E]�Y t�sC�+�5z7�51�z���ȺjIZD�0�����lOB~��X�Ds�17�H?����H\��	�Ӧ�h9��<f�'��h�;4Q�5'�#�>MNI�����^U�:�۽s��$�HH��tp�(&0S�3_��5��_�^�ߑ�Z�p<��q��}����a%<M��$eC@���x�ѭL�WGl|��Y��$�T\z��)���c����\�$���Y�\�Tq�D��Q#���X< ?�0�"�;~��P~��ƕ
�3�Ew��~�s��j7��"��@2e�.~1u�<}���-x�������f��x�̈́jO�l�П�q��K�f����V ��ߑ��xE��m
}��_y`����l���a��v�����3��E�@ƺ"�{�����L�����^+�X@������c���6��9�W����Q�G��Q�j��07yXl��[K}��	�����F��@C��|M{�U���e���8˜%?�db���2C�:�U�"���Wl���ɶV��pL��9;��ڊY��sɈlV+�cN����(N7&1g\��1ك�̶a��������gi^t��j����U����gQ!��D�� ������u�q�"�om�~i#y17�M3����t�r\��oR:�?]1��k^d��E�W'm\��{d˚�h�w��o)��@]���YIg��.����`���fr`�X��Z��~��
y�:��y
��3�V���~��0]u�����^��a�ʨ�$KjKD h8D��u�� )���1~�8����[śt��މ�E���X�	��p��(�|�(E�i����i��p����!f{p�k�(ÌU!B�[�@A�_�_�W�"�[��S u����?UH��ti��@�K���Ej���BjD1:��O�(��\�a��{��i����mދ���� �\M>�ʓm0��aD� `�ҵ9����F�ۗp$%8̔]$?"h�b1)mY�6]/��sG%������iD ��I�.�
��%t��o���.�@�Q��Y_�yOy��;n���C�S�%��%6�hkm��j����by$4�
��!,�D^O(�S$6�A���5�}����f�t�x�ӊ:7~���J��	敏�%wʦ�ُ��}A��av����\��O'�_.6��K|����Ѯ�'Q�;)��Fz��J�c�!�_�ũ\��MT���_N4��M��F�]3��������,�����=,qӌ��2���;9;��	�KB̅��60<�xX������޳�t���_�0Z<��Rq�V~�y�MS�d�����r��� r}K�$vR>�����4�@���l�f63��B�2���w-+2?۔��"��"�\��D������DhPԮ�P��%a�ؿ5��o�ZJG�T\v��o�j��{�l���J�j�3��CYA]�_��\]j������gٚ }��Qã/�PA`G̻:v���ȶ��8�;[���FW�ԏB����Xs��մ&y�~��j���Ca�aq*��L�γ�[p���%e���`�l�6,ĢEeAO��`��<�/d�Nr�'n/_���)_d�!��������?s�԰�_�鞳�!������}y+O�X�����+ar��W�Q�{�PĻXi.��\��� ڟ�+�^ߦ	j���Ϣ�#�R��P�����	s��I2<�?^*ꄶm��ïw��C3��C?<qfq3>�*wGd�Z��a�	
�z�)v��O������	.8�A�7r�(��Z�ndm��$d����&�DB���{�=��e�`4B�0>���%�}�{�1��奄��\׬&a���%�.�W�.n�B)�w$�8I�_����Ƕ8 >�4w���/��!�� ��j�g�Uud�ϟOI��)�O~��t�0tj�C]dh�	xq+i�91�݈��0��/$���c�ߍE	�Zx�����PĽ����&�������l��b -�K��?�����B]8��D�!���ז�E7�!��/�잘����N
��\+�J��w����O�-���ͻ��/<��G��_t_H�U��O��jK�<��M(W�R���񄯙�f
а �I� dh'���%�|�o�d�_r�g4H~�A�IKQLSB��մ\��1��=��E���uc�D�����f����L�v+㙖E,ĦZ��d���=L�`�����IB* ���:�05�8qFNkd�|,q��uߟN�s���� z�I��CS� �N��J���*�Km ̧Ĕ`L3˫��hE��( �y?b�ͤ�+Ʊ(�Zta�7�Ҙ"X:����N���ې�L1CK��R�-�C�#��F�x���9̈́HzX��є����1����(Q���Ȝ;k�3����L�{A�$F�������wz�4�ʌE~+r��[`�m�T���Q��ib/@ρ�-z���+�xN�_4wp���ҍXV���m���ơ���-H�d���NC��3������[�C����/��PO '%R��$������K������~���I����F+�(�JiD�c}	J;m)�kC�ǞQ����rO�I(�5�NP��S��(�AB[�V���}EY3�b��-U<��n���P/ܐ(��v�����w�Jz�[xe�I�E9b���w�?
!K����G6/�9�8�%�)���$���] @�6�I^�g兙?�O�������h�r�p�mJ7�r�ӳ14R��} Q�D�pOKk��Yg�9������u�g��m܄ښh�t}3$HQʦ�=�C��";/'ʞ7��B�]9q۾����� {�5H,zref��9�z�#�PF�%�����:��+�-H�u�m������O5��Z-���������S4}������edL���f�$�� ɔ�kMX�~��{��Ήw�PO��3����b�	<W�a�1H/ߣ���r-�����1����������:#��C$�:�_R��?�>���$%<��}� e�G�lfQ�8�i�W;�B�s�� hd�ED�xM�w�|����F%��.6�_�{��R��D�S��w�V�P�Nd� ���8�9��"���IΘ�P���l�h�ߎ���WM�Dz|���J��7"@%vJ�����g�y�F;�e]>ν.�8�2��(/#y�A�}�f���o�����<�DΚ��˖����w�
K��~=C6���A���u�p� ���H�SYA�8�'�����s�<-�]�CL��C���I�\��㠖&A�gbD�78�1��|�/̀�m�	x/ƚ��#�=D�������� q�:h_��}�a82:L�?X��hN�e��� �ѝ�)�zg�Y2jA�n^���Ni�+���dp&�>���K��ZGI��&|_7�vȐ�N��6b��x|<��I�o�bo�U��Y��x�3b
_�wO�k��B��[/kd>�â�̘؏YB/�{�<H-�l�"4'�#��-�L�s	�żo�Og�g�Q6d�{�i#x�r;���j�3s���&v����B*��l�+sYBa�I�<�&B&mY�m5�Y��Jw�ݙQ�_ݽ��������)6`��oz����A�k>�ַ��h2�� A�+RC���ri�}b��EJ���ѫ5B��� �oo!��t�(�; ����lZ�Pv����!� WvIሆܢ�6�7x=����JE� T+��Z������!�P�D[�h#Db����Y���v��ä���ֵ�i��JY��m���j��ƚa�Z�'���]�"�җ]�*��O)D�/N�O�G1���q~pF�]���}g�H�B�Rޟĉ��+���;�|R,��N��XB��g
֕�ɜ,��1c�����N`��Ds.�4�����D���X�Z�����5ߣ��|�_#�MvhQ��_���"�"�%U5��"Ű c��h�'9W,f�6�t�G�l0+�\�t�'����7��,o�$�Ĕ�l�⊊+3DA�|�8���s�g0�7�S����7�M�m�7�r�a�O�8<���mű�S����'(jK߈����YD*L�G>��/�pd�]~!��ͽ�3S.g��Ek�-`�1�S�Ch��cxl\cr�೤F1e��s y�L��TA��e�ԏ�9l5�CUq%7s���f����E�>f H����G�	�8V�i2%~4�+�3��b3a"�Ƕ��΃�V�'�����5]�kH�`�+�$�I�̍��h$~��ʆcqp���S�vn��e[�Pp�TM���M��=1����(�4}�K�����,���Ɗ�"!7$ ��4�~D
��=�����I�da+C��S�j}+������8:�ëY���2J�f��o��l#�bc���e&[<C3���SP��'o��?�F�����Lڂ�h\�ե�u�~��+��c 4u�v$S��G�B���M��|��0�)tRP�̺�����Ө�\��MoՂ9���j[�Rf�A�S2V�O��Q���.�;�aea�� �]��D[L�-�e�RxGY(P�q����[ �i��[�e�^�N�I3쉇>��3љ���|�Bهt��H�y�i0�J�_����\{9'fġӵ^\s��XZ����JF��!K��z�8���1�����.�5�H,�9t�Zy� �J��'*���ӑ�\�S�������V�m���JG?=��m����%�=9
j5՘�>A��|	�����8�}��y%R�V��F���"�Q��*�����T�b�9��k��?�����V߬��	,9��*�U�ܔ9�ӥ��$O4~���Nj�+$��gw���+���w|�����uЗ�PZ�x(���0�=}izkS�:��S�d�˫z>a le��HZ�]�8S���I��jɾ[�`kʠqJ�|��&Z��|�j��b��		<�����ѻV���>zՐ.e��fR ~�rJ��U�Ml�)I���� ,��"�4�Y)�
��n��oŴ��_�-5��C5ZLe��?OV�E`&���ee7k���w.$S���4ak>f�l[���&�dҕa�I�=��qQk$��G@��i�xB���M#��s�r#�5�<aa��w����L�H��=����i+ �.ܤ���7�@�˙Mn+H��������ݗ�ﰶf�e/c�@P'��3)�[��5q�� h�����,��.k��d�RwB�=�t��_J6^���R6&����5kp^cG��)��p�n�=�|�jw�z)'sqP`ٙ����D�������}�m+N��_��+K�Щ/�U�C"%H�Z���%�o�Rn�sv�Z�����'��f@lt"�Gi�2�� ͸DU���9�r_��Q��Mpg-mM&3�X��x���z	.�X����b�i�>�1w�	�Hc%�YLZ^ƒ��J
#r	��	���t���ߖ�W�� X��������Զ��b���f��5_��h�.�T8s��yW;>�^Cl�m������t�KN4�#S�e�_�M���n��p��-��F��e�6=��3�JVG���q�ظ��AC�V^;�}">� ��?.�6�s�(H~._2�f�6�b�<���[7Cv×��M���;��zm\���A�`�_�[�Ovq�c$A('�ނT �"| ����558�#<��s$��ڴ�x�A�_\���l��b�nXj;,�%�q�d6���54�b&����옟
���^Tx�B2��Hg@x^��\��xO6��m�����X֐��h�}�b�M<�y�+P	����k��e���9e6H��!��������͊���g>�_=�g���Hg醯���,�E�d��<50.��sg"��h��񿁧�L�{�cm��.�4;%xk5�C6��l9��T	u|m��ϸ��a���Y\a'4��Py�W�%�Jo����A��J)����)3�M�[�_yn�w��bZ��i���\&|��+�x-&��ˡ�$䞌)���ț�%��1�;���]p�X�y/��ԯ~>�to �;�9
��l
�5�+,4|��h�N�OV��4�0 ����j��|
�E{�e	�Ԍ�χBv��e��'#l��"�-�&I��sGz:n���U��z�X�_�Ζ���G�ϲx)�����6�]ik�Ї����;D�m��G�tU~��|9Xc�­�";�ѭ)��35�_��+6�#��	�G0��������A{Y��]�y�����4�o�yx"�[��E�*;��:9;0�qc��������� %�q�������&]2@������Om^ɑy�jG �GM:1����1p���̋�"!�%9���o/�?����k b;��*��Uf��1nr�T�bk����)�U���#wĭ�����r�n6�[@�ٵ�.�����c��[,���t=��1�V�Xlf�:�E�->�����WZ��=�O׾n^���N��|}�_(@�E��6�^U�����4r5����~^{�hv-�z�͉3���Іݐ��]�E^�|�__�9��t�|�}��}�g��'��O��#ŲY�>yn@�-��˅!u�G섕���ɀ�G�]�dmߠ��ራ�Q$F�!���9�o	�Y�N���ӾPOzSţ:�B�w
��4Z���t!�I�
x�ɷQ�cA+G����)��{1�g(V��}N�����_u^*탍�\�qNC0�^�{�Ӎ��*r��s!>~�WSzt�0Z�{SR���jd��"�-��Wm��e�+ �|@����ԣ��[�0Ƴp�^��:j����8wl���=�Y�k���� qlۚd�x�pݯ��ة�a������Q�S�$Z㍑-��_
�-�>ț��u69d���z=�L&����b?L�h���(u��Ss!F��d�� �J̴F�Mg�%�Q�=�$X�W:Xv�HE;�<~�gэɤꥭ�qp���P��#��F��3��@`��:��3�˧��6$xᱣo���N���^��|�)��Z� y����̢���G�X��T������
�N�-����\c_�i�#�³��q߹��0�I/��ٙT������I�~*��n���~��V�o�L��\R���#��mfNi��2[q�/vo���=�%$>���/͉XZ\��	���L�R�g�~�>9��C؂�#������C@�%ד���
 ���G�%Y�dH,�}nN��Sɼ�8'��Z���#��ڡ�0�����\�G�̡����e����k�!m2�w�ܴ��e���8�	�P��l���{���@0��1_P͍qI	$���j^`}L[�5��G��NB\俹<d�#������4'�=wp�e�D�j֢ں��wX�Mխ�G�@4&��<�k��Ri�r��][h#�����p�<��kd�1���W���"4����^i�WqJ<Kْ��T ���k�É!�=w!��c�WX���f�̧(f2��L����tPP.n_`��ËL۱"�4(O�L �E���3��>���+���+Dt����4�F6z9j�4��-Z݈L`V�D��ܥ��8@.�	����/4*j�CC�� �I�U���b�)'v�-Ր%�5�1���mΨJ��3p���J��M7x.|���俶L�Wa����2���\|�`��4��N�y�R:�Co���k�O;��À����#�����|�fN��}^d����3v[b����]e$n�2m?,�*K���мi�c�5Z�v���Hē��Y7x��<{ut^�L�M�p���;a�u �d	���Y�N��#^ڏ?�(o�D�tky\���_�k�нPV��B�K_�~�0�@�f�4��5��>{����R�[���*�e������=�#����l���,?\[��Z���d�F�M�n�mL�k9���zơ��#w��7Z`�6]̸P�f����(���y c��&|.Tg�My�����Ƚ��~%�����cCՀ�R.56��<M�.��5|�s��KjM�X%���#�r�a�^k�鮲�`����كyxE��q>8.Y	�q���x��I�1Se c�?&��o7߅�$�1*�~	�����#ßua�*�ݲ!��n�z��7G����HAŔ���[_�qJ�X:�ic�Y�]I��q��+Q��Ul��]̟���pR(�s�N�_j�Md��xǮѓ�^�?,�I�W ��ntN�͆�{�i�m4m-����
�y�$Q�`�j����+�DJ<J
��E�d1���F_v��w�j�J��A|�ڈ����;zYU�kd�*�(��Ehtݜ���bD��ȶMq��8M
�)��dQ��Y�.3h�����*��헁=XݦQ6�ƺL�87e}��^�Q�J!�-�}5[�m��Q3�lh��oY��-R�	����_�,����u�Aʭ�6c�Y4Q>_�Tθ�c�E'��!�3�����kW�k]���5h�^�b���%*N�X7xý����gߒ��8�6�1G�-q�/��Jc/�R����i5=���&&��#�C�2R,/�@/,FN�⍎�"��td�G�]!%��_T��{b�L=�E�����=q�;��S_|D�zn����.ږ�FYO�e��S���sҔ��
���b݇?+2Y%�p(�����U���S���!�h$^�/�}�}(*/���c�o����$���p�HB}���87]�vac������{uّ�:~�����
X���a�_)\���Z4�Դ��ݵ`��
���~����*u��͐��a���W�+��OȘRs�G�G��Iɠ9�Ԗ�*Ezt�!���O��)j����G��$�VN��I��[�vLQ�L�EIa��2�+�}�V������wu�~tXAv��M![�bA'���˺Dw����ݸΏ䶔�@(��pĎU[����a	��A��o]�i�=��	���ɣ�ke0���0��/h��g�3�/�'xK����dt2 u�l�R�L�D��:�	8,�aZڻ&4�*����T�Х��(�d�a)��ﾱ�ޡ!�XWB�i�e�M�cC:>Y}��&�{Z��?�Ӱx�k�!UK�r���&�\Gz�!�� &���lv&5�)1$��������@��p&��[��M�dyz]+���;����|�j�?�4�?��]�[c^�(�R�5z��uIG�����@
�z�I���H�MG��j��gF����3��
�I��&�q�+X��t��x.�k�- o�$-��>=���[6���D�r�s�prD��x�~�>�4i"W؃��w&풫c��y]���s��oM�ON �q`2�3c֫DN��m���&탦UgK�
S�1��ld~�k�w0h�6V�S��9q���6��sp`��M�R�'_D�Yf���KdK���.�KO��]�� p�����iTsc��!�Q\:��t\��ě�pߍ%��;l�Z�h�B�M���
g}�l�T.7�4x?�~W� ME�.�����+BRɟ=Ѐ,z���0`�m1��i��/b��& 7��� X���M�������G���!-���o����*���hUw���歷��-�$X��S�9`�^ڰQ�+������93�����YZ�g/����V*���
�wЭ���Cw\A旧n����x/T�.z�lFQ3�Tj�\�օ�CG���f�4�b����!xow=3���]��|c�e|�4i���/55����ػ�&�"㝥#Hs��MnoYSl�cq'2W��3j����=>���ʖ�n�@�դ8`#��~����}�A��Dkc�s�|l�
�B~�N����0���ADBlMU��X��.��r�ۂQa�9����@A^����|KV�|���Y02��Z�k�!B�N��oi���
d�=wn�3}l�5�GjԸ~�0�A�J��4��ʿ=,��O���V�	חU3($}iPQ���Y,"�6��
"әr]�VP Α�>�$33~	fzQ�X�ݾ,;�̧���ayˋ�2��؀#���_���w��R�K��T�	��}�,U�������?BWS���X:��'~p�s�hM:�_���:h����k��O`�Mw�8�*#��}"�B�崀�ԯ<'%[ �e-� ����rf:��s�M��x�E�`w������RQ���.(�sXs��҂�V����:8�l�E��]8g�Y�}�u��" ����]��0���G��|�й����cM���S��Ŧ��$��GEP]��r&4�V]�x�L�WB�;�v+/+��0P��w��e�������-��u�Rc�:Z���V��O�yV���~��f]^()w ~l2~���Q�.��qo���ŽrI[@�#O3}�^�↢����d ��Wԟ$�5��p!UIE��>W�&&}��S�J/�� X�r�$]�K��S�s_3�v����7^�Qh�O��
;ׁ�¢?�ʃ&G���a��/3��.��=:鱾�̨ŭ�F����`V���﯋�<��azr�γ��J
�`-�������&����OJf|��Y:G�D
�/w�&DK��cT�� ��G
�W�©�����臅l�8;�������%�Ű*12&:��k�siA�[�����W�����Ϣ��r�5�t�d�H��v�0�{�ԉC۠�3ya6�)@I��gY�t4���52[~���}Q� ����kc^7a�-H���C1�Io�+�����~�j�¿��v��J��Y&[���K��sn����޿*��`@��K��_"l��Y��:�/g����]O�J�Bi����-��"���E����W�Br	�c�[�A��bĒ� ����:��z�M6*j�lU݋�Ϥ�3�(L[8�@/���B2�-��y������7���*(��?�V
��C�tMs�=4�\��e���UP�Wۦ6�1���=�����jC��x�eč}8��CՂ�]��̺~�
��S���cP��9�v2�v��`R.�ct��:19�D���Y��eo.2ͭ�G	�����������~�՛׶�a&�Z����PvU�`��|N�<X����my�S+��Ү�
��8�
O�d���~����������S�hk��M	|���V��{OSƺ<rg�s�3Y ]�k	����"	t�X�e9��:��i���S[0�be�(�(�l�o���=hU>�o���A�P)�wW%|A$�����R����p� ?Li��=��/Gf`�F����H�YɅGn�wI� �=���M{Q���g��z�Y�^�5鷝��w�p=��wP���0�K4Tz�ƽ�'�U��-?Qy���ʛszj|���Yzfj�t��~͋|o��<E��8���TO���|��d1�bOLOn���Y��5e��?��݇28W4�V�����1���X�����ķ۱������c�N�Ud�K?�3�
8�/��A����?����!=�=�q��mU��w�O���_J�tJ�w3��$Ō4�@��	���u!�\���z����)%SgK4t�d�H���pẙ�o���HP:�*V�������8�Z�?[]����C�@�f�Zq�Z�§���9�WGj�wcGj�@pz�{4��3}�'���9S���LOR���w��6� Q}qR�(��]3�p��9~7�i���rO�^�)(Ыa��@F�8����Y���M������	��耪��Gݫ�]	7$���{�;t�"��כd�����	���{��ѱ]���[5�+[�<����I�^6f�w MU	Wr���6Gy���|�\QN,�W�� �P�J�����j�Ҩ�%̋�`6`	��ԒQ3c���ٟ�Ôp<S�`��pYy�]dm�?r\���8~i���;��+�kNO�$�~����D�m�
}���jI���^�y�ĿCg�E��:�nE�wx(P�c�A�۲[���Ή�������& �l��4p��ג�8�N:�P� M&d0?�f�fE?�w;V��z
�bR��A�(-�bd*-4<�6f�+�.����_2��T��'��@,WWeIK_���3���^�`�墸 ��T�x	S�:٭o�� Y�Փ��>����}Ȅ��~� 	&RV���d"��!r��6Ӳ3N�p��'A7�����:�BD���O�ʿ����un�D����lqr	������WkFY]?C�ʼ��R��^��@ V���i`�v�~"����Z�G�$ �Pl{�?��f����^��B��=a���%QYr��tE���.r������U���d�M���|J7�n�Z�Yܪu5��ks�?2�>���"�D�O�{��"�$l�Y�a�ƃk%g #�:#�S�t5���a�/���A���z3x�󯾼_tV��̆�Z�۵���
X��Az�o�K��C�0E�C�ͫ�/㥸ZO��pu$=2r�������24�`9j_x�7fn�����2K�
k��i�
)���Sd���&�]������=6p�tF�#�BE��=�bB�`�Il���\��{��k�h3|��b�3�kh��V�Q�0�3f�F�����������g:M7�z���w�&~ �ؓԙ�w'fV��.�a�9���D5���P�u�Z���V�J76��2���lף�ed�V�~IԹ�-��>J�����}��r����^=^�/Gf(�J!1,8'�ْ6���g�K�'�?�W�M�!��Ɍ�x����J;lA�1Z.����d͉.0R�e���������NV��K�5�I �ضT�.#`��,�E�k���������@/3"����(�l��+wչ��9ZMB�X=k��h��qO[���Kq�fy�u�].t=&��;���o�*T��ĶQ.x \�����ۥ��k!3��C�☜:��Kv!w�9�(A"�ͫ�/�c�Xr$�\׀b/B�������u�׹��[cI���tM_O��Bx�(D�N_�G�7l���:'�P7�ȑ�$��w�5�����r1OFw:�(>���J���j��4bJ�n�!�%��ńof�Gƛ&�ۯR��~k��bh�Ɂ38Rܕ�A�����)}CT6���8P���G�����F�Pf�/��ф7�>e�� �r������j��ż.�	XU�ol ��==u�~pjq��J�n�m+u�'���r��V3�ED'�n����I4?f��W���V�)N���7)~>�Dy����ԛ*2��+j�W �"7Ȩpr�\A<v���/q�i��I0��ji��Ku�a�_�%xY&��]�p��-�I��� n��,+]%�H��F���j$��<]���f���!ظx�}�!���C_�b�x�m�C�L�l� ���z!,�g�u-��]�r"�@F�:�G	��p̈́��(�Z$����b���q\��drǌ��dW�aX�]�`M��Y�.��1{�]��?�Ø��C��ɞ�f���_�}}"�R�,Gf`��B��x*V�bn�v$Xٺ`|a<��Q�n ��3��зTh��\'ۦ	���hcވ�,{:�8���M+�P�b�6s�o��}+F��v��Jz����(�C��ĨQ�9��hbz��G<�ռ���R���uF��7y�?͕�j�6W֎�x2��m�,�}د4w�Jì~`�P��#�>�`��E�?}S���X��"��q1J�j'�F"����a�(ɟ;�q��Te��;��QC�$�s�UR�e�R� b��c��5�kї�>=��.Gp�U�6^p��/����.[�ކ�%?+9= �D���M#���\����ev�!��1��� mgh�*�,0���s�����Q8���J���gW*�����Ud�a��l0��r�`s2����mҤ��^(q�lf/�����$�*�fލ����`��L<}��]1�;����*�,�Ylx*��tKՍÅB5�\�X��7�)1��L�� ���G��Q�(ӡ��e=a(��bn���g��b��o3�LóJ��'��;7�a���b����=.<+L+w�
w��`C�ΉA�pD�`!��Ϊ��v=�fsbv1=Z���lH;ϵ$�#5T<����ɣ	\(e;e����͌��j�������S����z��F���L�
?,��A'U��=q(�ʈ��u�TQݑ��7�е'��Ȓ�{�@���IMl^�M�<�S/'����<u+�y�x$��%��T�!�M~�X�e�]E�`z��ʫvTw�v�lY^;=O�LI������ ����4?��"  �3��2IɌ���*��A��(�����g���Оq2h����.�!�I��
St��:=�on��:ܣ�����h�S�ᦎ7v> 2У���m�/,b��5 !����ç �b�4��ֵ�3�n3֋�Gz�;�_�J�v�ԉ��KHH�U-Y_G(�q����Sۻy�N(%K�|u��nlW��8!	����z����c�`+BC?�i��<��S�Vj�����#W(b����Ŕ�	�����(	�=U>��5�2���Ғ�(��چ['��S��*�����0#�s��\7,8`�_)%�#Li�=���:ͬR�od]���%P�۩nHo�ԓ�O�<��g�= x�H���������ȋ5a�]������ѵ�P.�*#��Fn��=	w��@���!�i�,/vת��&�����	Jj�WGs����r�]�0s5g�DR�8�%nI%mDf/���d-b�K�^''(60*�K��#�H\�p�S�����mb:lw�_C��/��!�?QAwx`���3�I鲁7̣<�F�S�V/��BKi5V��wćïDgl��%B�]�X� O���m4&p�{�_� ;�˺"�fb�d)+���8�ȍŀh�[#�?�Df��z���O�����
_z.�&�_W"2ԤL_��dZ�\ǜ*��_�м`~@r�y��(4'BK��IOe����<���@�JQ�e��q�$فK;͂z8�l������2N(F9��5>�5 qs\(៿���g���@��3	��Gi%�A�ފs�݂���7\�jW�  �b�󭠤j{��Wv�^ x��ܴЏ��+�|���h	"�A�9�5jԘ�$
��f >YI�I[aw��v��S�F�#���.��]����.)��?��$�]i.݂��| Č�C��m{���o��#P�pL�ͪ8ȩ<�9��$V���Mw�R�%�
f^ǯak��V��M�o26���kdT�
TV7V�����;8����+���`���� �0q�0҈S���=a������FFs*�:��/�Ƣ��qI�S�a�3Et��}j@�>�~0'V�%O-\ewx
X��D�_N�&�u�CǪ�}���-w�ۋ�<�_�ˡξU?!x2\Yp%#�5:�\�v�_�|_*vj���=>�B�ЄP��(8�S�R"�
*�oe���S��A�~_��3�v\�G�C3#+D�HFa��s���X�&�;��
*�2�h}#��eg9�,|���$���$��U�k��l����=}��ڎS�j�Kd��:��_#��H��ܗ�BE/����:�r�eL�H{�!ʲf��:b������>?�Z�%����b��{��@K��{>�՝�����/�$�J��Q ;'��0ڊ���2*��`�� Ύ\��y��Kvd�u��>���V�ٲ�E%���HN��%�V���y�lˮq,���1,o��!���>`H���`�T�ճ�P2"8�5/��N+@	�!����Y�p��@����5�'�4��X[Sׅ;!Fܷ��[�]�%��$2uΞ6EmE0�ڼ
g�!{� A�Q��@�zo)�1lO&��_�(�:���n^I���9���T`��*K0O��ې��%�10u zzE�I�e�k|	���b�>���	�O��G.��o��"��bŐ�H�I%�0α!����C}םL��5HRx���qz�m6�W��4=�R ����Bu(�)�[��2>�k�1����ueB"%F�עR�8u/�D���r�@d���(6����=�@c�0�a3�9U���U�헸��5V��BB��#�g������e
�H��#tk��Rv�
T�L�e�8TJp�c���ײ�m�QK�f����J��%��o�=4!���q0�zY:6Ĕ��=��;;*�h�Y7��	Z���Fzy��8j���R1{Ȍ�6��b���@�1sB�����KC�{#�z__>K�i�)��ⲷ%��q���r|�Ha��%�NKBBR�����R#d�~����N��,Hp�'��.J�a�d`3���ja�2F��������סF�Ԭ$����2�}B",�г��pf��}T�3�KD&Y��]I fOt��͏7�7�b_�;p��ƣ�R�Y�s��[���/q	�W���{M=�q▻���+��,���7��?�U^��>1w+�-5�Ano�夈���8q}E�2%��JÖtЛw"H�����������*܆�o̗�̰��:k��#;�@�_���dt�;j�/�l*��1���A�	�]��y��q��P�V�����ƾ��H�oǥ�n��K�ƫP�o��v)$ԭ�u*α?%rp}�E��-Х������J��9�s?�]Jf�_H�E�u*���(�������j!��֕ce�h�trQ��{��v%�J�[rgpy�h�|�h��˪`cq�j��3����{#����Q=���8�L���1�ɣrzCS�q��K�z�9���ŧi�$6�!��..-m����6p�5�p�D��h&#��7ΗV~�/���^;��d"\M��"�	~%�W��mF	%ˢ��r���[2��=�۱�uy��F�]4�%hν+J��Q'�$0��#�8���.L#L�	�J�xYi�e8��n��pmC�Rc�oecCPW�"�3���}��K>Ԡz���p���4�RPf��?�����]}6w�^pv�'�⛶���¢������c�9�ѿ��޳ބpE0U�mY!*��KE��-��?PM�1��H��ac���iU�+�Z�y�	��w�NY(�a��Z|��
wKw���X�*�P
#�5��-.A�圵�]���@9��(�e����Q�d�7@0G�|[�������>����t�)J �1u���p꣆
��J�b���I�^�ƸC��������CcR'�+xM:��5�~�"|k���sC9��)���.l'�y�q����ֱ���]%-0,GT�a��ҍ�܇���O�������ps�=r ���SWsxA� �ђ�XO�Ǔ"�1*�O���*T�=9�����\�e���I/�a�p�P>������Ħ�牎э-W�f���maJ�w�.�7i	���l��v+@F�~�1�RY33��ek���
fF����_V�yy*��!$��j�x�֔�Q��|�+s�l�t�e{`��T�tF��<,B ������� @{;$�?R�%x�}�A�v&�_�Ry�o���^��\d�'�B|)����R@W�����L8(/������T����Qs;0K� 2�	�'f������J�j	BQVU0�)��?���JÀ�Ο�è^*�h]<�S�A)�[΢Ϧߧ�π�:�����^���}[L���b9�ȅ}&�BO�S �E�g���3F�Bb�g�q6�bק��Ca�1)0O�Op�Dt�⡆���lyǿuF��v�۠��Wcj�}�0�����͖�ZZ�<oFڨ��?Ԑ��R	��}X��C��
C-%h���&
k[�v�����K����Tj��jsoI��Ÿ$]0C.A�!�gc�滨׀g))�w��:�!�7eх�t5xa^�yA��;_�X�<I�6L��#����
u="�e\�ꕙ=D�z�	��
^�ө���5��$~{I��=uoDL(�	�1�F��K�e�л5���!��UZ�"�E�s�
�H��}�cxJ��.Pb{�6�9�>�u�=�Fҥ�~:-�G	��p�N_.)��{Ј-�d�����\d�w��S\ij��/�a56�$�ly��ۅV�~N��Tx�Uvqe;��`�TI5��}��3x�(�0�[������l����Z����Ȕ��6�ߟ�wzx]!�P��K��Y�����+Ľ����P��]��$���O���-]#��(i�:).!��_$�Fͯ�U��S	�[Wb,)p����-]%�����?����.o�>o*��D�8y�m���7�i��\j񠢞���Ջ�&_��<Soq�A`o���;M��e�ajh"�ȧ�m�6v��GHr����<�%���+2�������,�7�͆4x�J���{���}1˰w���թ�7�$+���%���`��>4�&��Gֹ����<��-�D��O(�[���A��ᥖ\1+К��`�c��Bfv��,֫���ݐ�O�(���5���!x�_:��Pn:���5SLQe$!�ВZ�C��KpS��O��J�����2 q�}����
w�b)�Hj?=j�r���Y��Ww�$�x=��j3-,/N��~
;�|�A6�42�*�CT�	�
�����RW�I��/�a"Y��Ut�߶���ڀ���XpsQf�M?U<�B����a,�J1���X��a	Q�Y����~��랹a$�R�n��'t����G�v�2]���D� ���K�a�+�g�LFO�r@��ͷp�<���<7�D/\����ok�~N
00�F�m�������4�9��}=ͩt����CQR�/�U�R�`b���,M�����,�������M]�8K)s�s�}��߇�5պ��Oe}:������t71�ߝH�/� X!�}����"&kS	�y�C\��s�
�S+M��3'??6�m��2M�)�K��c�vgd��2Z�MT:��GiY08�S���-Dguu��;�� j�U����D�p
�s�љ�j�}q7Li�h��3�#*Ѵ�bZ��{��Y��m�]	�6|��zZ�B�>^���:
�`���#���c���d��|�Y
�!�!�sԃ����LH�/�	���U��C�Cc/X�4�edy6�	[an��/fH��`
&��v掹N�1��V�
�:	�MyAT�2��k�W��C*lq+�=���|o��Ԅ@]&���.O=��ȽF�������U4�� ^!sh��'/ui�~��/�[:.*܀�TIT�z����qe�E��#��D}��ѱ^���nf�G_��'�(_j�Q1��v�7S�}h<[���X)c�a��'���4x���ǥ�$�z�o%�D�Q��qIp�}3����	ϖ��}	�&�y�ͩ#�j����&j�Ԯη-7%��Q��C�%a��`+��0\�^e�k��Υ�2��'�w�e��r�������k�˓�`�i#����û��g�$��E�1��OLU�ʖP	RPu.	���M��mP����?�z�nU\�h���j�bfz��)�˦?-���5�9�Z�W2*��̄p�c��R	�E8����AR�F�y��J��u������z��n���S&������DtWh��DMƍRob��ծ����Ԃ�aˑ�'3l2K���tXe��'��^[7qw��/h �V��D�Z�k>#F� ��.�fُCAf��vCm�� 3#?�R�WDl���\�9	���@�|п��a�@�+�J�Te���@q�����f���6e�qLEÈ���C�8������Y�����NZ�H�a(Y�C$.5�%�{(��T�v�~#���4��Utk��̸�iנ�#\~�R�5��ް}�z|���D�5O�΁��%H���:Z+Yy@�=/��4��SC�r���Z�׉ڏ6�"MEH�?I!@ͩW�q4�S��w��>&t��dx�~��R�ק9����^�]XP��������c��7�b� ���5�C�<�X��s66f�.r��GT��owcHT���3$�i�	�Mf�
 �bŎ �9���P;��o�n�;#y��/��<�c�%�2�� ۢ3��/�l��K����i�6 ����i}�w�'�� �g�g�/*���(�\������cF�&����I���(sܸ[�@i�Һ�j5�*�Iz�Lx�����D��$۲�7��c�I�y1+>��d���]�_���`@?u�8@M���g����[�TQ[����%-A'P@�g�/|�J�υ���J�}���g�LmTFnc��dsS�9���k*��2�Н���+�%�/��:GR��L�B�k�aC�ݥ;��cтH]�e-���}�����KM�F��2�os��8E���+�I�ĸz�����wg��6 �ow�ԇu����T5~���ht9�u����`֥������:7���](_��Np�H>�r��S�+7tRCrev�QL��7����^� V=�o`K��ѳ
b�$�$�(�yrA��]��I2+b���%#��;��'�>1���1��kr,����+�0����6H������Hw�A��	;�}4���I:;�U�0�d�@Rp~G*jPƯ�q��,��Y�7gO��GF-1X�#
6����q��8-�D�2��|�xBB�=wh@�Yb��
v�T��{��0��|�k����k��ɚۦ$ވ�*+7!��΢�)����.Y�O'0M6��E/�"$�36��a�)UF������$�5��%�A�j�@��B'V�wN�ٲ^��L|x��z6B���$Y� J�S������;�}���ʪ �m�D1�n��Qx2!p ��4�=�#^"���^�l��^44:�m [?�漮�j�Y+��}�"5q�]�r�^7���P�e^59.�g�y��D��n4�Rr��2�e��0{�%�t�n���Bg��؇�uK�qC��w� �� ��5��׊�c�u��������1��ŋc\�k*P�p M���uT����is
�&,D<�V8�1	a�e �]ݮ�~B�!2`�g`~�Q�j�ȾQZK���ԅ�ۙ�lK{�M�v��d�����YGfgs��� $. �VE�jj?\�u"�葜p��q���O�$��w�G�����É%�����hi�\â�S(.fq� 	�O�SdF�d��-����K
(_ٽ}HAB�!���" ��آ.��E�E��Z��Ś�┷�*�4�ȫ����	�s�Pd ��`n�����8v�=�y.�2�
��B��%B�=ql�q��o$�$�q,8�q��W����P���Gk���[Ł]ʓo�w��a�D�g�*o���,!G�/?��2�1�A�*~N������2�]A##�SkJN�(V�,�}oT�B|��^���U�BB	�$�O�3����pG�
����9`����t7��;�lL·�71����m���L���8N� V��q�e�j�L�0�D��G�$F�V��X1��34~��]mB	�)�~ ���F�ӱt�W�t��[ ���|ԑO[�Yw��IR����H�6g�u:�	�L�X͏9��n�`�H�O؞�C��!�7����M��tf��wy�v٤��?Ki���r�U:�`��˱s���5>�вh�G��s[p`*k�Ph��ϥ�&���<<ǣ<���&ٍ0�y
Y���d�F�SɃ�z�;�B�@� ��@7l�"!��p�W�!�Z)�;Fl��3�0��="���T�ȶ�xb�ۺ~(���ܙS�ڡ�qY$\�ى�6>W'@��^(��>�]-p�Ja�
�I\��ĿUB��ڲ�4u�w�rZm��ӆ5�����������*���c����ϝ��6��x���u^H{�p�n��IN]A�̒��S|��qk^�Ri�FZ�7	nt�Ue���w:��s�"�	���k�>�;�a�zل|wPei�P�@NO�7-6-{ �t���U��_e���-��D�v;���^�C�5�E����(��v�մ�#�5�!��e��~6)�T��&KKA���������i�����N;�,�c���0�N��Ʋl��t�zKպ��)��b���j�fG�͂���OC�2�S,*���9����B�w��\���K����5dVGC%��51�jj�n?z�T3���=U��Al�#���+@,���b����x�v��Y���k��<��f�K�Z���^�L~��f�:2	2�dE���z��G�۝�x��Ԃ�W�s�taz���d�Dt���Jm���$���o�V�|	�U���l�����ת*TQ�f�s9V�1�x�/iBA"�ώ'�M��<+ �L� �6��s�B��q�y�H�f<Ľ���p�%�3j@�R� �#�m����U���A�����2��݉�6��A����q�@*���kX��6I̧�~�.�����o�E?��%�������m��%��7�p��h�aUW��@������yG����`�C-$��U�$ۅ�{(��%�� |�Hj�	�?�,B+�Ǚ�s ��;u����i�)?T��b���b��Q�49���Y"���¡w�+Z�B^������Q��~d����Fw�z,e�Kt�N>�:�d?{��$Z�?�����Yq����ͽ/-~�i]fa(���?e{�>��C�� ��7���|ׁp�k\n�j�S�ĉ���yY�b ;�&��(��u�
Q�	'�l�,��l�Ѥ�9Hu�6r�a���
o2&ß_Z���MXb��c1 ͜*A��]����}2�2���P'� ~�橦���@�x�e
�m��������*KJ����黐����M=	�-����X���,�XCI^�n�/�=�{��jǵ�twV�t%�4o�͘g�вѩ�ʫ�R'�MEx�`��(���Z�e(\�CB��@V7L�딑����
}q�8W�	?n�_Ta��P�\������?]�5��~Frw
��<�����Y���j&�m ��	U:;y��!~�
2d�Tc�-���Lո������Z&'�Y^! pA�\y�L1Aw�TZ8�Tf�Ѹ�S��W^�8n��9�S����J6���\����_���OΌ�En�bh�8q����J���W�-Z���`�v�������'*�|4��3��OQ�h����J�fc����m��#*�8[C8%�S�����O�v%Τi^��i ��b�7���V1�٪���q�E�p�������6?X 豎�p
�+<22���yJ��J��NԥF�5��Wis����hݙރ'�]�#�?��VG�7�^���<�\!��!�J,/�m�KǙc
�w�#q����\$�?�����]����6����X����Ӥ�)ٙr~�bsɤBI��⠐�ICT*���7��"��ٹ��ܗ���<�ev)G�O�P����n��"�����\�[i�g;po�hk�����%�������k���B�X.�wIL\��y,|�0�s����4��;lG'�O̬�mԤ�+ʕnF3ֈ#O7��"�`��@;�=l��k�F��䫫p���r޲xvr�\�<�T�,M �Jj��7�L��1M��Z8�?r��݃�<����e6�U0�2�)v�u�aA��\�ˀ.ă��o%�ܻ�I �-�.�L�u�(=�����ۄ{��:
�?��C�XY4��CQ�I�K�\�}Jo�Ec�JL����2A��w��n���+eT.��-��������j�CQ`�y��ZR�N���aY���)�u�St�o �Ɯ�
���bA��[�3|���e�-j��NW(�>�����L\\[a��Wm<D��]ۆ�q������U ��'��xv��
���/(�}�f�ܓ��2�y��L,��n�\��^��^n\�H�ja�@�����R�y�Er$�@��Y��<�Mx�eQS$�,\����Q�}��8P�����֬�d!ʫq��o5L���xS�q�_��������#9��-f�S���u|o]��M!�g���ouͬ�6\�0i���=w���Z;�����j�5��H~�}l��`�d6��#h*ᶩ� uT��"�v+�\����6����ڡ�Vx�Z{FDO|�.y�Q�7T�%�1>8_hU$���Ҩ���:˿ycy>� I�" �q\�ө	�q7s�����<���I7�*U�u�Q�qO(-��g��͕z���#ee(����\�o�� SR���2h[6!R�J�N?��&���C�lAλ	��<S�b訽��iu�
V�z<Y�����UeKa]	�_{Y��r�r�ӕ�,��C;3�f~V7� �8�6%�&�٨a6�;�.;F�s�-��[}$6�xPac�'�O��S�o%!��u�AD �x�쀍��A��G5td $p1B�!шޅ�4B��3N�F͛������$56h�0mTv�����:��r</$�M#�>D��'�1���J�
$���z�8j���O'*rfG�������3{���7PP�\��Y�斉�C�*E9�.^�FǥQ0,_]}:rh�TӼh@h���kSP�^�lB˖g��>�$(1��W������P���0���r;=G��8vR1̦�*��Q<�$+�����$&;*�#n4�T��������z ��xf�z�av�S�b�M"����i��br�	$ �>�w&�S	��"�M�=+ygr�6'|P�`�xŹvИ�!��;�hYዒ��'����������nG��-J�8�{�+�a"�a�r�&���ѥS]�yq@�r��<�L�ɩ����K��J�p�h%�p%
��@��=i��t_&@i3��#5H(�X�
�i�y���B���0�|�/�4�#���"U���2}��h��A�\��o��b0R�r����e�1�I�
���>=��#w���F�Г[A��}�6�jL}o��@G׾���m�e����q7�NzW����(H٦)I?�1 �'�����Ian���qkXb���;�ˡ)B��,�K����q�_m�Ό���}�;�+7*ij�6$���c�F��7�ڂQhu��_�ȸq#��9 ��<Dx
X�IF_#�n�t
��{�B�-��!EG�<4ۯ_Da�&��7~�Uy�w�bY 0�e����.W�]��0�K��ؐJ�ў"J�Q��
��r��6����ГT�����&�i=c��� ��^�.4��X�^J釛	�&0�[���B頽�'�k���jW<s�];G�����\A�@�Sl����k{#U��_ ���?���<��;���h"DL=��7��¬8��Љ����?��8t��
ҳu�)�N�N�&�rc~�0<; C��/hG���.T ��E��h���n�֑'��hqL2M���)m���>fp�1��0���N�ڱ��N�6)\�⒌�Q�u���G�/K�jJ�z���_���+�hn��*2n�ɚ?6�$&���ϒ"��ֈS�D��J��\8T|Bi�n�`~������X�%������*�9�Nrt��e����v����?�.jk�W��d:|�q;�$��P����﮴����@�ArS k�&����v��@r'�@A�
ٱEM�
nm���Xr��_u?�M��C��+��w�B�_��Y?�zV\J4-���I%XDB+:ԕ�?[��)1���� �0�v�
��U�~�� ��_y�<���j]K��!�`�?���k��ĒY�~�3��_2,��2�WM#R���!���/L}7�@2� J)E�:�	�e$^�J��n�� qqC
F2:��&�Jx��y��CU N�%����X���I�5��[v\�q��7팳�>"��Pf�)����u	kP{�!:��^�4=�m�Tȿִo�w�t���O��	/�7�5��=�D7�}��ݴp�����w=<��tI�T��[ڗ���h���`f��;�f'�ݶQ��h �Y�5�b�+��rK�r��G���C2��a�ȿa�
6�(R��όL�A=��6L�h����n[�8]��𮓭��ڨo�l��x����P��Pk�&�u��������i�D�����}���`�ex_�R!�8�+dq�2Btؿ��������`�e�wycW���O���g���]����v�顁m7c*Kf��8'�f'ƽV��@��F��4+b�^���&#`;\���f� _�������
�����u�~�unг=.hF�5��5>=���}���G���P���=<.) ����R �Z��MJ1��X��`�xe����t�������J�O���t���}B�f�f!t�Ҍ��Y��cvb����R��d�J�����op�J�'nȥ�ӗ�����cY�r�.�� ��[��#�藜��U��%�ALM��(J�U�rY��^.��y�EQ]�C���?��Ex�[��5��艼��w�*��ѡ���,�ɿ,L�� "G�ƦNY�LQ5�P
����l�'������A�I��t��|���c^JI�� �����Er�e�s��e�w��D��&����=�N�n�C���G��C�U��i}����Ͳ�}b7b �yh�Ƌ�oZ�~Ir�߮b�S����9\4ׯ�$�w�ؑ�"3s!GJs	"ʤ����DH�M(��GXq]��( e�nA�	I�uͨ�$�*?=D�1/���(7cI��H��2��Fo"q��g��w��F@lkD��A����׋E�v�%�f_�!4���ါ �6-o���.E�s
C�U���Hϰ�aG��Aᡩ9���[�����py,����� �6c����Xߟ�`TN����-�/`iM�[#|J���X��#MZ-7P�&�T^�Y:W�XHqd�3g$y
-u����_k�O[a�I��x�'��'/�N�2Z�q�2�^����d�0D���y s�2��f^J�R*�{<����~�Q�dR��@�<~o����bI�h�����7��W	�C�VU/*rt��ol	X\[H��g`����Hw�b*a�f������-o�p�ZG���ğ9X}R�闼�иFC��V����Ԭ��1�����8�V_+ޔ��c3J0��$+��3o:�F�O��o|�eҟ%�;�;��孼ύ&���q�K40��b�&Ѭo��|:������MvIQ떱���iz���� D��%�I�҆c���QӠ7� �]3|d�Y)�Ƴo���}1��go�!9GD��$��-B�S1����a'�.���31�.K'�}l�0�O�at~�"e��7Є�I������ ]�|A�e�}��ahp=ʂ^�����n/B����5��a��֞�ȓ�0f���YH����%]9�''��B��C�u��\�N�)�cS��^��;k� �VQ=P��e�QE���HS�g/�|��f��i��h8�����'�����0<8(�D|i����ڸ���O�*�,-�)5��z�	���X��SG��c��]��f��9�Q�`�%�=�O�t?S�q�?��K���;GH���;���I8yAC���"����V�F&���k��s�]AMf��޳bN�� E�}��*?��.����4 �����;R��Qݴ�uJ�#8��'�qAx��mt�՗�פ݋��j�aڝF�Uԁ�c�Ǫ��M[v͂�IE�ni�%ќkr��]m8�������z'�À�U�,avp��cICu@������9oC�%*}��<Q������.����y΍��Z�Tc�*�PM�R�.}�τF��K-�~I�y�js&�d8oe;7���0|v2��<3�21-Х<U<�+?�]
���ɼ�8pj�z��w"g,��yO�ca���3)ƉA�yϡ����t���ۏ��Ӥ�禾�`�g"jx��~�ta����,(�д�Q�~0oKf�n��\�a��y����4�w�I�/���VKQ�u{�=Kk�#�ߵ�ד��� \�0ݝE���-NV�D<�E����o�5d��efe���:X�٠���y?�ܜ��Ŋ@�x��%�%��4��P^X���T7�����(�� ������~
8����~��0��\��ɼP���Qk����j��igg-$ב�O6�ρ���������P�Vüչ�A����~�ac{�F�����z�K�)P�,�!"C(�z$�)�f#�P�d��zI���綥��nu��
,��6VA�b���K��Ğ��1��ĀI��f�OV�g�2�Y3�*Ύ���䐓SU���n�|7e*�,�l
��^8�?�n��^ %��*֏j.�kz�G��k�[�U��G��ך��U�~�ak�xU����ۂ�9����2��$�	@��`&��$�$�M�D�D��TC�+��U�+������xMM�S��'/x 3�h�����o':�>3�-<I��FY#�#8on	�˰��&��W�eH���T���S8%!<�$�¥Sd{6>�n@��׿�X3_�_����f��y"�'X}�p���K��
Ơ�Ϲ�?=Ti#r�Mh������Q���[������*��57��@�:^ݣ;s%ɠ�? v���A  �ND�kS�*�;4�����8#�z��y�l�iT�<�U��h>���WY�ͯ�ma=>̛.g�7Lc>�&��y(%�?�%�":Q��Yd.��������o�͕5�n�f�?�U��l?.�����Όo�#J�! ��<4�����E^����l����c�W5���tfh��q��^48��'�&w)ױ�_~�7{�p��7�,K̫M�`�U�Chi�d���$���Þ�T�Q:1�GLxd��M�1Z{���M��&�Ҿ���Ҧ_O'����!��>^�g	������űta���-���M=�'�<��<S>{Y��j]� ����]N-X�8>��zضg����_!d�,	NHN���Y�@��(/G���@"�F<O�LP��J`�Sݕ�
�{܋�qF1�WA� ׳�r@��W����N��^�L������.vYN@��&�:�f�$XO�Č�k8�5���z�$����w�1`���A!�^1"�E ����h=�~; D��@n/t�9�9����S�B]�{і�y���h{p�U:,�6@����Aq%� �<�%���S���K��q��Vfz��ΫYJ�K�|��7��y+`�M�H�k0wT����Jɳ�� �^4w@����k�0������@�N��;��K��Pu\R�ڠO���fဵ����]��أ8��]ػ�7a��>[��j��ܺK"����*\?�Aӝ�����	ܤ�������/��2Q�;]]Զ��W�B��آ�
��I y��~ؒ'�$2d��kn�V�c�:Um�JO'_�
��<�RV���	Ox�`r����X�o�M�I�Z���4k*�f��yp5��n��`ր`xȩw�3h��B�R��U���e��;Aq@u��}C������)�bg�n6;qp�!�ň]%ͻbx3�(�׉�)ľ�X��+ݽ1�墳��͟�l4��s��^���m(�N̺��=���79m�l�;%R�K��HԺ-6���J�:�1��[�E�-K���jDo��b{<g���<CT�#Q��}!߅��pɹ��.yI�;��OHl������W���e4�Q��=�D7U[Tw��	x��+.���֡�TH�����LxG<yʹ�I^(]$u��N��Yn�<]�%\O�Ϝ��k7�{�M�2�Q�f����g��CU��6{����6���|9��^(UȝȾK&M���nT9f������=}�y�.,_��%�����r����N\A3΂�A�{ᚰ���(y���B%e�#ŕ��~;D��0�	"���w�ŕқ�7Y�v�xu?��	v��4I�tF'$�1>(>�WkQr�_��a��
�F"��n�+�׭B�0	��D��S�٤�����ױ�۳���*@ޖAa���ldx�'�#�&k$N��=�U��z#�t��7�}�v�� �4�H��͜���"��>o(p�{�EE��s�6���[@�6H4(My�4�a[e�EL?��¶I9�ѴD���ͨ͟�x�]Ѭ��#=�+�M�����s��,�'�$kH�&J�s?V@]�B����u�M^��="r�bj�������7}�<�Hb��Lc��l8~t�2$��:_�u�����w��P��cwv4����+~X�� �c+�_9>��W	�Y���I�і�{� {�4!��]�	�N�:^��Ͱ�;juv�����h��8��&�V��e�]e5�!h���}��re�D^ <L�`�;��,6n�/^��s�CHL�3����*�d$	�q� ���(���F��{d�E
Pz��~�Nq;��koM��d��(�w"�D��)=�vJ�1��<�y�`ɝ���ʿ������LpI時���';3v&B�r5'޳>�o<)y����H|�5���N�;!�_%���������b��g3S#;gl��r����0l�H�3��R�RQ����q�(\`���@tJNe]����� n�Hg�'΋����W##�~�]�3(#��kӫRqvN~�n;�\��KӃ\\��F��Ͷp�\q�e �g�����f?�E��r����U$�Ґ��Yu]"#y��]}�g�"!�Y�P�>�dw��?31�9oFVw�S-�^uɩÚ:��"��1��n��z>��o�{�Qq��;�PE|�g�.� �[�1��P�,-_�>��7R��V������jpR]}c�7��Xq:����-��T���0d�qQf����|�WҵW�]�|�_��K;��\�;�:��P8Z��b��h
��t���
=�g�-�{��hl.��$F@%/����H<���T��Q��P��\��q�7��mX���F&�|2��	x�����d#��#��2"B�R�5��£p��_�*J����hpCG�_��<��e$����CX�a�Y�Ą���\�\Ѣ��'T劗L�K���	�����'���ӮJ��8��a����1Xc8���#��K�x�r@���[oj��yMѭdp�29*m�~�w�SiY3N���#tR���b:5q�'��
]���Z��T��H��HK�K'��D$����U���m��� n�]��5�����s����	�{������)�(��4TcX���[��7�!�x�I�2�n��$�^��G7��R�o��q��X����G�'I����!n��$����j-��]o�rγb��=�)�=�)-����G<6�IUB���6���0f	~":��<�\?�>%MADV.cm�c;+C"L��A?�#OS!��RG�@�mx
� 􋔮�~'<���������YȌ�}��CPV�cv��Q��n�v����l]L����Lk��&����`h>��y�P�1B��3�6\z�9-) h�����B�����8�Pz�[������׋�!��G>�Ț��~��@��+\���'5>c��u1rH���Z��y籛k�.p�������G�Xt���'���\�M��ɫ�Ww�!˸� 9;E�¿"N�n�^f�&'�r/.$Qk���`��� O�0f���O���g">_�&�V�s�`�T��y��	aX��'�n"���%=��_�+���6b}���r�ؔEZ2��ÏUg��Ƣm.�ҬH�o�:a���o3gJ�m7�_cE�b_ﳿ��b	�x"^B��o4�������{/&�k����i� ��nsŌ\�߁��pFV�!�
�̍�Mu�=��f/��x�i`�Q�	�l�Q�O��i4��4�g�@�(1�Z���୲�Wo>��)Ie�
V�C���`� �B�+fģ5�x�F�!�����-gn�*�
���`�|����Q6vބ;���xd���L��'Poe����4�Y��/�^��0K���2��PyS�Y-�~�+����~��xEhC�d�a�G�d����%r���ط����,�	����tvy�p%,��(�
�e�,�s��l�7Eʈ
O笭�C����:�d�Tw��8R7dz�|c(�Ż�͜�~��~{�g�`� ���v]g��.�T���տ��>9ed2�t�x|�b�3�'[�+J `UNh2w��� |��<^���3�xB��ߤjo��� ��E��3�Kh��C�#_ up-�Td+�0�3��<��^�M�9���3"*xTR�����":�QO��WQ�h�7�7��	��RS/U�ۙ(�g�
�x���Y����"k$*��VQ,Ź����T��w��kOm���^>�͖�^�Y�6V^B�	�#�qKk��%�a��v>�
�w%2E��$��y��T��0M�W�s�#���o;�`A(ҰI-!�pSaQ5ӏEƼ�ɠXT�*��6;�m7�q��}�W&��d�8ؾ&aɢ1����O��Y>�n�W�2��BK�y�t�5�c�xB��>=�	���~y.\e~u*|�V9%���%ӟ���,NT��~5��i��r�t��<���t�C�٩H��94�b+�Ď��[
H���fLaM� $_�j7����X�����]߃�����ё�~�E)�@ HI��]<���/�:a�$�� H�A
!W@Fk�kG����3�U�V,�� O������bN��aamM)���,p�H���[��|�5AVEfë,�;d�U�l����gG��K�&�B�b$���Ġ����櫮t�'��mP]�b��_���}Ea:Y�<.�e*C�y���6nn�`B�;�������zV����Ϸ��̲}b�g1�'σ��c���QD� �}��E>NY�R�ю�9�P�ۄ��2#��ZC�l�ϥ��ռ�b���'j���.��`��%9�f�"���ͨ�^5�'��h�ր�����Ǟ�_Ҩ�:Y��ŀܔ� ,���_Ԭ���xd﯇�qA�H몕v�����Yr4 e��e^+�i�'%^_�KkQQb.��`��I@T&D����f!��Ip�����&�����6�n�!1�K��r��&�g�S�k�CbӫG@de���	��-����i�>ð=�+��u��'/O>��2Io����'�,�H������,x����ho�v�M<���@�O���S�׾Azm�4����5�u���ݸ��}�Nf��r�z7s��"�!�(��j���Nd	�?��t�:���,.7�x�gE���]pHlƅ���&�HPY���x*�X��ۦDv�"�y��<�w^��ޕV����A��𡫌_��~ῄ��@[Jo��%̎��/p����a"S�R#�t#�`	�&���UT��,�v�?{�5����,��!�ճ�>���^/�E���·�=o�V��ZX�KN3G�b� g�����F+��W����K\v�އ��@S-U�m�@��;����ߎjq��@�C� &����>5r�9�,M�XBE��(�.�v�,���*����ç`�3�#�B��g[E�E���0�PCص
!fi��oB�E�*�w:
2=�m����;B�B� �L�:��i��m�eC�3n�r��\�����7��Ն�EE�����n�"E�0��5f'KT��q�s1��r5�D(�����.�J;��t 7&�:�x
��FC^�M-��C�6KG1��pG��mT���h[Q	�ߍ��X��}�/�"cK�����,���9x�" �R��QK�*d䃹��=_?�.������\[�	'��D%Xg����7���JD~JH*9fm	K�kU�*۸R9��Ub��N�>f��W��4��TҼ=NЗ�"AÝ���/s���1N�Q�]D���u"����9�bV7�z���^
����	�7�V%���Z��}V1�*��l����eF��۝c�7�;�1yn��CyE���{6���/��#�*�ֈ� ��jK���9P�)*"u��Uo�B�,��ȿ�)�y�֮Ŗ���˿+;`���`;B-d��VFI�:N��״��Q,�m�Q�)ϻsY^�����G��0�n&��e��d\�ۛP����;;�oʈa��z
2"�6���,ɷdsY���*�����/?(Z���W���f�]�se�j琵w?�vܑP(����ٞ�筭h�:<S]��(:�2&�/yOM%�9�zI�Ɏ��oܮ�{L��Yv��)�*��xϖ�1�@x��;�����f� �2��z�a��Uk����2 �.��xN�*���i�7gf��FgO� �`�l_@�ͫ���m�J�����ј��=�L/��,�U{��-�kX*���
�;m�*�ik�[�y"j������g5�+\?��,��,����<)[�Q��9�z�Y/�ݯ%`���FYɬ����o�/q�����u�	�zA�~(�ՙ�(�B����N2�'g���oAɩ:a�ښv`I��T��VOT����@c��m���qJ�L����k]f2C�������V:�M4s�����ky��C���7С��/��t1�v���ܬ�����x���*��%c����BA���"Xr�8��F�0��R�c���/Y�r�p7�
J�
��L_K_Y+��#K�e�nV����e�����i��D�.v���PzNn@���Pd[QI4�Z|j�/����C�
:�2�f���d��ol����6�X5]�V"Y��OS��q��m�	����e�$ue������)wzX%��� �$�VD@��Q����
���Č��1�� \0r�{V�a\����v3��1�BYË
=bW�?2y"�ǑoK>p�s}�T���W-��./H�op��ݦ�THeO�pL�<��ÀG^�GUG�=�mw7�t2k{'rDWc��5=��-I���Έ�u�T4v��(��E���;ͻ#�!��z>?�ʭG�-���i���|v@�;TDl������m�:��?2��U�;��I��dX]U	�}���~��Y\6���5���7�P�)��P�pv��7�����% ��_�_��~�0�rϲX����G�g�r}�W)3�7�
��A@��ur�� ���c��@�ș���}s �t�ת�,�J�L4S=h�	��8�ze�3���)�.A���
	��[�_��P,W�Rc)ç���v�#�)-�/��V�� L� �.0ϵ H�{�Գ�i�K�����sD^��;����Z�? ��}գbԖ�"m�
�����F����ljy֏�y�%Tp*)V M��^��G*��w�������
�ٽ�P���.E1�Z��c$v�vF�X7b����|�a�ndw�-w�R�V3˼H���ұm�o��
x��O>�,�Q���'E�N�
/B��Y�	(�Ae���ݺ�Vy9Mm�O���<�`���)p+�^'u����k��A�oȀu�'�����$�rUG~�0���)���p��>��@����c��+�+P��i���l-�,��@p��	���v��I&�jC��zF\�1�㎱ ���t�;|vy���D�DK]���O��i�7D�.�5!�(y����K����Ri��Q�G�W@��ypF�����q���@Ȁ���?��u>�ղ JY,d�����uİٻ���NaS�lC�rS�*ua͢i�W
T�5��h@�U���$p> �q7�\�V�1��Hm�e0K��S�!+���.8wJ�
]>�͍��]!���K�qP�mZ׿\VJ~`ʢ ����򿗋��f�Q!$�b5�I�K�e��{�A2i���z�d?�	��R-��)j�-��a�`x��1���xj��1%���2z����K.��Kf2b��o�j�\�h�4�n���6�AIf�D�=�4����u+u�q�`�R׋���U����H���X��LW��k����{k�P���'�Z�wg�8�}���pE�ԙ�W��I��j\�jI
|}�8R�,���a�&�b�-��`�x����$텺���@�I�	f�ļ
�ީxfx�ͻ��Ri���_��P�WXd�3��<	�xa_���'���Ls��p�p7T�a��*�MM�c�Z�ϳ�7+خ�o�F$ؘ��A�*�M�LΉf췪��;�z�$4E�)}����V3���W5��kԯ�"1�:���#�B�i+��k�w��_�@R��^v�'0��<�fp?�
��P�P>��}F+|}��ou�/�,���y X���݌
hT��I\��ƻx�^�P�0�'�����-��Kr)7��E��vpʝ&Ls
%�1�{��E���u*�yYn6����{=�;B�s�H��IXWǚ�E�m'a��ҹ�?���'��6�\���K����
�M�sz>d�7E��\�;>�F�YӋ��!t�o�����ST��s�L�ը��4�:-����9fጊ
��j�4��9\Aw�z�����/w���v�!�SL��ߑ�z�g�ь3D�(��xF����>���\TD�-�ԙX�m��X�o��څ�`�B	ɿ��<Q7���
�m���k)׻�9>�$w�.�V(�P�IRG{�I ���ZVt��w�Q��)y5�����EfO����L��/�d�,�3-h|z(�:X2�*��ޞ�/��p��	6�^�9싫��.W����Vƥ"�z�'C�x����%	��y�l2�����e�<�d �<��'M\v�6��U"��O��U6��
BHx�TF�v�}��\@���2�I�@�GO%5�7Q�LYӹܼ�mc3�����!''!?oC�9�����Z����vtcFhj���Q�V�9[֥.>7�엟��]���!y# ���� �^�����D�㤟��_�L�
q�8���-��;	f�a$���D�y��()$>t���7'��M$�|s�-��(n)T;O�͙�T>�s��Hs�u�0p�oM��l�ZPP���K$-��GI�����O�Dc�"���@2L�x,1q�ݚ/���	�4�] �@��S�\=���2u��c������1�i���e������q�29=���RK�)hNn�*����I)�����A3��d��)���K<����E��p��/hA^��0�.�@�V�/\z���	/*5؉ �V�ɬ	,/�˔C��@:g/���Β�� ����o%��[�,�^͠o:�N��>��7���vNA����VK�蹕[*��NP�O"_b&|Eʻ�"N�,�,�.�SY��IX6U����wX�������C¢z�^�Z��"h��P _��6g�_��!D稟f¦�CV���*�oiFGi� ���$]ͅ�gO�PE�>��#(�/=���&���/PG��A�69������X�������G ��d+���;&G��Sr�Uj�ՠ�*���Ζl��ݦS�j] �O:M	3�����(hS(ڬ�����c�vJ��$���,`�v���-�X�L�&�l����$L1Մ$���e�zx=�;��e�F1	'�h6s:�i�(�RWV�w�b����do��'`h겹�'4�k�=�N�����yx�W��)�3�tU+�J��U~��SV������q_�ӛ��7�"C�$g{i�k��/�F�������d�J�L<��.�����Җ*�Rȅ�J^M"�Ke��9M�:�ϼ�_8�t���)�u�N:ҙ���ƺU$�.t��������x��oy(���;Z��PҀ��(���F��C 	��2J6+[��A�
�1��|7!�@)��v��DP'���ૹ�� d#��Z-��g��ާf])%1�B7z]�z]{�,�,z_���p��� ��2��p^��OBK ީ�+`!m3�����0B)�J7�x�"��^!?0Q-1~����䟽yL�]I�C�������;�����Z�c�Ai�+����3��|w�Oj��?����A��A�}��V����,�TK�1��%=�a�m��y�WH\o������t^��%,����Ӗ��c������s.J�UہS!�3U�R�Ϳ��?f��A��|����A����}	U�B.�`��#�ܮ�V)@�"�e����w@RA*$��F��	V�o-��s=q��5mC؂��Iå[��.��^�6�py�)��"���8`e�ױ�O��n�~���F��2�����Yr���5,3,w�rhjd�;xm[���
��jKϔ1���e�2P�c\+ųN�H<
�'���Cp=؊`]�o6�2�O� 7�J��ß���\(���we�|��uD��]�$��AڧP���0��l���@3&��H
�Ο�Q?t�'��9�o��S��U��P��f��P^�zWHۮz�n�p
E譑n���鵣���&)��lp�1��ݮ��%~ܺSH�->�[��*���7,a�D��C�Ll�!X�ﷃ�<݃"�i�s�
��X��(b���i�A*�K@��/���c��Ȩ�����a��5,P�މ �Cb���P�bҋj�0�s���d�F����)�������H#2��oXB��vG�F�e��5���fN����+�:��"�_�BL����?�_Nj��I�!��_���ON!5 �j����E�@ݿ�c�#���8�ʿ�m��t��O�_r��/2�;~� 'P�l�r��l�V�0Ć�[��G��c�Y��S�P�4���*�,L�����c<�79=��DݕO�Z(�ֵ��nk��=ĉT�D��KU�~נ@d
�ۺ��w�`��#�۲Z	%�0�[T^��iM�o���Ղ��آ�`DS�+=���0B��ɦ%#
�T�lg���i<�s]��\�xv4�^!�(O�p&�N�s�o;r�߱�/���#�)�e,���Gޯ�g�����*�v"��w���p�4�b�L۪F@�D}���br]�`��:Q)Tڗ����U���P�3��_�.��`X(�jڏt��x�����ۢ�PS�v�����15�~+��s)�g
���b�2�F�g�L$<�jN�~�~�����b���:�
��4u�ы*�K��lN=�ܗXo��y����;��Y��7�<`5�i1S�j|���K�����J d��k�{����ܗN��54uT��`2Q�NSFh+>��RiA��֠]�Xp?#��6��;�v@�"�ǯ�\q�7�%���!�j�Z��}�ݿ�~$�}�����}��S��=k�b:I��w�/A�9:lr�+y�sl�P>��S��xF�d�WBU�6�6��]��"����D�-���;��)	��(�Tzw��������t�&��-�T���c2�`�b�.��z�s�1P��v�d��z�hT�[a�qDq��CX�`��u�<�-y���BU�u"JnV@��=��w:VcŰ��~��0�ċS�1Z .m��W�0�ꠈ\��t�w��1�ⶪT�E�J��9��O5����Eв���<�r/�T����MG��Բ�b��<�ZD����1+ �-�:��t�(蚰�W�#��xx\PtV<߀����U)��?����_1}�/e�J>@��Ԕ�8��f�WC ���'��u"�"�G�׸S�bX�W5��M0`�Z;�WuϠ���(<}��<�)�RZ��?��Ұ�f�ȑl;!�N\з*+��P�1s�*��w�9}x0�<ˌ�f\��<'��?קő|M�˧���'�d�6h���A�)]��d�,�וʵ����~�vQ�m�#����'�SZ)D�6�F�ՐXG�i�<X�=�H��ƞ~�ы=�u���>r$�����G5vr�0-����κ�zN�\1�9.��+��6���'�(Yz2��wp:�t�`H{��Ɨ�u�g�oB9'�ǻ��W�c�h�S�Wוֹ��)S����;����v�-XGᱦ�ʍ�"��+r��v����`��"7a��sTr��*L~�'��i'��_U޵��I�E2�^�q�d0���m���C04��9o��1�d����#ؕ7%��Ժ�ϕ��/�D�],5�ƿ�&P��L'�ڱII�0t�� ��!ꎈ�t�E��Lx��H[�n��8
�A�,�w�Y>|�"c`��p�2�Uy��i�Vc�d�~�fp��ř�w���P����$�+���)�<k��<�l��O��}�ABp�tғ��\
L$s��i��;��
3��c(6_$ß*7��B������ţ_͖ -d�Qn�u��B``���p�9���D�z��1��k^��#�����Y���5� ��b>��ʸe�{��t���hH�g��>#�l�I�ck���[_��N;���O��h�Ey�ӽ��Λ��Ĩ���tty,2 W�J5�[�@P���Ű�h�uC�e /A�$T���������H��&׎��������1J��` ~��"�oz�%v���-G�e�چsW��p�;�ԓ��?� ����|�Q�������ܸ�wiO
|��'�6n�>�@���'�t�?���ke]�ʞ����Ђ~>s��M��m����2�肁��4VPɐ�is�gQ�~�?x�Ta,�4}L��ŇYBw��r�Q��<+_�����<�$R��F�N%�X���-�k��̖+]z��L*Y�n�%�>�@�=s�43"����(1�����T���g��������4����3�f�SMZ)zV^��Hx%p�L��]�6�¤��<��/IX�����R���g�cҚ�V g��v��>���k��`�BLv���8y<�IY�ue�1OCx�2E���ZL�`�4�՝r��P�|[ɟg�l��J�C�ԁ89�~/G���0Kb�/���q�;y�k�����+��1�X�ڷ�M�5��.��6��Q�;$4#� ��ʔ�����?R�8�T�F�O�1���d��,�q��g��D�y���<3�?<���`��JU�I+�Q/�ݎI�C�9z�u?on�~y�a����{�U���_���Ŵ:;��Xz_|��`�#�V������B���6��dE"��h�U<\��ߟ�c� ��6)bq��^�b�+|���4�g�iRbN���&B R�����������|ɓ��Gaz_89�?}N����н�uQ?��U��ܘ��B��&�������|���%�0h�]��p̡��Î�B��)њa1���KV�g���b%�������K��^)U��
�.	���M�^��6��/�2z+���I�����3ۨR�-�6\t�`��0�pI�f�|�ڌ,%E[�ˉ�h�r�~T��l��χ��{؁ܝd*�
��	�%��	��5=�󘐛h���+���ć0�ƍ����If�i�6ز��p��;�+���ˁĨlb��1�H�N�4��Ф�M��:�(��y������Iz�������LJ,X"���$�s!x=�n���]
j W5奓�N��W ��t�i�C�Nw��T@z�^�*K [gPQ���\��<A�	�#Ki�B������h�����Z��D$�]7u���C�q�;o���Z�"�|O���Y!#8�N�n���/��)��i��*��MaQ�_�-]�i�ʢ\�°�8cx!���@�2A�A�V�*X��L(�e�|krO�H��@�)�#��48$4�Cx�q����D�#�Z��(�9�qGq�H�[S�{j��27�~MIC*c�l9�5 ��xz�@õ�I���{�y�`^��WX�ބ�>
<������,���R�sDZz����W~�qy2���o�|�^������Uh��?�1��f��>Y���Ƚ0�J-���	D�]Z9Q�+XP�η�#:Q_�J��t!�;,n#�����S�3���g�[�We0�IQ+3���*�x��X�^TUh�E��I��GX��
��;���*�[4n�٢=',�W5�`9��ߴO#�`VW��V*���]M�י���x>�D�\4�ל�g�Y|$G�cY>:0�
?U,�����'q�S6�C��A�?Sһ� 5�I� ��['0��_<gM�*�9�M��}��c�Ƕ��<H&Q�8�Y=���82y�0.e9O����sY�#�d�����>Y|��T� ���wI����*[���Q���Ks�̠;�ͼ�8���(�>sP|����b�Z{ǣ���.��"�}M�/�iI�3�y+�*��^	q6@�wY��.a5�,���B�ʷ��[�d�FO<q4�>�s�9P0� 8+�k2����O�bo���6s�ͭ(�^� i ��,͡ �9�ʊ����>="��Σ����Ew9h Q	[Rߪ��é��Nx��R��m*�r��	��'��Kn��gK0�k���EبakROI��f���U���suI��<�C��_��)\)��E���5��~��\%�2\y�9���.S`�z�+IJ� �WAc�������;ڷ��?gݺr���*ݱ2��Rw�6[LD���g~w��nLp�[cƫ[o� usQʨ�a��=�r��߂Q�X�^�&642� =��eL��z�@�gv�tU�f����!7��B-�T7 
:����v8?���wE۴ �,�#8�EdQ%�9ٔ��Hp�e����z��f��ʯI_ґkv#Ƽփ��:l���K^�bĩi�EZܮ��o����{��A��2�s����7�v�w�]LK�WȪ���k�G��#>[�Y�q��� b�Z����Ճ
ty��C-$z!>B�$K�#��G��~Fk,E�Vd��p�������S��mc%�C���H��ڰv��F�95+_<R�m�R�@`H[T�|���36��-��5����p#���'�r��@��8G8 R+-��|�E������ɓ(�2g^��CS��K�O��p�N��e�|�I�
jg'԰�8
��N5�i�i��h[���ϥ:��+��i#��iN�i##'�0$�<����[��7b�ͺ�.�~�:y�h�$aH=wyG�]+Z�עC%+������9��__�}�D�5�P��g��Ծ��*����H�:��3�|nÇ֋Y����vR�KpʹK�D��F#]�e�N����;�X4�h�ކ��q^�b�����g\R���c\���r��C�7LF��4��R[�σ��n+X'���������~�Ի��f���V������t���Yc��&�2'c�� `\��C���k��MA���l9������3�X"�	��gz� Zx�G��v��>OP!���b���V����K�u=�%|>恕.0[��į�q$8����4=����m��Wm��wW��)������N	ȧ��o����`yޑ������D�XF�F�d����ݛ9��n�����r�++�nB��o|,��`.���n�ӑ�*`T2bl�����y�;�'��;�}�;�Sw�T<�~��V/��ecܕhO3�Zvg�W7���$�.�[�~G ���t��Ԫ�1C�.�7D�@w��{�T\����мB��>n��I�/�-��+2�5���i�� @o���\܏���%��ƶ�q���}������ܶc��,�t�+&��?Eq���PB
��V
gAmN�v ��^��ԇ�s/�kaq�54ϬϞU�|�E�}�7���g>�#�⏲3�V�tt���}�E��.���pi�ܟ����;<`��wEO/O����1�u ���[#�qo,dy��^;I�O�tao��N�Ck]�Y�N�avG� �������^���,�!�y�tn��?n���+��+�o m���t FAm
�{3#G��@"t���Q�/��+Js~��Y���>M�37(L�c���R�#��*F�q�l��{i57���}'d1���~��_�F9�l���ZKR.V�FS�����Z�5�����/�1u�	Aָ�p��擖{r*j��{/ߐ1lc�A����I\��{�0h�1��<a���	{�c��D��>��C5<�[�M�#ń�Y�xr �w�K��L,X�1��;�KS��3{�� � ���4~Xn��w���i���%�P��]^�*��e(�]'�ᇸ��KD���o�n��	#b����̏�`����i8cC���'���d�v����r����-J�la̨�w�>��%��Ќ��f��y
��o'�~F�G����H�"�.|�<c\]0\��H�_�Nh��N���"��0�j	N�^�d����M��v�k�뛕�������5���p@�Ⱥp���9�~�����_���}���H��ڳ�YOC%z�I0}4�ӥs��S\��R��J��2�%����ZX�����%����U�ܚ�Q��Ϋ�����C0���@��J@
Tx���F+7����ׂ":�)���<l����]*[8p���!L�%m����:5\e(����ǭ�Q�=7�+6�qa��#�\$�a��U$eyKv�'��B|���6�q�E�����������2$� m��C?�}�3�w��n�B�a`��s�^O�=ٙ6i�-E)��b�-�OX�B�C��=�d���DL	�`�+�Qʲ� �yz���i���M��,Ŷ<��W�qV����7M^�N�p�O�U�Ym��d���$@�K҄s�9M�L'���/qc�/�\j�4�%�����x;m�)fg��H�C���He����_f������8��i��
}��X�Dj��@���=��R��D]����ݏ�^Q?�0XV�����L���`��H0��H@��#,/H�A�c<�S@r��QR�E�1F��8J�oS�C����<2���VX��[V�Y	Ie<߭V��*�5��V����iNvj:�)�*D.Zkѵ+��m�chL^��(b��H����U ��%�1yE�in�nS����n�B��5�e��P�W���=��C���"������#i����k0�q<u!�������M|ߺ�ڌXJy�1���;V��v�m8��
��֨��]qz�/��ͥU'��F٬������Jdl�l���Y��u\/p���Lu�A|���D��� 0<h�%�2x`�>D;9�͂CR �՘�K��V��1U���̈́b29��k��;���qz'�֝�ܗ�<��@_7q����s�� \#J̛�B~�U���CA7-=!�u�DJs�7IjG��.�.Yu#�?����w����JXoO2*j�JЃ�}5�E��Z7\��9�zF\ڰ�Ђ�>��P�؉�׬��=�f�wy]��]'GCK&E��c
�D���=q�9�Ұ��;d�B)�m1"�C+F��o��ԭ�i��m?��3F�5}�����V% &Z:�GZ�g{f����-M��7 h��� �;��d`w:�i^m����[Vss���<i��ob�H�]�7�?c�r�.##�Cp����LZdĕz\�`��GnGHP}"�Ռ8�����mԯ��H�V.��*ƾB�o����`4B2���$�����c�ڞ$�|,�.�-:��m6�P���R��H���J����I��:����K�����4�׼��4�y@�=ZV�j�ۦ�i�)3���"~��C�{ڗ�����b�/@�a^�A�1&㟜��	�
)��Qu�̐���2�	�I3��T`��0J���!���˻�q��&�:�����|T�%�dym!����2&?�@in����+¶حD�|�v\"����W�"$G�-�$`��{��<�-w"6h�\.�?Q>�Q��F��e���� �ҝ`UF��3'!J4�	�ۭ�s~��V�JC�������5|� �λ�/�p�<�P؊ћ������U)�9�(1<��"�ڒ���߅)��3Y���L�q9�Q{1iIp�#��ϔ��M�z��ȫ��i�nt":�C>G0K�i陁>F钨v�1ё>fQ��}(u�}�5{3]a*�5�>���"h�L�w
a��3���z�a>�� ��+�v�����k�G����+���ý�+�'�^�?)S����~ǋ��1���TZ/� ���N�F�͌�2���q�>o5[�!O�� P��T�H|�4/�I8�+� Y�{�{.E-E�J�0�](��4[��7Z{�S|�L�����* q���K�Ɨ���h��H����8�*~��%��	��;O�A�j|�w-�m(4H��^u��R�"�_�XSg�tBE#Ԅ��q����p�ܯ	�UD��풙��H ���[g�H+	�C�f`[V��1��Bn��S{sYLim�{���̟PZ蠠 �ǰ�� �B�c>7(j����HLýN-�f�ɩ��2�t�)`�πw�G�|�)A��"D�`��SC%��J�+9���s����0`A{;�w�r^䫏��,.�-���wX�6������xd��2�ԓ��� �����qDv<Cl�M�D�%�ԝE�ҁ���0�@
v�������@��&���QRn��9m�w�wCXQƹ��(Q�Z��
<<�?�����<���w�E݆|�/vt{y��+q��7�Z) ��$�J����Y�}(�aQM��5��"�\��$���z6t������8�A����x�,i"*�1��i��J���N}#��x�ԫ�ٴ
�\�&�^YyTa~I�H��u.��e�#����d���⠏hX x�C20uϜ�輝_�!���L��������U0��Z��tV�v?_l2l��4Z��k�Gm�:6�F�Ŀ��5��~�ONo�Ч0N�f�$u� ��S���HS���6�+�3�)�w�}�����N�B�B�>Q'��i=�-���ݚ+��"a��H�je���:��H;WQ� �O�i���q����}�v g;�A�~�������.ңW��r{E?A��Z���ٌ�gx;�Sie8��Oil��=*�V�a�b�O�0U��`̦󓌃���Ww�1�e+0!8N�:x^6&�����a� ���ǃ��`��tL.��T�^;�\��F|�O��I>��by*�	g���ulfSW�*��?_�G}e����|{˿�85c�MPs�`�N�T�!�)}��!y�1sX$�4C��Y� �gX,�к���3f���N?�E0�L㽱�������>X2��S����X�A"!�z�r�fۑ�w}���+����%��[�1�d� �k��	�|��+4��<x���q��b	�����q�ң��C�S�ܥ�+Ś��t�͙M ��n����TX�*����,T�̥�Bm�5Z���!)/2
��� �~Ui��0J�}���+�̈>ȲZ�ݮ��E��B@s	�����Je�,!����ؔ"
b^�9!�˙Lgh]>J7|!��"X�T�����f���*7�O
H~_�o�Iƻ�d��i��cϻ3�}F��[�Vw��|�s g�aОu�r���?������
E��M�h�0�<�b�ȶ��b�/�I;��s^l
�2j�C� 	����=C9�`,Xd�������(Ep֍ �Q����D�ٹ��T���y�����w��;q��fn���mi��e+]��Ď���[�`7a����++�'�$�<���l�[c(N��Y�+�P�u��;�B�5dk������Cg��	��ptx*4�9^_{9嬜�
��4���o+݉UǓI������a�{����/g�Ggh4W[P�r\�L픻7K�m�ɬ��{q��D��-JŘ�|�[�Ŭ�]x�{V�V�T�vm�Wsd�v�{�R����)�=uʗ�ٝ;��k���>�v��Whj8X�[�
��;F�>�LUz{b�����W4nشY�18~mD�Nv���Аp�D�#��]ظ�����,��#��dс?�gQ/T��b'��T��k��m����D��c"����4�|�S]�7�~�w�����nV��IT�a%Lj62]��N/]�ޡ�lg�¥DfJ=�k	��ex��/��A�T��~h���T��ly{��a�v���"=o���=&��3hK���}�-d�A�ܛ�:��(̌M^�R;b $�M�&ˁe���s
<B� *�$|�@n2���n}̤�c�{������6��pJ���4ڨ�|��k� �@qE֤2�1|��y��`G�7W6UYE<^�oX�`1����`\o]@��nt���{&;���sx|2���?�n��]N�aI��d�׮)��p�d2Z�gĄP�<A�B�����Jі��i�r��	I.e]t�{�ap�UX�����vo�1�94��Na��@��!�r�1��r534��]���e��Q�!���.�A�{�׃g�<Fڞ40J��8�
̏�quǘ���?�,T�����R�r8G�eL���	���+�n�)Q�B�4�
��Ot�wd�������%�&ń��m�p��&�/w�D)��;���d����L���<�mBA���Cm���ynr���SэH�/Qm�y��;����C[��d	������"NdqX���i���	�����h���'�?�L\CW)�����r��Τ:g޲�F|�$���؀��P\"�׊�ݗ)�Ht��5�i5e��vG&��q�W�5J�8��y>Yw3}p�4�M�[ށ�95e�E0�Z��z�j�0�W�t���/���F>����$c����U$��b/)z�*������C<�M������h%�^�'�����9�*@�`z���U7��ݓ3�\���ORʤ-EƷ�ʸ�)hs�!���� Po�����~�L�����V��4N���b�3������(���r��\���~.|�i�J��A#�����Ѣ$u�I��s�L����e-T�e����O�ώ���꫖��kx"���H\�[8���ey,V�+�?d��k�Ds�j#h��Gd��H+ɏT�g�0�I���8j��f��h��!�o��KFX!�|:j�A�b7J��� �Ol���~�����0�(������f�2*<4�YD�g��rӪ�A�
��4!ȁ:��	'/�T�l�TBd��h���퀒`.���aR�o��9�2��z�l̪�c���R}0[��jCU>K�E�LJ���h2�u��,�J���Ys�5��O�Ѯ�k�J��G��؂`���^hP]����0���Gd�}�sĊ�<g����i懫�{e��ֳ�;�k���5�T�p�oi$}�B+"TO�B<�ޮ+\qOJ[8�8ŚM�����Ǫ(��G� #|��Ǐ��K�O��#x�%�?��d�/cǚ�5б5�-�rF��4S]p�<:�	��%�X����v!�[��[;]Z�ڙ��y�v�lj�Lis�rN�{���}^�z���g�bG5���;�c�������0H�.�2,ԉ�|�۬���M����ݑ�7kd�h�K<�h�4��y[>Dp�!��F|��t�z���4���l��ʏX~H!J��"S���LBiq��:s�<�VsL$�����4�o�3k	W��O.��5?�;i0�|�H��LE<�.�p�W��%;��=H�]{m[����%�ļ���Ȼ�i##�-LHu���rd�e���6|v�x�;��G̥t/���h�F��\�p���-��6� ���l���wį���S>3��7��e!�WV�;gY�J����(Ӽ̧����O�D��4�<��߅�n��CL_XR��.�mYv����x�� ���L$ ��`.��8�ckn��&DV8��hF�`�`M�9�n�]��)�=9�U>~T��qһ<�'�L��
�3=�+��EF��Z�ko���C� �������;��e���G�g�Gِ�ٹ�*�+`���1�U�u n"�d�����OΔ�Y�����(�YpN;͍W<��}�7��T�2�*�q)h�	q�I����Z���!K	�S"�.��9�������Z;W�4��nڛ,|�A���^��׸5n�鴺�̯��_\%�Ar���&�3��/�1�s{.�7��XS1�^iV�?�'Q�����ʴ�����l��;����}�a<ʳ�-���#2�S��I��:K-<xe?2�1k�7�OҤ$.p�a�#�Y�t"-��"�ة1̍�O���b��@��E��Ќ����2��q���習�R�6�<]x֋�x��^�`�_��~,j�&��|kEL�@^PD�5���% 4����#��F��;VU�^���������k/�%����s�2!��
6+lg׫�=�W@M�g�)h�.1�"��"@��un'���3Г]EU�u�it�������� yGo�ג�~7���- Y�y�]z¹��b��k<*H΁ �}���.T�H1
���=MP;!�}�7�6�M������#ˡt����c�8��B��Ig��q�QS	�����"�#(	�`�]��y+$�Dǻ�u]y2B�8���|'(�Xvcm��T�J���/�j�r5#�]d҈����3��$Ņ�&������{�GIS/j�O��u��tD�Hvйٿ*5�@4G��ޅT��ǀ���>^��`ԨB)\vz�e)�n]��^(�X�.`WWX�V6V�8|����A�l��.��,��/'��[j�݂��N�����5cz/'��C8����x����"��������}s~�g�8;	|<r�r}��Q��zW�'p#\l߁��Qd[ ����u��C�-W���N�*�?B�2
x�p�y��t2E��\
X�-�@�����,/vx[t�0r�$���1��n	&y;qȌ��w�����߶pM�X��a���M�7�L�ɨ�n�vm�pQ-�C�,��@Wb�}K���4_A�-�-��W�V���`/�h1b��s�y��[��/�O���l�b�g��+z}1Fe�(0�}lgMߣg?��#�g�8��~(�B�9F�D=�q��(�f�a��n��~s�3���؃̌)z���g҇����_�Z�X���@}�g�M��+�aG���>���wEX;J�^�I/�M.������2�:��0���(�ەC%%�l�Oz�?��3>��>�,ԬS�iNSb���E��B�SU�E��%>�����a�3^���*�؇�u�Wz���	���z�i�s��M蜕8<�#�Ja���f�Zδ�٣�U�,Y��Q��c�;y��¨�]*ض�h�pU��gN��W����L�H�I�`�Bw��^"4�<����[Y�m�뢗t6��"��uw��Yo���%a�!/;v��;JM��˽Ӏ���N�O�~���5Br��J�u
Kb-ol#[+Xl�첾�>⋹~x�2���dd��t{��� ��2�l�m�r��ft���,
�h1��F��d}r��P�^�����U�B�3!-?mos�)v�?y�<��Ρ�D��:Mux/�8$L�o\ sHC�_�!&D8/���?��J�B�C�
ub��m�\_�Ϲ�E�u� �إ�=�*6�M [ 2����������(�y�Ks��#��V
8��ٲ�����n���������A8�����1
�Jf��H�P}qG�c(I��$�mfb��(gdKn��ߏB�R?��sh�s	*ˡ&��8��Q>�A���h�`T��_�R�(pG�'��-u΀�|�*P�4�u0�҉���d�~B�"k��5J��F�@?�g��������$k�1�����k�G�P��B̊k71?�Rthj�Jx�v�m;oJT��E3\��~7V2+yޢ��=��(����t��i�� �m��2L��~��h�Z�7���C�$���tC�0�տg�\��vD�����_!��Q���oc�F��gI�7�Ĭ�E�b�a�{�6�v��|\^L'�1��M�=�@�K
})�W�������g3��z�9 !<��:�W���˴�E��('LB4O����@P��&_-��s$v�1m��P[DL�M�c�UuB�*�_�n��Y������C�Ӌ��6�i�5u��uJEON��{�fR��p*�Gr�!��fY�������<�v2���t<�lD��T�E�R�[���H��|U��f)*
*���q�W��LH��)v�x[���'���@4k�����a�h+�����&U��,��/�p>#���n(����	O��(�f��l>�>���P��2����L'��sW��i�e�=�V�FkM���4��秱�+	a/�æw.�E���e����$�	.#*�u��.�b$�G���Яv��������)~K�Q�ÁV�Η��]�>Q�	��F�zP)�ղ*�D���^R���S21R����p�����"� x���!A�R���D:�`�5���c�R��p��O2�1��ym��#dmA8�k��>K�?��c+�� ,K��cve�G>�_<���$�v&���F�OJ��{�Ap�?�ZV�-\��u�9m����\@m��( O���]^��O��v��ĀFn	��fb��s�BS+	2�Um��>ʋ(fC�i�9K_ �Z��W��cD��~:aiN]�$d�xW5nٮҫ��k��m����L�V����!I� ��?�z�0�}Ct��1S!n̸G� 6�Y��Q�����^E����$W��y2l"b�)��&����`|�h5v���G/�G{a��m��N��d8R�.�S�@��MZ~�r��+��T���c��R�pG����)ՆD�s1XW��~�ƴݍ�Ζ����CZ�A6m��Y���T�9��>�$����29}L^��8R}*ؾs��`�0jZ�03{8��g�@��
S��/0��(��y�8��O�UR�E1��3�����M0��N�Y���_�-n�qR�M�o�3-���8o"��Cw>�A����\XB���@J�J����`�)���y&:���wD���в/SQ��C�TC^HQw�Q0�B�,Ru��Rz����r�T�2T�a��.w@&R���/�������n6��H8�W���^�*VɄ�?����B�(��>��.C¹���	"5 ׮�3N1�HdT��y�V���9h����e��s4�I$&#2��0@1n�ۛ�#iD�Ja���_i·��Uq�ԛ�'�D���K�)4 %Gɿ��|� �����{����O<s�jĒA���&��J����"+�����߱s��q���y,���q)��g�'��3++�����?7�:��z���H�}�Fk���N#��{�G�t�>��ť M���ZK�e� z�_��2���0�RF�f8	铢 kO�~?M�,����Fę�%���\@#�c�������ft,���n����쾆�J����I��|Z=��"F;f���� ��ڎ�_��M��Bv���eɆډ��x����p4�0�6x{.�̦Y~���)���y��{z���7�~��i���5�d]����q�
�/]�۩4N���Z��I)$�h��r�C�4X|]c��X�����H�	h��Nu&��Q���{E|yBO�OÀ��^� /[ ��SKR`Q.D�����{8/D���}�?=jS��� f=l�`�[�3��M�ɶoA�I�ʊ� ��>7j���/�'�2��+�P�34
ڡ�Ԛ ����QQ/J�>���e#,}�ZKy���<��
�[0���!�(:���v��u���D4��4|���OpEt�_2=����n$�}����e�������j�Ѡ?����Xյl/ju�շ��:�B��aJ�0u�A�!�S���z�.���'F&A��Q�>}f#���a��ֶ�\� Cսٰ�=]�Tx�̓����Mn��:�K�)=c�ķ9_�{�+����5�(&�q�p1WM������G������b�w den��5) ��FOZ�j1�~U6H�9��4�_�{>�����&ˠ�$x6o���8}9ej%g��4���1���`��y�칥r/(��\a�65sr)��S�UYۭ�g��Ү����[���Q�b�:��������L�mY
�hw��Y[���))����a�3��\O\۴�e����1�67�'��1}��:v�#~܋O�n��1zYD������9����ް�����?�`�	t��Ã�~��t�t�Nv\�P�w��t\!����XC��]��FD��4Y�f�0_��Ê��o��wK:#��|���P�]�{��?b�1�6�bA�n����@d�����ޕGW4���T}��j~�ZbD��C����/J$ �5����0�R��DiC(���¬�!�����Ѭt(B��Ґ;��#6*x0�).B��SD��$P�+�!�v^)���ZΣ��������}(�&�������zCx�B��n@����*��;״���;*�Ԑ>�s�\e�f�-±l!	V{�[���<��t�Xa<��,����Mږ�b�_hd70�+u��(פ�˻����I�g�����"
�£fl���'0�? ��:�dh:��( ��օ��NʑpI����[��]A�n�N��w���jD��ys�u����O��9P�4vePށ���̎#DACǰ�"�����Dm6�w/P7���>[��{ j��>�^�dlU�pӘ:M4�m�.��o�
+�h��c�k �׵# B\������q�V�@� �c�a�pW�PY#�͉7�=N��
�TЇ?���Hc��E����8�	��0��G�P�=�i�k�	���|�a9����I94��������6|�B�-�^K	���]!�^<����ե��զX���u^��/�Y-��\�)@�%_�P��љg)�Xo�"�Qʎp�A�kײЎ�|U�Uo��y�圠��Fw�)�ܿ�(MPZ�3����9�h�m�A�",��Y���)!��6�h���[���C,�N� ���h{g�M}ql0ηй�F<#ǑV]�l�F����l�~��$ z���C�\�;�'˛8��H$��ܣ���F�#d�27	j_��`��t�q����<��	�7��}Ƣ��#�Xے}�x��a�Y�t����- j��P�
/�dD�fҒ,`�Y-�z
���i9�����s7|���Z��?������.��Ц@��	�vB�7��E�������*�Z���9��
d���N��ĕ!A3��I�.H*��� ���:l��@!�HoP��Zf��˩�K0#�L����ڡ~ݴ�#U�G��l8��W�X�*�*f�}g'����>�����R}�<�.B����Sy�%�C=d֐j*�vд䶶����"�j��0��tCoHԼv��d��t?�D�p����XE(>0p�\�m��XE ��Q�]3�eS~L��)�!�K>�HE��z5���~�h��K{��<t��H������h�l1 e�,	?�@b�⍋�P��Z�U���'��Q�gW��Y�>"�_h��vڱ[�Tsa���d�l?�i3�EU�+��9�՘�?�b*צʲxDD�ћ�Q���u�vT������ �T[v�J��!�\Dz�0�$���0)l�
7�ζ��*[X�s1����D�4ImpR���0y�46�K=U��ٚ[��9`�T@�.��u�P���X�<OW����x%�3��oh��/��-��F{:u�s�s}'%0G��/G��c���g�k�B�rA�E5eX�Mŕ�mΆ���-55�q�Ol���@��,��a�G/4�'u���2�~O��%?���[��O���Í�[�$`�R2�a�h�AT˾?&1*��*��(d�&��G0D�]J�}�� ����	��� �=��<���;֩i�y�Ot�Jk̗<CeG�~�B��s춼�����&�[��`��6k�C�K��Fc������Y�Ƚ!X^�e�} ��u�:r#�؀q��"ÈP�%U����O�"k\�+�d�[N�^X�?����&n�Cֻ��o2�{fkU�9Σ���R�����,��@$�w���!��A>sJDg�}�}�����ifPh�� n��5�9U��.�m�H��ưa�,�y+>�p�o�_��e���a�*�Ÿt�v�!ta*���s5o;��H:ͺ'}�&cYJ�u@��1O#���������a6;�3C ���?A���#�+�����)Ɵ�ڙ�\������{3�(��ϝ��M�qV�12��hf���X�Sh��jk~Qcx~+AlX��t�&�1�h�U����T�yx[��=P�"_+g��w):�o� ���/3Ύt|LK��2�J0�?���T}p���!�͗���>/��k��Y�/(�D���-\���0.���NڹĿ����?�\�.�Ss��+�D��QR���^����?��w�-�^_ �7�B?�S>QxT� 5�7�x_`�\# �Q�Cڗz�i���
���]qs��l��^�@���PK��Mb7�3�F��%�i;�s��Ҫ�&f�������G�Y�q�B��U��T❋\�Z�Pg�m
&T�>%�Ld�!����%�w�C��XT� �UN�?'�3�M�i����9�1��}�}�c��ƞ �|f�l�U��1�T/�b�<N�����'=BWB�{ʓs�rSd�Ԣ0��QDz�LH�pA�2�q�"�BJ�kC(�9U)(�k��
f�B���s�R
C.�q�bm����Fm[��Ձ��Vtu�sZz��͎ JNwej!�"!����[k�byjˍF&E1���I�Q��x��p�H�� @Q�5�����5N���=�f@����� ��
̜|�QgF�TH!����.RuE�T�7�C4�c�|ʈ�)�Y@	'It�~�4޿5R��TbR���7�=c�;�ܧ)�U�������)���'�k��6@��I]4x����3DB1͌� ��ǾUP�4�0��{M�hJ�F��׺]{�����k��C� �g5�r�_S��E3W���`��!�Z��LT�ԗ ;����:��J$Zu`�C�64=XUi���1Elc2�>l@IX��XL@=2td�Wj'�������'�V#��.��O*a8R����ڣ|]���]��-��Q�mV���=�E�o���-TBB�T.7���d8I�d����yYkz:Z��S3$���-�1��ҞTI;��'j}�k\!]ӽ��@��H��&�!��W�}nK�*�+[�S��$���V\�UDZ�W������	���@�I~��
9�T";���P���`�o�@�U+���!4��+�y]�=fg����A��~L4�!��-��1�⩢{��U���t S�]��֤�	x�7�ܨ�/ם* �镭brrcׁ�!��.M[r��?x�����n�?���5	P�jȰ0i�Y+�ݗxʙA7�X�/M!� �W �� ��o!�D(�R**PG��0=���gx�.��2	%9*]ϋ�]/�!������a��H�{��<�>��>��	eͿ�,&������ ��n�C�b�;s��z��'HZ���Vثi�K������}{���)��ޤ�]Sb���6{���bCo��=�R��.N��/\v�m�����J�nN)�뻦�Cc�� �̠Mp���H�j�7 T��o{t@�˖�,����[�3��������()�ښ��nh���Wg|KqX��A����}��Lp$��6^Dy[��鰤�Va�x����yE@h7��I) �o1!0�}�f# �P3�� HI�|��!vS���L5�<��<4��|T���I�/"͕���Ǥ�z>me�)>C��ָ_	�
 �0�`��"&3GCxGC�a+kGNrp���G�$��/�����F+�ʨݔ �ʺ���JAӆ�?�6��j�� e�g}"��!��)b! nRްC��|"6⾀M���ǌ�ɝ��X�W�0bO쒢��I�˙��� 8��IY�>���P��9�urZ0cm�`��Lhx�Z�R�6�%���V�ۍ���]]K!�LB=��#3r�c��U����&���W�.~���!L��j2�W�n��.����*\5�F=�/��6�DEl51�@�K.�1]Q���L��)��1�b�U��u1.m�y՘Z�Y�����<i([Q ������	��a8���)�/��	�|���n7̞�X�3_���=rG��I��C�u�q��b�9a�%���qHl��������S���M�Z��}%o��L�/�f����CB#fG{���©>��^e@,eǟ� U�� ��I�6���Oi4*���Uh��������+zܤ;I��!�Gю$*�h��Ba��R�`�i��tnxX�(�W�H�����$�D_�}{I�ْ.��@_9��@��癛o�Qk��a�No��\���]�Fǘ�^�)��!3ތC;��������1G��-$�Z�|�����Ҏ��q���F�k��L;G��gaӐ at�e�O~Ht)aΪzN;�0�#�V@H`��׷u� W����;m+ej���/yJ�>4�3_pW�Tv@�L!�Կu�,���\�Ȏ�32j��3�1�i�X�!���`���QD@����M�PIYcAA�-�]��!���MA�j���K��[�bVt���3�O��B�Sn���m-?J���6x����s|�s�@G^��Ϻ?|zh/��6ã��n�4��&��zr=zӴ��B;�/�`�ل봚P�i���A�_h`�?��Vd�k�8�N�Q�g��VfQ�z����1�~�Ҝ����5�戁N{1�Q4Ɔ�SiI�p���#h�\�wr,	7��#k���;	�ek�Qӑ�旕�}�ql��ƣF�����Z�W}��/U�Y7 K&Cի9��?�K*H���qk���Vڬ��S�(��0�+ӑ����/Ƀ&��ݿ�NA�^z���m�%�8&2󈑚�v����Ww �&k�A-��L%���.��7��U-�q��;��}�(X䋀�E_��>�Ʀ�t���hsOK�D�<$�����;�	@�a�z�+k,(vZ
�mA���W��uF�ڰ�+�@�פޜ���7d�y����ho������%:�Y9#K���xL�� �Q��&��SͣگTk2(Q��O8���X�I�m�)ܼ�&r+M*���Եa<��V�/:O��[��^M�1�X�r`��~m��"���>�����&"O�Ȓ��9{�i�7N�u��ܦ��ͬ
56=����c�EejkCy�Z�����N0���f0����w����^)�#���҈B���󊒳1d�Gu���t'm�[��jf���Y<�ׄ��x�F{de`<c'�����M#23�)m+�l�S���dCy��r�t�y�ʌ�������H�Pı�T���k���>��)����y��Ir����Ί��3�C/����6�X-��Df�H��d�� PW�������|҂:��j�
�8����a�����%�؝D=�b ):�W��h�fp���s#�`x�}�$23�H̺�%��[��G�P����3�b�̛������e��7�H1l�co�Ҟλ��d�Z��~xy�:����J��+a�[V:��d>>q�+�:3ޛ�M�B������s����J#]��fe �E�s���ٞ�����������dI�at�_Vg��09 �SF�����ɆW�K�^�`�Br�k�������@��F�H�"���en�K�7��#��F������N�'���_�Ax���`j~�r^�#)ꫢ��/�/����:Y��y	''��b�b�P9�����œ�Dd,g�Fv,f��h/������m�[�B���
�`��� ۿ^<��{r�3[��C��28�+�G5�J�3�`'J��iB@c�z����fe���c�T��}r�%��į�2dJѥ�v��h�� V�$��0���/ �)�3]�V�}A��o!������H���o��d2Q��{���F��Z�g�Րb�h��92���⃠o�k���~���*p�6N�'��������c?H�R2m�sV� r�	|WV�l���Z���p��y !�Ѻ�d�ǐż���*O���{}�@<���ڪp�G�74|V�h6�z�u�<�!,�j�&!|t�}h��OI�n���ȸZw:%��&���Q�Z�Ը��⛂PI6�a1V��]T�{�I���'\4��0bu��=�sn�<ŏ;V_���L�e��(��(7a8[UI��Z�c��.��y�a�&��
����W�s�,4M�{۪4�$d�wl�̜����M��ck&w;��I9Z���׹�����Q�k
��w B�zI�����ug4(RV\MmTܴ̫>����аH�|� ����Ƕ�Ƿ�kۭ7e�d�@2��=�F_ؔ#y��W,Bi=p�	��A���Q	��ČNJ)q��i���T4��Z�$���]JkV�zy�.�ax�z�N���#C���6D����y��7�Q�����̳Jٕcynb�ƃ�O�=,��.��ߒ*� 2��+-�xyW��%Y���#K������W�����a�}�-���i{cT��i�v{E��r^#]��mn��@肧-���|Mg�ګ	�Z@�u5�}rN�Ɏ+I����o�L1; �@v\@�w�*�Ojm��5�!�8�M�Խ ��RWGH�u�ĥ��/��<^x�4g�e&��p��_4�p�� ��>ر��T9�<���m6't��[��x<!��}���eYW Ͳ���X��H�����{�^��-x���ymv��%��q5+����7<���]�p`Y���V�"Pr�6�ح_)�s��M3)�A'�)�K�.��8f�k$kiY8�Rz��Y+]�O��YԯG�v�50[4��G]����xK���~��}&J����m�+��D�&y��XHf��������`bczh|F�x��Q���+l65L�IT0ٹlFt%����]�=�O�q���>�Q�S�eK���O>���w���n��;/z�rd�}���/������	6�&��G��'"u����M�"@+K���,_	�~8��ﺟ"W�hĪ���_V�Y{��Qm�M��`��s�L��+����鑇�gI�@e-x�-U�
��p��B�c�`���
y\��Њo�ͨ	5����X�ޏ��
���kˁ����:0lI:��4A3���םI�?������zMK�����:��-�区Qn̲�tF����!r5j2 �&Ց���T`*}��YaM0Ԅ3���Z1�iR�[�82,�r%`Zd��̋Kc1`3������ږhM��gE�W�_
kCP�n,�&���u���3i��ǵ�}�BC����e*:iPtRW;;�;X�=>�׹ԩ��iㆭ�-�Y���T��@[�.���8���$ִXX0m��z� ��5�,7܉&t�������$;x��=\Ql�����Ķ�?ReX�%(��#�^D�ȿ�=q&Ǌ����F_[Azl&'��: ������#�:��p
�&�qظ7��Ok��f3�`!n0@���x� �sp�\ߪ�uM��p��~�rT�=p&Ț�^-lE94�$��5���8�D���F�10#���O����1UI	z[ٜ��\��jk�Y�u&�aV}GJk�,e;�r�*��$z}��|���ݷ"�E�?�'X��� �(��gK����QE[�Qxs�h��5�bE�G)��rN�E���*�Gթ�A���,�jJvn��x�J8@�h�1��yβ�8cB���)�5n�C.������x�
|��gNli�,�p)`�V��8��j�|M��^��m�f�R�a$+�Ĕ0��ҥ=������.*xu��M}��(���LF
��-��P3�3�E~��\�Eԙ�ytr)}իҌCmʄ�p��XF�>j�fnB����_I;���D 15_�?i弋uм&����
���Mcﶁ��M���C�7`��˘���]<UW� 3�.P@Wm��iGYm,���R"k�<�1S�/�P��5 |�(Bhd�PY�i���5�K7;o��5��14⧒$����n�Д}�Z���>:f�C�q����>Bߟ���򚈮@y%�G�Z�xP�=�Kt�i%��s�������>��gӗG�Mh3Bj�:�F���(%��QK�4o~z���\����v�