��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|݅o�@
�nI�֛TU�PP.�����+���u�Jf]�ϫ(#��$�r�jO!�Q%y����m����T}�R4�?/䃭0����AU�(�ƾe��������f�7�m��v����of� 6�{�
N�m�H2
��j�Y�?�:�@��;�b?�f��^�����M�f(p}��&~!���i�W�/��>�d�(�j�2r�L���QEl�	�зJ���MBj?�e�տ7����d�JK�
�!�M��Tt<:<���SHT-D�	��z����X#�sY�$p`A�q���li��+���g~r$���Ikj��|��
��Q�1��>�Y�����J��u��ի�gU���	���>�D�����&�d��͒�v���*A�tG*����/X�USQ+;I���ʊ6���%�D7�9�
��0��>g�z���	�\���~���A�(�{�R�{�a���oh{���u=3�� ��ai�������H�"`&��2�G��/�!��]CKZ����S�X/��lHU�s?��|eZ�����7��o���m��(�v���o�d��,+��i'ڱ.�{"'mu{�nɡǼU�
����W�?���N�\�{A������ɢ�����lt-`#x�ȽGT�=EE�zv��fi.�tK�~Չ�]�t!��؁�3آ"b��VR��������������BCc��H�p�[�B��8�U!.lv�%^���{?�I�6!��ar�j}(2���ˣr�>C�c����-�Y��H+.���\$�����S��������:�O���	@��`)6�_FF�d8���1�J�fBU���0ǃnj}p�g�����@�I?-��� ��*E���"�+5{6�"u!��F9�(R�`��� �MU�e��Yq
��jn���#H�j����hyk�Ieʯ��F��Tǵ��RO��@�p(E\�G@���>O��mPЏZ-�v�m�`A�q�!��v%6{�a��z4$,S~:N�1w����mtpˤ�{4�S���Ji�p�����_�_\vH�U����؟����K�,I���*�Nh�~]3��*��!n�F4�A2���H*$ִ
&�I��з_�6���)8�_��ǂNH4���p�a�s��q��I4tM3��a-���*�J#_w�_�B�3���$�D�;<��?MԺ׏8���Ta�sc���h�P��(���7T���כ�
�k�"~�[)6N�|?��̂@��_��ɦf���dL�"�D���4�|��W��J�l� ��|���#8�i6b$��N�7��0��'���4�O/��j��w��n؅<�iȹ���B d�`���R����(��bᣐ��AH��b�ڴ1+zJ���R6j���5��>��F*�Y5Ξ���ף���(����v�ju��ͥဠ��e�)�@��P�s�ϐ.g)8���S}���P�aU����"��&b��49�vmX�W���LQE��k5��錌̢�O�]7���$kZ��}����z�Z �c�� ]�����}�%���CI#w�2�r^�_Z���8�un��S�y�3��/9�ѹ2	���?4�^e��x(�?�K����6VL�P�Q�5�ŝ�n�B��W"�9W�4�݄{�ۆ�b�W��n��P�q��� Z��h����7F���*�x��,x8xt���l8�sH4M����]ʡ�i'^�� 9�*�Du�����b�'�]�����a�(���&oK�rA��Q%@�D�X]�D	� ��:zʽn��)�|a}fQrZ��5��5��r�{�PC��HNma!M�	X0��/��{���?B�Z�o��#��5�HU�������2�>tZp��\	�b��X��3/r�E�1����\S}5R�ת��0XQE ^�eV
:@ S�>���g�0�TI����Ź�����|���j_�ەlgA��
ǡ��X% �.{{�����6D�C�*�*2�T���ۇ�sB]�wv�x!���ը���e���r���5^�mXx�����?�� E>�K���z��~#Z���&%��->jn��Cz �۱��z����n��y��3��ٷ*�*���ѣu|� �K~���N��h����*�<j�,OJt3�Dhw�Z�~�~��-wj���(b'w�7�������X�*7�����>j8y���v��P2+j�' ����0_8H4~�|����F�ܭ=~�%�tn^_0N<�2���\�ģ
�!�d\���|OX%�v���È���|�i#%ݽ���|U%�Q����@�_��|w-�g�S�sx�τ������^p��%㟝is���pq,M��1!H��KdAM H9
�ǖ���[�Q=?K�"��x�u���tcS�|�[����>��4�gm���~wp��|���Mу�܁F#a�g`�?1kN(�p�ꝝ�q��	�F3�Hd�����a���y�\��Q�h�����I��=�N�k:-�l��,� -"��ơZ	��d����gޔ���S��ie8b����Y��n�'�f?�:b7��ZH/ȓA��mG�y=JK��8;S���?A/�kȠ��b��Jxg��ȵ�e~p�-���h��|��x-��(�%TW=p�r���	1��[3��c��vﴼ4�=��-L{�����)����j�;p;�,�b.�w�i}�E�� ��6y`�૯k�z8��"ד__���7�6r�}��Ǉva������vAc���/0�@U��h�*��xˇiCԃi]�J�9������֗(-��B�m��T�����P�,�/ޝ<��Q����"o�[	�!����q_���νv��1����г$�?CG�Q�c�JFp�J@NL����i�zk��P��0��������ce���-J���Ί����"_[��^W_�0��jc��P�ǧA��[W^�GM�Vc;(��_�f���y��5ᵜ�h?��+���F|�����Z����>��(f�����-B�x;ז�]�=E�1���=0�����V��Pө�o��&�����4$ef����7��۳�d�3s����)�jH��)���n�bì���&�&BE�ٽؤ;���2):?\��+�Z��o� ��h�C�W�ߡ�|c_[x����Y���1-�����I��D7�f�乬6 ��a��r/'���Y�0TB�?�o~�*�R6�d|�O�| �"i�%�8����M��Ӛ0\��D��&y��������#���1��+����U5lw�-�.(����`��_l"�e]��9�n��{�H�@B>Ϟ�|v���׎�&�����k�{�x�������&�1uS�F��ZsF8��X�9�)�.���ފ�lg�[��d�4�ɸ�.%ҼX���`u�N�t�[&�Đ_���VFX�C[\�KW,��w��P��!u,�Y� ��͛d6{��&� F�66�#�*�1o\�Z���UR�R��=Ȩ�Ӭ�n�����P�����Na��Ǵ�8�cK]��UO0�ozB�v��4�:r�O���	���2�߱��'�\���ڲ$b2����Qu��*=�_�{.�!��8Dc\�V�;57:(��`�������5�=?m+����~�2��f*I<��}䃝�!eש@�oc�U�/�O�Հ����pdE�Seo�{ �COcs��c8�3���lF��Q@1_�UA������b�(�F-~��Z-@�g< &��w')K��%����,�y���=]��H�ߑT� �y�iZb"˶�xf5��~F;�h+` 2�1�o�#��_1�l+v�xU��!Z�E�*Y�^n\TE-�t"��
c�F�h�Jj?ϫ�b�}� L�ꈜ}��n^
�[%`l~�55y*�����#�`Z� �l�J݂�����":��O�(��:^%fe�l��oO(�8z�a[��ђm0��,щ��ǃ
��*������Fc|@k���gǮg:O�DO�\r<;4�n��u�SEӍBk��6�m,� ��٣`[�i��1����`�I�ʝ��l��H3�
�+�֧5K�$���&��'�#����(T�����n��Kw���U���yQ !�+�&K��VӍt�ؗ����G�x�r�-P�^��9w\!�%.�Ϧ�PI����ҳ��ǫ
nF�=*�i�d�b�0����$��~P���x�����hǰ��]s]��Bl�U���8,�x_��;�+�3- ¾&�w�5���ѯq0�I�$�6MBF��ʙ>��W���A���8��	,���Ph��{\��$��;�X�n����S0�秓ֶ� ����;֕��_S�*v۴[E��VB���8�%2�E��LW���*��i��]	������ހp7�Nνv��xQ1Ԩw� qG�����s�������|��v7��1͟3��w;�-���O�zU2�JV|	v����M�h^�q�p�HX[�ʼ��Ĵ,sp��"q�Y��a�;�8Y2�S��$�"�͙�BhḈ��A�{�B_2�n����?�־���E��6N;��Q(�P��&��3n��d�]��暠��O�],��= W[��PW��W�K�V����sH�@a��'�pg��x>�>���t]�'�zL�O���e��A�u7-�!Pxa��pu���۹r�2�$�^{�y��hh
7�bv#�:�T#�nna����=(d�A �bD�������W�]��2���i�-��M.��6~��+'t��X��y'���L*����yw��P��O[ߺ�T�;��H�3oyV�[W7�+�,r����B��O�'�4�G��Al��Y#�E�a�	�����o��ZJ�il<����!�]a<uY+�FNB���L(��ڤ�N5<�K������9ݟe	����+
l�~;�^0�`p�ę.[ά�f�Nr�%�WB�i�>y���X��e�E�E���$F��PTq͡�b���*�o��-b:E�s�����aF�"��6=xt���M&���ȷ�^����F��ж��-V
�/4w����TBU�D������9]���<����t2I��{��U&�\�yV����In���踇�?ba�ݴ e�Jp��ك��Y.4�JB�,9�R�e%&�b�l��i��m���"���⡰߇X����[�g��:GZ7���h��4��o�l���.��z�cR`v���I�cJk���}R]��h��D��gg�bU�9]����@uh[���Z��0,�t ����Px\�l��z���
�pw���"�iĿ��՛���E_KfxK~�r��~J��^�(��_c�d��k�^��`�.��7E]eP��aӀ�����)�T�u�)�hǑ�4
=�������,������Z{Z�L5dzJ�U��3ת����/[���"�]�&����s��/�Fn��޸dР�����e'{�ުQ��=��:���S�I�i?��V�Γ�	u)2�m��!��V�cSh ���j��?�n}�J'�$Ɏ������	v>����#��fH88��f�_!��,�#0N��##J�x}��U��_n�C��L�0˔�5?�&����)�ԫ�hW9�$)p𬘙t���BGn���
���6>�'�e�@�3I�Q@� �HG6X6�`� ��`��3�<��t"N/�I����zQ��9��{Y�]:�t��߹���%	MbnoJ�^Zf-�Sn1Y6?d����� �>��G�굶�pC[�	��ı�r|��ǹi+a���M�&�atҏ�1Z%o�`
�ķn�]����$�K�PB��
&E���=�9(�P[���˒H��ͯ^;�G{�o�F���U�q(��Z�EK?���yH�a��Dm�#��*�9M�xd��U�Q^���}	Mj�`�0��o����%d�g�:qTWV���a�	�C�f$T:���TQ_ ��g/�9:�GHl��(i�o����믉�-���*a�dd��c��xxL�K��Ů"E1�<��1褸�V�'�"urf?���#���V1N(�n�׊�r:���
�G_k_�iNX����.쓥��)Idm),����	��s�O}�3K>iaL����$��_~���D"p>�䏜W��������~�Z�j�$���� ��7�o���v�"/{�g������(�����+�. ��-�	����R6��=��~�Wb��d��f�vV��b��:cL��i�Qy]>l��i����>(�CA(��EIV�I8f�,߮G3�R�1�Ԗ^�|��ٷ<���W���[TV���&�/%dw��B�J?Y���wf��?�� �ԥ��!]��9�?*[I��"$T�j��!�_M���^�_CD�ם��T":�7�c_��2GNLX�K#����x��?�kʶ��ӻ�7V4[�a�Ɯ!��iE
���9�q��B4V�JY���J�[��c��L�B�S����?O{�Q�x���K�<�Ӧi������Қ��Ϙ6_о�#����W(��~�W�h�4���)^�z`MK!���H�R*��9���u�ew����ڇߛ����
�
>%=��ڿ���a��W_;� �܋*��e���)T4���Ҽ��L��;��'�*4�`1�
��*�=۪�·đ���Wg��h��7o�+x'��J�Ws��:7���J�3��69(%�x�����'D�עlO��U��y1מ+����ϷܡE^��#�f2jn���,��XbIWKXX�����C�r[�*���hl8��O����DҘ�&4]�|�z����8l�3���4͏�#���}$��l)����8�H�w�R������>�.+��&y����h7tR,"�@(����Wp��y>6n������ �qd�%:RꂧtU4��@����|Ƀ�?vϴT-Z c0os��T����X�T�dD���Z L}��D9�iM���/��'?���f�#E�J��%�
a7���ֆ��$o���U���/�Kzc�8W���C�l��,��-㶄�U��U��K0(��C,��4���\_y��C���uS��=�\�-"���X�h8�x�iH{cn���.��
�͈��ͨLe���0��Y"��x��(��ϗ\Z=z��z�[��{&\�a�*.�>n�ge0u��h (h2��v����<�F�8R�r�L�\�%L2�S
Lj�H;cʸ�}�/˨i<ڮ�:�Wy>)��(ǲ!�U�����R��h�إ�c� �)��Gb��c�TQ�ڮno����^v���
KA���Ft�ٽ���7�����j���"A�� #���U��Q?�y�*a}I>u�ƞ̰�,����xY[�M����˕c�ʹ=U��s�M�jR5J����qț�x�FY/:�3.���q�|�ht���s��R���ɟ`��3
2��*:�Z�$��aP���n��B�B�+��	[Y~����(8h�v�o����zӾ���e4��*��g��-w]3����S�. �ݰ�&��~u/j����Oi_\�I�vِ�H~e���R�-����E��M��%����{����x&,㓞�����xE�D �6���X��	+���3���la6���A鱞>\.҇?"K�X��z���=We�w
y�c<13�����V��� ��*YO��2�� ��J�X�_x!gW��۞��)�|����u/��H�-e�}�x�=+�\uλ���@�F$��7V�G�������~���	�v� �L;ǫ����J��t�T���i����� o�z�^O2����U'�[As���о��@0}6 E�����~j�w��'�>װ���Y+��s�aT3�I�ѻbwq)�CK�^6K�A�� �`i��ӈ��Z2ܲ��7'�b�Ζa6j�C�Ugt�"����T��?�3*)�'��n�-B&,��r��+���NְaO�����%���k�p�I��G�b�'�9fp��<�6�p�_��/� 9&���<���$���g�kVrhX��T��%�&)Ǆk���r�_�\bY6�r��6��5�D26��W�Ur�
˕�1P�#���f׳g��0����V���pK~[;��V�P�>f/�Z�"���{��ԏ�T3�c#��t<-��2�I���޸�^U��ǯt;�B�5�ׯͻ'>��\m��G���)�a�7*�n����~�io{B0�{r�v���3��"�fJ��t)�u��r��ܖoZ�P�ඇ3�������U�j�^�%�[�>	�.�)�b����5e�)��]����"~�p��ӫ�.�QV�[7�_.d4A�5��3��i V(�Ά��Ӓ�P~�h�B�� ��w]�>������;J�8��t���ݼ��!G��@��ط�
r]�@���0w�Z_;v ��ɓA O�Ӧ����IU>Ѷ���M���ڀ�#b���b��
�#��1�?���]a	��CW�M�+��Z�^[�$�J����G�g��N�=�����S+�}��q�$��i9>���$c6���m�0l���1oO��� �R��%���_�4?���x [$|]�
5ѵz�o/аC8N��s��_+1����%�o�`�X�*7�i��d �C��^�rd��|�:�5:d^My��ҍd\00������r�r�F�k�/�YAs]��FIi-�t_C�~�g���Vq�+:�%��\��:޷n�b������$����'���b,��Z�����;	S�}�0x+ǐ=�bmH&R���ũf��҉��T|5ϱ7�ˏ�bF»Y�Æ�����W�u���#���,�@ӡ��_0p��w[d,_b��ES18Ǘ�%ͫ�" ��W1O������M��18�N�X?���[Z��8�w
�XhN�$����g%<LIu�`�swu���q��+�lp7��6dj<���d-���u(;�l!�����B��a̪�?�s6��9�.*�X��:�'�����)�lU'Q����R��Kŝq���c� �9C���m�i���E
�v�s�q��qb��ɥ\�8��vt���	��xC[��|D�������c�P��~�0�:W~��xJ��0����{�CRD���50�qb����nn�O�-����#=M�:����[����}���b]�6�۷ݑ���\�Y2���=r���Z��k�G���`�x`�H�? �0m������k��n�=VP�(p�
E
R΁xh�7z���/ ����\B���æ���(d��bP��˲_�6I��	>�G��+�$���n�zO&O�?�H�Z��e��`5��� �T�(R�1;���=����ְ�X�\���7֪$��uL}���D���8�Q��Ζe�Yq�}5�&�hB�H����d�R�y�u Ұ��@�蝓��4�7Mo�?�0��Z;����u�@���sā-�?�[�
�k�֕���N`R�����Ƣ
y�wOP�:�'�A;��y��|Мm[��&�H|TC�wR�W5Ö1.;Z&�e�D#����M�e�\�7�����g�N�=~\�����&E�@�m��U�N��{��͒
�%4�3�~a�m+v"�+x:�n"_�n����J�� N�󯢆s�P>�Z]�H�\�)�'�m��"d'p*C����T������D�	�.#zgo,� ����m�ɼm�(~Y���T�42�@��:�E�m��b��� /��>�v�jX��@�W���=�9K�ZIl��j<>���N5H�9�~У-&m����E�$�жQ���VF�O7���VN%�W*��AD}�>'+��ú�����B-��6>$D��C�Aw�(�~�D��*4��0�q��� ��!K'�s͖�bЊ�d�0���>S��=��}xuݤ����z�SSy5�K�_��V�fJo/Wt'�ؚN�oV��е$���F�U*��1��}�;��d�GѼ���ׂfr����I�!�m,ўԸ�h���r����ÇM|����+5�0�����`9��$���[p�*N�'�>Mj����͠�v��&�Og�dE��wWU��eA�[���_�+ �1EhW�C������ͪ�po��V/��fBB׳7ωѼl�sяs{V��]_L�7�D7Ϙ�ʳ|�j���N�;�n��i�/
�U�G��
��5Z�v�=~1�?Ie�,�e�&f_qƉp�C(����I��/=Q�NEz�9k��L9��rO�qC6!(l�Q�j�C�`y|�<&\W]"F��0|�.~p�j� 0"υ������`kh� ���f���d�~	�	m�e�� $"-�rGJ��}H��$,P���ьN���1P�����z�ݸ�H\6�C,b�$1;��*��u?L\Hz�*���7��hej�pd��ܵw&YXv���a+���)���e�S�j�f�VcF`F���X�&���؇Z�mY�+�D��d<gɲ���&=�\ނ7���N|��\�%S}�W�TD���I��O�+r��/?U�����[�������zԬ���R���⒣�k��­'m�1�����
��`S��V|��s9C�p�U�d�b�(�@9���R��=\D�TLxRl�DE������tg������S�W.}c=���P6.6���t�bpZ��cK�3�7(Ls�u��*��d��\r��Oڋw~�ǘ�+י��c���o��Fc�d)��m�4��n�wj���T ��J�dTx�dE���ۦ�~Pz�GD�G����p��Ճܚm�$h1��3J�z���Z&vd�j�e_�(�}�6Rŕ��?[(�ߡP���YnbW.Sus�ӵɭ��w�J�<�Z#��h�L����hkG���� =K7����9*,�]ts���r] |ɑ[_sIW��(�R2����ێ]�s J���*�^F��AQV9!�A�/��,8�
2���0��.!��R?�p�� �n�*�)�ҫN��'��|R{�Ɇ(JT|Y��=b����ŉ�y:sҲs�����(�F����"�J���cA�$��\��bS������s�!��jPOa�����Y?P�it����F$�qTk�(��Y�]������*�,� `e�R9OU��L��`a���FZ_�ě��6D��+f�$�3ʷ�ƛu���ͼ��6C���qi��~
 �� O:�C��;;�aX.GL�^o�>�1�@F4|8`��S�.�l/(�Q�qj����T�z��Hg��t/!d@���`N�4�e��|���|�RL'',����/ `�o�F�`iȟp�?�W���T�p:`�n1T���P�ъ���m� gp-�>�����V'2�_(b��q��j�Z$���˟*9}���(�TN�Oͯ��q�n�)(9m�j���c���6,�,�T�5�jM.Q}-EY&����0y�i�[��}D�&򤆔T"R%�\��q%�,���4�'�
D����F�m�$��O;8d�<!V�U��0 �Ko M�H�=��O��\$���%�EФ�[EP�n)�z	[���qke���,��O��7{i�H
��B4�Ԙh����W�1괋��ӯ����^�ެib|�*߽��L\'ԏ���5LV6���ܰ�U��?��Z�N��'�m��P��r��-E\Y�)�L���G]v)�����3'Ϯ�@H��N�.��{���(V~3>T�a�e/�_�(�>) ��'�E��bIj�am٣[>�pG�e��� �e�*;S.��=����rq���hL��"B���x��w�P��ع��������,�iE`!�/��wC�h��jEY��oů6��z�n��3�l�,V�1��>�S�No�Z1#`s'���g�0�mkO�4=A��U���@E��4�S��W�``���t޾��*��φN(��܇^��TWx�+���\���mk��~%��\�t6�H*h_[� d�V	��M��g���VW�� g��E2��1�R������CC^e���ΰ����M?&��D������7��W6 ��o�'�i��r���ܔtb��d������:���9�';�ņumn�o_'����X��t�-
+L�=ڎ��iLT��3,�Z��:�j&���N@#��]j��/|�a�?��������0���%Hi�Q���Z�A5�a�+b��
H$L"��A�rK�fb�I���<�x�jp��A]R��b�T̊1���Щnc�"u��K�1z+5��?��l����%9���?�1(y}��	�@\��`B����/#��� ��K޲�  Oz�V��F��2����_����zޤ�&���)��ʺ��a�R�Qph���C�ʀ������!��8b6� A��p@N���0U,�r;���O�%^k_�V�I�)��,�Gh_��q�wAf.��.4/d�q5v�waW�-��WߴXw����-�h��]`�:ݡQ�7������i8���W�N�u�܁�/���ϡO�7���Vg��mE/UR��y�z*e^�l���D �V':O)�5$��͝����d�c��ĭg�\��0�"b��^��uF��b�f�?C����Z��7�3�D!��nO�b����n]�;AJ{L��Q*O�5�J��]���#��Ɓf�h0�k@������d��1D�.qI�ՠ�<\�+�/���?��U*�.�")��[u��	������B����}y!}p����/#�+��XJx�߱���N|�����'�o�c�&}�1FDу[�~a���б�c:�R9��W���Kk�!��x��1�"�=7 ��G��q ��"��x��an]	E:�lPV�6ۓ�:a �16	�,�F@���ɄKϐ]�ԯe�������G#�A�n=Ht�ي�T|��*�/|d�����q%���֝���O9�ɤ��f��k�ƨ�[C,z����3Қ��,1@R�?>x0��*n�D��	"dR���~ra�k�r  d�t�u *0d���hv�Hz�֬2���+���%�=}f�l�48�*Qu�����ϬY�+�lx����q��7��J�٫�ީ���Sd�v���F��/q�Qܭ���}���q)���O����~��g�C$4cE���B�u���W�B�H�/�������t�]V��<���0����ܳ�aZ�Jzg *��ĤX���ފQ����e)� &f��^��u ���^#�z���dd�� ��s�_�n��q/�	����R���a���yv�_͚Bm���(\�[�S�}��>��NY��Br$��/2���>�i3@I}ͿUN��x�t1����:�&��۷�gX�g;hQ%�T�l\�ج�D)A�,�L-v1�/�e�
og�R���X)�p�E%�c�c���a��!�p�� f"K;�>�����"�.�a�ƥ8j%���wi�9�g��� A�by�{M'6p��m(�y��6�%�/3
�]
�\�t��È7�NX��qsOr�*��ߐ����[:Ր��gP���������V0	-�0b���,��@^���j
QD���i��~i�Mz	uY��-�;3�ș�g��5���pw,~��tԗކ�܌򬉶�l�@�	ot���[$��j@�D:t_����w�4tv1��A8ݯ7�(s�0��y�SW���&���Z�]��Jr�r�w��k�o���J�5�������(���z촭�eR��T5KW�ɬ�9�S6�7�hm�\)�5��fB��m�^p�4n+��6���Ӂ��9�7��p�����KR��h$9�}	b�V=
�̖���f�)��&��d3'������+*�����e0��ϧ!�)̞F&�˻�Ϲ}+�w�>�veW	Ҫ ��8���xU�5З�R�d�"\=n�����\qv�S�ٯ��z� �|�Ê�JJ��T�ۆ&������1	��*]7� �����-��]H��#4p��7�._`�dtMo�6�ث��b������O�wq��C>�j�Sz������$�Q�5�ٍ?&���Qb�����h�Z�J�����g��+!o�e� ���>�����C���%����!�&4BE�D��@����W���ǵ�a0ۣkB�L�F��VB,w]��jv� `l1�������%/Mv��à�rU�,���hl��oG,���F����"���m4x|*����18��#[�����X|��*�뵹Z=�oC���z\ƕ�9(��A�
�J��k��3L�?s��Y=�ԇ���>��Ybv�|r�Ȕ����p"���OӘ�K 8@���L �;�ȍ�ӕ�9Ў��b���馹���f ��@��a�=��O+y����-��0-��ʦ-e^W��6�i�kLJ�Q(isNO�Ua���\E0dsPN�{�Ӽ$�0	�i��D4>�XYM j�Qg��RO�@�x�6�pJ^��<�v��D!�K��+�;���jI��2Y�J��̱����إ�x�Rh�/���k�19��9C�eH����1)�z����^�G��ْ���;,.����}	��=��ה����F��`)�{ߊXG��t8��`�mg���P����m=p��\X۔�u���v���P��Ł����Se����JO|���j:��dDJ�E�As$�D��yP�T�gdh.�#f[�h��GD����E?�f������c�ۜ�m.A�����}W;�	��ܞav���/�q�Q�g��E�!SM������3�\t9�Nm?�gҿ�]��%��=���R��dOq?i)y>ą5�T�,��3����X��bL� �)����s4 ���9;�c�27pñvYÙ����]�*/�0v�5Q$E�J,�g��x Ob�ه���� �B�b�&�?T32 ,��>��E�d��a��a��U��\<�f���'+��84�F2���-}���YqYB�=u��k�e3p8 �E��N-�Өm�AA�'��G��N�&�"�p/=�R7|V����-Yʽ�jVkVf��X�G���:@IJV�cA׬���?"�o
��g/2x�=�2h����[�/0L����`<X�$敋��&��PD!���Z>g2Ьm�̝��sb�U���	�b3BD�����Ϥ���~�W��r�I���R��	����ɗ��n���|���i}��eK�*mC�}�����뼾�3�w����[�l��xm��^}=PK��b�JɸUl��$<��	�H��x&>z��Ɛ jlK�dMϩS ���cs���E������ɜy�p�y��AR��礪+���y�7?�+H���mu�w��	��(��EA��ɸ����}H��7��1��R�-�I��'c߄ž���/��/����P�j<����)�4M������N�i$CT�����nZ�F�A�C}��By��àRЁ���iCYů�����8s����u_#SR�_�]�-����Z��sO�Ո[���͝��Y����&5����X'������j����̐�_Չڻ,�;j�l������}^�B�X�C9�\1$^u���z��|0ŎLq��:��f��4Er��dߑľᢡ��Z��'�:�:ʬ:�r��:!)�啌�7�*U\|9�M�����iԥՇxg(K�]�P����N;�bi:;��u��U~5"�J�0�d�۩�M�%<��.+z�)�u��;���{������/�������E��Q�%Jk'��Կ�:���C�"!�)����K��%�&Zc*AvB/0̩T��T���@<y��M�jN�^U����X.X?���V\�?S��̽k�����𢡊�jZH���������%F�6����z]��>]\�����T��by�'7uձ��u:���~!g^�<>=��p�iOCN�&i���k�D�`��������Gnuq��	���aB�S��bpS�U�k���$j�@��ޱ�f� ��eY��M��r^E��5���X;��^4A���|_�2_��
 �x��[�֦M��m"�	�\��"[��)�e�\�sl�|o_|����UmH��w�Kl#��L��sm���b��4��T���te�=r��z�*ֽ�
���Ӊk��Y<�Ng���+O�Ó"_|���}o�P���`������㡤ŋfn]��C�����I��@|���]�أơ
�͌��|��+���-�ۘ N�E�8g�M��7�8�;��q?k�A���b/ح��Jn��������G^H�Vt����0K�M�Oe�5!O`�XM9��:?��j��
�ʏ�;%J}Ւ.�'��H��gÈ�n�U0�}��y��>�`�y�2� /yقU}#��v/�3�9f�hB�3���I����� �a�iRyŉD������:)&?׿9�rH���2� �;/"�X��
G׮F����\D���j��X�)��>��C���o���qn>75|~��&��<�J���4�6�:���~[@u���}�U�}��x�
�0[�B����Y	�¿O�F�� W�@��<T�Pl0�[�\I�����d��@��A�D���M*b���F���ɬK]���b2V�������G���4hN���P�.zF�f�7`�ӶwM��>��5_HԷ�B��U�n_�Mm݁��+��%>����V�$st_
��RG��p�Z����2��w�;5x�������qnh��r��G�oo��~l�z� |��,����=��@$�wKWj����ꃞ0��zd��]@%��Z)��jcvI����3|[����9Q+3��P�}�F�I�Y��osaz��ZШ����2�9X�"�v�la�G���4�H�I4������%'�ښ�B��E�D��Gl��ǗM��]�ZuJ�h��BE���}>}B����	$a���Ѿw+�B���b�ƾa'�J #=Ia)b� ġ_n�<.��,�˵��a]�:Kxv �����yś�s��E��N
�i'K:��M7���4S����F��|�e��$���_O��D�_�LS���Y���ŗVKk[̖���+�<v��L6�sL����_�|l]�WV�����Ri��-X�0����r��@��d{�� w���M�$����ѐB���c��Bd�^��fS�T�z��6b�9�����4���~`Q5ې�8�]q��׸E�`�m{u���N�%�� �������48�s�a&���$Г8��0�ۢ+0�cjrV�k���yPύ�
�mK�����Y4:e�^u���5���ı!�����p\���Q�mG�5�vU1��1tCJ�ܭ���<{_����q�+���Ȝ,���
��?��?��]�(h�e55i�@]���^�Q%�\�j���p�����e�
2�����l���G�o�S�6x�tz<���K¹gѵ&�4}��;��Ax����"�Ceg�ܖ�~1|/V�{|2�t;�h� ��2�y�X$�y[_+��.�[��ߚ�{�0��K�'`j��[b�sa��:))Y����@k��e��ȑ����F��&y�/����Z�
c}�������D��	�/7�2^vA��ޞɴ�9�r�N��:r���d�ϒ��5���J�
3����f�)����z7na>����Y�a<ֿ��	E�r@���)�Cu�5nχoh,	}5��l��x!�W0/��/�˹+���r5�SHЀX��Ǿݣz/�_"7���!����S��:A�3�����2h��]�y\G�B$�XWWߦ��p�x��k�R�>��'+M����"��@C����y�Id�#d�m�<�v��{���Χ.XUgK��7%�+�皃���ֺma�����j����po�ӌ��DU�Bbz�禋r@b*f~���8[,[16�(78b�B�ֵ�H!eG!����Hq)ƮR���u����x�9L�WLY�Ӑ7#Ȩ�����0��P'�!��|?%���]Q�˲�LR��/�
�A���2�z��1���bD�^�	4_4$����IiCZ��{�2���ؘ!��S'�ޚm<��k���#3\T�Y��fٍ�MGR�p�LƖ1g�Mr^���Ábę ���*ok�sf`��sz�e����/Ȧ��1�}h�4����ґx����F��C�o��mf�^2~��9\ǋh�5�دb���r]c�+]�0�,A� Ԏn����ە���&�1O��mGZ.3mʍJn}���s�����.���xC=�����k���N��Hޱ1bOPcd���|�0hó�*Q�U3�~��g&��S���џ�e�E��L���������������fW�JJe�/��mH��΂k��.x���y\�r�J*�S:���^�7k�/�=e��Ɨ=sC�K
s��n�N��_�$@��0K�Ǥ�ه��X8���vB\gŉ�0��!���Z�Td
������A�\���i�����b�l4�����%��G,�{�n��璔ҟ�aq��lK�����'	�'C�ү����t&������>�|�HOP�.��\�T5�m���Q�D��
J���%��FW�~*�ꡤ�0��xoK�{���?���g��P�U����	�eI�1}��UŬFg*���_�.b���)��Ò$ G���(0�j/2c_�?4̍�C�F��y$Fn(Ӽ��〸o�j�6n�U�Y,!��h��_ԁس����$F���6�Q��zv�Et�!�X���$����tLkLϐ�}O�S�+p_����u��qq���Yt�[��m���O*|����螠�$���:������9��~Y�׹b����#AU��i��g2�it4Qt;�I�C�:�����Nq�|��%G�Ѫ��w���)��h�]� �{q�f�Rq~g;d*��h��cn,h�/�B�8�g����vW7�cV��r<x�}�[�V �PD '��J��ϊФ�w�9D��)��X�*Ӳ�YQɻ��Tj�f��ECa��
��n��C2�_!�zT&C3:���Y��H���<����{�3�6�<p�����T���B.	�u��0�MM1�F�&���`RĢs$�� �ɢ�"�y{��T,n�M�����8��P4yZ��^��T�&����yY�n
�JIO_��{��6!��i��gXˁ7�??������5=GmP�p8�r�P����@���ʩ�H"0��$�Kd:�Hz_��>�v�%4���{M��V���`M+�2�ِ���rD��ZZ?��)?I��@���u�S�(D�����-�Q>��%>Q5�Z�
����0򢎑�ow�JB���^5�>�N֝7&��ce��-�D�<�מ�`mX�Һ���.5� (��ƌ����E����P�l��N5-ݪ/u�����ٷ��?GX;�R�8f�G� �s��$����6H�O�J�X' ������A'�)�JK'��,�!(b~:.�������NA�t��Z�*|�*�ZJ��h�d(㰦1i����&B(D�
����6�%3�Ui%���m�`�&�,��E��׈D��_���f$C�RIצ��t���������q井��퍽{R�g��� ���*�rO�ZC��aO���s<�O�� ��8�I�
�Th����T؁�>��@�dW��b�u�T���� ���"��R��f�͌�&�vu�3���9��kv���J>�?�He�t�_r�y��b���|�ρ��$n�"��a���[��no*��͙���nЃ��b*N���nis�B��쯤#_��[�@$��Nl���Qj�
��'��T�R�vfc0c>�^ߕ>��頻��vg��5�����d�0�?�ٽ�jnʰR�tI��8��o��j�8����$��A3 ��WlGC�#h����㎿�쾹a�U�e{7-o�8^(��p�l��# �K~O�^' 69`S��B�|�����9��o/ѭ���.P�����E�(g���{~kː1��WO���l���S��R5����/RC��l�[��#{�wꠏ�	5=)���7ߞr��I_s>׻Z?]����� %	��ܧ#A9�T)ٓ\+�Ayd4r���IJ��u��l��<>��_�D2zv��)A�}ϒ��0^7�F��F�ex:�D%·����P�z $���n��_)V3�����y��2��x|,8Iix�<�i]�t�����\���OBp�� �NE�X<"��
O_=�V���o3^� X]Kg5��jn�hh�I�p� 8q��F}=��<(��z�C��K`���;Wr1ZM~3##9�!���~�z�ރz�����G�H�u�0��,��jT�ji��I.�߇�w����8��VIB���>yЄ��E���^I�Fjca����wF�eGW{[̺iG�Ȼ 2�%z�f�j����Z;�Y	��f�ep"1zt��hǇ[_Xh�83L>�y��\��k�����47ʗga|�0��DB�� K�xF��c�H�
��n�Z6��Jd��Rca��x��֗!���z{5w�O��`!|7<����䩶-H5<�k^�� T�ID�vb������1P&�8�ʻ����Ct�#���%A�r*������^��4�M�^LwL��]}l*�H��#9wK)�g_���wbr8�V��YJ��+�	�(�i�f�5K���3��ӧҲ���ec	>J,x�-V��_�)�̡��A㭜w���v�i��6/ݒ	Qy*�aEx�a���؟�S��dm��Ҏ��莱��	��_�$�n���(��-p�?��a߭�?�%��h��l�^*��t�=@��EɪM�9��N7���Ǉ�mj"�B��t���*��s0T�bU�R�Q&w�&��#��C��[�f�@;�����ut�q�Ȯ��\���e����1�+{�?8G4������g�'ϖm�U�o�l�D���~�q񅁇�1f�<p� �3R�����--OO�8J�B�W��r�m��D�޶T�uPK1Z���q����HT����GQ|Zδx����=/����i6W j�