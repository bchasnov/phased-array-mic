��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�tڐ�!��Q�����xZ�H������
��(��B_K;bA|���.-ƍ�B)�wr�q�h1�oDu�j`�3|�?l�d�U�J��%��{�.Q~Ѻ:��E�)�֪�3��g��UvT���F���ћ�2�&�7}C{ ��e�9�W���Z0bnf��*�TS�sR$���| �<3��5�oO� �2VBndYh�h{�l��
s��P�1�eS��"�&�xδAP�P��E�Ġ85����z�	d������CV�!�ft�nj�#I����%�{<�G$�=`h;�Ka��L|��N�r �V0��w!I .�!έ-9;]��A�۵��0h��e7�W+v+��rr�$�
wx����>4���<�g �}��9������r����t|�k�ŬWTn%5�H�~�\��e6�C�܁�D~�G|�:�L�O��;1�vs}���p1x���}G�GzY�R���Ei�"�x�T�b�ǕU���sd���j��Z�!d1�ԻP�	2jq����"�k�g�����1x��'�\qefX��]!�"ì$Tȝz��\�F�b�+��ă�½��z���@d8��v��]U���q�pg���̙a���QY"h<�g����DRi��T
:| /ðY (����'��Jc��n�~�y?�����|�����%�~�c6iݲ�e[^�&��<�ғI�ɲ��Q{��s$O?��P�2_n.���LM����Drr,]��V��<����l�S�b�����m.�E�/T3a�x����j�t���<LXP �ij Z�N1�p�z2���0�����W*����y�'��狘w��;�N~3���d�GSYhb�7���^���=�ci��m�؃�-��d��Pk�<�lT�}WL���D�mad-E�g���]J�X	�mE�FSaQ_s=l �W�@b�1�i�)�Y{1-d����j�����h�fT�U",��f�rw��*���*c��ח��;Ȟ0��B�u��
��e����
|�^3��cǁ��LV�E����G�S`��ۂe���%�P����/������������HHj�#����w5>��)��L�{48��+�?�_��%�.?V��m�^[�ݥ�.mADV��D�v ��]gF�{��/��h�G��?�-�#etv��2+'z���}OƏ3
E�u<�O���y���{����Jeja.ǆ	5�d��J�%���bqdG��`J�}J>æG��u�[�Ž>�
���]�1L)�ҝ��2�[<�
Ƀ�zF�S�������ud|;��(����v�^��Ђ��e��J�f��h�"����_�����%�*9>]��_����D���E��li Rt��Vj6��xu_�u�sA�j!���k��4����9T�Z��9!om�R"Pⷜ
_�}���uB�c?(>�[9�g:j�iE� ��k��WÛ�\����������9�|���$k�ňi���������!m��[{yl����"�<%���R�_0�0��~3�s�^��LQ�x�(: |�D��<|I���F�i!|]lw�o@<e����{G�R�����h�� ��Ґ���@�Y���ʸ��Q�������g'�,>oR�����zb�Y��R�w���6��Қ�U��p���f����?�E�bY���j@��zI+��K��,I��g���Ӯ���� +�)�>a�,ǒM�Ψ�V}���e'�v!�ՙ�I�@�r4]0~멌�ă�:%����Y���T���E�!*<�7��LF,m��`h?�f`�ȏ�yf��@�p�R��ϡ��)�}Ğ�9��L#�����������v� ��\,�z���I���J��c����z�B�$�E��	�x8��E�2��1�[�/�c��o~h�9Ɖ�/�k(���z�pep�7⳺�wO�����:[���X�Ll�_|���z]F���_�V�����3�&U���3�C��xD����5U\�Ϫ��/��CXܗ��s^~I�`]�${Y ̀�������G���x���ޛ����RSc*٬�Zw �T&J��18/'�Xs�'1��5�\�J��N!�:�E�8�c�%�xZ�-�6)��?�Z��bň��������io��?�O+�