��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1h,�mwG�� ��q�
dh������n�5ӫ�2
�e?4�K�����ps�/)k޼��������a?SrL-j7%�"�1�z忄Q���͗��2��B; �/^R[����wd��\���
A3W���w2�;�uhs�SE�%�i�6H� �P�6��v挻g��Z2
�*UO?���d0�0B5(5��������\��6�j�~���%�W��Arx2�n�+I��}�6}����Q��Ч��]�7��x!*�\�-��Ǻ������>l���Z�T���	Re|{�D��+B��=��3w�(��Z�"v6~.���Q���{y b���n��R�ZS�L��ѓ⫅4�Z/�T��6*c�מ�=rs���ޡ߳���W�76t��_����B����X����?�Z皸H���K�>��_0�w��k��&3�t�b�����>�H��c�y"��Zk�l�scsA�E5 jC�V�R����\������eH���o��N�����Su��ǆ�(�6�jUa�2�����Y�f�����s5��B���������\i N\�R2�q�-N�������X�� 6�>pWW	%���O��:�18K�h$z�D���ڒ( �{O`dW���/!(qČ��Aϰ�qe�O��s��:�So��e�'Kٗܤ�Q1/�����mf��E\�u~vBh�z��!_�w���L4�R���g�$J��w�]CT% Q<kʵ�t*���@�[�\�47Y����dBa�<&��{���2��dr�1k$0� �&���6��/�����c���l����^�HU���l�*�[ß�I�����oẲAv��!]L�`߱8BE��4�
��=
�!=��o*E}���J�s�%�Lq�U���d]�>��7�:�����)(�����q�\#�ZTm"�E{k�B�Y�'W:겸T��ͅ��ݗא̇]�0�ː߶V��; +��)ZZ9�Q!݄o���ս�+����vͱ��M��l������]���xHu{5K�'�p+�:�..��c]��&��K��K	L��3i%�I����LBܚ�
zk���UB�	�)�і�k*G� ]l���'KpL���:��b<υQB��#����TKҙti�D~b�oԴ{�H4g�	[.d�o�I��>wr�82�;0� ߢx02[�v���7�=`�
*��cln���
>>j0rΎ���!��+x��ޞ��v�tU���*
1���7��GO�֐���Ƃ���|C%D�=��$r%W���bF��Pa�0)�geu�c��JA�,�뿖�ǞP[+p����I@�E~�1�z�|�/�gI3��<�񥂂g��H<�~K�U����.X���h~��6?�M���J�`lw����W���[���n����2,���y����E��k����0]��ӷ��

����4uO�n�������튇n��#~�Uf�����/Rj��k���p��a��1%@r�?�L�6ͼӰ��i�v�:VmUDNO\�7�����l��{ ̐7[U*R�`��Z�_��xh]G"!Nl��|������L���}��<�����Cr��g�O�L�[��O�n���w�-l�xUB2���?@�����&�j��j��F���h�Vq4}ˎ�p���d��2��=0��~�2�^��~1,�\l���$�"PE6
�5�	#^"���'B�~��o�~K?��(��b��C�*^
�z)����Qq���T͙gh�ܦW��S�U�Ҿ
�L'b��WI4��q6x0��h��f<�H�[�D��OD[st;�$�Z�y��-w���DyQ��� 4w�Gk���p��]bN��|eb{�xn�
?�U�q�Co��"c#x��:���q��q_�%(x�M��`��}Ӎ���SWl����
�{�U�t�mr����:j!����]���?j}9�ʁ)�79ޱܕ��������)XG��E�m�n�q�64pS���S�`���Nf��N��C%�D���5�A��e�)�z���<yY�uX��L�cpt�e��N?O�f��{?�c���i\ ޒ�����qb# ��҃C�\��BE�#�~W)}*��YϒY|��˭r5kzĸ�Vo����{�\�dz��#J�Ej��������ftE
"���2��9�(BX��B�޸��2m�g�����u��3��[S
��t�\��&��SDd�׋�7F��87h��h��� ���PP��6��Ke����U�.BdJF��c��#`���MX~�К
glAL{���2���/�Kd�/������G���b�]����W��?����ቱ�Ş��x�"�^��!/�7fʱ6� j�����t��|�*Q?7}�0d�f%lmn�%]爭�
|�rQC�1�nq��R��}�罈�i@�)W����qӳ����=�/��6���0���o�dE&���*e!�x5~�d��~��n�ZB�	�8�Ӹ�'{.�xl�|&2�53z��q�9�Տ�|}�ۗ�)ܛ6��q�g��dspVΖ��A�O���F*�B�}��o�˗���� P�'��j߲�־<FȤ�#Z��0��Gz��Y��u�A��K��HOQ	lߜ(��~��p��I���-�u��+�o�����Vµ�n��Z�>,�3�0�㯚�>~�W;�O{�a�b��,�\�ta��y :~7[�nf��ف�W":m� iZd([\����\��Ep� ��tOB�7v�/���3tta��E�u��u��qC� G�յ~'#���r�(���\�������?ؼ3q�t�wU�JL�k�}�nC��eo��][�v���������P<��jd�l4������8�|����ĕf/m0�ɒ^��gD�:?r�2-��_d�o��҇�Tpv7O������9� �����ʇ���j- 0�F�9�\��I)�k�����H��py8v
hH����\Z(gt�T�ϕ	�ֶ<����LҚ^�C�뎥�4��E�`�d��7E���<�Z���w�d��/({�3�}͜��Ց�e$��7��$�kŕ�T���I6x���%G��Wn���2"�,�nOڄ��m��d|�0 �6��"����H�c�~�p��_pW��u���X\�G%�+���\��UWb��W��l�i3���AZ-��'��S��]�:e� n��H٩�ԭ �.Āp���UNw|�c��i��E�����;��ǆ��m�Y�������I�Sژq�͂R�q��r<4�bR(V�O��J0\��R�Y�tς�*$z�Z�ʒ�����:�0q�$p`fc��)m?�}8)��@�NM�S�G��zf��mIj�޹�-��a�� &Sq���,�YJ��be���ǒ=�Y*��֧��߲��7�
�~#%/}쬯��Q¼h�
�VG��H�k��G��b�	����������P�[q�,3Gƪ�@�>�ӵ�[9��Mؿ�k����7���ן\���yj�	Iŉ�mE����"%C�}U�-���M�l�<`|�|��{]�Pf�X�`u�4o7�d��Q, �>y�ڦF�Q�3]�������������XJD�P�u\m���mJ�;��)ܸ^D#z��1�y"��w����I�@�1�%�ʯ�+�3���8uosm���$5�ez�V���h��FWo>�^��"�F]�R3��5G�nQ ��Y\0����W�j��]4��a:{�M�xd�Y����֛��.���Wb$�v4ε��[�fp/�'��)3����j�K��� �RM1|y[u�CA���?�]���ZB��/������]���\!`p��ɠ_*��Ņ� �w1|�]�&ud�a�b��BR�3XE�%"�4e���oJ\0}ZY��[l�g�G��[���S��|�U㙙n���˩��N �7��Q$a��BN��3�zo�*�A�{6 ��͇�D��1����56n=.�g�~Q���O�}褻��[q%� ���{�~�[g�֛6)�L�BF.��a�D�K��Z�^����J6�����
Z��ͻ��1ۤ�*�(��Wl!�����
x�����S�}��D:]��`��:?�]\��]v_p���LH���cO��%X؍��)#g��� ۨkR��y~�ݘA�ꊷ*)_��á����.�wG��mr ����;zf{�+�5F�I]��͕U����&,���@
��"nX.\V�L�2�!O]Q����W����s��J��e-l����ѽ�4������r@6�ޛ��i����Y�7�~đ6B�,�? z���I��(}a�=�z�nP3�~'ْ�"�V�Tt/sGM/�����$)�U���&�� �ַσ-	�YE�Td§�G��#�Dv:Y}|ُ֭�i���G>�V� _p��O�#���z��C�6��G(N$:�V�!5����z��g�rS]���;��؂���"8��Q�5�x�I�d�*�!j�Xv�q��i�ya�Щ�#d�����C����o�^^sT���>W��%�5�5"G/C�ݰPn�צ�{L��
�X�P��|�͂�2ǳ��۩4��M������D�+y
�H������`lԔ�����Q<��z��Te3�b�n����Dz��F��[ti9��Ck�ʡ�����E�:���.�hbނZg2M�$k{2���Q!�<�X��<	�ϧz����5޽���p���>�{h_�.�����53]YmK1J���<d�*���&�� ����w9�Qpw,��B-�g� �ID�Q0W8��-M,��=F����;3��)�~��;�ջ���9l��&�'�j3����md�z�D��җ
���1!���GC_l��\��7�m����wd�T�/� �qWbw� ���V)Cg�<�$US���6=�E�V���,7.��0J}S�����7���G!����jC��5��7�n�;�T2W	c�o<VqP�
?��i�yS�f�M�IoSl����q��~P6�A���9ɺW��<��*:dGN���(�UR��?�g�eP�$6qQ9{����ͮ埽izZ��(�[ࣣ'�Ϯ���v��va�$��d� r8�$O�߀ܹ7����C�ks���hK�7J��2�[e�k�Ov<g�{Հ�?�F*�~�5��0N�[�݈4�W	�y��S�1Ԁ�HO"jh��ks3�L5�j��Zl��pJL��S�b�A��	�����e$��)���َ�$k�f@�p�������� ������ _�vC�ճO��F3>�q+�5ED�a�z'�׼������YEJ�]�B�7ԚQ�������zm!�mڽ��Vaޥ��KVT�����wc��D�]�������f;��_�X���t>�������_]D*h'���Ϸt�M��J�n�����6��)�J��'OZSs�̕�����m�%���.F!�Nsu�����gԐ�6@R߹ڶ��������%�_�DzF>��a��Bj��;>�[WzB,���r��|S�9-/eɥ����ᵸkS��������<|1Ô`{�M*��N�[�e�t����P<�+��f��%+���S��5+҆��Q�x+�+��p�U��Y�@f]!��I��A��R�e�c8�����=R��G���D��:M"�<qE䨾�(c�#畬db%SE!$�09��}�r�7�cw�Ф �Ƥc���D]�|�D� �����OU1|6����"J��A���������|J����3�  	�#�(=-_o��z�+\�H��R`l-4�ݿ�[�'?k�q-_�T��x0O��0Zˀ��C�>J ��So�<ѥ�#&�.��Sןr6y�٤׍;�U�ʅ8~6}F��7N�,�_T6.lz�3�} "��Ҫ�F��>ҨN���2��dޱ���3�O���7�E���ᡛZ��F�E׷�(ֿ�ڣ������j�<�f[���LE��Lp�/��[���?Kէw�Y�ET�n/5�LM�;,z��~�+v�m?8���������ED�-#.X^��},ꁶo4܆�	��mS}~<Yڌ���?=-��K �+�LS���u��9ô�"oXl0y�X/?��W�O��ɦ�k�?�52�	��X��� 9ض���J�*�B��=�&M���-�hձ�E��B<��ɀ7�rp�vRD�$,����`#Z�Д��MWQL�ZQ�آ,N�'l�&���s�zV����3����Iz���T�I�W���"��w�yx�8x4�$du�1����7caE�hQ��&Q�g)���}�A�s!�
���~Լh��r�h4�;o�69hє�F��L�ӥ:�I�!UE�݌�t��n�&G��;��c.��|�H��\?���i0&_����.���=Li����ChY��:�p���>�3�?��+�a��ݦ��uB\GhЦ�y���D$��^o�yV�lzꐢ��Ppſ����51�q�H(RӍ�l��%^S��-'�� �?�������xEt(51a���V�B��̔��V}����Ƽ��.�ɑ�v�$"d�`��E�a8�4�T�@��}�\I������Һ����ݰ�]9m�{��M�bЕi�^O���,����L����܂$���g���
���o�ˇ�e@��d�6F �	9|_�<dL����o8���f&c ~���[q�`����G���"�,��a����- ��2����@q
�TZ@�#��b���"i�P������򝌳_�d��]�P�:���1�m$�g��UG�n�pg�G`�e�#l�?�3y��S��Pt�������
��<�R �U�K5T�Ν�$x����K:p��\�-4F^g��+���f���?��l& ��|(��︎�{��7P{�ȵm�N�$��5{�\0A	A���'25� �L`lx�"(��;��dq��)2�6c�	2v(�yy��zXa��tְ~�pM�W\-),�����ssB>����8lT��C>��� ������m��b��6�tu�5��a��Q���됡��//eI��g3͏���\�ȅ�$����U�<Ov=�QP*�\���;�59���3�QE��$�+�f�
`�X�̒\��'��I�L.h�)�����is��B��{n=jV�d���G�����ؘ�;�:�2����c��+��ϐ�s���ȟu� D{�M�>R�'F���s����%(`�%��h�`�?hv�̷�y�X�%2!O��Du ��l�ᣚh7h�.7 $04��Y���X��\�{�-��N�
�
/�����9ɵE?�����������ꝃ�O�L�|s��Z�F67{���#��L��{[�šq3�)�vp>d�:QaA�7���8�c�����I�┽�}Z�܊ƈ:��|��?����_���Z�>�N��`���N��%^�r�#gNF�8�.�$�W��~[Q)����J���BVd넒��/�w�{i�D�\�z����*g����JD�!��M�S��U������~=�l�G�b��c��P&�߂\(A�6�H\s���j����qG)L����~� ��qg��%on�)�W6��+A����I�r�)��Y�j�7ZJ7�����y�aԼ��
ס�����8_ҝ>�`�`�M}�tж�^J�(ϸ�`^2�0����K)9���e�`&������E+���i"+��'�1ϒw5���a���HU�t�~��x�3v،�\~ P�Q��s���j���v�"#bgޑ_��4�=� �jĞ�B�X�܃�`��_F�/�q?����9����+(�sY�t�~��(�]��_iN�b�聸�
�@�t��g�M���� ֪vM�3dS9��
9�vG9ĕd�s���1�xw<:��8n�)��G�+
P�"�m<�`�O���J�c ���m䷕��ë� �ؗ��
��5�X��_��,w�ַH�P��W%�����6�sT`g��ΆUj����*��Ri&!7��G+19;�{�1�0�cU��Q��&��t���̸��D88�[oo.�%�|��c�T^x&