��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�P�;�{��3�OT����n/\�@���V�F�	G�V��]� z�`t���y[q����a2�QG����c<iU���z:fj?�?��	1פ��s���$ɍ&�oD8-��\����6 *�+�I���LYx��"qJQ #��\}�; ?8m�)����7`���#��'���9��O�y�bs}���횞��bwk���D�|����l�8?����He�Z|���jo�㒝��� B��HO��bE��۔�=���)�k��BW�Nij������%&< 5y�Y��	����τf��K�V�R�Y�L�0P�S�*]�8EK�a���P�J��6�H����v������E	����}
3`�ge �d��1�$�ܬ�\Z�tRO����U���g(�n8
�8���K�y6����S���Q�,zͰ9J�"eP/�}F#,o�4�c��;������A��2Ҩ}�S��s�d��*�W{�-?OF=LHWǨ��⴪^�}c�=���-�
mӖC�е0��
���.X�>��ΐ��v0'�yɃE$WA��$\��F~Ǣx�c��"#H��- �ד���Й/�Ci��J���������^	P�`��XBn�ݽ[=�������� w�#!QQ�DhK܏_tڵ�V��=�H(B��V_]�K٪%��a7HL}�u���ܟL���<}ݕ�]1Y��&pi'.���|r�煯ܚ��h���D%�����F�bg�S1^�Ү&~H��1>��W=n ��C!�id��2gZCeւZe ��Ԥ��K�������A_�����np��uf��L�k|�Q]�tI��dPt�v7�q�Ե���̭��)�C�5-c.�П��(�g6|g�RH���E��_� K<*R\VoN�Ts�r=�w�FEl.���j$�N* �M�u),�A�|9b��&��ǒ?�ى�<eH�*��3��'��5������+N#��Kl�a�\ܛ���?�>��3�k�[�R�'���� ��C��z��!��f=�ّĀ .F�;S�ԉ�O2��]
��ݦ��W�E�M�$]�gsX{:p�M�8Sf4�9%%݂��*9���`x!�-=ФE�Z%>p9����u7%O�)�ȩ��򹯡$Z3���=ѥ���V�ҩ �D4�bq�܎�ӿ�x����Tj��xfȮ�)HuU3���J�o�3g�=�w��SF H�T<�B�`��MG7f��-��ʾ�b���1o��zX��!w#*	��]Kb��_�}r��xg�r��OtdO�B{����њs����S㍂֧��v���GԆo��RŨ6z�*����,����
��zC��V,�� X��T��{̆���gTmYb+��9ʒ���y@��&���j*E_5�,Gz돀2	4ԲM����u��ܩ�1�!o�h����D"��ˢ|B���K���7�k	 �����V��C��OYߋ���	�>�/[�M!�����rD��O}�
�,BQJ�P���	��nTB�蛞e�R2�&�׭��f����\��^h!0�3ek�)����~��h�e\Yk��5�3 &K8۵1���4}bh���j�����ou��^�p\�4aV�>� $Ϝ����N�"x�7,b�Q�̝�%4���$����1��bI��sCV�HL�%�<�?Ҡoqy6����=lEW�Q��%���(U�J5��9����g�k�]lk�*p���W�+މ§[�;�; J�,*�k`6�CNMH����/�2�Ff��l��%EWF��7�TZ�T���I�������^��H�:��e����}GL
�EP�L��V"V��z�7V���7�_L�I��И���!+ �3%���" �)�]�`|}=f^����V��`'S��k��I"�(�wR��5�	�K% r*E�Θm�5��/¬TqxL�|G;���L3i�������߁PEԽP2��~犡������Pa��y��'R[�8�Ņ��}�2��$X`�V���'�u2��V�Q��/מ5Z�:��dF~ɴO���s�b�I�s��ߛ&�h��Z�"�����_�N>L�ym��A_�|�)�!�6�%�ku����"�NM$��\���p�jJb�n�g.Y�z{NQ]ԕ?��& ��@�Fn�<�� ��Θ!���9H�w�ܔ"ˎ���5�������`��%;��h����W��J�����W"K]؈�f!$�  ��*M��OC��g7�k�6ݘL2 ��{ۊa(��=D�`�,�����A�3c녷�@����u�%��p~M�?Xߺ���S���TAЋ=|ײ��
�=~X���	4S��d�ߌ���ψdL��g�1�ҭt�m*��ғnWǱvejOPL8}0��ؽ,A�p�\�5�AiܶS5:;�)<��>�OF�b_���US��F��ű�Y�J���&�[�Y��T�x(�@�# ӌA�ܖX��)���1��|u
�:���&�uu��ގ�,\M�Q+�lȖ��|ÌG�<�F³/������{Y¢��\���˚E/���������̇7�2<�5?�5��Y��V��r�G"~��U0������e����o<��I��,*d�=���1���3W�7Ŀp*Y!�(	�l$DWA��x�):L�Z���V5b�bjK�
�`���3������k��C�>;�.���\�^_c�n�q��T$:-���d�8���Q�AWw��]?3YC�C������/Y,��O�a �z�O�y�����5k�W���V������$���q\�$�O5C�Pө@�QWNw$J�w�q_r^��2_� ����[�$I4�@-V�B+��l�g<Az�����K��<�#�u7�#DM����R>>}b���*��]��������_&��-���iv�>� `����be����
��=b�x���O;�p����4 hA�V��}-�������6zR����n��KI�3ꦺ��
GҹG^��zJD�<�?��0p�*N5OZ���6��!`�\��%s���H6��|��������Vq�<I��WϘ����Î�΁k�e��.��9�/�B�[eW(99�r|�5��3+��Y�74��=y�'&�<��]�K����E�V9=i�$��&��x}dX�/��>����7޲ ľ�@��T}��k��8lB�i���uv�����i��TK��<��1�?j��Ɉ�����}���r2t7ɽE��%�#�W�,��D����
[ C�dUb~�� ��T3�l���v&�$�<n~���?�DK��؄�e.y��tV4��U:Q����5�\%��ɐ���5�^Z�C6���e'�5����{e�-��Bj�Pr �1��B��(*h.˟�o}�-�W#-ܣ��/�I�
�p���_�oI��w�A�?�m�ъF��ArjR��oG�[��T!�3�D,��칹^��/kzR*?I+(���o �N�@5��pd(rV:��뮧3�� 2ٱ�ڽ�.� �0)n��;�Bpm��K�Ӥe��>زa�v��Qwu���]kWʔ�0Fة>!f�\)��yE��<B�Yw\|����}3��M(���&ϛ54��f��#�_ =�K,�|���Z�X��4�DR	%�*�!�U�ɞ|���,<Х�����0��|C�h3 )Zf���8��n�ibU"���f6����)Ơl�4�E��j����\yMBT#y��q�=@��!a�7,��,=�k.�B�#}�@9�LhU�#��Da���0u�+/�ks�,�BR}����k��?^�Y뱉K�i����S?�6h�lIBC��7��qPjw\�t��OJ�����w��l��b��] ��w�ʣ~���6AO`��~G �=/�הS�d��H�*E}���ס��B�T��]��	�<���������el1[^���z~/P{�E�Z9�X�����:ʵ��\l�'搓4��w%aa�j�3H6�k��ZR��]��O�K//wI��8�x�ܶ�Po�/<�>�Ŀ������jE@���,�n�C�d���f�B���
��ᙋ�cǰ.�@頉����6f�����l���J�x}M,[���ظ� ��mL���^�gb?��[��,�#�ϡL�zڪ��kTJyy�{~��&��pV�J�x�N�ܡ��|�x��6�J;�!�a�h�߅��N�IQ�!*W���T��Q�;�}� �Dހ�s���#�}�l}�?_��MVB&�j��yS��B"�ed�i�� \nL6�d3���|�7
E����K�szt�-�Fhr[u�~�����M��2�f褆5�_���b}M���dŘ��2�=����AH��O���L֥) <B�I��(~ܓ��K`$˒}�F����L#Kvا==�g9x��+�}�FH��� H��l	x���-��x,{������D>���[V��ȝ��p�X�b��ʳ[��X�q�uJG��S����}��j�BF��b�x#t�v��M̄04�c.��`�<�l�$�Bv;}�$w�Q1x�Q?E��O'Z��XNQ�0��ژ�����	2ou��/mf�O9DS=���y�H�n��dCN��7]�N� �	�4��
\�H�"�\���|�'��� z�q��� �7�bF����Y��,ǒ����	ys�:�C�G����g(9}Q\U�(V.�?��Ak�~�$���N]z�u��4��e�	a���G��H�ө;�d�'R���!��M2��2��?4�z�G�G�7����$����ŷ|���>�chZ�6+#G{kN*�yˬ�����U@��>��l�8�E��j��\��6<����/#ק���^��2=~u�iօz�0���`�Ɵ<А@�Q#T��m�˸��H㚒C�/��}]�}�@��";�`Ɗ�!�+Pr�
=CQ稼k�:Dȡ��X"U]�Ze����Jx�@E��2���=���X���Y�)a��u��:��ǅ*���n7 ����$i�L�֟jr �wr�A:�\l��:s�N�ź?,�K~��lM,�m͑�8h|�@�9����g1��^

ٽ�l���hg(�-t��k?펯�L�Z ���<N�G�6�:}���9�tb���|F���?6���J���$@P�/Kѻ/����3�<W�0������@�=}�#8m4ۜd�}>�_A�>E�2�ᨙ�pg��<*-K$��`��+<WK�������"a%��PĶ@�ac��DH�N�39Xzo%���,箇]�<�s��0x^����81q�Z���2v��� w�A9���]'�d�]@6?�u�. ~�]�����޺$~Z@,� ?6���B�<��"9?�_����_��"�w�e��ٙu�C�/+��A�"�K1�fh�"����)E>%j��ޖ1����'���)��n���%G�c�' \���dQ>7��$�����E)ɛ��b�"A��]؊b������Q�GU��F�GU�����:�2���'T-��(8�J:�Q�a�1�|�LR�H9�	�/9Z���<�fUԻ՛>��-��O!��*�����*X��u8|�����|Єi�_?$MY�0�&��W|o#u��0�$�l�o�q+s�ʝ)s�:w��w����L����gw�a�A���ჲ���@����FH�b�3l�äO=��1�c"C���P���	���;�#����൉��ot�A������#�IuǱi=��4}���
Т�_j�W���{w���<�Y��V^.X�r�FQ?�(���
4��S��p��?h���^{�F
|�k�:�+��Y������^f�㮀��j���D躁�ك���@-�77��5c�:��@h�w:��џ��)�Z_X�I��E�4M��ᦻ��e#.�^�Z�	|#����u�{��~4)-��<-��t�9��M��{���p��V"I� $ss*�V�+l�:E��"���5*����P�M����Wq���pF͹�?,��6rw���g�Q&�LΘ�\qN�Dʴ��im����2N]Sv�[o�gT]�N�l��əG�N@^�ڂ�({�Q[�.��OXxNw$��`@��-�9�ܕ/�>V�����E��������n:(�`�_3;-�?�N�]�!+�y�mzB��i�K�k���D�Z!�܁-��/�\���覢2�J���a��qye�al6Ȫ{k��u[�2C�~�����[O@:ƍ�M��U�&gA��߁����*��C��6�P-2�43V�9����̥;�|DTO�$+����9uQ:��V���,n#1\�J�n�*-C���;)
Ho�E�~�&6	�MԸ��s��㏀��c-mi�% ���ws���h��M�P�ۋ2�� ����Lz��ڵ�=~������!I�V�V�����r���[b\�i`ܜH�A�:�9���*Ɗ����Ri�}t+�Wv/�`�&���eS���L� 3Od=�y&X�;z���4���<��l��	~����
,��ʜ�K�k��3x�2��'���U;���Y&j�W<Q�W'�CV&�(!����k+�1�q
��vF�u�.;w����"�b�i<�������D
E߾�Wk�_�Dc��v�t�<��c1C<�4aI�g跿}3�y��e��R�M �nB�ˑ�E�C2%���F��
$D��"D͵6U�NX�c��ϗ�I��a�&F=z�b#WZx�'�q*ѨVҧ}�h���_�=���]�;g�R�XU��^<Ɖ��a���;��Yv��Pu7ӧ_ ��([��MԬ� ���l٤�qq�3"h7E�f���Aiif����@�����j�^�+_�h�XL����:�*y��W�P�G� ��?���L����"ti���$ݡ��o�y�T^�2oђ��k��H�J���#����� N�����""~?�1�P'kA��8�5&<��}���=�C���P��9�����b#ph��ȝ�)8F�;R.�]���A#�xχO���j�X*�����-��W� ��Dc
�����m� �Q��底7��W�y�^�-�qy�F1���SFy�܋��CRvO��H�8����"zf�Z��M�xK�& ӫ[��~��C�a�1Rk[��ߍ(��r�ו�D�3�p>����HPq���=_ӵ�J��եx\�yf���{J@���,U�m��i��g
!T����v6!�`��7�de�n���1��"����
9�,��.
��)�zˀ��0�|%���t"�B�|4ϙ�>-D	��4���XH���ͯ\�.i��^�h���-}�_�Q NĒ��u�E�dc��i�U�q �1f6`��O% >篊�3GEJ����t�<�sҹ�q;�|����b���([�;���W�8�id�w�>�Os *@�)j_����/m�<~��YV���j��OlJF��U��{�2g���ą��g�	{��d���ۜ扇����X��3�[�l�)�4W�����>~��^ܗW{��z��|W��l65�Ы�#����j~�m�S����q��Uxj�e+"�H٤[,._(uEj/�����3���1�31nȒK���ƻ�]����(�Wk����ȴ��.�H������V�v�NIB;� �nPo&�X%N�WǻГ�$��)g��9��Oyx���3��,K�1̿s�K�׏i:	͞]̨�n��f\�<�x�K���u�y(��fZ~}렱���90���;��!��3 �����@��J]�H�|��C;���]��>�)'XO�i�ğ��t8����Y!'m%�����ܡ��0vUVxǙ/���	�V��á����y<�W����]W�������=c؎��иJ!]�u���A(D\� ؔ@�z�g<=!|w�ۦ����$�v��q�I�C��,��U�P���jQ�
f���I�rя�oO"B-���
������]�̦�jf Wr��@
T�Ć�#��@c&�3C}�rE����
���|L}ՠP���F�^N�&bU{�MC���g��f>����0f��{�d�*���Z�l��~���05�5���{^~ٲ-���:��~�#���ЇI�4�u�ϦC�a��;����Bʞ��6=F�'5Z�>'���UyЕe�(+�$��8���G��H���p*��M���������P��W����;��a�M�_�	�Q)vq�/���W\�������@�P��}�\W?,;��@�DL��y�yu����țZ�-&���9r�B���7��;��Q����̋DV��Ե�t�J�[�76hQ������I�B�s��I�1��!����Dez%1�>��Rv{r���k]��;w:�3-���$)� ��Xl��ma2-����q�����l�[,�%�,'iɩ�@�r�����X^�g?�Y3��+�"��O��Q�<L��؜|�D�3���GY�h�فĲ�޶�a����~_tb������d���@�M�v`�^�ԪN�׶��?�W��-����`ɻA���5�-D�-��>g��H>�z�a���٧Q݉���s���,���=�K��.{5�E$b�������B,��b�C*�E��	^�	֌x�)�j8�(Xf�h�����1N�'n����8�}�`矛-��C^iY|��*"�_���Q>�濋�2��.ajE1qk>%G�u�N��x�N���cѣ�b��R�S%PD|�Cmx�����f����u�6z�y���`�.����9���T\�}���C,���`��󂜧j!J^֙�W\��J=����A��γ@�^�{�&0��zu�z_2�ܭ�`�z��S`c.�~z�^ƨg-d'gc�0��� �3��WO�L�������D1��3Z�����_��ȡ��qʓ�¼2����p\̞~�#�9<�<���~T�rh��:�N�~��'�9��j�Yg���36Y�R�f��C+w�m�<l#{�iJ�iY�R��%׷ɪ���"���:eF����8~���P�O�~���;2H�ɟ'���b]ݺ���R��$M�ل3[���N=��C#�(��`��X��A����5�!Y_U��0��S(1�km��ׂ�xgC�|���5I¿�+2ٍ5��;[۹�VLjm�I9юM'}!1EËLV]���U�qM��g%a�M&*m�v���Ә�~��B#��^m�V�k� �37�C��RR���s��I��'��%[��~�~�w�:�˗(n����}q�@�!�d��Bbwz�Ď� �vƼP,^�2��zف�W��.�<k�e�p���OO$ˉ�����53yhV������}<��E���_�],6�R�C�*����ͣ��uH+������V{I�1;�R�o.�SMT���C�y�u��<F����nd%�(k�"Q����,.#_���z����<�D�| ��"s!ᄔ��Y�h��Nx��%"��Q�/՚Y �j�H���fNP�e��<Ce,ȿk����H�/_������2/�5fYI�OYr�f
�)�o���F.�lD���w���N�v{_�xot��y�n��j�S�u���N��L_�y;��ݸ�n����䁑�g�T�3��x�fVV	��=Æ; TD����,����a�Z�ɖ�t00w��3��d��V�}����#o��U�|^Y[
�T�Y��hJs��HY3�Y��	��� p"W�:�G�����cF��ҷ�v?���pR,��U�����
�]�D�&ͪ�-��pU@�Y�>��@���s�����is�]���K!�K�0�x�C�j|����:�����{"�͞���p镜��y�̳�r%�6�3X�]��Ǧυ�,�o��U���u��M��׵�-��.� l�B`� *�R�\��bjӧt/"��9� \N�d��������uD/�Α|E��S0җ�F�q�g��T�7Ǚ:$;9KN�r�3S������s}�ܦk_�Ǌ��7ԟj�B�Y��&�Y�����������c��Z9dU��#@�H�$-q�d��զ%:�Ćq.�FFk��U�@�Z��l��<����'������V�U�m��Ѝ>5U�u��Č�A���)���!~��[���o��K&FJ�� ����<w��Μ<��i�;C�"8�e���	�ݿ�##;���UYr���9"��D:U��ۼ��v�8k�&@�'M��Kh�웾)n��*�lFX�D��m�2ۗ6�N"�#�[z�{�J�E)�7�*{]"/[X�ƒ��Iq�vVEs�0��K{츬�<��&�H ;�:`,ºM5����)�E�_P��?]��� �g���m���G�i��g��u@u��H^@|.(��P��n��q�e-}������i��D	ܣ���J� ��G �Id^��ā{�͕��{o&�ic��~0aKR�m-Xj��A�qh�W� � 5�Adli4�i[�>��Z�b�(�D��K��8��������W��?�73��3�g�+���G�9�s_��8��2yZ�j_:B�3/rA+�4KaZT�-�����xh� ��D����h��5�j����^�l����ݖVt���N����$�-�ĮR�����w:u�]��٬����o	C�Kd�_]��I��"��������Ay�I�W���EԼ.����d��W��ڥT95����D{��`9��48��y ���..���"-S{���*��(���\C�l
. "�R!�@ƌKMcq�N�4�Ee�nEah<t(u���|�.��e�Ͳ{��B�Y�<�`��+��N�㛲b��W. L6�B ")^A�S�q��q���#9ة�gʈ�Ǻ����w���֐	YUǒU�3���˜���i^�h�bQ�g��+G��e�U|���U�am��x^��$Qf��S�e �8Sp�7 -;o%'�*\�UV�|��F$�#ך���XT%J��ە��qH�<����Nh�?,�)ri3�l� 9��t]�IB[!~�
��/I���<�/T�4�k��w7����.�_��H�%�~���;T�.�G���k���C�͍�A$�Ku3�ۧ0�S �c����?Y���/��^���ɰ'.$�.P����(�M���ts��Џg29��W�uw
����pT}�J�3[�Pd�jd�R��ݞE���P�����&����*��_�=�H�
��C��r��!�Ħ[���$)+4�(psX�� s?�';-G�d�i�D
������(��L�Q%O����ٙ�Oʨoc���G��ݭH=4�r�f(�<�Y�zaFQU�O���UH5���1�Ei2Ď|��u�;c�/	N��' ��H�tG��ʉk�܌�uY	��O�x5�O��w�\u���E��Ϭ��m�j���)(�ӻ?�$M|�@ -�a�8#��QŹ8<��n�?H@���i�'Q���I ]Pi�JbU�Rj��ڠ.�����d��E�џ�<af�(��c ; O�週a�?"ִ�:ev��09wL?�Ԃ���=��	��r�s$�H{֕fc�!ޒ�Zs�2�R�N��֊F�j�6�-�J�D��dk� U0�r�P�.^%>oG��/p��N��Z�������Q�=0���G�M���_v�\��J��T̢�}��`�B�r7�e� �U�U�Ī�U��R�x���ߺ	U���	�+��XE�8��i�]����Pc�]�,փ�c�K�ҳ�#2�7�\����6W��"ZR0�^M����\������l���ꖴ�Ǖm+��
z鷍�D�����yUCɘ����1
��@	0�����a>�όɤ�v��vs�{��$�=�J����#�����c%��Y;����C	����� �9��vUK9��!�c���M%�����?�V�W�%9N��s@���`_X�!��(/3Jl{�b�ZcGp�x��>�E��mu0n�����"Y���$�Ֆ�dR`��H(���j���T3�"�Z}Vy�[�U*�)���`=���>�D=.��mHݨL����A��'��R���lr�.�UAU\KYpz�9H�> ut�����p�/���E;�j
/A��9���蟃ő9K�.��\A*����YUf��Z����Z�,;�}�T}]bh jE�l�O^߀���J�� ���!������ވٳ^]y&���>��]��80
3I�����h��K�w-H��T�\Aa	��t�A�r�	$9�lL̥���	���6�2�Lt�D��<�S�h�v@ �[(��f��TO�[�,�d���C�k��*p�B	�4fC�V�� j�����,"�0~�#.�7��P����`~;�u���%��8�q�ջ�����L������¯��N˴�+7��%�nAP.�1�2�������w!�|x�cn�-n<�o��m����Z��T	�����FZ_�4�3��q�<Ҕ��Eأ3J5��ۈ�0������ŀ!o���"G�i�`��쩭�J���t�H>�l���(Nh98�ځP��S�W�t��n�h:9w0�m��se�h�'3�[<�Ay��L*�4^X;g��N�rlH�LH�8�A�����c��Y<��-z��W��2�/�Xzw��b��v\"�r)������l�x��;>(kǫ,�f�Qa'����ː�hU�HO����r�|��ꢤ-�Z�S�	�Xmm}+<V�#Ѷ
LF��P�_��'4"���nO��ՉO%�5�l�O:�)y��[���6ڐv�^%P�1�-�O%5���qsenʭםN�����n�b*,��`e2Gy��N��.�WC)�?�a�u_ا��D�YeC�0��y*?�qe:7�Y�����@}��D(��T·G�m��}!��z�׻��=����<Zs9#����w�\���W��ܖє<���{,�+z�C!�%�z���0�jly�����Q3%4Bd�^�_
���Q�)��ݽ��<���T��
���怠BN�+ٰ[��8�D��(4&v�� ᰏ�/���Z�R�N_بDGAOLu��"�y�g���,����k!��qh��Z��6o7��!��sԇ@Z��m�dɎ���l�v��տ�_�9�e���G��#S�B�i	'����3��u6��z���*uG�����'���Q`������7��Ԛj3E��nr�&���z�G�݁Z�P�q�� A��R��=wb��p���_����@xtqs+~�M�Ѷ=��F�%
{ϴzU$;�Wzu�M2����ǚ���$Tӿ#A�1��æP�+����b��������k��\�nh�!��יз�;�(ڲ6�9�p��z���h�̂ݠ��x%o��]�v�> r]p���FJHƾ�B�e�	����M�	�ոT��֎�Q�*�nn&�C�����/����3�Dq$�>
��[�$�΂В��k��(�fyȔB�����M!J�\I!	XRV�<V؀L�@P�3a
��eu��+��Rχ�`�^**.���׽ �b�go�z�l9aBϻ�%=̂�~�I֢W��
�%1�*+�Px>��v[�%`��b���Ω,�C�uV�������+�Zg�����b�a�K�QJ�����������v��U��B��K�p�����]�0���Bޢ���_��%�$KȺ�y�OrD�S[M���H�����E{�> �).$�'Kp0���1n�H��R�&���U3�+��C��HjL��g��^ٵ-�,� ��G2s���[/qø�4f;ϻ���y8h����E/V�H=8!TՉg��4�)����f׸�&I`]h6. �9XE�������Yi:n���)�*[��w�u��<w�W�sY���`�Ą�f��{�w)�!M{6鼃�^8Rx�r��R�I<�>|�� �i&0	���J� �>�X�ʉTQݫ���%����,$�-tٍ��,:��*�ٍ��� 6�\S ��
�������E�a4�^��f�s��o�\�Y�o{:ؼ��}�ۧ���^h�!�M�~r)،��ֿP�O ,����F����"����T!ZYlxI*T9	bkD�;��e�k�A�,�S��O���6?3u%��,��G��p"��b���;�㉰3�N����b ^��+~��58��%�����<�9��"�&sE/�o׿��x�kG-�5�3	��Q¸�N;�o�I��N� �]J.�Q�o7�n�E��E�?Y~}L[<v(N�Plt� �h��'=0�~4����?U�x�j�b|��GT�����	�Y�,`RU�����V��=����]%}>$ń���c�f�*��v.$�? ���ٞ'�>�Ҁ����������{�_���U� ��=EװZ*E�w6j�*�pZ�F�_�cu��E�
,��^��!��������H*jѷ��R��Y/h1~�Y�Z�i�J�'����_8
r@�`�1��:/.�A��kK�%��6r�y���\�����: �aO���^d��9+�����tF��$E��ѧ z��E�<�գ���y�꩐��������h��K�{1w�VL;q�F��Z�r�4@0���t&U���^F'^��
���q��>9D7�n%o���\w$������)e�i��������Y�Ñ6�	<0k SM;3���k*�;p�[Xl�ki���
���T�ӧ:����ηU"�,*r�^��Mj�Wk���1fٺuA�mñ��y.ɞpɴ g�WkΨ($E7�Y�oiuX�SU�(�L΅�A����@�	��S�y ~@ ����A�-b�t��i����-*2�l�(�\~�ScoCC�@ɭ����:S�D�ޖ �?C�"Xg%��s)���N��״s8��F�1ƒ�k@룏�R��P�	�r�zv� �l�5��6���+�s�F�I�3z昷�=���ЗU>8B����ք��D�s�J�<�6�Y6�"�>f��:|6[n�N0OK0�}!Яy�.��M�CR�ⷎߞ3�up]���pf0n#0ܮ�D�g+�-B��`��D�%�O����Od�94!Ǭ��M*�!�>u�������|��r��PX��dz�ʖ����7��&'�)��>#D��a)�O<C_)7�gknw�����n�5���|�������.I��b����K�^��v:��l9�B�G��u����~.ᰠ�ͺ\��T��׋�?w�2`@�*�� ��y�g!��2���+f��`~ڠ��/ȍ��a*��r9s�SLj#��H9,�&8�
��s.�tQ�9X�oi������4�o��wH���*����w��B�[t9H&��� *[*�"S� Vh ����bS����2��0��A%����yǍ���X<��at�t��p�{I�������|��5�����g���硼6�@G��(=��?!�蛤�����5�@4	����*'�W��8�wg���dI��n��������?;[^�k�*}ߨ��$'���V+���I�OYxus7(R9Pk)Q #�Js(k1Ĝx^͂�%��:��a�~�j�ɂ���$�!or�B �U��`�-ē���*��!�VZ��y�38f���6i������2��@�;sR̛��0�8�*�qc��5$�c�*Mnvf��B+� ���#)�B`cq�vaL+��!���6=�z�e�y��|�����ҘA��ίrd�1�/����␶n�G��ٔ0�v@�JD�q1�X�	S���6�]ۄ�c���ϙ��^'���;�RH'���p}ic��Ӭqw�'Q��nӣ-Vy���
�d�$UT
�����̘z^{-|ZŸ��X%���'���c��1���iH��3@�����w���OѨ��Q-,��Qh���l��N C��x:�D���:98�	��'m��L��3�YH��h�1с"5$�d<^]��ݎ�͏�|$��b%ZV����5rq�(�9 �t N��1'J���X�˻�tŚ��.[4�7I�������4��CE�/7i�R9��F��{�ٰ+��0��]�te�c	�z=�e�V�%��CXB'�qOG��	 ,3osYr�mJ(��o
O�D����׊V7�P�d*w�^�Z.J!���C|w4m�nE�2�������=h���� �C�17��Ҫ���d��T�{�(�sg��a���&���K����,�TǪJ�NE�Ǔ!S�� @����w��VQŠ˰S?��nC�X�<h�sd��(5C"���ZL�����`�bc���E^.)y#� ����e�����묑3�i�s�A���G�XNH磯�Ӆ��Ih��~=�,�o3BD]A�����ɑ��a��7>+s��@�����썀[u=�nY�&ț�n�������BH廲
o�)��,Zbf�w��&��L=� �㡍ل^dŵ�e3�3JPm7J�'W�K� ێ(�b�z��p{������b�2��7����2r�K%�{|��q�O[q��I��E}Y�ఊ''9ʔc���]t����L����r%Y��^>��h��6H	�F:�9�����I�}���Dg~h�aoO�v��eGe(Ӊb}�+M1�M�<��]"|{0f���Yt}���@D�$����SL�%�TzKxA��eG��l�j�B��=+����\��1q�0���hn��)?ד��?y"Q���}G{��Y��V'|����f���� ���H^E�2Ǐ��l��F��6��+�D���0�e�5�D;E�j��k�
�.q�؏���Ɔ�Q���^�YP�����n�4@�� �y1{��on:
�ǃ��~q�������'���iW�M���E�,��G2�!6ê�6�!cg}�1(BC{����M��� ���}��7X�����g�0���|������5�GEQ| O�}�'�=�a��[����쮢%���B"V�4�l}�f6�-��>i:�_���0m��]�d��#X�YCŬD�ٿ�\.#7�o/7�'��d�F��-�Ӫ����ӯ��^���,j�S�VI�����1�"���<;P�H� A������,� 1_f�C��3]�;c�$�A`B�)�|u
nFyE����j�]BQ9:�1`]d+��*gt��c��=-+:�Dǚ�][��m�_y�������t��˛��K�q��Lw�Aή��@�.��Aۏ@�u^��Gɵ����q3Q���
�1I�%A�`cJ#��ڢn��CXH�&5��@��N���cl,��"�gf�6e�=��諅\���s&>kr>q�!*&��T��=���Ӄz��Uctq�d�qy:�o�9>�C�/~�Y��K簁:o=��ƉW���Y��JyU�vD�C�)(o�,�\�[����.7'~��4i�qUQ�t]��_�.�]��R���-*�7�	��?��[Z����y&�PΎ���%Ȅ
u�sw�����7h1�%�W5Jԑ��p�͂D(�\�!�J�j��M#2Y)�[���c�2GЙ�����rC��s��[힭@1˵`�]�G�$�?zj�� K�=�{#���A�X��ٶ������>�7�Md��6���{)+�T�l��YmǦ���b���cR�.�>j�.S�Y߈�rv?�·L~�$ȌW��i��q⸷�M]5Wsp �Շ�����I�O�b�PfO;���$wȁ�<�>��]	�ӵ�<F��X~[�;�2R�[%Nc��M���/Hf�sh=�,j�,w���޲^��l����&���e=�����!5r+��v�x�	R�4/�� ��5ܙ��^�����("q�˹T��*���6:d2w;>d�'���������g����*��+U^�r�c�����F/ ��lP%���E�O)MOM�Q"�-��2C�OG�|�,���
>�*�lr1�����H����z�W4�ANVS0B��dY�䄸Z�N��� y������yRq��5�cx�=j�s<���#����t[���6�㦷�v'�ӣ@q�I�Eϊ"tBXI��]�w0`�u$�`N����0�?�� ��4�Z��Dʶ������$�.G��XDQ�+,!�;��Z�Z�%�i~]J}~���&%�/�4<*��;n�c��b� %�lm�נ�c:<GD8������a���	�%z#��7�sZ��Ϟ�.
ر���8��&��5���`x�� ���r�W��FIU�<i4�@O.�o�}��.��g������?YrƯ�G�X��5�䫭��"+Wo+���W�h��8�&/����)���,ϼ��\p/9�p_��}O����x��{*ݯ ز����;¡�D�/(Ʒǚ��X��{]E�uJHY����`��Utf 3��ćȘz���Nx�ހ�P5
.V��Qa�����FM��b�o��;�l<��g����'D���H.!���=[Qo�Ғ��_>�l�Pĸ�Kp�����=gQ� s�(��Q�E�K7h�;�f�Y*<Z��kp�,�n��:����s�-ධk��`�^��鋇�Iu^f��A���r�ˉX-��j�C��j�~���Uf{�����i�\����u��L��O���ܒmb{'���]ȹ*�ʋ�-�Ƹ{v+44t2�	���f =A���U?���=�����;o;���B�M��.B�0ݭU�}�X쵔~��[���;���7W�yj�Ϝ��s
P��m���(�fs�i��eq���qP}����w��y��C&+�|3O�$�%�ϥDי;>����qq�X��Ego�:�/�0�Ƹ=/�t'?}���e�zWjrIG�@���u��cl��)J�<�"e/�vo���GP��V�#w<�	�\��'��"-ʌ;wM���"lg�7� .�%I��
>���+���N�D�	���B��w���=�Wt�gGݶ� J���� i��-��[)U͹vl!�ߕ���vPċlE���ɪ�����c!|xI��S��@"Xy"�d�~��Bߍ7�����B}�U.&�/p�E�Qz��Ŀ1�\�t=��c��\n+�fw5mE�*jj��ڵ���D�g�݋�0b5�r˱ˮ����	{Y�?���{+
�S����36��Cf��CĴ���R�Y7��u.� ����X�L��Ac��2��3�V5p��LY'L*�D�b��Nř������)��L6�a��|�@�D}���e�x�!�������o�2?��aV�V�˔�]�㊈�18�$��F�c񰮫7�l�>�ĺ=���)��	L	'�O�]h���-��w��0%�#���bĺ�Ң< �i�B��8X�6�58���2�u�s�6B����V(��JF��{�\�C��`��'�ES��F���p�F��@%���c_x"D��q�A��8>�<ut}�ri�`���%}��B������ЈY�1������w�̱q'�����(���0�14W��B$b���Xa6��� Zkw#��ܩ:��h�_PB&��@a���ds
�d�}�)H"��_;0K��p�D����Q7�L�2<���i!�o)�ֳ���t�[�=s �]���b|8 ,�a?1{�K'?hψ�^P�2{ro�2n�d�Twl?�ĵ��VN�q�� ��Y�����z>L5���m��>OOY-xV�{ף��ě&5��e�z��-R�5��ܥ�u:!����K�7��B#gAS�w�B�xT�ܡ^��������[�JښZd���Բ�{,�=,�4T����u��2��3�>��|��z��A)fM�����%��N���z��[����B��D&��M곗HJR2��y~}�)�xo� ��i`�c�Fr��$��r+�	����z�/�.)gU޾��B��c�wn�o����SҒ�BE[uVӅ�(Ec���?�!��=K�����ν�
Po゘�\�QI��Z"���LI}�M3�3F?S���\���Ȏ䊥�5G�E<���	�[��Qv|��ͺ0���Ĥ*P� ���]��u��93X��Ѧ˙�oQ&��!�k��p%%n�b��Z�w�q�%;�Q�,ȹD_KJJ"� 't�X�.wq9M���	�|!�?�le�#��p��:�6}�l�3,Q�"Q&�\����vb��F��FeI�&%��)��.r�;&sԚ��-OKF�ƅm_�mܯwM��H������Q:����$AJ�6HZ���𿍅$r-/���P���)Pj;m��� �H�Ns+pE,DS��	��ᅵ9�~vR6�0���T 
F����t������x$Y��"<#F�T�MZT���vO������D��?��'�mP�4���Y mv�����nh`��׊���Ϡ%C�#f;���j�u��z�
+�*�T���������F*�"���I�<[�T<{X �Y8�h.�AV�c�P�ëY�q�³�E�&Aa�"%�G [��C�-�a��^�1�t����bz39=Ⲡ����*��v�նk�J=i�
��ο~vh�e]+�����L6����b���:������uֻ�@��s�0G�(e�6�r�yz4'�ėpJ�x�<k�z<|��}��	ɣ��s�_��.��yv���L8K����R|�0��G���̯�D^���#*��u��]9�R,�h��+�+�^s��)ӟ��L������	�].K14� C�w9��(��Y�o_tРO�^\7�迱=�(�V��x1�v;$D�ib�O	�68�A��h�W�H�I ` �KJ!�HC��0R����E�S�:K����ps���$m��0�ʢ v3d�� ����#�7�$j�`(��k ��uգ3��N���+U�댸h�0D 7�TE尦��2���/����k߇�i���ZG*��y� ���aNs�%����o� �t�s�f��I �Ô�Η�,�e�Y^�]]�{����pxqX+#�Ӱ���at�EIj��<̛��\��X���$<5+"t+=����U�6k6:��f�-!�*���pE��"#�m��~�� `��2n�(�OAڪ�Fŷi�?vH��W���6���#AU%�M�P��'ު���^��=q�\,`VO�% nxf�0EN��[\��)�������`�ǽ��x�vj2M�����>��jl��̹�O9�<��!^�g����\�xK�)����l���#ݻw�&��{RNsS���la�R[���C0v1i��{��!���I�� q����4��j���� �]�2L6t��Ӄ�.	>f��GH��2��<�^��ܸ�6 n� 2!�t N݀��ܫ�XtV�/�ic��jRK����Ym �Nd�9Ш��X�g�wP�Y��E�?�(Z�5����lӁt�e��.�,d��o��@��36S�x'��öHaf	;���O�k�ҽ:5=��{뒗��>xe�xoʹGV��j<b�s�׉/v|��#���4���e�w�� ����=��L�G�k�CDڪ�jj�Y6�җU���v��C�1wM ��^ ���"�
8,
��-�u= �4mV�����VF��T��8��v�S]�fx���2g#"M���:��|Y5��z�z�4Zʜ�8`#B�JW��U�p�����5������>��Z}L?�������k���
��
-���ȫ��[Cμ:/:8;��f�[,�l6T�����6�O� ��:�d�0��}2~gGjB�}^� ��}�@���U`P�U0�t\B��"&�JE�vYXaԘ��P�(�C� K��������㥖Z��GܾZ��X�S��ᡠ�X�oK|5M�="�篙�Q`x��v}okD�g��My\^�t�$�����ˎU���@K�`zBHTTد���W�F��Ђr���S�^�xȫ�s����/�����d����O���o\ ��ޖl(�u�^�Ż'�(�]�WQ��at2�Gz{5n�C
���fzu�0�M��~Sҭ浛��+��$���a6��U�s �`OYךӐ��h�3�����iX��坠���x7�l+P�T.��
�dHh@�
�o�W�k/�Jd[��çV�l&�D�������[�c�zɓ��E�sy�!��I*8Vȕ �F(ŕB�h��T �����D�J�K*T\�� X�Z0wKT���!�FS�9ϰ=� yV0�&2���`���ʵ�D�*�P��F��(}��L�"u�95��^r�k�Q>A�.y	ez�yQ��]����b��h�2�ψ �@�E��v6�!S'+r�C,FM�?�/���UZ��,��p⣦@�;����wK3;��s]�^sj;��&5S	�8�E
�V��?�{������,���K�k��K���.ܼ�BЗ���x���zc�a?�;LӚ��'WƲ�{��N",���}���ѳ=*�!��<4.$O����H�= � �7Sq�[L�Z�ۙ�h�D�ܵ��N�a8��̃m����81��FY�����q�"<�9v|��#�e0|����c7�u'U�6��	��U.���ȏ��3j�'&:�>.�{���
ž[�[Um�z^=�ZG{1�8���c#(ź�(]���ݡ��)�v=?_I�!L=�XYqF=a����/k���#��N>�g�EZ2W��ޕ|�=_�qΦ��_7T�������k���	֡ԋ?�9���8�r�t��"�O��o�+�c���B�asP..Q?��bC'Nz4v@�Z���P:��l: 了|~?�2`�j�377�R)�r%�$�3J�x'�d�<�����3F�*+��UD���RS�߂%X��aU�K��aQ�"-�Q��MW������A޼��0�٥��gt4����q��2BgbtP���H�]�f��)�5�J�?�d�++������#(�A����N3gA>��nA�1�D`t����(�����u�>�)i'P�Q��a�X[F0I�s��<��V������z�c2M�`%lq�T/�V������ޘ�D��R���Ĭx��.~�nE砻�E��`���?.��FT,��Q���x�Ȼ�s�/��z��MV��E��O8�!���b�����3�I"�W;D:?ě �*��a�}bL�?�5��)J�F�BK
d����%�&~ݪx�+P��!k�L���O,:��U���k�i�$��$Z��Z9���C��bOb�����cFt�]B�o:"��$�Y�βښS������C3b��n��A�a���bOyz��S��WE�QS��$,>����~��ٓ�Z8I�����ѽ�ǒX.9�O,�}�z��c��=b�B���ˏ &����Q/�F\����N������4`Hn�-
h����SF���6�}�r�O���%�&��w�ܧe�G�"9�{ ��>�F*�V&~T�8 ��9R����>�K��D����p��ť��kM9��Q� �6H8n�(�*�c��[�I��+Ԗ�������'�m�������>�4-4�/Sl��s�(f9���t����MRP�����NX��x~kfv�Jc0��SD;�:�ˊ��6���B�LbEyES�d��A:�dv�Ċ盨?��&��nrK�+r�����fX]��'ٜƷbpt1�3B���\�~m��e�]�nۜ��c���cJ�_��j�������q���\e�6}G����0�~T�PT��+
Ey��B����f��Ѓ4�m�J�9""~7z�W�@d��H�m{��}'rOj9&�l~qM����[�����B<Z�Y��ٜ���F3:��		A��]dLMEr�^5g��Y��n������U�2l|a�Z�@���P�J��TM���;Ur�,�t���輷B�)�5�_]&5��YXy��\~�Ey�<6��j�:ݞn�w�@~l�{�zB�͝K7�߰o���P�ײ5�Z��-M���-n��0�#&"֕�_K��w��ng���K������ ��p	)��T�y�V{B��&��G>�A�O�����o����Dw�ْ^=q߸�Y)�r��ԣ89:3�7�s�Rkm&���Y�t��0E55�qApr(�>��G�)'<���[�&�bz�Sv��)��k]��OK�L��m�B�O�u�ʝM�!II���z��U�lĀu���f`/�U��ԫ�]ᄐ@�){F���R�K��vj��Ajw~�*[*�JuԒ�����)�-󾠻�s�Z]�0�r�(�W�|z�������ݠ�ʕ�C=$^���iѴ=��:�Lg��z�Y�ihw���~��]�d�kgb�&Lz惰�����(�/�EC��W@�=>Y�)h��� 	��V%�f;]b�"z[ӷe��yu+[����$�J'g��7'�;��A�+����Yc��u0����CX������c��X�HG/� A��n��A/�U�0e�e��xqI��f8��Y|���z����b��I����Z��۟fN���3�&!���ɴܨ���&7���k�{C�Dbz��H��f��&t�;�m�n;�����\�κ�x4�R�5�B�Z@���� �A�F�_���Z�� ���݋����h�J��26&�$Y'B;�	W�J������\q�8ݥ�R�v	����G�.��w���x�;�"/����\��Fsƫҏ�12Qŕ����W�ʌ�ou�����f�vE�u!Qר�t����t���.�"�a���*�-��QQ�W� ��ab��'6�#�����03q΋�3�Dinٸ���]��ܗ�t�� .M)����������Z%�m��"J�aI5hH���4/
OqO�0s{�f�_I�Sd[�	�u(��Y�J�&˯l�����w(����|]������t6�M�j�<a%X�/��!LJ�7����+��M�i4w,�g�w�5ݜ���3���R��u�g��Cu\�Ņ7��+%�܁"��d������L��T��)u> *����R��`��-5�>=�5�[NF��f�����΀����nZx��v>��kI/)3�0�����P�ì,��T%5x��k6�&d��M�U�
��d�Λ�����%ș�8Ɍ9s�ٌ5^�'?F˼�M:�:��<���v�pU�����.2�R�ի5j�5��׿�w��h&�g�D�f*)o݇��Sa�J#��S���|ӝUM�1jwXA�����t堈�U��O�t5�O�������{|ݩE��sJ��󺌏�R\��~Q���r�\]�4�	6 ����
�p��:kиF3e�<,ƞ+͒��#����3@�o��&�w�0t�Q��Z�]}r=�(��[(X%Z�huV�kB>�CK���\[:�X;���#Y�#\�1���֙�%����	�k@���'�n�&���$:v����f.�/��{\ÒB�+SUE{4���ك�B�	�t�q�N�����|��}G"�Z,G�ԼH�ۯ�]��'<mg�f�t�3��b���l��0�ӥhD�V,E?�A����#ѹߝ	<D�J�	�:��o%D���2E��������Ų*�y��%dV���`ÂnȺ\�Rn2a��3e��h@D��_��"�2��Li�+�'SBb�`7�ꮼ\��/����s��Yax�u4;c��A��`��YO@�N��4W�YP���=�::f�s{�:�c>��B�u*k�w ����%#����`�M�5F\a��1C����d��6���Hg�>c����5���f�~��F��ɧM��vI�ϛ|�m�"�<��g����kQ�sїGͫ�	N�!|�a��M�d������{;$�k��s3�k��>s[i4l�gzB{�:z�C�%=��ċ�p�Qr �|[��<6ev���Z�w�*- m�@�KM)���,~%�qA(A��'���b�� +i�I,��Sxo��'}��H�ط�]�����mV�)0�r�e�[BN�/�m�0S����k�$�{�q	���MK�F�)������g�r��6�Xx�)Q��� ���v!+>�;8�dM�����8� �|{N0P����U��PӬ�Obc������)��!��Z����]@�3[��d�θ+�=�&������Ξ ���� y�����Ӥ~k6PX�^��h_гE��Uģ�V@��L~�'K���!i^RIl��keL�,גl�4�8�����򖀇�%�߃��ep���YȱC�L���G��$D΃�Vw��u�{�i�*=�b�b���)=�dVɜ�q�'�HR�mi]��~���\~KC	Q�K�o/ ʁ"��e%U��$���᫭�7���_E���H���B.�f������ҵ�i��xE�,��:.��ۙ��l%�Y�V&�#�u�����#�MG�i(�k�>:��>E���>s?�:UМ]X���j�6�:p+gޚo���bi��Ƈ�lp͍�+����3A���\KXs�_�^��D/�b����Y��Z��`wE�Y�����~<T�p��#YƲ`f���veoҳTY!L4Pt�D3b�a�������
b�cC5��A�Q1���r���o�FƬ��n:a����S��	��a��ZD�`������>�Ό:�M�σ�t��3Q�x�~�@��l�8�������9�j��܇�ɋ2�P��G ^��ë�D�C8�B���Nu�di6�k��+��v[l5�t�+
9��1�AJ���7�_^=]�K��q�}X�ұ�)�,�Ȧ�R�$ϳ�H����<��e���v�(��H��	S�zU��P�u"$�Xa�9��5�bO���#��h�;C�����^9���e��Ϥ��P������*3a�SQ~F�ŤW1�=�M�"2w�9 FO۲��S%\Y�h:�����a,�F���<mC�z�$u�Ȱ���3o\�f{-��u����t��G����Qd����W�EE��~�X���9$xO�W M��ݐ4J�9#<;4N��iq�XlO�OjJ�S\��(��ydH`%sIB���^��T���h���O�vyG�-�83,��D�W!���#Z�s�3)��L�Ӑ���a���"�`ʕ�&­��^r����A�-�7]�fo�A���i�����= (9�Rf�O�w�V�T`�d���A�c��a��$P�����-PSK8��i$�j~���,��`ZU�}�bo�����i�^�'f����U���-�?���*8�q�#!�
֋B����W1�`�m����<�\{��!�����?��:ÿ5&	��hi`�Ut �}�5��=�h��t̗A����"N1 ��v0o�| p����(\)�*��Bd�+�0f��}U+N�O3��/۶D'��u�J�p���g�2�-�m��C�!�9Pu��<�$ݾ��Oq�hd��{4��n��־5Ի@S���n�P�>���%��Y�F;�F�tX��&}�U�������"�W>1��up��Y�����]}��/Ե3���'��n�$�W֕*�gQS�8���y�B(W��I�.��S�*��,��tq�:-��#q����T��8c	�\���L�xe~��f��`�7&���9����^�b��.6]�n�T\r��
K��R�Z�J�Q�-���;����+6��b�7�r�����H�Z$�B�%����g��k	��F2[<T����OCt����z
�Z�r��n/`�fz�#�ݤ�gS̞�2-���Y/�	�̘��?�L� ��|��2�V��x��X�2c�՛��H�׉�~����*\\�_��5/Ɔ�p�u�X"�|��Pz��&�K`�tC�q?��&�s��ݩ��O�js���ۆ����WPi5��S�lI��8�G=��)��_?݈��'�.e�K�q�	)�b�t=�.��A1�����WA�k���a�:�q%z����S!q�C���M�(�q�Xsa�EÐ���X��,��������>F���
-ţ�CZz��S�P��z�rR�=`���DI�7$�`J5ޓ�%1[�T�	�p[�}H]�x�<i��w�~6��L��k�*�)��\$v.m#01)�Z�����|���V,7���eF����o�FyRVv��`��)�"��9@:��fjvV��LuF�W>��Ǵ���>�ǋ�(U���vgV����R^P8�����1˴9��glfu�\�%�}�}z�LQ5܆�Q�Yo؉v{�E��#������ń��}p�$vD����~́�Ш��9����?)&6�|)�g"�����2|?i�hrC�L-���@�c>�h�ڜ+���U��L4;�S�/?��g��\�������"-1\j&d�{��c�	���u������c#���O�I�V\E:�ƞD�� x���@��gPp[�����~Zp�1N�\�hE���6��L�Z�IM`k&����k`����4$�?O�����l�up���=Fy]a�ܡ�H$�Ϝ"�F������5r�3dF+�����x�p.��`���s�keLD��h�^^��փ������C���{�('�\:j5������<ewm�T�Cgy�~H�����]o�}Z�wF��9����j	��f�9�Ӧ6�
U�0.׹X��"�x�#,`HgD/��?��&�iD�����tbm����
��|�qt�M��w~�3�#�[ÔQEYr��P�b^^�.$�B>�*�7tamTd7���q��2?�������w_�C�������;N0yo��|��:���wn��(�Yì�׊�<UI!ܦ����ƈ?�&�{��4�5�z�Z{�yc����8=2_�f�_m)1r��m��0P��Y�i���a:�zfj
��[���XS_�9�ȷ���WJ�_8$Du��<WD���X���!��5�����B~�bF�2q�(u_��~\�q��hx1Y�K���d,=0�N,m�Y:�|W�c�hT#�l ։̐o���`��oe�r�l�H�uԐ��VHadx�i���{���6˚	n��Y.��SO	���ס=p����!̬s��@��_ƍ�J���;�%�s�dv�����\Zp/&H�cZ����Zvuh�1�[?y
��{p����Pw�ྑ�َ�* ��T{@��c�2�v�	n�o����X��|��� �+�-~pk٥���k�k�)P�
ۯ�A��?�Z:}���%M��^ֲ1��<�02h_�.�"2}�D���|F����	;�%�lYh���E1%��gVR|�J�.�xBVΔlh�,Q��&����Dy��i]�U4��Q���"���[��X��>i�N��=
���x<T]ű���;�8�=��8�>Z����6H�V���������&Պx_��A��bo���'�L.5�<��A	F��01a��9 NiAE��\>xrT$��R<��q�V3�v{@"$+s!�,�5SJN�nh�b � K��}�����f�'f^(�Bʦ,�F��?�9z0l��G���Si��)��%٣���|�AC���~�_}`<
[GYն��ѯ���!ǝ�l�Ʒ8�W~�j��������%�N᙭�E�z*�?9N}iW�?�ȫ �>�EX�:�#�&��ν6���AE�H�-]�h�Ð;��D��x��/\ְ�������+�,-nB�����{�a�~��BCx�HPD�^��Q���N������v�nM1Hc	�������q����R-��|����L:(��$�eX?�=�H�J��@��tf��K��dY-�vD!�4���~ѹ�
��N`= W[J�)����c��T�5�����!nRٹ��8>�^����J�@8H��@�Τ`y�Z�K�Gx{[�B��i�[�3�jQz�!��YTY��8*@55�;�Z����p��F�$k��>.�	���J�mB�V{��q[�_�J����o#�ڑ��7��D�je��~���e�V<Vn�Ş|���R��g��64�AY��RA�	����
b�@�̞���c������d�N����H�� �*�j5�@mN�1�E#���k��Zӏ]����]���^�� ���&X3.��p�`���0q؁s�N� �'�c`ζ́Rf����
�l�/f���+�>�O�Ģ� �=_��E}�8��L�*�����I�e��)c*d�%��ʹ�mt�'B��x���ȇnޛW��P��e�;�#K���>��ƕ�w�L���L�6��ӻ���Ǥ���1��siq�g�>����9vl�k�ܬC1�eC+#��DS�_���a���E��Ⱥ�dr�>����}}b��
��>��(��cn���x��K
I���a��*����{�$#�X1��j��Ie��k�5��TÞ������y�Ztn���4ΐڙ_�{����j��vRX���SZJ&ڧ9��M��=1���br>���=���]?�;`�T_��Fs�]f�#ȥq�p�N3���l�q�Y[K�����O3�UN�|S�;K�AF��'�t|'8��8�%�X'O���}���z:֠��1���{��`��o�@U9}�����ʄ�7Y���?C?$��^���L��RH�UX*B�Z��)oX�9��QZU��)+�*����2ב�Z'b�ĩoƮ���;(�R�����zIǊ�0��8����76bE�}��)���O8��~���r���aM��q�{y�*�*��*��ȟ��&��)�]���{��N_z�gMWc
�Y����,І�AG�'��˅{Բi~L��+���3cI�.�2Y٢*e	fI�dfJ�v$£v�Í^��Sa^�\�[Y�^�P�s�����^���섬�����6��`�;1���aҐS�I��EU�1�l{�}��2��-��/��е�%��~�~4͞9�$T�N�@���c�P��K�۷�ޙZ����-�G�^Cd-pm:��o@z��Θ*����� �^wT��/?�b�Se�E2`�F5��@(2S�p��t��^��� �s�,�b9����9���w����1�!���!�Σ�i̎��],�4e�3�>��BT�]��8����>٥^�>2b�#y�uݡ�t�U�4d�\@Z�����&��\���/F2���|՝����Z�| ��r����̭GO^#]�Ֆ	ba�}�?I��]]0_)��f�^� Ȧ� �,� ��>�Ixr���9�E�wY;�,��Ǌ\>�1P	݅߹Jj��7*�ӟ����T�?\�K�tG�r���SԽ�]�5�Y= *����O���c�����?���p��Jw��������Ѹ-B~�O�
����I�b��-'�����#>��T����`��}X�('�\*fr'���M��ŗn:{��A����_p���MS[$�Ew��D���L2�I8woз.�5�F��;f��s�H�����YS��m?�ݸ�'�PD
t/l��l�F�Z��/qM�B4݉�����a��L�u���M!����a[��G���~J\u%[�&B��,7!QZ�H��Ϟw��*��H���u�T���2�ú����	��UHB[ܹ�IL�_JT	K��b
�j�*���%~�ޡn�+W�2)�M,S
��jq'ڂw����yU�v��^tJ�nw��_�^���*9~�'����篚��4Ӵ=������E}�:�ei����1ʽ����p֢��+�8�F��5D�� �=!37� CqD���5�&Y��������g����R68�������7�_j{y?1��߰_'@5��cU�Pn�Ԃ����eׅ�3�s���l��? 7�X���g����\�O��D�w&�B{��o�+�b�A4b�FԤ�B{&.9[�.���Q�T��h���.QP�;��)������a���#�&��JM`w5��
m�9(z&���ꝰڅB��1����)�n7�Գ�����ӊ"]hP.�D��T���	'`��G�B�	���0��0�5}fC������P��~�9��zǊ�e $�����׈g�|�Ş1��Y
�w^0��/|ņ�X��]�
|/�WU�,�+���Yy�$�$��p��We��1�=�(���`!����%�Y����0d�B��`3�Y��5;b�r�~G,h���r oĚ⒫�1$؂��"���*6^-T�|�!��랁ڟJC�����`�L\
�8��H<���F�p�=,(&���Ik���լ�Y,��S�w��#d��c���OM��D�?��K��uU�\���@��\+�'��jܖ�m���҇��ۘ�+������ȡ��
�noĹM�J���h<���^&Ajb�C�q|$I�k�Q3:��ʡ�o�hԅVeuMB���[^:�2��\�[����r��O�+{�0�{�I�f79X�k�J[%�T���#�tUE{�-l@+fIΐ�rs�����A�&$�j�B$/����H��T<�Z�������.�VAy�en���W���������������\1d-d=S��݆��#�k�k���U�]�jӾ�t��>���;ȑ @������υ���S�X~�M��W���G�>s�kG��<WC��e��2j�1���������0&�����*=�`��0�9)�ؚDy�Rl�r�˙��X�W�j��w��Z�<I��ԋ/�q�3�vDAov�����Р�'o ��� н���*L��W������x�T�,���1����~���R4$]�:��2���<����T�'^�9�Y�p�m����>�
�VU�T	c=��_T���l�!m0q�u�{��.9�J �u�����o�C5�Isx�#�ր��ò����CYL9F�-�p�@ˈ nj���\1�l�oB��T{�O�K|T�I]7�7Xj=�-�B�[	���ǆ<��y�|N�S\���4���?�d�>m]��o�t
��u|��2��G ���¬ݬMY:����c�����f�O<~�6��W4[pf��u<W���٢*竿���~Z5����p�s;3�3�q$8�P��^���ǌo�ׅ�� ����Y+��mC�5�����mn������jw�w�U�����J��r�5�%�kL���^{4�v��	�*ܟ��|��͘&����Q>�֫��@YW�P��~An���6��E R�bfV�-�/U*FZ�����"ꡃgX�F�l������d�n��8�B�w5�cE_.���xwAPVj�/�3�IMv6Tܜ($�z�N��K3����1D��y$n�qt|�K(�����;z^�k[�XB6� ���C��K���+-�+���܅۸�j���ү6�Jr�?[�`0Q���sX�<Ή=fj�I�����cw^Jf�Uah�;��_��eD>�V;�<�f<t�{��cp��&Q��+;A���'�nޚ����9���uJ�ّ�u<����iZ�WU��!r��7Ÿ'�Z.#Ԟ�$���j|�>���_�A؏�Noh!:��@�g�9e����#ؓ�?&Dv����2n᷆U�E)�!Нt�.�#e�T��<��jӀ~�L�bC~�~ ���%Z9f6��8�@(~vk��{h^|$\��\�;[��X\#xvP���G��sP-��Ֆ��["�n飫�ub_wM��	���B���,3�>�W��T����;+�x��>�	]:�n�p�A�<�=�t��jpme!�-뽆�P���TOU%��f�\y�*�UV��'��&I	���8��`w�r	u]��Q��`�Ф�$XE]��0�ef	��pD �ZXp�+��:�Z��7��܃�;�~���
�������`��%޺Iڪ�ON�A��%N�T���_�'�"]E��c������[��������c�O��i�Y�ʬ��N@!$�|��)�$���.x~�z?+'�cu���6l�/���'.��׭-��~3��¶�n�S���JR�mпA÷}it��˛34_����?ZoD�������U3-e<��NC�� [�7��"���.����Klيt��D�N_��o�셆��Ko���Ԙt���%!�t$�܋�4q�G@�@�����0��?�fY�S�@,�,X��K\
��D+S�N��ٝ��#�x�J�*��-�_{� .i)
FzH���F!��u+٨��*F��gy`��[-:D��P�JLA��L�A(m���jb�L�C{xR�}�V��ВlFJ�);��M��-��>>6�x�l��* ��=�֪�v*��Z�|S�����@�Z���{41{kv[�R�>ei�|F
�y+9	P���:�8t^��2���T#�{��Ru�qAT��=����_$�s��c�����v*\J�q##%�|�#���R1�,٢��b��ý֗���0%*�RY4�!)P��3��]#|�z&UP�h���O�l`��W@C��N'm�_���|w��=|ϸ�f`��byӈ��Nf�`Iݚރ>��f�����=*E��}Ǭ5��e��s���c2����9S1rbg�Tk��BS�؁;������D���t��0��䧬0�0EW�j����l�7�F�=X��oL��09DN���(�}� ٸf�0P�� �r�������#i�E�&�YmԿ4_�����l���B��B�x1כ�O�v�
��A}���{~yE;���p�S�I�J���i�V����¿~��d_�����Q���Ѣ6^0.���cT��̯0�~p]"�2s�	�;
�h��36�4P[�V�q3�F,��S�?���י��42#�I���ԓ>ZM�1������\�U�_]�J�Q��e�6 R��5��q�#IS�<C ɲf���h8vt8��=�>j�؋f;g���O�����3p��~^PT�� HX!��ۊ:[���(�6��U�q����^����/��ɚ�)��pH9Y�H����s#Z*�*��j?�����jS z~,����� Q,��wnCX���LV�:�����)����7hv��%֥x�vSQ�r��٣pS#-��ey��8����;2B��6�B�i���3�a�▘ѣt<�}�[R��a���6�}�ف� x��ԅ �܎۵��E�Mg�#�}���.Er�U��0F�J3Y��E������R�w���:/�,���Ҹ:�ӭ��"O�s���D���
ת\~L֢D�B���$�g�>����<b��/��k�)�^���"qbfZ��f`j�Ax�O�;���Q��3p�ү����)! >��Tx�RCM�����醬�O��9,Ӽ�c\x�%R���ͭ?�(5i�;~�⤼V��C�Z�N��ާ}3exеC�<5A�H���1�,e�sN���Nx{@����P����'3��Q�_)G̘���g)����5r�[&@}Р����M�}�t��w>Hk�r�'b��D����,�i0��%3}�6��YE-�>�%$(��)K����N�� >~��s�C 2G�5 B��S���}),���p.�����Q��r�x�Yi_���2c��BJ��<��Q�u/#�'cIR��$�;WMxn�Ys����>�F��y	ȣ�1�oM�t-�j&�U��EG�̋�WA������ͺ�!D�P3��_]A�ￇ�"9��BrG�H�u�_
?렯��"o�#Q�t���坟�۪��tf)P��j�p#�a��z��q�H}�mX�<��`��R���S�%�^^��-��a`I��yX.�A7�^�'���_;�@�혩K�=�r^��|�G+-�j�r�ddЋ��<��yO�;�ž�0�B����R���ai�1<�طI���+������\��C���@�x���L���N��9�^�a��o��;�[>��
��7�&��677^�tMk^ �.�@��x�����z�5�Lv��=�4BT����(k���.�3o��)����`�Vw]���1š�N�����uc򶧲���8�OT5�;hT�Hi�5ف7ñG��shlcD�F��޲���z�����&���i߱�M�zD�Ԥ� � �sm����[���q�H����j[�fZ��h͏H"�_��N{e5�<�͗?�%Nv&���B*<6�A=|�z�0�D#��@-����M�[?>�  &Ź��'�ҡ4���(P"����?�-_���lm��l�`1�����wb4�|{��
š�"�'P���z�(�ȭH�؍�
��"p��]P4���� �78�T��c�?�t��N�wv���L'7�$w`�q1�<��M�v3�&z��[�A�S��o��\"\U�f�J�nKFjq� ��DG��rE n�M2)y�*�=���zA���Wd��i.y��Bu��5�뫨Zӈ�AXu��2��@��Δ�~ɚ�RNn=���x\����"䍶z=���ͮ�V��� �=(��q�j� �,^.!�� �N'y��Z�F���z��i�nF��-����i�N 	�(��I��8@�,O5�<�.n��g���f�*���T�v�g���<�A���e��SqI�W`vˣ�ysu��!��N<�Ӄx�� d��"��ZB��i����z����dm�!N�~
~��"�;G���V������)�5i��"��4�KNĪh®��+�*�Ӝ�D'��`�=�j�ԷaVx:6F-� kh�w��j��8!�K������x3�MBW3Go`y�U݄�:���ܠ���lH����Əz�d��2�T��c��q�K.�@����9�q>��m���n��7��
�t"Ń<�5����!,��3i o�ޖ!.�5N�xO�g05A�R�r;^v�z�Ս:��q#֘��1V-�+����_h9!�G��)��ɇ�P�Uw�t������9�"��&6�$�6���};���]C{ʢ��n�K��:�LJ�z_��+���P��.�`�+�qG����p�:���\��&�;)Yͥvz/�q*SR�,�.j��o���Y!��R����x�/|�Dݤ)� ?��ae�����,T�x��[��]�E읠�7 r�����l*�� q�^�T���c���5k�Ћ�6j�[��a�T��3J�1�*�U�1�r,��d�j�}%G�&��.�J٩����Ĝ1�r0�k�z#�A� Q�cN�4��i�p}�9^��n�nT���'0��g���,��S�G�N��N�;p嶧|)>+T@2�s�V��2��=*��@�0�T��f��Q�L�����`e�e.��5ҟ�y{X���qt�v�{�j�j�!�Q�RΞb��;�Le5!/1��F�½�ED`=�Q�d(ع�'�R%�L5�0�zEڽ��zop��uzla�$��g��Rm�z�C�����t|��q�{<]UaJg=i�Ǖy���
{cԈ�"��m�B�����.0��IkSH���{D(�0������B��BRyS���g�e�
�:��G�0�����P�V�U �Ǔ�|�w�CJY���P[�ݟn��1,���WR�w3e^��K^h����
��ʔ��(�\Hz*��H�0�FN��~FC�Z_4;�o�=_�ޖ�v=� >4�l�
5�Sfj�w�o&����>(�9;\�LU-r5#p�u�cw,Qa���h���w�z�W�9�W��?l�Q�Ra(?����)@�r���W�H91�>R5�Y8���XC)�����X�2����],��+/uZ������κ�ngٕ��w����W�p��Z��G~���	�)n��ܔB@�%S���f�����2�9��/�������W��&2J�"1�#���Q��~EA�0��>tD�������|������	`_���G^��<�S�����y;6�Ǚ)����2BaT�3~U&���H=���i��g�A�^��� ��N\d���8�h�D�wݖmA�z�Cdڙ��jC�����s5OO�b2�������t��n'�����g�5<0�Ȟ�PW�"O5�a����fkh�0i��D4�K��S�v�� m�g�v����m��Ԡ���g�t���y	���e��R5$}6��������:� %*�J��|���ޯ4��o �'�L�0q���V�1/(Sq���T��l@��U�����r�$�Qڣ�Y�y8�u��3���	{�ϖ&SL�J}U�Q~Hׁ�S���bgu��N��k�|�Ųr z�B��m��>�����YW��8�s[�e� �O���z �	��ؐF�hF DG�}��z��-� -�ȣ��0Y��B#�m82K�F	!������=>�;���Ò��R��.aD����r��M�[x�n)���-y���pάG���\�K����Uop=j�5��2��_�ߓ�#`ߦ;7g�1�-Ia�L��dHE9��u����'y>QP����I3"�/ �s�]ϡ�mGt���� ձ��{�'�P�:��2=�&QY��6	W��d�ki"p��%d��t�>���|�������u���,��	:}��-3�b��*K�����A;�ߵ�LJ�����p�`ٶ��=����x� e��TcN�*�=E�<�����*tɷn�&���x\�����/��+�r��.�r�ӟ;�@�������x�WK״]���B�Y��t�Z&��r�m�i�U�:w��~08�(w����&��um�yk،�΀HR�{g�DҚ�3Uڭ�t��vx`c� Y��y��3�|��:��e�.�ړ�}+���Iؔ�w�27�]�f#s�m+���('
�Ve]�n��F�0mO ��$�w�u�7Eu��3:�<��Hg=RfM�����FؔB�L��b[ ��T/n��g]� �]�G�<1SD~�UG�)����.���sf'�bi*U��4�;�~�����s���HIp��g�|J���qH&=+�aH44�f�b��:9�������{��$ʣ"3�C�-�C�c�*�z�'x������{^K�pUN���z]��(��&S������� ��2��2�����C'ʞA�̹9����������Q�	nA)v~�C)��20���`�3{�i�D1Ö"В&5i���`x�2Z����ڄ�o=��L��ǔ���]�ߘx��v���0��*��+�'�9^�0T|,�t�R^X��W.���VE�o1��/>jr�Pfw7���ā�x�'I�!D��'#�YB>|�7��?"�m��{U��HEF@&u�O*}WJ7)ؠB�۹9�rm8s5�2�B�q qΆ�垥�!���0�Z�}I�/������Ɉ�;i�e�O���4�H��Ti�� 67>�;���{�vmv�Fm��C��΅�S^���ᗚ��kz|�:b��fZME��3sG�<�S�+�:44ڸ�!��
o2b�.B�[�U�0�Zj���wՎ���8ĕ�:�ؘ�z#aʜ�4��GT/�8�n{Cڞ�MK(r�Dy�iT�(_/=jZb�Nhȧ���*\8��2��*M)	S`��Ok{V\�n̒j�k���W�[�[?�x�'�?���)����*ӊs\�	��"	�c��	|z�[*�l�N��*��G��DrԕZ�������t�m�0��)'9&����d�|��@&��5�c��������<�P����c�~@�8)����c%z�
�)�.y�x J+��Ds>a����fYi�A^_���g�g�m�c.Z�6ZD�1��1��_h�J压��\����#4n[q���X�n~�Y�s8�l�ZF�����&�06��܇�j�l#�'�!��9�̌9����P��ν���l�f	���/�CQ������0;��y�
.�Uf����V�4&<��l�`f�����~1/'s�}g{f~��/�d`f+?C��Օ����K�z&.s�`�T��i�bCa�����Z�Q}u-k��������H���L#��-�h�S��(J��>gf{	̤�WhX����G0��EPA��Y���n��2%҈��Zv-v�7e��+(�0���ո����?�^�/�1�� DE��+qs�Y��yA�F��]��Gd!��cZ�θTDli��e*F�^칤Yi���\�#<����d�7�����'�^5F����Kڌ"����3Ĝ���F1�����}���Ig��.J�p���f�D':��.	�&5\jL<<� ���srڧ$͸�','��~sKo1���%8}���fX����]� �qR.TK^�j�76�c�Ay����o#��� �R��M&wÉ�G�����a9�;��j3'�;S�j������S\�;�������hX��LQf��Ga��/ ���o1脄��\��0e�v4YXO#q_&��g/�v�O����t���܃��\�=����?��o4,�8�K�eD�A(����qT�9�!��5�e�{����7�/E�y�B�� ��c�iC���������(}�
ٔ��v�d�HTJ2��q�b�f�Y���(�E�z��Õ�&9�,|KyG�*Y��ѐM�����ϵ}�e�Lw,!K��a;��v���XGyِ��1`�%
/�ML��7��V���I��C@�Y]D�`	F�'�@�1���!������B��Ij������N�4fpTM�1^�+�E����=��!�o����=#����=M�f1�~�J���q>>��J�D�̲I=���)tNX^��4�"<�����l��`�/ȴB{��X�_��:O�q�k<�z�׹��J���>���L�-�p�eg&�(���n �'o3��МG�������耪�������i��Ee�E$q�k�\+�,��G�L~>�t�,؋r�γ
{䧚�����,��2�t��Kv6�<�<f;�lJ��0�Of$�Rhu3����!�&[*�{�� �AG�	�PI�7�37�����c���ii�L�^��,P�����R���"��