��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\����q�?��e�I8�b�Ǽ$��"����ׯ1�V0���g�~����ⰼ����I�u_��M`��}�u��̩a�}���1"�Cd��G}��n��"�9�|;��W�[�+�k)̤cG�A�<VѨ��f0���i�'��k���?����z�irqC��R���V�)��m*�f������T�o��<A��.�G@���B,��@��+�Nc�0VCy�T��sӻ�����_��?b,@s2�/Z,���R}�}w���5?�d��a�%xg8���C?4���zAZ~�`��h���&���"4�I�_/��c�Ck�s���`�0񞝍�+�⚝��u���
�U]��O�Z48X[5Nz�K�--���Zo%c<�ӹ�so=�׹Pu#� ���O Ԉ�Փ�6��ې� ʎ�r'��u���P�]
n��A�53'�^h���kuj����l��@FV'��Sh6���-S�1/��s�ϩ�B7U��]��lw���%��J����P�92?e��^HE#<\�d�Ј~��{�Ʋ_�]�`��hK$��Ӎ���*<��!Z��ںa9�*9��|����;�ڟ���Yi�AQ�/���0J�An�"��AK��ad���3��=Y��� ��X��!U����8��7rＦ��K�q�KkvU�~��ޙ7+H`%�d�t���dQ���մ��Ɓ} �:���]�cH��mj�Of�OM9��.�^D�u���o�W;N���+�`�0L_US����̯(,��V������%^��r�&������a	I��X]_��#���ƻr����5���y�V��W���c;v�9?�*�5¹\�*��^��
'��Ff��Z�B�\��g�fҎ9��m�a�RR����v-4d�Zq�i�}��f�W��Lj�ѱ�e=Pv�n�G� �9u=���K����X���)�ؠ\fs+]J��a�j]���'.л���(��X� $؟�ݤ;�~Y�z�����_נ6A��G�|$�T�N��׿��~ 8zn��`�c�!2+)��2H~ˇa	k;b��mV��4��9�"��,E�m��&���p�^��g�%_iB��h�(��B�St/��=aGU/�����
$qZ~�G�£*g񻏀�2�p۪�;&h���ƥ�9�9Ը���,IG�B��2��ˊТ�g����7"s����uG �4�v��d����f�	]Sj���
��de(��R�)��D�fM���4c!�@�U{T��!w��9 P��C��HT�� Iߊ/�
dO�@9}�iÞ%���j<�G��ę�SX��޾F���:/�5ZUxu(V���IM�z�E�D�)�T�n�����l˫�	?��^.#78R�.Y��R����������4%�N�S�t�S:J�����R�m��߫O��y�$���g��#��'�
37�Dz�M�;�kO�j/-����[�Fel�p����%�9�����YKipwK �C��-�#\����eU�v��h������ +���4{���+�	 �p�o'ƌr ��2)9�}�S