��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@���$U[H_#�/8�y��,��F��`G�m6f�f�aiI`������tC����dl���=eZ��^�٭����B�FYĸX�G�����݁�]}~�s�cC�_�V?o6���p!��#��9~̢z�x	����M�8�DӅ>q 6��n��  �	���Oi����P�ª�ج�9���Q3��eS�&�ʟ۹����:�V�ۂZ/'m}�Dv�Cf��)B
�n�ݘ�I`���e,����i�����r���+=���%{��V�ݴ����{��L�����3,{���<�@�3��N�0X )b�t��~����=����y��(�l\�m\���?��B�*"Rߎ�R�ʃ��t�6
dw=y`j�2�e��J������^��ò��-ƀ˘��yqXy��1Ȓ��h*�׈��.�T	森�y% \PU�*AH��i����Q��w�YH�#�k:����db�s叢]����8�Q�
���d]�5�h�Vr�(��C�c���¸޽`f���Y���#�:D?��.Ĥ_��5c����D�Q�{\l�M3�r�������
n��b�������6AZ3���r���%���Ly����7?i4p@�tƛW "�o`α����n0��dv�qnh9!��П4��[� k:{��ERS4�ۇ1"5�E:ԄxDL��AFqDu ��b��e���6ϛn�?;$�=_�t�s�RL8��""#�Z=vv|�g�t�嗻CYY���m�n���
����|�E}������aS0"d��*�q��h��a�9��Xy��1uY-6��Af�����F_���Ԩ��|�Ч���_�y��\ g��H(����|�&�D��F���Vv��&Y�kP;T�7چ>�tH�w[���W|��5u�S�p��[
�>���B ��{�t� и~h�j,^@0��Ƙ���(6�ɉw�ި�Q�D�je������g�����M��i �©K3��䜕��1�S(�_?���Dk&Ϫ_b}ܩa�r��7�xNz�7'�:�����s�����&�L����R� ��u�Ϳ��ݡzPҽ�&�x�����.,l���	=�3�ԛ�� e"tx�>y"lC��8TWL4T�@���璘��@��	����A�J�;�yz��>�H��>F�SA��d�H�=����e�
��;��R��\�|wo������W��?C#P��[�/q�e��g�ZIk0d$�(ԎQ$�NRwVtY�C|`��>7\�p;Uf�ns$	J����	AU�����w�������7h�^a��糇 ���+����7_��f�1^+�
durV�HW֯{��<����I�h鸰�I��EP��E�LIY����m,���1�6�c���SKŦdظR��	������iz��`�˳�M��DT�Ϯ�Y.��o��ɛ����2��;���ק��j�k���7o~"�zh�g�,�M��D=ȟV*�hf�f����_Cݍe���pbֱ轼vH�Ρ��:B̆��Bg��t��X��.Fz��/�K��(,�9��h)1�Tn�x�{	��m�X(SߏW'�g���s�>�K����ꬄB�M
�F��<���������7��])N�Oa�����ӻd�綐ԪU$6c�0y�c��(�hÐ����7�7���H��Fw�8��t-_�z�P��]^�9ӭx���v��=�����4��r�~2�W�ih��*o�/E���.�sH�Dμ��:X�J�s� >���la�0� � =�m%Ⱥ{�P��x-t�F>&�Cs���N)L��B+hf;\�{�I�k�KD�X����`�ew��,q)#|`Ѿۭ"�]752�7���?���`K��]�A��_l�'I��}n��A`J@Eo�ݙ�#�>.k��FH�gT�=���c܈"BF�~Ó���L괫#���┤3�z�5Z���(�N4�����Tv
�a<U���fR��?�T�$k�}��G�~��b�1-�t=�E��# 4+W�/p�P�{��QcL�WѲ�Ї	,�P�*$<4O��**oug�(�S��]��#W�5)�q#Š~���X��y�U��Ws��������
Mzo�i��+�k����"�Q-9���$��GU�LB:&��[���l�_��1SS�;	�PA2���Mu#�̿�1���Fؤ�Fe�#�R��)��,��o�W�ċS��Z%J��W��Z������ ��/e�MY����!�Y.�]0����(@�E���B x��u�mh�U7����n�?G�9�mĊ�D���!WaT¦��(\����!3���b\Vma[�	 ���rO2F2icB�yR�W�A���A�����@�j��ٔ�]an��vYu������X�|tvi�d���V�J�)��;�R�ų�1$�Y~�[�ѣE��d�7���l;�S����F�O�F'�(h�d�,u�:�qm.i|EЏ�z4����-���<][�ʗd�}��8����D�-8����x�ń���ڼ���w5 ���L��[��}���p��S?�,=�g�Z��Q"�0m�khJ@ ��Y���ޭ��k[@DuF�:Cx���W���PM"�O!�wy�|�Kx���������:$T�=3{.�P��rqA<���z�Q�1�C+YsǆoT����U�)T;C�/q�� ����|�+�����#-�d'���Hu�y�g���n_�H�����A�%��pO�O>�u�ʱ�;����PH*�ĵB7ľ[����-U���� �Vڒ�ӀJ+H-��f��+nG�S\�)$�g{��s����<5qe�8-�ۉ���Z����	�
��	N� =b�9�TҮ-S-zd�Ǔ���T�Cďp�Sc�I�O��L2T�a��|���@�y��"=�.���e�o�Q�����n9u��'�$��B }�.�%�`���޶����ڬ��^ɲ.�AeF�q��*���5�ַo�p[/Pn�����L�G#(����O}�̊�η�D OǍ8�㈹�� "N7\M��_w+$i�b�Ƀ<�.M��	aD�4���/���+'[��H|���"}�����iK�3K�2i����H,�Q<�H�`���n���t`݊l=,$������"�1�e�lO
2K�=<PVw4������MT2R��bHtb�3?΀4!
�H�n���;��R��������2���j=$Vj��pAH�r�A��P�c��@?T�)J�s�� �$
�R�J������J 4��������E�~���ʒ��NغÑg��b�%פ,������q�[Y��u��^P�P��nE��҃8%i�s$
3t�D��=.3T��a9���U��2�񗎡U��g�2��e��<!z���P<�.7yc1��_�l&��$�ZP��G��]�cj�4Ѿr�����qV7_�L�S��L���g�D��*�q��w�ź�_������|�H78�˖����U�����5<P�~��ڨ!W����b|8�2�j�Up.��`C�ߨ=謂t���`�5���"G�N7�����2��5[+)F�D�;n���`}>�������0<g����HN�$p.�O�՚����Mkb�<j���+9pδp�xr��J�W��&�<���n�f���ֶ.�k���{d1o�-����5��@� ii|^�fedP�� ��	}ΰ
ijG���HJ�i� ��xi�]|�{I{����$U��L�A	^����?��Rg;��7Г�0^���5�Y�,���1��L�:���������Ә�\�Р��|�� %�hW�d��_~4c;���#k�E�(N`0,�6m���~�Ӆ��R����[��"9����Q�ct�+٪S��Yh�sۄ��^��fV
~XD�&\���819����?e-H-��F��_|�
%��4�E3�HX��Џ���P{� ti>z��"
"�$_,�