��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\����q�?��e�I8�b�Ǽ$��"����ׯ1�V0���[�#_�;�]͸��i|Od�cP�NÌ�X�jW��!`��8Ti滨��Y�������MG��uV���pGVt
����h�A�#xM�J��5���֧H[ᘁ��f
E�	�"L��*��Яl3��oxa�H�>��E�o�(��TܽBL� �f�I9ˮ�LK��û�)Rd}�(NO���T�����`5�X_�=�<��F��;�8�D,μ	J�i��_f4�$H�*���l>AP	��)���X��W��Q������SÉ9�7ü^c��L�2��`wϩ�4�Q k���fa����\��!.�~gsm�d�5(��j�!�nqM�CU��-x���!�`۰s�0���遗�CȂ�7k�?�\�]�[��KM��ف�׏C��E����IP!9?E-���9�j���zF��<��Cڈ$�r,��9Z���ј� gw�s_e�)6f!j��=��9Ɠ�s��OҔFS�.�V����"/e
��1s�RG��+�8t 9�\��T� _I4D�j��ʸ��G�Fťzyc1ֽ�
��@��ޒ���+Zy���uƒ��=��0tg���2.׎�� ���m	G]'�6	�)R} GB��!0��d����Eikj�&��1��>D��ؕ�����%�z��J�G�Z�
�
{�����G�@�Ev����@9l�#�6�ơ!O,?��2�2g/Ք`n��]no�� ס	�,ݗZ�x̓���E3�RS�TkH^��HA��9��g�5�M��Im$�i�Qs���W�T�d[�go^
i]�RDZ���oY��s���/ލ�@���]�
^�Ǉ��H���R����'�b��0������]���s�R|V`H�~�����c�ղ�1��DƋWz�j���}��q:"���|||4�2P�}�X��G/�n��^A�0R��z��(؆��;����:�����"�;u1\�y��
�P����H�+96M�0[{l���1��E��qN�x�f�C \,ʝ����o)&C�' J��JQ:D����Op:�?V�,��{wb�FM\9�%hV�������*vW_��\��x5���K�S�O��6�{4�A�X/���p�����>2��gsirH�c���x��ϋ��-_K��`��ӇJE�E�L�ݓm2���hBxQJNs�R�9he\"���l�n�[���ٿL���^8��V.�yW�bɟ
M㳡���t��;9�k�w?�jӍ�ޢ����x�U]����6�d<�%��2�UH�Ú7�c_?��!0@���wEҥw��z3�c*���r5�/ �R��a$˴�a�	(7Ɔ��Ϋ��~nK�R��[�v����_��[���f(��9�����;^�^��L9#����O������2��22�.LOs�����$�Q�M����5��d�!��HW�Bl�}9ջ�����td�9%Np�Z��p�&:�? ���Z71�Lh��i��?�3Бmu�5��!��@L���mn2�6o{& '=�#�i n#��A�3լ�9W6�M]��W�,'�5���rQv"M�B_M���ڹ�tE����3Ǒ��Z�,���߆�����k�����~>�gm��ͣ�0��KYACav�g%zg�7�������6l,� r��d���u���:���Ga_k���E8r��_PF'�C��[�񟭞���zXtg����=XY��d�_���~����%�{�:����.���q�-?�C jۯ��hDZ�f��ՔR�.�t�����(9j�zVS#Ҁ�i4�Ӱ�td:5	�4��&���e�w-�'�>=��L�r�%&�۞��� ��v�F88[��܁�M�I���}�]5u>1��Kz���t�?+- �������l��S%�������s��y2�G��7��̵�0}����V�U�͐���S�M�252�j~5��g՟�'������s�DJ�>ji�c��y\�kv�Y 0e�.�'C;\����s�a���3�u��E�8-�ƣa-��o�u�Im���<F!˞�\��C��O�G@A��x٦�U�i��/'v{���)�#q<�#H���g�������}l�dT��S�3"f��;���JJY�U��o�>�÷�Pu���~��k�q�8~���� �	�?�rg�ss�� .K�f�^���w�W�o@��,�;L<�\�ys��>Sk�5ڃe��ּ4�K��������{��Ւr�F"t����$�#[���߽J*�?T�@]��� RB�_��[��a�H�v�j$+�E`EF���cQd�5��dE4�JM�%��&8�� �	1��h|�87��(&C:9mX~+U�0K�"g49�ǃɗ�.�;{�euȵ��PJ�5�I����Kx��9�D��{Ƹ>kك?
�Թ�>պ�7�+�-̘:�����шO�&8�:�������J+E�i���pN����@@&Hd~o��`�^��� �}$H��"\K��W꼋�EP�[h�����h_z˶@��ac!E7ת�kk� .Y�	�����8��$�ȉ�2�m��)��;T���e�ٸ~�& l��d58�3^���/�|z~��n���K6�g2%\H�����5T_�e�vh�(�` �3�E����� #A�a�+A���B���#$o�-�]�}LN��WcX����xQ���u�jTd��~c�E��/��iN%�
);�PNA�g��z���I����6q�ͭ^wǉ�5�o�ö��׃2�.ȫ&�wõD���Y��Õ���w�%n��~OB��@G��*M��rj��U����<��)45~Ѽck�4�Lw���m˚E�m'�ߵ��%�����G���g�F�d��|c�D���A%����/����+T�s��B�ң���|B)y����[�?K�l��Q��y�(d��k<Х�]첕ȣ!���Y����)������C�|�L����>�ӬK^=;����~�GN�C��@�O`��C��2�y�T)�>~�62����/�I�.��B����Z�V��5�æ�\�)#$C�GT0��Jg��K{N��[��0cǔ�X���-
Hp���F4�G�O����_ff��wL��ߋ�5�eu~Zf�#{v��ʬw��R�p��~��]���-u�s��71.��,�Ƣ��0��	���z�~��k��"�AbP`V�f�4��va�R�mfc��Q�Cm�~#��bB����k��hЌ=��Rf1a�R��ӖP�6��i�N)�O@�8�_R�"��[�u��ި��ِX0"���=]qReb����������bn_4���l���u�Jm�ĸ"�ř;��M�r�~e}
���]����<T�}�A)$����`��"�W��v�nד���0��Ua���:Z\�X�x-Z���9BkN�}��j��Zmج}��!e�*�������[��`��/)mx{<k|c=�e�]F-!��������ŇY��� zt�0&OG�X�Zi!n����+�wh�|C�2a��A�-��s��/��L���Ix䬦�K%Nb�1�+�e����H�J�����c�Y8����������ci`�Eh�f9k��Ofՙ��֭7���1xU^�1�mp�F)�����*Bb�,99��l��^9�0.#pΤ�OӤF,\!�s�O?��}#�hy�`O��Ƥ���D���x)���-p�-�M���7�g/�뛩|*u��D�;�K	d|7�~��:��x�����7v� ������!O��b� ���ؤ�e�,�R�S$<[Ph@d�oё!�!�xx��m^6M��nRܨ��������I=I���bn$KZ���I�z��[���.�lH4��,�ۻH24���Ў��VޖZ������̆Q�l��j].�<�e�J3~����a��
�R�Q��Z�,L�<I��OQ�1���su6;���c��~��ɍ�? l�o<�pS'��Mg�� �$�+�c�a1����.����ކZ��Bk"g������z"ϭO�$Y~<T�R7�C<��l���=���|؈!��k-�IR7�����P�kkf)Ϲb>]Ez�u�� ����6J���-��"�w�������ݯ�nnQ�٣�G�u=?�r[`���kkÐNX��zC:�������3�2�>�P�ٍ2 �Փ�S}�d���s�
�r-pT�7�y�t�8��3��9㙙U:D�P븡0�Xx�rU��7��߶���1+�y��8!�vx�V�WM"c#�d�)��)I{�V���������S	��ۼ.ccWba.�����b�c[�HQ�����,��Q�(.�{W%;4 (1(�F0��%I���,/7���ݬ�`|����_-�O�Ǚ����t��g%�ዬ�mp�����od���D���l!^�H�8�$��dv��&�p_�j�x�뗵h�0턀 � �<&�ɱ{U�7"ku�ݯ9i�%�[r��|��(����N��V������薽����N�:������`������6	0�C��P/L��[�߼U'\��A& CP��x��Fk�6i�e�
�Kj]Q�s��>9'f�R� ւ��և6�[�x]V=�S �//��m����XR��$ڣZ sݴ)��&�%��%�}%�"��&]�(�k�S���l78�OL�هGN�kY�f�aWk
�μO������������n��'�?q�\�'c��� �_�7���% �p��d��K{�u�B��>!�8�~���A���5,��2M��b������wb�����{��_.�F6�������=�D�^�=��Ύ���R�$��<D�K�a돾��lI�]~F�b���tN�K�!DN��.��{
�E�\
�Ƌ8��0���
��!Ⱦ���w�b���N&7~�"��	M&����Q�iزՆA�1�[�NgW!ޣ%T�ݶ(��m�0��������u۳?���/=��"���Հ�ۺFoY��	UW�M��1�E����(�+\Ӊ/$ܻ���XS�5e��d����q����]�p�Ú�9�_L:������c��o��D����1���1�C��3�xhp�,�GV�����N�9�LnzR.����4�M���%2�Y�~4�q��>G��z �7�$H�'Y��K�Y���.��g�MJ%?,kT(ߜ��ϯ�}:��,�>~r�t2��&d��t���~�ib��ݺ#DP���ӝ���I��;4��c�c����2�ER<���Ǖzg��m���^�Zy��)҃�7
����YWoԨWn>�:X�٩�O�N� �>�~5�a�����׎��Kj�*Z��#����Y����a[� *��3P>�>�=���㩯qV��`ȴa����������pQ���$D -�E��s�%3i0ڊ�QSJ����O�{����$�l��O���8�0�]!
t�������\�m���ߙA�Q�ϥ�i���+o5�\�x�.��6\��	��F+-�syp�|�㼡����;�Т],�=�c�� X�!��s�����Mx�5�A���	�? �0M'V����5��HX���ʾaHnYX�����}�������S��XUt�?��I&��W|�KQ�ը�E�*R�O�5��VX&�QȬ�Dz�/�|z��Bh36�I�3c��)Er��2 ���3!�2f��(5�����;[�u�x�q�+�3ӬE4��?Xn����aݓ����d�JX]I6F!v�jc!���cߟ���'���+0�+��`�[��R����Tc�HFLc�b[S�|�L��������O���I�r'c����d�V��h��6���];�/�D�+h����ڛY}R1��5��K����j��N�w�**�H1��Rl�1"�ǟۺ�5��B8g3ϣ�z(�\.���]m���l��)�U�
/]j3V��Gk��4�\w�E���+���l�.M�{y��E��nW�qRӜ����VLίs>,Rb��q/�#[4����o��v�}R��u a�[�v T��A�A3S~�k�Sg�𸧹��Δ�t�D���aɥU�ga���Y����c>e�b�^�0u9��s�Gۙ�l	�g�.��=���Q�Ў CUĦ��س����GimtT���(΂3��+�� pc	Z0ϭEY�����X�l�H&uI�5b�p��#z\�R{R�iӦ�ۙ;Ӵ�ۄ\��_|�ih��!�o�����M�5����Kk����kp9����[[iip�K�k�O�_V�,���(�Y	���M ����<;���\&g"Ҡ|�jiN� �dN�"Ԩ~��R"���q{{�" O^���	��J���bT���dU8�)�w���Zi�kJ2��04��B�	_�m�K+�Ǎ�e�9��*��@�өO] Z�:{�" dA0uN��7���7sF�
s"-z�j���z�6�p����
1������>o��6��OE�4iK�h�ygfo�X�oE�D��%&�\�y�T0���Y��Q�Uw�}���`5R�谗�?�����(����E�_\�U$�l�%N�)x��ʳ9�	4�h`ܑy�9_��z���R��k��b�+���_4=�5�+��G딠�ʴ�3�1{%s T�L����j�p�$�(K�cEk(#���nJ�@�1��/n�eL����Ս��B�
���FȮ�@��"ɖ!��ҟ?���)Aԕ�ɣ4{��U	$)��Go���J����c�}k	��N��t�<�&�aft����E�mH!$⟙����u)��&��}~<ҿ���=x��ζ��s�#�w)$n���$�q}�"<����+�C~ADt�g ƣsp4����]}�YL�7�u����蛙7�]��[�{���Kv�u�>T�~���)f&��5Cw�7fZXm0����UXC�BNg.�n5��m?�� �	�TR2�����g��MX}���s�E�'��Ֆ��U'�N���t��c�_����G��|�mӸ�7#b�T	����O�2��r�c  �U��+"��@�Y�
�"���#���@�����s �:��N*3Ę뉃�s��s�|�f9��qr'�CD�<�uAk�1b��P2�&X]~W�fALl�ai�L	Hv���bA�4d,78~Xnj6����B�iq��x�\�?vr�S>˄"61#�`%�虡G�d�2�p���:\�3a��յ?x���:':�:��z�B ���'(����ݥC	����o򧶲���~�rR��_�)�UБ��S�Y2�9S=��n���������G��9�	��{#{���"�X�R+�^c��W=�qc�¿�f�o���/yeN,J��u=�ֆ�;YWĵ�kI"����[�ACz�W�u�nm$��W�\󶏈!��D��秏���>LL��Ƙ�tV�_��1�t
 _A7���a���u�P5� �$6 Dֳ���%S�B}��c�vd����q�<k��[�A81sm�, ���Q��SH�jJ��h��A���#�JX�XMae�}߼p����u��CCݴ�bn�z�B�#��0`L��)��'y"*4#�8�ȥ���!7S��`�^r�_M50�AIW,B���1�?���+ܴK�k��~��ۤ� ����U?� !�&�N�/��B*�O�^�H~�(��X�"^n���2�}���X{t���F������U�B$��O�{�Ӥ�4�gU�n���X�<��t�J�L�%���5�hϮ�#�&T����)��J�N���ʞ�'�1��"?_ovN���C�mE���t��Gc��ی�2�`���C���eWb�0�4����د8�x�t�Rj��g����u�t�fD���Lb2/����@�F�w�\I9t��a�0aIP{�׻��/��V�@L'���H��C�A�k�'`>��L��o1N��e?M��
�����6�R�֗�_M��B��*<zy�G�!4�&��z}pVR�c�X�~��97d�@�t>&�X9`TJ �Y$��B�I9�п�������p�z3�
"e��pַ<�>�	p*˿W+�����\������ ]Ok�ۿ��5�� �cb:0��dz��h��sDbl�w1W�.�nr7�T��}d<�-�i<6(�ބ�	[`7���h��SH
F�����ݑ�N�����;���4dW�4�3��2\�?��JUV�R�Jza���v([?_A6H��̕��C��pw�<�G=��>	xȟ oަ���7�ڴv�;-B�d@�� �"�
���<�Z��U ��ry�[���<B���hYaʸ��&�x�J����w�ǵ��}	�`2x`��f[�2k�:�����dY��g�d��P/nH҃�<���	���Z��PJь�̉�G�d�,���`+���]���Q�ӯO���W�$�S��t�oˣb1hS!����H.�j*����E&�o�u������/G{8,&ׁ��w.m3�_���1��������o�̂�g�7�b�2�4�@��� �9.�ן7��Y��T[�{��R�k�sԌh!��!�:�[�+׋�!���4�Z�E���t��\�s� ����Z�3�lO�K4d�B-�q�
+�x�7����yJ���|0w���]i�-#�7:�����Z3	�\2M�׶��E�S���ܚ�n�B^_�6�=��&�F#�;��`����u�'���u��1K��q
�,G�|9�S�J�$>\#[�l���kz�8�a�52�W�d����f�Ȓ>�Hv�<l��f5S�yJP��2��c��wg}���4��NV����;]6{	��B��'O���
�w���d?��P��$�����,Do�~��n��,�J��V��S &
e�a�-�P�>�y�!U�`y��qd��H�Ā>����ܖ�er��T��Q�"6z�+���^�m��"\�G;O�J���M�&eX�&�=oj=��m'���co$8�"��8���H����|�[6ğ+
J$5��1��`Gb�5� ���R�E�0��v��@YRK���9�_�
�6�AJpV��h�5��I@�¿�֐��)��T�)T%�[M*=;E�B8&y6�&�À�'��#�p�2�&p�?�$G�ZWu�-Xٸ��.�ߝW����K5�I��S��R����D�#�J�Z��v��>g�G�QR���K8�C,d�DQ/x>��_�x�~֒�RF
�ʭuq|�q#h�
][!�T����ON�9S�曲��A7�F{�s�jэͨ�\�z����Z;��S�V�����n�� ��5A}�oZU"��+�	5Y ��{�����?l�'b�}�Ǘ��9ݼA�7�R��M���G��"�:��`�T�h��mCm�RJ�����	���NST�{O ��V�4\�/5W���-q�}̮:5�,cR-N��-�0o'Љ��-ZI?�aH2���a�����-��xU'מ�q!� [M��Z���|WIt�,�X��ڜ��7�	�мĤ��(��6��d՗��2M/�)�O��[�gr�"��� �g�M��U@��E��~UV&2�����;m1v�u!�a&�"�/��}��c��I`�r*�7�ˣ���j2�m᫫���MC&a� \��P��x�,��$/7���0��d�T�����dۿ�dO�9�4ۜC�1���
������*+��B ���s��@	B�Fs] H��k��h�&�jF7l�ytNa��TH=J�~k<8���ɽ�94��c���Q�E^i��
Fe64�V��P�O�0�����×��6�2�.D���=G��7�ӥ�����h,�O5n����r�7/�����$�UՑi�`Nr&� �OՁدP��²���)�<!쓅}��fA�Ŵ��g9±��ZE�r,GǱ�/��<H-:uw,Z`l�֤Uؔ_���~�G���
��N���*e�]2?I*'��#f�]�6̈́'E��BXf�����#���3G1��
�Шw���C\gˋ%_�-G$b�����a��Qk�E�2���qPd��|�r5ҹc����Y�l�:��CL$��-��9`��M�ڝT�tl�庁�Z��0A*�q����pv���v����q��e�+6���<��ܺ��!�<���o[l�-���o���0ˊ[�[�� #Ĳ�,��6G�,���/Q���-����I`�M����|����z�����������@7��:��.o_fb���r�%K/�@����58�^��<='n�^i�ꊭR��mu�\q��u]��?��]Y@�8��	�,�2�Sla� l�����LP5F/�1ϥE�_@�"J��lN�:.�s2R��� 4WRB�ux0�� 
��b�_:��^��F��)��j(IU���b��
���<>�ڱ��@�l.�z`k^�_̾�ќDk���V�,{�ă/�c8\�{�� ~�@8~�~��2U�mrνP���w��I~�`>�`S�(�u�����!�,.�����H�PO��\/':��.f�q����m���X?;y��U�5|γ_�.��Gw��cEPb%'L*l�6�w	����� d�ٕ�5|��)��#��S]�B̑q��z��Q����P�}(�H=�7Є�ln0ڊ3�o�2ò�:S�S�b��Ah��u�zZL�u|Å���T[}&Yz���~�o��M�o��IL_�`�H�$�h��ª:!xL Qmb�h�.�^!�G3	�kls��5&��T`��& �l�@��,�]���̪1z,?����b�OKH��5�GՃ�b�2Ո��m��"��4���ܯ�*��
�6>�����kZ��p÷X��_0(��k�Z5|�m��,x���`�(>X8���Z ~H�cO���׏DsR�B��@�/�=o�$P�T��S#����aۚS�])�Y����\6�B'�\�g����Y?�mۓcܟw�'6�� �L���K�ח�ǴDӯ?�M��*!r#r]j�"�G�;)��TpVg�x��T�[�	㓣J��������a�P�����X�U�V���"��-�G>�h��XSb^eU)�x�D�p�O��l�¸I8Ge��VF
j����#�4I�͝)�E�Tp�����$�:�6upf����.5~�@{b�C5�2����r녎{5��F+纾!k�δ��� �P���B��0(05�Ғ\���'�2�`1~�!��7¥����hv��:��F�~��%(4J ��J�O%��u��g0ь��_ebo�[5��?�xl&F�Mˊ�Ԙ
q[��;a�������۠�a"�fu�8���{���k.�6� ��\H[	)�@�dh������AbV��������!�S
=,��P>�q�?N���B�,���xQ\E%o�DL9��5�b=��*ż/��tI.Pەx׼	B�ٿ��Xb��&�v�	Y��'�e�h���N(�?�0��g�8馳�wV$���I�z�Sl�^މ��\�ķs���mK���4�KZ��=/�a�\���]E�~l:u�[��ٷҲ��#~A����Vh�3�y�ܴ�I)�b׍il^�[G ��
��#��G������D(���I�rX�i��]�q�N����֖p���;E~�̦�G�W9�n6�'�%X	&��qf4bҀ�~�����n��#5!����i�t�_��>�I���iNT�����rl����]��Ft�\ME��N�¥����E�����odUrbOS]�r�96�a"�8��P����_�#i�l\ M��85��1�����n��Q��}v�N�r��8�p����]�`���Ժ*�>���P��4�"�,Ss�].�`���t��~�b�v��˗���/��� ˎ�9˪}���C��a�Zi�OV�7_ ����ĳ�d�\3��� ���B�����n��{���̫^i%��y|p���$���Q@�`;�C���c�	�#�$И�=!Y�rt�N��!⸖�ob��
k�5����w�R�&x�y���ֺzjkTu�+���>|�j�^�7��Ū};������'x+�ET0���o��`滨�'��GV#`H|VL�F��SW��5�ߘ���S4�S����Eu0)�P����˭'j=�B�9���z>O�0�3�Ƭ#��o�}��5Z�3�p�Ľ���t�a$��D�#k�������Au3Aɩ�n�B��*Z~u�ζF��ZeB��Y}����Y��#ګz|��v���U�8���^F��嶽�?W��ʹ	%�";xVy�@�;�e6oR�@y��z
��!�@�Ppɯ�_��G�'nS,��^��΍���űaJ+&OtZ�u�S�	��vv����H �W�M�V���O�\!{m���y� S��&m]�!.эhޥ��J�W�* �9��c�v[Qd�����ˣ�^�7��۶�x<�x��m/BN&%��Y��b�Zt�dJ.����ߥ�!	��?�K�i�@��}z^p��v�1�����>r��"��X�Հ�!aq2�L����ĞZ�
�c�G�Ϧ�=&�C�$5S���j�%1���;Z#��|�ӆ$P~��|�8�J�²���q��FZ&L��9�.���)�ย�g;�5+�h���,��/^�R����đ�0"���#��$'�"�_ 	����|	�	'\���D�$f����6��V|�YW��ZG�r�k,�Sm�c+1���Dx���#�N��!�i���WT��F���R������nXP����2��H�v�1Is�W�������F�]M���ʳ���Q�{A����g����9$ĵ��m�h��3i�^��k�x�WΣ�����\F����ǈC$�mH��>Xٿg�u����C!��5�l������j��"���v/>���OBw.��tpA!H��oY8n1�-+$h]�XV��+�Ƕ��?�g��ůD9�n�	�=��4kV�8�����C�~H��P\���id-�`�E�-�aK�  �����s��J���8R� r���v(�������^?m����Ʀ=�*�5S.�Ň���j�����*��bBuL��Ǹƛ�_��;R�����L��[��@qdx��0SP���SĚ^�ü�8���B�q*e+G���e�{���LYԖ���k��n�-��3\$9^��?����L�B���B���5	\���*�]L��]^�͓�,yn�b�憨�8K����p�բ};�6t)�}pO��*����j3ʝ��Zi�?(]Z��I8m �b�5��v��A���_��z�C���ߍft~��#+"�s�]a=�&��������?�=mYm[��H�I{6i�����٣��yXu�}^�-4"�T����c�t�­�_h8.�Jv5���W*QA���]\���.��_XB@0�&%���e�?�,IT�IrX�m3)�ah���&����RPH����`;�쏋��%�3!�7�(�x0IX��_^	A��N�m8e��߬(f��p�g�nV�]z'J�v|�"�x�K�e�j�,�QX�K�LK���^-v��Tmg��}�Ԑ@�]MӇ����1Q
�z�L0I�ݱ���h:��-�V�#y?AT�� �ia�N��I�!�P|p��U�{�~c�(
u��e5��hC��f��֢�6W[.�X#�h^)�tH�슧�ŉ
��w�(k��I�����f�#�������!��`�L"+ؘ��;��^�/w�Kj>Z$���0�������&M^���Ñ�T~TB���,�HY�7�n��&؞q4o���������8��O������5A��a/ԕ/�o5S'vM2�U����s������.����y���) �rh�B�T̊߅�����od�9ێ�ʰi�*�.I��m�4�^�9�2#����Ħ0�NcN���^��
S�(;����ɖ)Y�+�{��*�eLhG�%�e�=��V -a��(|��P�_�4��X�_"��G��n){a�Y��1ݻ�������9�v��º�矙�G�j����i'�_+L�>[S�ߠ��X4Ά6![��'\���j���\fGYKyo٭����-��n*Q|�	u��J���$��1��'s)	��y���A��0!��0Y�/\6(��Qfhs��38
��#M����ßY��X6d ]l!�[�L�B�r�E�v7�0h_��э�$/-�#=��q��{N9�r �,9����23����-���%�@�4��F@�~={G>@3s~��D�*��ъ�Kb��K�C���UY�/��B�&�>l,�л��m��j&?C�'��9�WR� b;|0N9$Z}ŜC~����/�粘5v��`q��v`�K��0�r���?�.�u	Oy-�h
I��J3,bj�e��� ���� ��5�Aaq�MD��֘�u�&��>��!*gX�NF�����0��h[Vru�/��{z���O7�	��
�\�G�l��w�t���d�%ߕ��>�#�I�c�W�:�h�eN)�\�5�n�}��6j��������&���Z��4�z*�|����G�>�
�HT'Ej�d�x�7%�6�M/����u�}����1Wux�74 �h`��/��!������������E#�,]�ވ��b���|m��(��5�6F��̾q��.\�<g�2:�u�륹lm��]�,͝ ��"rR$4R���a��$%O�W�*��f>|���z��h�S���#m�^⟙�YH�K��J�F�9�/����z����x�����ό������@g~�13�A*���\�Ï�z9 �qA�����z��Y�#D�11�5(�'��k7��/iwc�(�frMo����o1)��8H/ah�hFz}��;��;b�W���I�"$a3�a�,ۮV�&��l	ħ>���2�q�g�[���3�hǜz㒪�y>��O�
�+�,Wf9K�B1�^y�n���e��9;{.���e�F`�Z��
�~���ov��i�Fj_���t�q2�ɷ���X�s.X.���^D�0����r��k��q�6"
O���<�
���iaic�+�O��n�P���v�@�T7((y�	�����V���W�OM��}kWɬ�"�6�A�HQ���鐒]@d�˂�ʉ�%��T�^�gQX�[�=U��I�O��L}����3��L�n6;�y�0+	�9���,��k��N��;�(�u���7!ޔ48#?��؛8rLS��fv��3�3�ym�cF������/�xss!��)Z7���(��{-������� إܜ�\�TwF@���15º����V�L�ґ�y��d��s��Myq@�~��w�8�lvy��d�'1ˊ����D	O��4��$@W�`����7jH{��.4)����������H�ؠ�k���H�/ge�|��+&kjr�l�#�V�1��cA�6�B@d�j��,O=��]�*#�չ%�A���7����ɯ�]Ӕ~�#��zې2axlҒ��^骄%ߘN�%w�u�B����������N�,5��=�T��
����-���`<������Z�Q�	htsZ��h�"��/`Z�S�ѓ��e�m��L�uSn,ʻ��V���(�W�qE6��y�����B��qc�y��,���tTZ��N?u���{'�����yC�G�ƨ�8Ka��hRN��*��0��썹�4�D��4�3��V���VۙƟ,u�N���}�>,#x%�]zȚ��F��,¡�QQE�����`�$��vR�)ʰ�>J�ݹ�3�@��f��W�dQ���$Wr����d֑i]���V�A#d���ݾ�=� �o��pQ���<����j�h�z ���7/�v%Yho�V�7b�h"kclY���u�<���GڮЅ�Sн��C��2 x?���7W>, ��6^��f��  &Ӹ�)�u�h�[�]�����
�Z*-�#d�,��m&���U��y� �̙un�j�rb����/�i:)��;g[��m����y�0iI~L%��U�hy����%m~��^ ��hATDʃ��r���B�#���GM�x�S�ׄ�4~e����
�&y���Dc�ooyn��'�与�����ƞ
!U�&��4���d;�eL��d(P<`�6�t���*�6�t�_)H� =���z�K���ƣ[ ���.�=7����FT#ᷛ��ɱ�T�J�Qk$Mt�H^�z�����^��`���oz��D1��N�hB_7L�ߘ;c�8FE�N��=p�4�PޜA�lb��C��E��L�����8�V-C�)����GMc3��1�O��q����^=O�\������p��\��}�:��? �"R�a:�ȮvNG��$���	�a����3�$�a�b'��C��P0!sI�\Z�{6�E�ޮ;�-�^,Z鼂���wY���|(��ny�f�+��8��zĎ
��-��r�����b�Q�ب�)+3(����W���
����&��d)5bQ�����r���h"u�{�x�a���&z@�pH�X}8�v�K�Ӥԭn�0��=0���v�g�K|+�% �����U	n��[o*������t3bc�Ƴn�L�ӄ7�ϟ!Ç�{��C��^�!!�����2�ceC�o�!�eQW]T��Q����H�i���K�go�y�"ޱv��n�(O�Ƽ�V��}J�N���,~��:�Ys8lL�1%��~3g�M&�pwr�a��L��:اvX$���^�17��~8ZNp�1��(���.�������H3 ��"�����|NW���d �(�#Slǁ|���w�#}��w'�ϫ���A{�D��4��W�/�������t�x���"�����Yy+#D���B�9��-�P����Vqϵ�4�my���>�h��l�q6�ov��ԫ*>]�ب�32~,�5ۦFo����۔�}͍���q���^�_<d�>H��5Us��ݵ(t�חm�	�w?i���ȧ��d���~�����}��O>�$�[�z�|r��֕Ki��XW�!҅�K��u�*g1�$��=���W�'7����0տx$C�,�H^X���M�x�G+ÇG�h��M�����6x#QoX�%Ρ��w*�'/�4�3D@>!Pd8�[�'��o#|P�>8\r��<j/�Y�5�q��
pd���S.`}�H\%��T�Fđ��Ǖ��lZ�Au�)��.t�_�"Ga�P2��1�� B�Jp�R�Ѳ�X��حVdg�s�85Ǻ�z�����e��k��|*�]G
H�qV�\���)S��agn�5q��V�d0��4N�®�6��'�*Zn�ߢ1Z^���t�i�&w`!L�[�j���n=�P�%��@8��Z�YRey:�C��ĝ�( �����1��^��l�-�C��6�GӲ'����I�E���n�w���;���]�N�w@ɧAk0O��]�lFrى�x�q�	���c�sW3�: �KnL��:j
{M�]��A˓��жs��VJ��m���r�w_Fʢ�q��%%�dY��Vdg�U�2f��|S�Y/�i�gœ�������0�B�5�
-�og��/!i\;q�H�7lC`��xoQ�L�Q�����qs�w�G�o��&� �4O����{T�zB9��9XNR3���*�8���������7@�?�"c��>x� �;Q�x��v��k`�+&a�[x�
A�خP�}��Չht�E�2l�z���u�?��WT�_��%a���&S��ͤB�����c�&.���gG1`<;�
#�$HMX��'��ȗ�\�"	�dp-^� �)�� �s�7�5Se����j�s��m��ʏ�Rsվ̂���?:=�����"���%�a��`���x�O������+F��U]�f�"n-2�m ���GYǖ�@�_�5|Gz;��ܶLP��mU}�u�C�)��C�`-�d;|���G�y�m��8�Y�HųK���_9��:�Ԍ+�[���K9>|F���mQ�����O�����	ج(#����Xvҍ�%�z٬�={�ӛ<3�s����5��Sn�^xn|J�`��9�]/�/�&���V��A�����Q�?��V�����d!8[�\C�s)\�ٞ�������`ߕ�pp��Vz}���"R��<�rvh�p	3_�މ{���MϞt�@F��Zfvy�ħ_��ִ���Oy7F#��_%ygC����]�綂��N�,eKݩGEz|���G�[���3�*�E�u�[��W�Vy�������s_|���D=D5�kO�r�*��2��$T��� �~e�P$���
��Ǣ텈K3S��<v���82_�\�����+��5��&��Rfk�YVw�#hό�avBwϊ�w�~����{+2$^^��ZN���$"�@�&8�����O�g*�P�:���~��ŧ�]8;}V�]I�7o�N�����X�,ר����EL���y�:;���b���U뮔��[�a���3Q?�_�Ft��]�m���{FH��<�
�hXd�[4 *3������J	9�S$W���� �|T��@r�5���Lm�o ��1�\ɯ΁[諒��?"����"w���[(�VF��CW�!���Q�1���i�(���F�#h�����O��kFx����sx��am���1�A���e����?����5� ���ȡ�H�����I�.Oٰ��h��
\�x�v4��rg���vE� �O�%���0h��F�|� �T�7�kc�黻ھN�di�7ȚᗷXD��O�B��g_R�`a�1��z�;~�W�tۇԬ�W���r�*|��V��+Z0��};�-���~���y���&|7��N��#�57����dk2�:9��0&�����s��!Z�bcUN�A&b
�C
%���= -��
-�8u�T��Y֓��EoE��� ��e#חg��vwfy���b��+�~bJ������l�}�`�"������*��MIc�ϟW�3��
�I�-�!z�.2%�عIĨR���,�S\���� c���2y��'|�``�a0(	��Tk:�Y��ւ��,_�M1�_ɠ��$�,b���^�ŕ�?Ԫ��?]A�ju�/�f�a�m|Y�����\�a�lL�q/CzN��/��=r�ʺB�����&��"�I}t�W\��A��*Xj)�_�E�
i,t�x%��}2R:�<I,�.l��ɛ���[{Se��gaK�<|��tG��W�D�x_�0>D�G��M����ƙn9���!�H���{UW)����ɽbͽ��o&�\Jŋs|���ޱ<p&���g����.�Y�Y
K��)c�7�w6��_���I��/�%Tc��\��w|i� {_/��q���!����E����	iq�+����RS�ˑ5_��ȗǃW�u3	����)�@i-G<-��ơ���oq�0/�����E�WU���j�lM�H��t�Hec� �WTm��|�r��i��~�ҹ���R�̜��9r|������xm���\���2塈h�fK��#�4��4�/r'�խD�G�³l��k&u|�A�9�k��py���9��3i� m$����zB�_:XN�'h��ˆ�m�l@ǪA�V�}!��Z�'�EFhC!�w�1�TV�n�'\��[�ͣ;q�;� ���?_�)|
�+���ﬂ˯#l����<ϰ
wK�h?��5�۰4.������=q6P��9��[���rg~�����F�y&VNMt��@x���֬I�ԶlI�Vk�����:�z���D�\��|��_�I�7(�Mɒ�.�!۩h<�V���r�p�fh��Q����ƹ�심���җ*���V��,����;�l�6N�e��Q卹vz}�-C<��}O�e�zsBo�蠭ʀ����� 
v��d4(���?j�Num�9�D�m�T-,��|�~�حhյЊ�`:���Q����f_SI%ύM�-<�6�Zl�e�|�q�ǽ�@,�j�1Bi��Ow��/ �FRs�/�Y���)-�B�?H�'�gȊ�P��[��uR��ϛ��rtA�|�h�V��rG����IyNh�%FΒlzH�j��2�����2b������\)�Ѻ��b�W~�
X���3��V%���pq�������w��M����0���x$����6#i�����}n(<n��<CT���=��@h�墨��w��$�zD���g�Q)� _�@���.�c_e)��]	o�ҟ����?�;&�^�,A� �K.N�����s}n谝������
��<�Jg��H烘���i�-����ջ1{l���U�B�L�Q�w3F��uu-}@�e�ܧ�o=�S��}7,��*���~8�DX���_KZYZ>I@�;�#����Vųܦ�̧��g֝*�Pz�]^��G��s��H��G�Z	��s�d	ɡ��2�),?-���t�7ˬ�%�a����y<֒�xP�|��UЩ ���|̘��c��i�s-{���yF���������k�>�pP������>Z��^�*�몭Վ	�Z�Af��ñR��A�>��G;���l{�h�u�l>��^��4���T��f�����d���}���#��X`w�I(k�����k���]����=J�B������M ����3�Iw
����J���k�e�9�5F�ݕj�����4OP^���PjW�	9-���sq��YVD�~����L�&`��<�Pa"���e��yYɄ�Ꜣ�S�/����2Q�����i��T������.E���砃��n �db�͹�4�R���g��m��1�M����h���o��NQ��L�����g�����k��]���˯��n�����jO��ɹ�Pv����4���xB���1����7��w�� pJʠ֎��Yu���� (E:ͬ�cѮ`[�؊���G^�(ID4���@�|�]Q�*�ʏ��љ=ˇ���\��[�����;�+DFu��r+��o��?�)�s�m5� �0�w>_*ruWw,�T�މ<�fW�p;�4�t���6	J;m>���F-��K_���4ϙ�{��p�qrւ&p���%�׃�3��>ӭ[l���PY���I�F���9��;�8^>W��8,��M��Gw?R�w��֥�`t��"�!X�x��7,ڴv�:fp�Y�7��X^£I����U������]��)�A���v
o9T�ր��Є��n%���hxB�|%�-;�l��G�|{	�ٰ_��V��~dHj\�&ۻW�/�]��.@0��m$�2ap���ŉ���������s-1��N����be���.��$��3g�dL;�ɲ�/*^[��'{rJ̏�L��"�I���Eq�h�?aXa��J�۟�����	�HN�_Z,wۧ�ٽ��A���P���;�M�ag��M&�t�o�p�Q��lWԀ���i�oX�R鵦?���)eU,�(��Q	�c�����#�W�Y���LƓH3�8�^�ǭ��>�b�?� ��<�@6�<,Zy5C�c�u!#Q�n?0�-�i0���,(��[��R���kaTH��8�ke��2�,�]|��\�&W\��w7b���]��@���/@E�b8�[]����7˱i£��!��y�ܢ�J�dB�m���ev�� ���n����Ũ
���o�n�2'�*�o�H���ۣd�dH込��(.i����リ�]�
�vg�#�)��ojE��K�1�f~�OZ�T;����ԶF|��]Qa1���C�<��:�ǅ�>��"XC8%��m�]��;��c&����p�_=�Z� ��o�!��eè*k~���Ւ����̣yz��C�b��f�`:򹭌�(M��*������e��(�<�EK����I �%������z�$`��=��\���P�4�4q�{3��e�G튜�,�ĺz�;MIq'�%
��o�l��_��n1��0��m4FԪ�Io�
�[�R1H�ww�5C��;�tLs��..�F��3��rS�ClMt&x�����?��/���Al��0�1���qI>c~eM0���W����T=�~�ƅ4������7��֦�A��k�p��C�}A�Y�������"kM{.�y$�Ġx!�Du�L[91�gxBs��Ç����ө�z� �QjT&R!K��P�$
��v> �-�����-�αyU�r[@����m�䆼�����r�P��ҹ�����E��ECo���s�}F�7��bKF���;dD!n�
�Q���Qf��툟+m��̗!.?.�
����j��
�	�V3��h��B���u)Uw3�vd�Ӧ{-|9:���e-��n�-5H��<̯��}�~�Ae�S1E]�Xܣ�8��a����l�kQ���|���ᅣ8������@�E��E�O͍`�	ٍJ����Wd)AM Eh�OQ��`�W�6rxQ����Z1١�i `�M}�A��G��,�� ����8������-;���4��G�C�U�쎚�UM�aV���վ�������"�4~Dk��2�������Ⱥ5΁H!�W��f���Tז�l��+%���k;gYPRp��C
b�/G{�O}��͉�UgHg0|��GZZ���z�uH^�Ґ0V��-���k	.zh���n�4߆Km��3hAi��9�P�����_JKO��n��[@�2\��i�Xq����+��Զp511K��=p�if~A,u��/��*�^�t� �\�~�9��I�X��B��DK5��b��,�|�� ��]�Ky�%�,�v�Ӏ����*���-��S(��p�`Y�/X���"�^esU�,+����X#'�C1�J㇒�ǩ�knֻ�Iq#Yo!&,���Nb>G�|m��b7R�(�������ͧ��@1��L��V!�,�����Q+��{*n�7���9[�����\��I}���-Zr�����xtɷ[W"����":�W3tl�6�����}Ue��9"x�nϱ':�Sږ���:2ۧ���~�E�p��A=07	�k& q痗25K3̪���3�M���|�O���vio�
���I���|O�J���aF��<�<sN��>��[v��XL�@�E�/c�8�)V�R)���n�;� �3�N���1l�����t3Ȍ>�\4ܴ�s�a�`��JB2�a0!y�����݃V��s)�r�K��e&�Gzk]�2�)�֥�����}hB:}�$�6���[�O(�*b Y����ZJZLa���ٛ �rm! ��:��A�oS�>O�Cst(TE�#����*��7����ԐU.�z+Z�8Zsȓ�דߵ��v�KIq_pT���5���^�q���KB�}� z��%tp�-���\@1�)�f?/؇[9�����.�yg���u��_R��U�m�2�ċ]���ǽջv���q����;*{G�^c�*�"�F)��� �[�A^�����9�\����QLVA������P�-P�x��ؿb�{���"ޫ����(���b�`�h�䡯�o���P�M�a���A�}ޏ�빌�'$8�v�'��A���y��+��'�i�p�+����0}��,�˨vb��bpdkk�;�ʭ�.���(p�E�6!Fe��yä�Ru���H�Y۳lA�ks1��-��'�)��_��M(\��H�?_�a.�L�t��H�rh>}��r�5� W�`�}�>u�����,��L�U�N�Q�@�?�����H=^�x�>���ϕ-W�#��+�0!<ـձ�W��te��;�:ۢ�,��+_��:�zv=_N#�*Ń�@X�����ܒ��h�@���S�na���n;��@r9��Q`�0�x�J��[ɘ��4�Kʦ��b^M*�\e�Ƃv�w�/?]��t4bܱjG}�[�e���g����	UX�U�?��0̜��S2L�9��[�	$��3~��)g����C7�W�/]Y��l\BOQ����jԞ�#��V�v�3�J(�� ���ha!&t���oJ�����jk�#�����HVC!�2T}b�i�At+���h��/sSW����9�Vā$�i�js}m6A���pcr`
�jzҦ��oi��q6}�0��\����?4|�40T�7��AyG��h����Xe�O�iC3�Ak�T�EI�R":ګ�����w�o�)��o���д����3�ݷ�.��oF��`��"Kȥԗ/��\l�MkL������פ�$��/�R����S�_}�S�[]��+���C:�ʃ�mM/&4L��Z�NV�����jm(2D���?(�A��o�)�ő�V�G8^{v0T�r����~Ó3,<�+&�gx���Չdq�|���]3%C"�"�g$̼@�Zյ���?w��{Oay�E+��ʪ�� ��l5�F�<��C�>���ݘ0�H��d��u�!jwT�_��+ ��s �˧��	y�$�ݸ�������2D�nD����M���rP��G�+�2��'�W-jo�B��c��9��.�M`=�~7Z��i ��=N��^����{��>�qc�D?��LP9 ��桚'܉S�üZ�z��KFN@k�J~�"��g��,~�?�F_A,/��u���i�f�ȴEce�H��x�����Q���h"��(q�83r�Q2�q}ۚ�̹�V�~� �4�cg�9�nL�Ƽ$"CJ�56I-:���b���ӄ���SM-�,$g�3�)Vz(J|��(��vn(|��z׹b\�a�d��`�R�ZҵY*�8
��ؿ9e�e0�`EL��+��[��j�����Z�~L�)my��?�۰���qV����ڷj�0-�u���0i�'Q�b1$^��-��~�ݣ����8�H��~��U�4�u�w�X���sy���
�}��Й����0�m�t���.`�s�h�V�w�t�O@�㹕���1�����hX��N�B�D��=�2� 1�xD����p-]�3�&���p��[���&aB��b\Ә��^������3`��"�%��WP���ۈVX��K�C�� ��at52Yt�����q>�s��T�eˎ�	.;��.�}A9��'��m���>���/ʜYXM��b�(Vsƞ��N3:hc�〉qY�$�bۭ2/Ie|��pn�b]#�E��:�*sh��Gc����v�l�{�pdjY5������Z|Ջý�!7�������#[G��J�>x��t�5�C��;E q���$�z���_��Ћ�Y��"Fï��9O�<�59a����G؝�s�ov��y8��4qR�u�Qᯡ���Ͱ�)ZN$(=.p,O1A"�"0D�"x�6^��<�4O�W,|�ɡ�k$�?���Q�@�,AE䯨֞$�����������BꦇUq0�|���t���!��$�h�e�<>�7�V��2g�J�$P���.=��-?��0;@�܌=3:�����kLXY���]�Q�}R\�n9�6FI����\��O�Ac�Z�D`,v��У�"OY����r�1|ʂ��9�?p�6��7�nW�)���a���$�|i���-e�Ky7mw@�o�I����+q�T��'���KB�u���?�w�x�җ�X3-"<�Y5���gv��t�zk�n��S�*������#�́Wh;�W�|p~{D�����s��?��	��@�A%	E{zc�4�N�\�NѢn�'O���M�y>��+��)t����T`-�P��CL�����F��o;+�+���P�x��'���;��QD �q����7Py��p1!���!���ͻy�1s~X1���cK�$e$uKp��!��y2<�!G�~�u.�^yv�����)a�.k�k{���^�1�p!![8���7��0Ӄ�e�$����t�.�Ne�xh[
�q�b���5��Ȇ4���~�#�����͜�G�r��c���S7���4�%�b\��:�z�4��CŶ5}n�e�ɖ���82v�,nzʸ�.�,}�ꈁ�/��͕L�lg/)�&�,���g��jJ��6�l�C\�rJ6;�WCm
F���'��v/g3��Z\)}K�?j��+�����v�"7&6��N6ۆ-;�萴��-��V���#���`vj�۰�]=>ì"Mk�N|�%�4+~�SY�r��_:ax�&j�RI�uZ%#�
+͆���v�򌁢������9<1>P=�P��7#�Kl%��1f1��&
��n�3].�W��F��]¶v�16V=aJ��0,���<����d �?�L�fx�^+�E��n��8�ίXw��U�]�ܳC*jW>�W�IRB��%�S�9�����WN]Ҳ�vBd�/=\���S��|�f��Swp�?��钱�@�a����C�?G�G���<�+2�R���|��1��'mys�#<���[|��\�1���u������	0y|20ㅿy��7��#��Ϭ�纬�P:��J�����L�����_���}�Sjf�O��>GTgH�b�}X��9�s�ǳ:F�I@|"L1\iB���D��'|��cE�ְ-F4M�5��K�H�U1�:�/�.����a�FB�I�~NW����}�py/>��Z�`�ͩ5�6!�[S�3��@�!��e"	�c�z]����y)lm����*����x�F1<m����Oޤi��=k��&� ��؟���Z�K����Ztp�%�H�&��g��hz�c[�k25��QtSR�p�9��E.�2Ӭ���E	��u�^�y�^�]�j�y<]��J�D��K��S�S?=A5�^ Ց�/`j8I�x�Ϥ�5m�-�);��t�9�$8W�Pkn>�Q��ɍXyx$�����l]��]}(S�Q��{H#'�[p*>����G�X`��D�d\����1��?��z]�|���ꐷKgХ箣�7�����$<uq��qo)UV��g�WLa#��	#m�RNW������ؓr:��;eT��Α<�+?��6a����_�HWj���-@�˴��#�Ӊo�۟�_�A���WL��m3�13���É$�t��|���z�n>OpK%����O���"9@^�A݋ӏ�	x3�T���ϓ����&��or}�5541F\e?T��C49�q�}�!q��p4���tW?�y����j�,�#t��	~�2�K���wE�Vr�I?��9��3�&	xbD��#KSn���K���w�uCX$���x�My$���ab���
C���oZ���[���:Gv�f�hyw�Hצ�s\���+��,�������5�KkR�V��_��}�/���B�N��q���0?�@�R?��Z�E�	hN���a�$>��'(.��N�ݽ��E������yk�4�FC$߽�A9���;Dz����;<�����=^���	�<j��ګ�"�rc�59�{h���-%��q����o��I���	@���lW�9����\��pB�Vʛ�W���s� ���W�DW���pysu���2��6#����^Sߴ�Y��o�����b,�2nCm��ON��j	�I]�a/��R�E6��<�S�J�ǒ�l�ni?5����O)Io˵7��4��*T��۔k4j����(7Ǉ�6�`	�6JH@Y�3���.�w�zu�)YK��
nԕ������Ig=K���.�SnLa���/����y������;�Y͟Z�q�*I	ɰr�z51+P�t	]R�ׯi��O���tZz����y�4�����y�}3ͽ�j~&L'��!*�7Z��q�T����Lr���>e������y|g�[:hp������L
��*��Ә~�cm��8����o��KbEW=�6�B�_��uM��G&O@K�f�3}�>�9��V�)gr9����33P��{�h$呻y�X^n駔0���@c2��,�z�0�:��HU���2e��6`�����H*ji�P$F���=B(�G��ʌ�����	���4,yIu�^~�+�=����i�E��y&]���62.U�"b�Έ=d��Q��>��g*j*K&��xӲ�,vm�o �i�����TCׅhu�S�p!0h�5x@�5�ɪ�zx��)�/��S�?��;ær��ަB,ȣe�"����hz�-pѧ��Q�$�"� ՚ă۬�j�j�,����?��*&�~��X�и���>㷷�^v�-E��[<$v��x��-1���?0؇���Ƭ"�Z��D?�=�VV�ؔ�����>.o�7�� k�|�A ����VAa�bII0s	��'�+t��;���oc!N�lg�y��0)��Yqz��
J~,�S��_�\�Q~�k�B��$�b�L]�!�*^/��9Qb'"y[0�h�Ԏ�ӔY0����O���(�w�r욧�-�d�gx4�����&�Η�˷P�Sd��Wi�+��8��0�	䣒`�ݸ�JH�'�����Q��'��׌0G�}Fɜ���kw�Mҧ�����["������X.@μ�6��/�lC\&���:-Ͼ@����o_�!$�V��z��G�I�n'�E���$u9��s�Ή_�u҄���A��k'�\�䤟N�Ms���񪲄ֿ�5��3�wM\b߭�(��vV�+���ԩ��ou�+y �Qt/�ck`68 ��,��ݧ2����̞X� �Vw�����v�H���p������;��vƀM�lS[voZ��K�E.X}�Jh�w��/߻ZD�� ���"�K�3��k0-�g�?F��a�E̝߽� ��ԝ���7�ok8����S�">Pe���o�
>�'&aR�Y#���b4eb�A���?�,�*�����p(/��١hi�!�3Pr���|/�ܕ`����`A��$e�"N[l_"]�<&�1��W߭/Rϓ?��4�s
v�3ք-��mY[R�J�N�u*8ޮ��r��d{&�"���(����`�H>�$M5#*�QX�RO�a���ZTs�R>�|��m��6��5�qc0���@�;�
���H��u4��B96F|Nv�F���ۜ;�]��aX�m��b�<+�̴۹���ŧ3���>�^zD��v!�h#�9�s����q�驔���O���$��J�x #����|��)/8�RtT�O���+����茆ʛ8�����$2(+#,0Ў���-��4&/o�o�f��w$�FK>W�Ű�c׌"i�������[�1~��R������s=�=�[�ҹ��`��ڂ�z���b(��
{�34 	��I���ņ�WN���C��Y�AH)qn�؁�ϩ�7�V���������H�Kү�s9���vNG���W�!��?e��o��@t�6��A
��AZy���&sa�s[�����߯r�?^��R��K�	�9R���1 ��[��~��D6}�޷�i�r�*fW|�S %ՔaEW�[w�Y�� ��a�T��򀙊�ť���p�Q 1�b� �3�3m�jn�� [OO'B��"Ce���춶�V[�+�9��|���L��Hb�!�0��ԒP�y5ݭ�{R�W� S?���(,B��ݿX��=7�Q'-�jk��;1C:���_^�]ױ)��!K�F`_;[<}P�����Y�$ۛoxIiq���z��X<C�6��S_��K#�@��GŅ��3���E�	�Ԓ�S�-�S���9'�	P�_�����I�!K%nZQ �ؾ{Wc�Zƛ��S��}���p��~n�CTp�#�LJU!Lt��V����&L[h�F��E0cu8t��<(kֵ;sZ�h4Ҏ�R=��U ,�w��5AKۖhY�}� �����(�o�
�e!�g���a5˞��i���w�~�K�h�.�c��Bfmd��?&���rce.�DB��A���¤��W@����[�_i�zo������0 ��R�?눑_Hk��uN�L��
��@<�o�k��B��@�e��������J�5ȫlJ�� �g�=cX�|9iFg2?�Ae�o#`E��S���g�q����# &���uUe��{*G�7���Ж�>s�������Nl�:F�cD�k�3��5���͚F�X��0e�)�]:=ծ�"��n�OXa�r�UH�"���o��2@.�o��w�R5ig�}�Ώ����;-M��&�B�M���|�IK��j��V'3W�I� �|L��۵ Om4$� �x�D8(�FF�po<j������TՉ��x|��J]�ܴ˷�!o-.�/����3��pޜ�H�r����!��A����NΪc�I��=\Lv�	~�B��;/�U�u�"�o�����k_L8��,Kؠ��uC,�t��O9�KcH�>��{*Ѣ��J��B�9yKE���k�A|� ��z ��k��^ٹZ�)$k�ʘ?Qc����gڱ���p��n}�V\ٛ|Y�|m��/��a�/l'A@ru7sx�W���x��V�C{�J<?���J�����f��]���������Y�9���/{'��F'�<��?�
�ܭ@ޅ;�J��n1�\�������f~w�Q��u;|��gHG�3����]q(���6�-��@�,����2��	T��F�/���5�E�f*����^�n�,V>�u��ړ��2���|�&�)r^�;��kME�~=Z��ho����y�{;��sLb����E�s�J�F|b�9z��7R�?'?D>����eݘ�<������'Q��?x�a=�{�|�3c	�6��k"|�^��<	������Tç�J�yU{��T7h
:/��w�n���3=�-ޓ�Lʕ��I����$�I:�Q����%�X#����ԍQ��ґޥ�Cl�a��?~/�3�!��n�~0�!��Ƈ諈3�/\<h���IeY\.��e�%�0r�jJ���T�M��˖h�rR�j�M|E�8�q�4����c�Al�=a��@��R�mن����w�`�%G���l����/���`� ��H^�I��Ֆf@q�ۜ'X<�^\v�/ko���������L�@�"w��<n1}`�� ��ө �;ҍ�,f�Y�fBw��)v���6Jű��?ó�,HMo;C�"/P0�7�x`}�^h[C��'�����ڞ�o���f��_'�/�$a&���|��VK���B��&G^�N_VKv�䘐�>#lhv6�����3 r7t�y�R���Ci���:�i<T�8yYr��|,�8��T"�w��|'Z���4���c;��d��_�]�:Y����7�o['o}��e�y)#(v��+��ɺN*�����q����9�.�t���4/�/�V���{ϕ{��׈p(ċ��7�laQ��8u�E�pd0�t��ʴn�Ȝ)|�}��7ۭ��d�LTf?E�cIο��S��ǛS]K�;��b��(���{�Ò8����c�剸1��Y�a熜X�}�f`�Qh���>��nƾ��}}~��s��=���Ti��U��ܕ�;�Y��Q�����9�G�Q�ᷳ);�b�ր�r��M띟�8p����tAj�a$�8��G��;�Ϣ@�p?P'S�u
t��f�S"�e��2�r�a��/	����S�MW��K�d��+>@$�k���H��̡������V��D�9�K����Gq��]�]����n���TfTX&�9f�����r�yZ�V$rƶx漘�G;�UпS/ݬ�~~�Juz)�!>X����<�х${o�1�C	���q{�F'�5"ʕB��g�8�+�*��Ə�J(h��V}��q�v��?�v��'ˆ��j;O["�����D�CfuR��ŠO(}�=�,a�V���FZ�6�g�wu/��֪DA��Q'��O>��]i����B�������)�~tLS'��	�Y
ڔ�)�N�A.x(��+MvE}�� �َ�}?w�g�9��Q�N>�2��h/_�dh,26�&G�ƩM��I'9`YWr䍙OX2z�`r8�"rd�Y0{����`��Ϡ*G����+=X��%���p��ʹ�R��hE���2EɎ�C�Iz�����jH��R
���U���W!��k�䠒w��:y�t�,G���dW~��A�-���`��h��fTt���]���'��kb���u��
����X3�x9�<|�i-��xL������	��J��<2rS�BG@>�SG����inC���w�2L#l^�eA��~,��H`��\� )�i|�)+1K��_�t�8��3����"Z,�
�= �EF��W3�>Ͷ�_�=�����H�h (oP��2����:\Z���ֺXd�unc����VY�wn�,Z->���ÜýluA3�F-�#1�%W.>��o���)�_泧�@����Vg�kf|7�Su�<g�����Ms���kڧ$m�������+�ޙщv�b� �����;Lw�9�$�%�AsH�(��rt����lEz�^m\t"����A�������	J���/�\��͉��'1��������x㬀��W*n� ���M%*hJF�*�#��f��U���#G-�&�9����UB�ES� �d�/^Ǚ�X���؞Q�+I���V��/���z�qXGW���2��eI�� ֝c�.��Az���039�m���?c2���̰�XMc��J�Cl����V�Ҵ@��hQ@H� {�yǤ������u*����(�#m�������HoW����M�^ij�e�u-��7vAϟ��&�L���(�Kh����%]~Y�>naV�ZN����α�e<�@)���IR�D���,��2��-�=�z����� ,���*���k�;��L#��!E,�� D"���O��74q�=_�	j���
0��B�\K|յ�ߧOl�f64��̼WѰ�٨wVH4b.?�T��4�u.0X>���ȏ�^�Ӳ��R�M��~FGN,k�h�%���On�\=^Gw�}A<m�P�������A����]=s�߷�QK�6G�q�jbA^����k&:f5X2�� �oΆ�.2���5�� ��|Y�"�Pnq�}>��Y�~�Q��{��l�0Uy��a|��%�n��qs�L7=���79��������[�;�4�ȫ_K��N c��%��{��U���
�+�0����qα�ٺ�3����݇�F��v�+�IH�.%i:+r#P�n@v/�5Tl$��𹠫J�K�������!��[H�o
�$q�;>$b�����!5��@�`d�3���3�}�k^�sX����{�T~1u��3-����oV3[�8��~�)�)���r�u��4ڪ����`^��/�
�3P�YLl���L�nןEjPm�̭d~��4�]��i4���j�h����m�9c��-�Q�ג.B%�1��+�<� }�?��n���)��M�%�c��z�f�u\iه�ChׂL�[��N6��!P2����8������;~�Y�]�+��A���&�k<�9{��T�Gi��}@���1���'{h�5؉��{r$@�2���l�:�UL���MJy�R��򗺍Y��f!ʪt�,��"4E;�Y3]���A��8e�/��q�n9m�C�9��!�7l�t
���dTC�i�l6�|�`k�62�P�"�$����P����.Y�Kt�	����ג}���q���|���U2��pi�b:M���򹆣>�~�Iw������[Qi���Q8�B���nv��n�WޮB
�\��R&�5b{�����p$��?�`X��B���3�2��Vα
R�Db|�dlϕ�:�I��=n��]�G����.~vc�i)��M�cO����)��K!��vw6%��jH��2�����������lW?u��zM�@u�DK&o�\��N� �����L���5�3�j3��/g2J����;�+�|�X�b@?�j�$�7?���F��H�6�oϧ���X��A�Y]u8`|��� �����̠n�3^��
�I���/���L̍�c��S�9$�+3xY�3�=x�Lu�e�vS��M]^y���.х�O]-��:�O�:�!��|�Ɵ�[h�l���)�7I^����"0�ӃXƧQ.
�l��ZT�WۓPH�{&� �>�;S���X�w��\�L�NÍF��}]��k����ߚ�&��/X�װ�]g~�Ѹ�Ь��
gQq�i�<�<�R�v�([�z���&�P���< ��kH�Z� ���XY߸���C�Ūtz�no�k�*}R㮆�˭�	�@y�V�)Ux�z$�[��M-wy�zMڽG�W��s�Xl�Z9���7��owC�ȒM�tMq4�t7�/F����|���f�ݐ,��Z�Ef_S$�*�͒A�O�����u:�#t���X�����2�TeKF�)8)$���*:�^�:sc.�	�H���z>;�US�(6!��ƺ�YW�t,T���i��y�#�
���/5������^�aF��X�������8��������r#�>s���:^�VCKL33��HL�<�4t!�Ѻc������w���.�>��I�<s'�"I�z`�0S��,�#�O	o�s_��nI��h�a$'h������-�
�����7��&��2*/�I2��Ѯ�Z�&�G�~0��9�.S��_0>��5C�JZ�fK�ۑ��ND	�b�[}&�`�N,����_�{a\��7��\�����uA���m����bFA:F)G�<:�ݳ� �w�;X�X��2`C�V��=�T���%�3�,���c�󿲕��.�&'�-F��������N�BI��K�*&�w�u�]����{��d�b} &�S�B��-]���y�S�4��nf����
�?�b%���\2�	�����&�X���c��{Jb�s�ev�΁5cy��@��$��ƺ��aY*��o��������&%�5!�&y��\��|�=�������u�����!T�������ǌUQد�`|�]�	�Rq]�<�.�&��H���%�|c�^QA�5M������$����Ü�	H���~�b�m�,�~_.!�����'I&�VϦjx'j8n�T(��w��Z?өT��(�^�V���#����@x�Ա�E�q�W�D��b\�OFH���6Ԛ���V�_%rPmE줋s8�WE֦
J<w��A`o ?\0)����ǚ���4�r;
p�͈����t<l�d"Og����9�旴�~[>����[n��Xm�a�" S#jAJФ�� �LNY����|釺�
Q�\.�.�c��`Ls���h7r,?7� o<n
���ʶ��K�Krǜ�@D�JJļqE�)Ef���w�T�4��G��Q��o��7�@��-�l�>^~3�����Ӣ���4{�&��<x�=o�Xe	}�L*i�_|mac�`�x�`m ��n!�����4���cvKOWH�c�6����D4xڂ	�|�e`)i��������
��%W_�˶h^���?w����mX�5������QGhu
�U��pu\���]{�I��k�bO;�I�{��g�Mg�K=߷����d�@�Db�.���]\�hy���\�K���f�\君����
b-99���8����0��!r�t�U"�g؝t���$�8���1}��j^� :��ؼPWS��O��"[��Jq�'�3��`��ぜ\��2?�09&�f�*#��V�eQ)��U~��NN����\@5&��Q�.Ѯ����m��.��BAK2h��!�]S0�v���sZva�b�"�2��������?���R����k�{)���vw'ey�E�\*�����y����@�;�9��@�89�FL����l��7��Q|���T������ i���u�A��$�ȟvd�d]�#J!D9	"}� �7)��0��4�k���8��m��&�L �U�s<T�b���G�Ҷ�G� ���G�ow|HJ!c5���q\x�2��yZ�*&�$\���Z}�Pxt\]~I: �w��ԱS�z���^������s��եRJ'@�<�d)�k�]U������Py�8��:}fk�H� ��rO�[�^S0>)f�[�Ud�,�䚀t��ϩl�|��Z��C~��Ա�ZsL9 z�1�J�G̬d��8[�y.��eND�9�x3
"z|Zh�D�-6{^�1�E�l
z�9��b�C.�2��OJ?�<s
��>p.���Q)9)�ȱ����W�ɠ?��Ύ��):9*��f	ј�V�'D��);i4��ae:	߇!狒�t��>�ɸfNÄ��y?�r_ށ{@U����g��6�B�|z�|��y�D������� �G�:0��&�����@�t'��κ�K-��t.��Q���ϺXn�n�u7VT�o�c���l�8>���6��?�>�(Y �r�O�Q`~)��ƤG�%<�[��$J�+u�Ӄ�H��u8��d	�t߂��T��62�"��E��c �f�VX���+�{.���B��9�.���Lh�!�3m�+��	^l1� ��v���p_=�0�h
B��Q<'M:�e�q�N�PI������R����i7Թx��cد���eq�N�i{�H���:xH�q��p�oP6��H�Θ���G�R�q�í�RN ��+�����0��T�' ڑ�0�lԳ�k���~������8�rf��#���� ��$��2(l�����}p���'��!�j������4Ԗ��L8�����2�Ұs�U=T�6]��07NlZ��_��z�`KD��U���:L�$b�Kdv�[@��	T.��� ���r�vmy����F�6��^�j��|O�v��ܞUH�,a�B"1B�fġl1���1���$B��(ꝰK��i�&:b=�ގ�Zѡ�D��dR�]XݟK��7z��l:l[T��x*�6SR�����ңw��g�Ъ9����s�W�n��mEV�Te�0l�oa��]v6^��DmT����9�ձ%�q�ޜ��K侐����)�w�y��`�N�Q�/~6�Zs���9N�J�[�����@bA�kn�1��$����;w0�Cӝ�����n��G3�t��V�n?_��e<b�6�D�xЧ���J��P���!����Zخ�7|�� ��Pnri(P��@��p��YsM�5\v�1M� X�P��/��	�%+�M�����5Ӟi����{�������ȊZ��h�B<zT|�;�
r�ޟ@_L����;�Nt����Z\����Ie�O����Lm]lOQ�}l#��/h�~h���ih:��d�}��Q.%7������n9��Rf�̆����˴Z��jQH^�L.��9˳.���(�b�̅MA��U��?Y����襷�~O�)�϶��\�AV�T
pn]Ȟ�����雑��7���U�b6���E� �����Oq!�i�I�[�־cY>�uڲ��!]#�&a�Rx
���h0�	���~�3Z��s������� [zm���I�������#,�b�1Lф@5G�/�rxb�#�������6�߯kᡕH���@O:���pq�����:�r�?%��=�k���0���=LP	�#��dN���yT�)�8c�ܟ�|�S��0��}��Y.�&�� Ak��6����%�]2�+��sC���R��B���;B���g�6����4������pٞn\�Ig6��= G�?��P5�,�R#���a���e�8�S�^@%;O��.}����3��54?�љ�{,a���*����Vr3ʫ��`B�k{�,WIF���d��ARj�3�Ux-�uۛ/�X�n������#�>��<�e%BT���AAsh!S��qy���sGPy��?)Ev�7W���:g���VI��z9h[��#2��1r�ti{�_Q��2�S	p-x�`ԡ�H�7\�wm@�7������i�,� -ʆ��o�k *>�/?~��/����r��\�;��yBKڻ��'��pD�Oέ�>P0}�f;z�Dp0�מ{�9�mD���$�m��4
��x~���󯌹~n7{7��Ø�]�����^��}s�ب��ٮO�0����w=+��e�w�%�1�ta�K��&I&�,�[��? �-i�J�N��韘V�{�Lri��U�.�:�.`���=b�b�M��9'�f#UN'B�6���u!�_�p��fN-�P��EOxr��Fp�Cb/S�����zW>�R1m���4<]5(ݑ��l������6hQ�����E� v}g]a�;�<&���vU���̆��r���!39���7���/��P�X����A����W�?��]վ�0�ȠQ�le�w������FԋT�;g�Xu��7x3L�1�kNɐ����q�|f_��� 21 g�=����B�Ċ1/�)�%���Ðbw@��.Ga[���3�52���$ܔ���WГ��� \t�H���tܜ���c\2(�j��2��rl���%��|emŲ�p�2Q�J����Pf�cR��e��� R�>P�.�>}#����^x���t�ُ�#K��>��fn��׋���.��p�,)ں�3i�Oh,�ǹ�T$�IgJ�7P���hZ9���cL��6ε�VM�������o�=���C��Ŷp���S<����Ƴ0ؽ�%1��H��0�^飬�����3&�i��o.�������fX0,QU��?r�S�8̢�|wRQ�7�p���;�_7�/��a��z��p��H�&LȚ�`���%�
�1wf�i�����9�u�!�n��Ԋt��c�V�Ҝu����n�"�1jŮW*��T�PZ�Y����w��JFSy�7�ޜ��R�xw�Y��8���T';��E��Q$j3�_���z�V	�]iR���ȷ��U#ݩQ߭"���!�hӨ���6�i6X�k��I��!�,�K (fRY�>�"��	Ce8�!���IN��F�����]o$�v`J5�'ٍ0���pK ��:���yx�|x�ˏ忧�ר���H�f��^���1�o"����@^���K�?�Wj��7د�VS��u����2x�3vKM��SL9��s'���C_�������!N�@Q-&LP�������������&g���s�N����"5z��t��!�D��H�2S:�K�H׷9�ojt�v��רp5���-��=�2�z��W�;���9�D�5	pA
;5w�2��x-v� ^ͺ��K�V5�e��W^�jd�[9<gYT�
*��}��"��&�"3�8�p)s8T(� ����P��X����ݍ�*��H�ߺٮ��bK,ǣ�+PE��5��!S�Y"C��{3ӨkX�h֡a޼��z���N�,�oJ�C������Oq�L�3�N}@s^�>3C��(l���l��ҺK���UE��Pn��IykE.sDE��ٴC��gZ��Wމ�V/C�QU7�1��@/��T��#����ǨA�Lޯ���]�Q���T3�)
��@�q`�H�y'EP^w7섻Ј�
.Xr��J|K_��t���@C�	H��(�V���FϚ6��s�iV��j<%.�b�>t<'�3\��0nn@��E˱q&��ӂf}�Tp&��@�9Y�7���Ƃ���pF*�@wy�М��V��}Wb?5Q������%$e�h
���U���adU�W�1u�����uyź�=��j��ɑ@����[�_��Y���r� ���}zE�L8�'S�i��_x�U\r�8�@���,c���Ɛ�֖0[��ʡe
�#�`*�H�M֒����k}�-}��yA�ȉ���%�1���ܠ��8�Y��p�R ����C����7a!���'�
�_N�6�G;���Un&�H�TFn��D<�Iʽ�^]�c��?)D�dx,p�p0����"�7�$l��Aճ����G �!0���X���������[�
 ����>OE's��&�%����}��uT���y��r� t?�����`�Tdw|�E*���XH��cH���������+��;;�.�/� &���i�B�o(�o,��{^2G{8>	��[��iQ��ZͲ%�DҝEV�������r����ᒵz1Tk��b����$h�Fۖ�"I��_��F@��ʌ�W궰��Ӯ��8����L����x^�P��ci� �V3���wZ�Ǽz�9��a��6	�[��6��ilC%rA=FWH� źk�&R�KN�!�#�n�Kfv�:�o\��ʉ��T����-���yKp����)  :�m�7��?�ר�{>C-|��s�ڦJ��<Ϳ>���Z-��ʟ���jQ!���G�h���
	ɣ�Yi	y���r0�/s���*��g���!��B�����v�*kz����q��얪a��w���� Z�W�3�qP�>`�H��6^�E�0�d�����~S���t���Y �"�q�#"����:�T��2�]���=��6�s���Ts�"��g�3��#�H����WX2���Gf�<�+�I���}���.�	�7'�E����?_�`�̨��m��c�{}��T(��a2�x�~�9�M�l��V�Z�LNRNi�|��%���'b�1�	{ې:�D&GI��g`���-�����Qj�,��op�Q���T'coY��m
H�Xv�d��<�z�W����a��&�0,;1�*�ǩ���*�Oy�H3ZȡI,�衳���|���C<�#6�+p���j�~��xdL>úZ�ix�okt�c=;>?E�)�d��jc	ك��A�u>a��I���R�n���U%�L~f�������9<@��>���hӴ�dq��^�DٜG�&o��4yW}6���_�T�e*>�~)��~�?����7��Y-�g	�-%]+�f�'��;c���^�z�K0����!�җ4
�����E�3p�v��n/��X ���|ytZAd�۠�cվ���%�����_�O�U������'�w(���s$����%q�8N�s&i��E������KOѭY��Ѱo�hV�Kc��bv�����WF)��Ň.a�GV�:	#ј||�'-q[Ge��FF��s�i�ȉ�	$uD��\����.OZ����4{��e���p���1������4ٯ°����N�[]b��B��xd#0S�r:/h٣LLLB�B�.���F*<+Mͥ\�gޖWLw�Y�$[�De��r�>�_�ARGrF�����0�ɫ��wU �ua���b�_���:��xm4x���Py3Z��.˟�i�K�L�Ւ��%�cE-�h���G�eoG流Ż_��v�����w@��<N~k%���>:�!�L5Տ�*�>�F��KkS4�y�M�@o1�T�Z("��X�����ұF�!3`y�5�7K\ 
.yH��4�1�}��Ӯ�����NsB�П��dMB��9��U���*Y��_��3�ד:b������%M�oH3^4k�EY��fm9Q#�Pȇ�7yu�Da����p?V�,}o��V�A����%���֚�� �Y�-<� Y�;N��/�i�w��d�~�˲�����O~����61�A��oG�d�g��K�b��$AU=J>#j�n�PQXJ��;#���!7P������6g?m�>��^7��H��s���H���6��T��ji�EQ�z�G�P�{4Ua�.�92�0�{�ҭ
kZ������6��%��W'D�5泟���x"�L@��5���*��H��eͤ�G�a�����%ǘ�A�$�E� �G-E���+�B�"*">���3oof�b�"�V�5	.B�B��q��;y�_e��]H	k	�C�Hz��@�T��ng��%3��(�_�a��s�O!�Cxz�c~��.q8ޭ��X)�Ш5{���v{i����� Y)�A�iA]e�5��%C�;�ſ�.~��H	)�{N������.]x��U���H6��'��p`E*����g��Ҷ[��ș���1�����ݺN/��
ɋ
����Z8{�o�����D3��\��㴴nV�k_,���!	%���]�&��*��٬�-�`�����;�϶�G�����Þ#%N}*�}�f�b�t}�/F���O��w&08�2n�L�f\�K�(��X�u���A&�W�"h�ز#x�m.�O7�pVK�R�%QB`�L˜;��_";�p��!3�"q�*Sҳ㍽jp==�8 i��I�@%����[泔i�4�D�u}���J�J�q�jD>$�l���;��S�ʇ3�V#�l_wj��c����~�1�CҤ��8)�J��Lݣ1��)��lF�*�7�,�N&���["d)i��]�?N�����0P����k�z�U(��Qh�~Jpa�,���8X̤�@��Dc���`�����q�.�-�fݳ��m�e�C���P1S�b��������hT�2M	p��m��͈0�Y8��C�[�LiP�Y1:6'9�K�8�������JV���o ��	S���ReVd���a��Ъ�0d�Lڙ�z�5�;��7bh������l}�3��LpG�)�vrB1q�{k,�����:m��AיJ��"-�N-��W:'ޠsy�9=�ʀ�Ł�a-Ì^�B���>֤�pm��B2R����{�_��U�Y�_���ߵoO��GC���3!��g����W�̫O�\�0�=��g��o�.�.I�*Q��km��)���F�ǣ[���c5l$��l�? r��!�_�����<�[��C!`g��v��x��}Uh��q��G{��M*��X�D�1H��.����	Vs�xW�}�7���"�G�l�A�a�P��$��2c�Bq��T<s]`��`K�*{((D���l��I^�l*�0�,��J���z�_�"�-����G�j��}&��.$�o�!߃���$��^�w1�t����[qa'i|YƟ���`�*΂x1���{[ g�pyG��a�=� !�
\?CE���|;�7��,�;��X�[� *=�w��9�2�x�������Y���˿�[^t����_�r�֡&m �Q}��׹��>�l�0
>y��t��E���,��e��t��Տ���o���lNs,f��w�-rq��� �1`��jȖ�
��#"Шv"n�B��u�U��Kv����%Uf����5��Ӕ��j��@D�����[O2��{�0g���j�З��>������·�`-'#3�%����G}$�Iˣ.Yn$Q!,���H ~��Y����LI՜�x�C�ȉ�T���=�@����]Z]�@e��Ԇ3���D�j�XLl:�ϐ�������!�8�'��ZµYlh�r��1xE�4G��?��BO��.��ҹ��d��/)|*9�2�s>,B#�yr���\�M��hо���w!����,��o�m�h���U��XFE^#�ʲ��W��۫�!P����6Ϋ��.�~��vK��f|�WZ�@��ͨ�#@��(������EY������'�$��*�]�����H�6L���8�[?3t��X��*��}m;�o'y����SΏ��i�ꑊ��vMXH��6^�Ǔ6["�Ӳ���ǜ��ӎ�r�5h|d)(��#�u�͘�ۘ���JN�<8ˮ���i&� &k�X�#���d��þ�*&�\��H�h�1)&o�I�MC���4�k�)���/org�$��dԈKo�]�����)󐙛�����,������hJ�$�`!A�f�x�K����%ZQ�N晬����� ��0���ᱷ��IGZGo��%���7S�a�yP�X��@���A׊����Y���Zy9y��et��c��ռ!�6̎�9;��e���,c����g�򻶇GA�d|��h��*�eWFx�J�N���:Fƪ�K�Ymi{�g���A�4S:	�Ⱦ��Τ�gX��9�\�F�����d:;>A>BS�3?�^�"b ���L�J�a��);h�e�@@!�M~A5[3��D4�8ml��y/ϗ����1�	�Ș�����l}��Zj��pt`)�7:����tYK�W�e�]#����"zs����#�Y�|�#�wݵ�w8R*Ze*��!�!���d�T��Kҏ�!f��Q$�q�$`����\���~�A�Ru�oy���d�TսE4�0��/�4���N�ū�l�1��SP mc�)����``{/O�mJT�Nc�1�^8YR���n{k��@���A�$��U�2��Л�;~r��Hg�}�tG��2�(P|$�
}�<�k���uuB�ŹX8�ԅ+�g��SB��"�Χ��^Hv(+��4g���BE��6�i <���Ѫ���n�j�+��f�eFk�m���?�>�֭��B����[8��X�^����A�4�� �?�e"�U}ޘ���3w[~"P���3+ƥ�2"���C��VN� } 7 ;��na7����Nt��ĤgUe��P�1��I�'�\���$��MY�*m�0^�^��ݿk�|���9)oZ�&�Fߙ�􂞇�O�F]̨��X����j Ғ���H�	�y��
�HɄf^��A-$h�o��m�ݗ-l (��<ʦ?�1�2�I�W�X��N8͛^�*(�,�1���ܻ}���#��.כ'�G����;�Pd�}�����3��I͗V
q̂�ߦ�O��Se��[n�]K����r���c��|��g�ı��U����ϼ�Kj�9�*1q+8�N�S�y'��ɣ!Z�Cˋ��ޘ��g�}��{2��Z�|�8v�z��/�+�_�����DM���oQ��F{r� �H�U�%?K�����N�P�<P�iU�0b?��wE\صf{�)��R:���['�[vʁ�;��@^��E�Aə�2�����ԅcޯ~A�|GB0�9�nsV�x5�ԚA$Fi!�����8ag���S����rG��Fw=��\��W�i8��i�Z��6���"2�8Y���6��"JX�:�X�]�5�
N�8���8ǰ��K�G�����J�(YaA ��Czۛ��=8PN��JZ��s��N����`���m��r\�Qc۱O5b�P
�l�Uq�*�@���=��������o��T��h��Sd��.�g�-o�&���e�}�9CY������� {f'��0�R�&��ߟ2��d	V�l�[�rɧ���s#��,�\Ʉ�@vB�9�\v-i܌�Hҟ�U���♖��\:uߩ;����L�	^�EP�Q�P�����x �	���\s,�W�*��83~gM�M�Ox�{�^��'i܄iK��ŋ"�k_}tQTq:ͦul�|t[�y�x��_2���V�p)�>S���|����h:�V���t\)�dMRS}�MG��G�gk��U���a���f�9���(ǆ��V�d���X*Dp&�\-�$�W-�Eo�Uڀ({�9�����Z�i`{��ź*jB�W���a]�a�+T�#�i�o��pj�Bz�i�=��TH<�X����ä���M����(m��KM;�Z����'�z��S0�ro�1�P����� ���#r�I��B�o2���kw����$O��{yV��tjLRn��u#'��u�[��|��V\�{hжHlI�:�f�����]��ֺ�����R��N�&���E��#�pª ֌`�~�5�ԏ���Un��pg����9�G��l�'ɹ H�Q@�$Y��(�^p������ڲ��C���8\rP�`;���y��n�>\IL����9�Ԙ���B�=��q�(!�������Ǉt�t�p����9�7�V��iެ���H�n�\E���:��7�&��nO�}I��Ɛp�PNyH�_u�rT*�lD�?b���7W��)||e����"�ϟA��8ȼ�v_5����͙ء(��(����W��d�h�́��j�����R�}cS-� ��z�s�._P-[�-�Jh�H����V� `i)��]����9ɓTz��V�p�p��t`��
Ū���'C��^n���2Sla��N�u�Mc�R
�.���ߦ���Ϲm����r�ߔC�!3~qT�b# c5�B��$h�����Z����`	�z<�ʔ��P��#�ޙL|n�%0-l�u��xl�_R��o�n�����fny���I���#22��H�_V١��g��)\p[A�������@�.�J��M��˱�B��A��d�#�!�
d�Y��(����Fd�����E��͐�Z�����=U���"R-=�� \gOD�V��W0��>�)��#	'̿I�ib	qi���0|Xzb�ГB�Y�i;����Y�W��@��(SXʤ�?�/�5I��n73K`�hp��] ���I����I["�t�3aγ�N��@�t�Xb�H�[��֐�,�P���֍�*�/h�����i����@&����"��E 7����	>�/w�E�hاNx�E6d��2P�l��d&X��jhل�"��S D��&�ܑ����;��e��E�qN�_k�[q-~�ͷTe��Fڮ�'rM���?����-�$�#��Ʀ���_AJ$��I������KJ��&�@���f0��a�1�'�^�]զ�����kkP�m���s����a'%$�	I� �m��C;&��Z�;>�N�5�K�,�w$_3���(�#��`�X�G�_�w1(��|�5�l���Hϕ�Wtӿp���|{��?	e����4-���xGz�*�0Jÿw�OP�@��'6\ �yr!QW��C}7:�g_`V��ƕ���M�:�>�l�ó����a� ����?�0��O?���EPs��R��1 h릨�*�7w�h�iL��ѫX?�>o��_/L�q^R8#����m���zы������vX �-
`�cf̃oD|�a>H����e1�+{���@B�p�)��r7�����p��O\��s�L�� ~�o���Fvwa�A1a�ޮlaRKʟ��2�]�aBN��,3� ȏ��AaU���=e\u]P	R���9-
{����j�Z�����P�ӥA�X�3��T�������H�S/퀌����A@���&xU�8�{����~`�bRA%��k'�����k��:��5��.�ȹR7)C<���e[	[=:��ވ���i �`yQ^��SH�
�e�mX��� ���I�$Vi�)JN4g>�Sk���NM����F��9*�gR�pޢk�o�g�Wҩ ��£�=F���5�0�(E'�K���uxJV��P�E�C/'�b�KQZ��M%�8eɁ?��D�R�%yu�G0oM�����N�2揖�o}���3$	����H=$��+Dʜ�a%�t��N��3O�L��`��NQ�{�6�1n��CՈ7��uVjc��]�h?3L�޳J�#?���4�<Ԋ�߲�!sF�;V�v�hѶK�p@���}�n@���YX$��HvE�W��"����}e�_:r�>��K��� ��`<[��~��#����E��5�x0����y�"
���n�ʰV� V�%)*Ҵ��`75B���ٹ�:�ae�i75hC��������ڜ�lo���Q��"h� �ǰ?uѸm��#��÷�ր/��G�i�P�f=p�)2�8}��lq��R�N�NR�B�6��o}���aT��݀n�	�ns�/C*+!�8<�2= 	AV�F<��0]���_s��0��oj����o�eql��d=���ߓ䠐�~�>��N���0��o�y'�]'��n����t=��{�b�wߓ/���N�b�����%5KW�w��֍7��� ��XE;b#��04{
1<ܨ̭�&�����N��X�[P��
�D��s;������t
��ޕh�d&C�"����e�ʔ:}E���X�|��-��$� �0Sh�RV��-D��p�d���q�y=�NvK$��A�A��[��hk�:�G5�"Xq�!A��*U���t�B B����c@mp%$�@|ð>=^o�A_�G���;%(W�!���:8��f�u���D���#pY�qo�¯\�L�O'��{�.T#9�:D;�n��@v�Iw���@�Nnt)etdX��K3�e��h�u��{�n}�7�]2BI� ;�9S��q�}�t//Ƅ�dF�
��}����
.�VgRic�@/����Kƺ������V%�^Ց�Y����4|k����.�=������hߖ��r�[��m�+8��j���yz�QLx4r�XT�eT�x���D�ܣ�wg�|*= ){#��#M�Nu�v���@�m��Sr�g�ҏWkk���V�mkqb�L�㝧���-��n�Wݑn�7C� �E���\���[%���ɬ�\�|k����˞����3�b���T�-ѱ�Dg��RV�f1�12(��(��<iC3���������A�"Lw?tkH=����e���%{v\�f#;\B7Ab�ϓ����7tV�&4���ӿN(�Ziu�SPi�!�u�H�rZ�.����|5�!0����X�а�cC�0�Y�gk_�/�OAG�G��lzb\�d�Z�=��k~ז}��C�j��Y}��M�L��1m}�aW�@Ķ�aC�\Ӟ+���}QG?v�v[�����d�%]�&���q�W�:�2�9����t�C�d�3��!W&G�k��X��oS����s��`�Ko��,���DU�p�	PS��]��|�'�R����t����?�d���QA�F�`�<�G������'k�-��р@C���W�2��ʧ�`�2�+Kհ��y��T��W9`.%�y��޳��AH����А�j�� jN �q��fi=4\~j�O6�q������LfJk{���9.ɸMzF^\}�V��[:cZM|CD�\Y��$�Zl�Kj7���r�Șo�[y�1�k��/�	�,��U��TXi���L�eB�6�j�__�\��Q�~�a9�+nc�K?���НΕ�h�������CY��������M,�Ĝ��M���>�^	����p�V��;��2,�"%�E�Q���\F&���-6����~C5)�!w�ESD���`r9S�$��ƺH+d�F����E�\��Ỵ�A-e��O��4�����2l*z�g�V7�ذ��,6��B=?x_,(=ӭ[H�'~�yX�F�}���X��y�XA����m|I�K��ɲ;;���X�B�ص�I�$ۺ��byO���C��0}��"�����K|u{1v��E���$	X3��1���o\�X^w.q!J͞�+!¤F���Z R$�դ]���.��"	#�_��U΁��np���'���zW+�k��y�:kQ�4˾}�r
��S���w>�*�d�G���:\aEo#��d�d�M0������#�_'<ř~\���3��<�,(:��݂�4����N��-yR=H�?����/8RB#&ƒ�����������������W� {��|�R=!��]a�J��ʯ!���I#�0�-��YҾ#r7�7��pI�z)�)5J�&�_�]"\��4���]0��^��33?`��{7փ-�'"�0"_�Hd���J}B=��3����rN��~b�|����.�
%g��̬��㭾�^�M�)t+ڽB1*��>��̬a��
nH�%����B�̕�>H�/�TR]��Z���T.�mqK!��@_��?!�=�c)$1����.�¢/�:O�-�fȢ����z���}ǹ^����}.n��1`�xW���Ay�t��WN�\�Y�dA�yf�Jd��N؁R�p���r9�̤�U����+��:[B��`S�2���D�$�Sߥ�fښ�Ρ�ty�n������Hh��k�l���H^CV1MB���S�O��|��P���dS[h,B���3���P�E�
���v!���]��)����\t���z�\���a$�ZI��Ε�ws<q��� �ce��rΊ7�Q.��u�;��ʲ�����^��TWԧ���[ ���d:���ݶA�2-��H�D�R��y>�ؓ|�P{��9ՆWjm�#��򘁟����S����*�wa#ݷ��% to?¬���X�n(��%�o
�x]�}�XD�SUn�n
p�D��i������M�v�¤��@ҫ�'RO���[�)�6���,��g��R�@�z��6ܴ^��cO��E��(`_�n��T7��]�����o�W=B`S[��{W�j,���.]"��~f�05lɖ�3���d�<�_���[4+����(�9C�A4<��O��l��Gݤ�?s�Zd�Hg�$�:�c1�����ɣf����62��y`;i�8�eK	���%�%�4MB$c�Z���M���M�QȨ���OYL�~�;��/Kk�5a���j�;3�%P<�;Xq�L��ks��΃����6��x�X��8z�(��:�C�����߯��j^I3'��o��J�R� l�]k�̚_.F��A�*ОS�Q��9�y�*�wa�$��Z�n"C�x�w��D�Ey�)����K�J+��R��o�;"��wP���	��꡼�@1`���Ï�����1���d�vq "�݄Y��L,>�j �LUd��fVʋ���r[�ԋ��F~K�UOT޳T�+M'��h��%�!����S�/����h� ����v���, j �<�m�c�H�2��=KN�*�Q|-���A�O�����Ѳ�
"2�f{bV�yN0�_�h��i���+Ӣm�0�L}��
�j|4��+�W�.��Z��wD��+$>;���TLܤ\$���iDAV�[x0��6Wv
�Jئ�����|ƣaU��$�rw ���z�b�*uu[�4너^��D�{���G����Z*f4���$�q��j���	i�&1�+���kG��}�,���;SPiC�z��O��PD�h������&]U.����f*���Tَ��Ǥ��֞Ն��43Ν��K�P��-.!va,"�-��݊v[cD!H�z��Q6�a
����0��񀈣��%9���y�(�u������d�ߠB词�V�c�����&��%��o[d�*���f$�sy�*觏�0'��Ĝ�1����E�����Y%�L���^˫Ѷ��؂�e�%�o�z��0 ��S���cu�X)������:��ݤ�"d�4�y]ѸO���~��oq�q+4����~�ι�4^��O���
m����jF�@�kc�z�\��CC�~y�N�h��K�I/�!*ӿ:�d=����9�*eҡ�������_�#B�GP�۵��a�2of�5b`�6�VJ�Q�>t�F�A�- B�W%�ːS��O鳦Cͥ���]�h�>�Ms���;�ޭ��~���a��6�ֶ�,p!
����i�	�-XpW��ź�6�ۀK��G�K�A>�✮޼Zu���� ���)n�pUȵ��$�Md$mk�5N��ūnP˹C�{p�H�un���1�h&�K��6p�ӈ��K���h�63�D�1`�� ?����yh6���BLp�5|�Ү4�W%O�ּ-d��#+�3'?��V�}�� J@�9L H�:�Q�������i�)��Wq�I2e?���v&S�2��L @b��~�Zwn��? �J�=!).�ᏺ��e�����y��Baw�M�	_�5V�G�Õ�IB�0S���o�R� ]�����KY�o�ʫ��X�Rkav��A kJ�u���,�����CK�>9��gҕ����F��_y���*rf����	�MY;�I[�LG,Ciph[v��(x^'�'�l�Y��`g
����׉ַ4�Z�����Ѧ�X��E��#9�p�&Ü����I���:�e��a��� ��T�6�)ȋ��ʗ�2)5�hu� �����PV�z�]��6.L:�p�{R����,*!�T �����(S�(`rTY�D����c�)�Oު��9S�whF5�_��X�rA�N��lj(����R�LmN\�Xu)p�������#��8L3mR����f�+W���:��1�N�x�8�����qt��Q;Sr��Mv�vA�ϏP���o-��v�`΋M�j���=��4j\�4�A:\�b�R�;ώ<�9�c ����Y���l����B��͖�t%�~X�;�{�G�u(IN���os��<��
g��������1��e󉡔Fȉ�ʞ�E:ז��:�w.}������(NNB����An֧��Ƭ<`��E���ˣgy�N��I�+�yo����m=x�u��5.��5Mit ��c�m�Nrnb,<�v�k��>�F�?��"M�x�"����K�7�I�x���5(�t�hFEΓ5U�N�km�:eE@Ы���J{_y[OOf[�I5��
h��< IZ�9o�'
ٸ�!�[�a��?�� $�6^����s`s�[9��p�w{�Gmw9z�ݻ��=�\��W4�