��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����Mڨ��˳0��`q�M�'���2&��Ȯ�W�4��д��|�6�K!b�'mY�`��L����T�7r~��<7�C��T��RLiо<��{P:��w�[�S�Jݖ!�s��?���� ��\��Y���T�eT�' V�(��>���ꁇ���4�M����k���͑�[��"Kpx�!6%�IT�W�X����oH��j �M��6ዣBX	�Rs��A4�eX�� <i���t'W��=�h�1����e(��?c����Hj�nm��˩�Ej�c��{�?���xm~�ٕCQlk�N�9�
|c�cb��!X?��?-i�Y�x�g)�Fk��Lx(�JaX���B�ָ���WF�{�(�@�hH��1��d�g�i���N�m2d"��W��o!&���h  :����
W�ra�Q~�����ͯ�jJkI�G��O�Bww&�F��T�\�]�\i�Y i�6ѣEDrE�L`����L⢛p5��/2"���z��� �g/deZ���K������.{�i����!G�t�SbM,��"������(��tR���a���ߤ�\L6tM�N��,�5O�5�p�7�@{3,�M�^������M����0s�Y���M�Z��˾>�_�OKV(�^��.9Y�o6CZ�~��U]�Q���D �;�M4�~d��?VW�a".��5[��!�K�rl��@��So�T��J����;����x���@��^��Vy��I����x�/���]$�O����N���e�P����(�8qF��p��7�|`�F~�}�f�a(�+`|䴞9EiOPH�jC!T�s��~ Af��ĸD6����?H�Ī��m�NnO��	�Z�\��<�w5��*]���q�:OJ��}�盷�>�C4)��4�t
�VP�$�p"�!����,9�3r��ч���7s1X�T4�:���cb���=f��h�!]c��89�ދl��=�.���N|�~���|@@�����`��a4�W̤^��(�A`"3_�QQOS����갾h�p��0O��f	�UcE�;�3hp!����GC��P��a@ ��>������c�@r�s���P���j_o��j|~C)7ŗ� �"����3r�9&�*.`��+��0y)h���OJ���V�U��D�Y��]����"���@O��N���,�w������C�ϴ�pd,6vY��`�]k�'r<~��X*��2w�X_|}�vῩ1��<��9���,���X��UAnfmѸ��*�z#���4��%�),�n���tX'�^�܁ȉ�� %1�8�ozi-�q;'!Q>�J(��I��P 
jD8��������y�T�=N=3'� ��,���r��]՗T͡����m|�����N�����A��܌�H3韬��9'v!mK���mT_ ��A/�	{�?x@��ȝ�-��J��?)ɒ��� ���])Mtg,�&�4�G��ث��y��{n[uU�rEtv
��Szi�c����"�'яG��=ZՀI3�Uw��n�&!���x�ӯ��Ö��OŹ@?��R\# -LG��h��n�`���K��K�5;�ytH�２��C��W���W�SDf��e_*�6��{4�|�x��܌f9��G�ײ�D�c�x(�����o�e2�-��̷��eʮ����v!u���kK���ތ�
3o�X�|�kj�c�� �w��
����d	�mښ��-X�Xe��ͺ1H�R׆d��ѣ�M�+�� \=�~��j�^�	\1�`�O��|�׎y�����ws(T}�+�e���J��>i�z��h���Gf��fB�������]�A���h4���tOa{Fi%f����\��)t�(���~q��g���G�9�%���>�z%O��&�k}��l�00
%%�YInv:��X�t�̊rY�x������jݒ��H;�.8?>�4'6;餾��83���jh����%F�, `�1×$��XN��C�8�3	R��+V�߸��,�/�'�o0+�s wo�>d�2����5�;v�Νi Y@8���o�B	b�7��7}�*x����\B�ey�V�/��3��;��I�N�;��%~�ѱ@{����W)�Qen��HK��_����v�c�V��^���4cl�zI�V��j]�T������tB���|gx�<�k��U�ԹY��գ�Q\WL���K�F@�:UV�-��b,B�����቎��/>�`3�Q�p�ͅ��~�8��إ����F����A�x�:˵�a�h���|)�c�\��mIX�r��$` ����@*GXP�=��f�}�ݳ�\�8S����vG��)�pn1 �}��g�$�p<N�(�Ő\ �s��(\�����M~�P���I ��NB{J�N�C?��1���>�A?a�g�����/��%���Np�a�Ώ�d��|*1�3�9����,��<�����ؽ���C�-؟#���O?�lc�|�-} y#��1/_�ۧ��R���!�-CR7+)�_���n#�gV�����BO~�D���+�z$}�u�<�B����ׇ%�4��V��O{��OU�G�v�I�M�O<k��)�`��k���yn���q��K�8N)6��2{�C2��Dш��z<?����7D��}���=-J㻑m�R�i��_����Ƿ22�^}�Q�N!]<t�-�]�X��nu@S��O���1�@,ቱ#xC�g����?i����+�H!%(]G̞��ټ���S�9�J#���_��`�E��}���2��tZ���t��}��*�i�kP0�F�	5�D9��3����:b�I^�γ�Z�Ɩ�وC���c�|&�m�Y�J��a=Y�Z���w����Z�,�)R�Ǻ��$l�`�U���黥 �*�/��`����*4�B���w*pc��\����pU���w�C9C�/�9�.2�d��_��K�G���nބ}v��̺Ql��elv��J@�e��#gMe��Y�����W^��4M�9#e�dnloȪ=��"�!{/�f�x�ۣI���������'CS���&D}��ͱ�x�m��B>-
R )���k'?�0���&���.��L8�pdh5k��_��ZZ7��mJ\�E>m�����}�}�BM�a9�ȯ[�'<��qI�j@,[���_���^,����~�h�hGT�6��\���f��<�]��u�dY������� ]�g��Θ�Ɇ��߉���_����D̋075?�cݰ�>����X!�P/����i�\_U�,����ß���	4�Ey'k�������ιAMhu��f�4[����(�4���+DJ%��1?ٺ}�ײ�����f�,���tO�PKA	�(�q]���U�mX�܌K�`g���D���-�T�%��̢��i�����a�k�^�$�Qa�\�[�/V��s-�
C��op@���"���Z{���t+4}G)[�ll�f~��[����jb=�'A��Mr�k���@��#���l����>�M���d����375&7~%'"�g�A"�hb�[��:�r�瀪~0=-����#}R�mۆA���gEc˶J"�}�p�\�lu._Ѷ8g}L����Cf�,y�vKn�O@�kgԝ���%��N��y�2�{\����ʺ��#l�]=�Z�ʺ��3'���\��(ٱ��|��3@�J��ޯ�n�)���
x�X�iM�&�ޘ �?ݮvw��!)ף�O��	x �S~-���j��=��S0�P`�&~�C�09��r
_�������"��ؚd�Xŋ?�&������L]�K��
����Mx�<Z��GТ��UtS���E�����9(���!�ݭ�g*��CRtn{$���sN,�8���qQx��Jt#��e���[Vp�F����ZB�� R�!�1P�2���kϵ!$;��
�IW�zq5�u޼rY(�j`t*M(-v&��Oi����AY��ȡ%:��U9_���%�?� +>7�^�r�/�i����;pG���E��v֭2�܏�����Jc��V�����*���΢�|ޢ,�������wȑXa���B��Jph���gиǕ���,��VBa��� d��.8a?w�kR���1��3>6��i�>���N7���d���.e��4�75�58W����C�7�.7�x��b�����(�攞K�{���r�c,A%y���Y(�7�K�����|���1֏�g�t6Y��0]¡���Ͷ%}��*P����k��c`�s�T#��Ч���(��]�tzAj*��r+��S2@Rg�:%:C]x�C�hw��q]�l�r�x���[�[�ŁKq�%Z� �g��k'���Z��Ԋ�u������i���v�5;���O�e16��m��O�6��G)5��BfC�ea��E���v֧���6��hb`�,Q�a��Y^����kc��=l��Lq����������[n����������6�a+�+|��
z�?x�J9׮��Hs��+�]�fq���yjvPߧpS�u�7kt���#��C�,Ա~=�Ͼ`��:��@�B�0㊥k���r����֕��'��e�Y��郵��eƶ�㤒΀���`|g���*8\�Pa0�̀�~�m㗔6;�\���B]-_���+b���<j���M�۠��]��Z7Q�(�R��ǔĀ�7�#���f)�Xzp����3A_*����Z�HH�G�p�<��ߺ{��ݖ&a7#�������UH:�,�L�%Uۈ�1a��Z����ԅ�R\��:��'�6�>5�K���TRI���vcg��Stj*��N���(�.yX9�*��:��Kg�b��
J�ŧ!�e��-��Ĉ[�Ҵ��M� ��:*o�¼��d-Ro}2p����OҬf�����)1S�_Qeݳ����#��6TqXkd����� ���cP�n��PF���{� �Z�<4/jZ��̧������,��7]G[�u�GBG�#�� XFK!p��AB��s���4Zf�߯����,<2V�C��oۋh��љNw�*��&��V��c�1����o��3!덻�0��k��k&����k�����%	I��
��A�ȯ���N����Z/��SUw?�
B����������L[ko@cW��wo�<�ڥS�O��!�qe�70�� ��_l�49��M��U�i]>C�%����wo���3�tb�#�9 #w��_���fJ�ruk[_����-�p��B&�t&�Ia7�M��oAQN�^;.��L_�$e�h#����������@hp�WZ��cw9�{L=����ؔ+<�yO|���|�8
;�iA�Ή���l�$��K71A�ů9*���v6磀)��&�VF���g UН�_�q
��S��!�i%�7uB��E�3#��~9b�.�SldҊE���
p�k+\ b�d�������3L�,�5�nj�b��h��:��g��.�W)�;���[pfԩ�̝2%���Z����2��?�{ϐj��U�f��D/YA�N�j�\�kX@��[���#��ʉv�Sr�q�������Cѵ�Z�F�$��2�+�OT�� >��~s�2�r�{��U�Ǘ�*u�yqm8Cx�VZNF�~�.����@�%�<��Ϧ��L��9��Hp�2����Y(�n�B�c����">�\/$�	w>c����N���˹�/�+���܊��h����	i�tҋ��� Y���U>t��ds�Z�tW� <���P	�q}�Ș{���1})���pEМ-+ؚ��*��#�;���J�U��ag"Ri���Ǫr�ESi�h��B����J�<�u����k
��	�5���ϺD}	������$n!��T2�nߔ��*:ݚ��.P)����r�����<��X�  "PM;[l0�Z�F�*�)��3'�4�)O�J�t���A�8�8L[e)N��L���e�������J���ȍ5�(� �ɫi�!Ww(~E�m�������9\Q<�b@|U��hWP��m����L�&�ڕ�W�N����N�tp��W�_h<#��Ѩyt�[�tL�ߣ7�7�v����I��s�&_�Y�h���u�V[w�'�&[0�)≔��N�-3�NSڙ� �6���n%K��H�Z�v�dF���(�?�Ռ��x����m��>4��I-�����Tb_Q���1��n
��F�b�S�`��pj�o��Y˺&�r�����Ȱs����#���YDBjCfB��K	5��_������Q�+-m�T���#7Bc.�T7�Z�~��f���8<7̓鶻����*��v�F�ǽ��΢�~m�t�C�
�d�����0J5�fuۙϞbX�v����H��ۋ ?�7���5����,p)�n	U���0�{�l�e��iJjň%NJQ9�3ނl�׀���W�l�z�0a������hK���l�lE�sd�O�{?y)gs9[V�?ֺa���5V�y��E�A�K���n��J�A�U��[�ڦN��}E��_����lP"��!����mD�xx����8�@��U���� YM���E��>:�f��Ϳ	T�į�_f�k����v<��;���֌Wt����2�#��w����8^�해�E���������������rR+ �#���x�J�T�FS��m��/���Ϧ�p_�&�i�s�z���3K�F�s!�����g113�|��	���k�	��Vȱ��=��C�;<�E�$Q�Ќ��jAI�n>�?�v/�\�ts&���-���cB}�_�)��Z�5�q8; ����U��r�M�|�j<��7�^�K<)��K���fڰ��m�I({�H=Ӟ���鈖L��R������]�y@�ED/�~}(�x?���<�[A�/@�qX~a�*�M�s�����?�����K�����*��s�y%�`�ЃN�>x������� |R���n��������=﨎��?���u�a��nsD�[��(���z�6L�C|�� ƒF���|h,�L�g�U�X��.F~��}i����I�ǚ��a+�)y�<�2�I�o��{K��86�eI_e�������ayD��G�Wk=���SP#�N�������@핢M�؛h�p.���ކ�0��pg8�iQ��^��*bq���M�5K�Q �8>���ᩴ=I�J@��ߓ�l(�u��Ǡ�tY�