��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�k�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������H�W޵α���N-�`��6����ݾ�FF��eF4��_}<�ےA�[,�|{�?r+-��]n?���A'xin�XO�v⨺��sZA�R4��g�psXdm"�d��Q� N�c���%���9��-SX⨣����jR8#H5�H�w!"�]Aļw��)���F�P�4�Ո������2"?'� |_�-�e�����-���^,�l��M۪��C���ĥ]����R��Y�AҚa��r��cF�Y�q�aA�����^9'y��z_���c�`�ԗ�p!r鯬�h�M���i�2�{�y&�x������?�v��[�
�/ǩY�|�����%�n�����h�fZ���i��*����[���p�F1���?oO:�9�\P}w$8@�@n�8Lq�|�w=�\\۾�I��YY
���Lj�h�q-��ťbUY��,���ѻ�_x�k���y�a�l��a�Je-�ߵ�P�z�V�O��z3�zﻬM�W��!aπĬE|�q��JRQg:^8b�ο�KjA�%�j�KVz���2eN�Q}����{��&u<?�7�L����>�b�	ٶ�����X�����nx�㾔ԑ&
�ͿC�"0�q��&N�/�_���r�G?"�q�i��7ݹ*B��9Y�4�b7�Ҵh��0 <8��,��rmh93�r�D̨���.��b���#�V�(�H�R�����(�Id�. ^�>�7�=����V���H�� ��,Ȫp
 �a�2M�W0�P��k)q'5U��N@�F�_?oy،�V=9 Ǭ��{�|H��ڃa�I�ދ,�$6�]N��HT�3k����Ɨ|�3�X�}I�ϰ
�	*o[kހӘM���n ���R������������	��>���/_~��;[@�e�),޾���^�e�f�͓d/u�`P�(��g��:�`W?��s�y��q�n��[����d�S�3zզJ^���=�&�M�x[����k�������r*DN~��:։lf�c�0�n���:}��̳�My�SX��dS�9e���$[ق���m�i�������ZMQޒ���񳅪�QqGX�*���3Ho�/dĳ�Ƹ#{B��1O�����8H��e�8C�ܳR��d9��Qd��cs<'
���))�4����bǬq߰�(�,�ǯ��J�Q)S���4Zu�=?\�T���o��܉8:�ԛq�/i�54�{����Xs�#VWﲡ��Yq���oǹ��"	���(E�YK��d�"Ҹ�J��oJ?� SY)����.�����m��40zP�h?��6t��~��m �<�,r:h�K`	U�H��n�Mb�c�$p��P�`�^���	������؄�ta��ǝ�Nc[	gӝn�^��Q%Z���a�/Z��@� ^{�Լ��;���v�"fŠ���ӓ�Y���@d��x�-���s{m�^v��t�۫��Z����s]"��y{�&�F�
P���7��L)��O��~�Hk��Y��m����TW����;�kH�;ڒ�`��P���:��=����z ���P�iT�[I�l����i�����}3E�?��r��(,e�gR+��W��-ťx������Ѷ-I�f)ٙ"��/�ۋ��w��o�ͦ�l�	�G�a���f,q��)i��J &N�X%:��	����B��zAt�