��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1���e}ʲ��cg�t�ϙ�a�:�KR�%���ݧw���ȼ������ :�8��Y��(�[�*<��uǏ�y�Ѹ!��+S�g$���Ŝ^*�Ϥ�0Ҧ�ǳ�ț�x�BpD%��A24nx_܉~�%�\���6&�+e?����6����/�N�|tR	V�r�^��ʌ)y��=o����{t���H<\y`����sPև�l��M���,�[L@�HTS���K∂)���(.�#�ʖ��F	���d
���}�_�45 �7꠸���F�:W'ߕ[�/H���_��+'T�J߱��J��ݦ�e���o=?ɵ2��y?�h�����!��ԉ%��Ԑ���v~Vְ<}���QbwĬu
4���)���]��䗪/�q�1ޡN?�ͪ�1Ë@R�&R��<?V;��-@���	��@�#b^�%yHM����m��o�����Ʃ���D��cx[�ңJ5*Q˛j�m�Z�ݲD7�V�)�p}\\�����A��j�FB���pl��Vz�$�0���/Sp.����lg=�T�C����k>�y�52
lAdch���m9�B��D:�ß�J��Ćq�8�I�WM�^��Ν�w�l+�8�!��Nt����ԢaԥU��p�%�Z��B-�D���»K�Q��m��aн
"�y.�uv��4�.�<���d8wY}�8���mJ8�C�|[�®���LT��5�:�v=�?!��%��_)k�A���[�W��/��9l�$��]�Gv��ufs.��N5 (:F�7�0gMBek����05�^[[��W�����gX����i��w��Mw�����Zypy綞�I�~�K�2�7<��0���9'R���(�	����%�?-ʠ�Zk8�|f�b�+Ox��J>ٹG�鹪p�K�Rg�Ϫ� ���z0�xN���+sm��J��f>_,KF�SC
0���nɗ��!�uꩁ�=��G)K
M͝��J�23���L^�$��Rl��˭$�,t�b��2	B���	�"��:Q�=5@��:�����lzc]�w���w�k%�;yȤ=B�߮4���p�#��Q��ہeM"r+�
�n�#�@;�K�a� 	ی���rS��n�֢����b�W�ɲ;�U�3�-�S�u[`���\n�m�s��EC�*�u��O�aV���v�w$k��>��yT�g��/1�U�e���?{Nf�&.��d�}k����b�M�L���/�����1� !��F�K��2#�GT�����7%��҈��:ڡ�,�˛�du=�rb���LOȆx�X�@
,�C@Ԍ�g��v���F��+���u��{C�U'���h��R:�Ɔ�����M��1C��{u9�!Y)�'��sk\��

�k���h �R\��g�uO(��\��qwC� >�٥Q�1����<�P�׺�>�`�����(�]��n��Р1���J+8ҔZ��$�5�5��֫�I��l���ʩ��p�7B*�h�8�����#B
���MZe�M�1������G���O{np��범54��Kc�x�7f���G*����??���B���V��+�ny��cTt���oPc2���Y'���Q��g�4Rf6]*����C����������u`���
������^{��M�t�V��ld�|����y��2i����Qu�!K��h	��\��?0���%��|���D4Gd�Y��!�gS�mXϜ���S�xq0ac�`N���I��t��Bqj+9B�mFÿ{���O��.|��
u�Ҍe�<��!q'Q���rm�Yp`c�)������b��l���(*��~���j���0�2 b�6�o��.3ޭ#�pA�`�H�ʂ&KQ�*o����\�o^(��/�+��T���DOC^L5�w#���U�\=U�oI%���w٫Y�}�
��x�^d�R)
ya��dQ%���^�I����B�Ρ:in����`�	ATNn~�R�7�.7��@��(DB4���c`�.��"ֈ����`؀��M� 8W��p2���S���7�������#ٿE����*C��_�����C4
��0����uCO�x�x^J��Vm'x��1������N����z��&�cL�ܹ����t/�k�t*��d�� ���Ν��<��0�\ <c}(�	��#��?��9:2�?��g�p�S�"����1v�=F��9e,H������^�z
>?V"{W��ՙ��x4�9yG�m��2َZ��Y]���{� !j�<���~f��.e�E�"P�B���)��/�ՠ|HG�G�e
N �:'��6Rf�~v�Ϙ��eC1��o�4��ԭE$H�4�|ܹ��S�1��R��;�5q��GXS h���
W��+����z�߰#(�$B�8*#���s��0&�z���	�84EvT�8�x4Q!������P����w��Q���`'�,%�,��b���~�y�$��?�g�r��6�݋1II=������7V�&l@����Y|�u(k��]^�U;�k�B�	M��]��s�,��2q3*6L��iI��,M���Q�b��MH�)T���Q��&4щ0S���?�9=ٌ��6C��m&h�c.놽j�4�䭴B�Y@�8`i�fX#�0 ����U'�U�7}��'E�(�%= ���U�R�$� 6�aZ��a����u�.+tu�J�G�Gڒ*`D�v9�!pA����S	3{I$�ZR�9�~t��뙍?�מ��a��^�=��5ͭ�~� U0 WAٱ�'���A��9�k���F���dic"�'{-(�T�~%޲Gp��k�>^]�Ǌ�!8�J$�� �D;�w#�O.l	�y�N�G���HB�\�Hښ^� 8�eDvSF1Z*�S?��L5,u��u�t�ve�N��M�t�:�jKy掰~��&<ih#��%^�����'��N�}O��*��0&���2$`ݗ'(Җh �
J7>�0i�u��+s�&�ӽP�V�����������g�ց�}��d:E���*��D��ڬ.<J�<R�$����p8�2�&#�;FҞ<��s�Co%'WA.w��ڕ�r���G�JMU��{G->U�Oݾ�6	1��Fܰ���{Y�i���Q �F���`d\).��~5ԥ\s����V�BPP5m+e}�.�d�X��<Dބ5�z�Z��B05�OH���`�z�_���&����S��a��H��m}PQ7؟������X�r3�&rߊ_������>/�d.}������au���և�v=��K�v�s�!T��yP�:)����G�W�P=bQ�p��PL;Y���y�"�>Z=�C"�n�`~:���S�tr�DJ�4��.�$X'�}���ܕM��iv�� 1�6��� ����Z����Ā$�/n�m�j.\�[����ll����|?�YqM|��4�²�{�%-�"YyW%
/z����/TL/ƥ=|���V���N}5�'`��°D!ԅ�d��Iu����?��>��pP���I"-�1��{���5Tw�?l��P�T�V�HE�t*��^�P���ڦ�e�z���1X0pVZT�X �r��U�b�{����X�]���b+��] w��P��EI��ڗ��~���&I��2��t�3'k��:���	O8�M�GbSn7VL��ě��T��M�zԨ�Ӫ̃K{�䙞ń�a~���~y����yj>m(��ܴͩ�2=�V���[骉�S�P�?�W����z*(S	�@�q��Q�c�*FI�Ζ�|	�����O��p�I%��2�rk
U���Wnhv�0!���s�D�W���k��O��Ѣ8�6xB���,Dq[��ީF�+�
���~e�W� .���D�����TpP�q�4nss��4��n��%�Xy�:=�2q��(6���@E������(�^������}��Qz�6j?Q�K��~�m�j:8q�!D;�����IkD�@3��U��d��>꠲-.�/ě�`̅ǥo�O?n�%�/z�-?̱?U#�1�,4;\r�&��\�����e���6��4���V�P�гT�Q,k]��bׁ
	����7��ޕL��E��%ӯ 4��\V$F�O���L?$���E*�:���t�l,h=A樂T�r|?%<�i�!�Q�:����$���y%F ��<Z@��'�	�.��ؙrS>�JLǟ�h����8�<��;6x��3��-8���9�Q��ӝ����!Z�Y�Aŀ��~]���]� f��g4(�'��M�Qi,E�\�%���F��F����lDti�W���VI
�w��C�S���q@�6��1}lW�E����(k�O��u4��g��I�:�ʧD�_�2zr���ʙ�xIF9:F'ٺ��n%o�'��4zl$P��E�hR��xXE�E�m@a8��C�4O�К4�O~��Lo��Ƽ�,�˻�x �$������MOV����"[���vМ���TS��M����;�WP6����tGO5.���h�iD����m�3��L6��<�BÐ��+ŋ��@�����
��-,=�d�U'�b�W��r.0cP6�a��s�fQ�P�C�\���S�ʐ�آ>�/�("����i�@��R�-9?�MA��M �&�r�ཤ���O��X���D`N���/�J��'A&����"�^�*1,Qɼ�ǌ���>���u}v��*��8OYL�0�OS]8�U�_�7�^0髚�����f`��_J���\
U#�֋�z���R,&Cb\.���EC�ί]�~��-k8�o� �Z��W�>��S�{�g4��6�	��J��L B�^,���L	�Tc{�W?v�q+G7Sk�+�Y��2.�!2 �@��G��Ӽe�Mu�.{1�f���h�WGP��xg�uab0+�*�;yw}�fA$8w�\�'�w��.�*݁�x3ZX-8@&HY#�}��-� �&��
�ϲ�z�D�3(�[m���Ƨ�~�OE�!���M�B�w�iӱ]����I7Z�Ae���3"4�M�/����@�\�%�0�Y;ZP�v۷Qy��jQ�R���-�I�1@��K�ca]�~�p�r9�G�Oj�~�œ+J!X���B�>d!k���L�������n*22��^��L|�v�.X�Ҙ�:0�6�0@�����a��c�c��>����,w��Dt�lT���ۂ�Z��B��X������&�'P~`�f�tI��Y�3=*��L��7��їPY�����(��c;�X9L�+��������I��\�0�� ��C�VXG������� l<��+�2�x+t*/�$��&���9"F��}ͯf����RԽ�&�ԇ���}P�	�Oi��<�ձ6ДX���7�YY��Р��b�<�Cغ��F�)v*�J�|Z�t�����������Q!�?�yR-�*t/O&j`v�w�/h>�4����zq1��bs�I0��Z&�|� ����)�������ߠZbV"���[�}x���;�	8���)9l�m��M8b豈�Z�p�88����� �7�lA��Hi����X��fSv��,�`<�JP[߂�ef>���`�߳���l��fJ�iC��%;�����2�α㎷uJ�	�p��k�Y4eºm��E�����<���ʖ�r�Q�Zu�-�44���$@ˎ�#,�"��1Z��&��;���/ǈ�5,ğH�Zï�3�"����Y|�L����	"�G&Ȫs���3%/�4�σז&@X�{�@(n}����x
Q��V�Pr�5�0 �Z��5�Vd���5Q�N���S��Պl�|�g��N+���t�X{�%�g�Dr�D~F�E�O6�l�U�L@Ѻ�+��b���M�T��!z��VZ$�^Dc���s��Sa�~��/��P��k�ܭ2_��?�:s�A3I�ܧ�r-�oy4m<��/*ڞ.�
���%?JLSYJ��Qc��7
r�tTQ�E�[j�ʲ+�Q���J�Ԭt�\W&O�_"L��=�[��D�p����k+�����{+�{q���`jc7��]�{ȷ�S��]�A7����0���yP
�3:CZ�f��ET�2�{���eֽ�P@��]���B|�q4�|��Ex�`3�,�Q����Z�&SW��{Bt���E����?�s�ܡ��2�����d<f�2I-9\;q��*�ـ��N�є��d��P%�p���(G?O���E � ��PV^�kW�5��쿋��lTd,��R��UFE���S.xu�t�*8���`�@���}
{���x�9������z\������͒�hɣ���m�%✞d`����{U	dO
�~�I=Z��W'��X26D�ѫ3pF�|B���V��t��%R��-��)�f���r��g`b�5, ;"Vޕ��A^��(+�k�8��ǫ�����Jk��m$1w_��������9(�f�� z)a�?�/̋?_]c\+�;6ѡ�JW�BBlfj|-`)�A��0�$��pN���ʎ/�c@���zMH�����;U%�c&�ޠ��z��^P��':�`_#s�Ѻ}�2�jNLp�4�d�|�-WB
F����Ď�� ��U��#�+`�TTb��_����J̟�V�Ny�<��΋�h�[��7� �(��;��T�ܩ	�i�C��>��}=a�#"���[R��D��c��J�A:[�Ȍ��M#����#��%2P����]���1����2DqBw���/�苲�t�6 "|�҂��+�n�+@���.�ɿ5��j5���B�R��UJ��H�����~�&��@N�[t@�� �`�>hd>�Fb��09�~��|\)ձ�[L<���f0Mz���:��䟬,r�	
��KYTiJ�-A"�4�Z:� "~_�y>�>*׮MEMn!�)ĺqW�Ƃ]���2H�[*I��gl}��;�P���;Z��JR�s��C�� ��*��-ݲG�֋�\��R���	�rǱ/fVuX"�K�2Ѥ/���Jj�l.��Oh���W�^t�Xe�m2a��Θ.b�=�.�X�G���FL�,�:(u-L�\Ǝ��L���e��/O��P�q�ȋ8_� �y�1�R1�f��F����#Aur:P|8�y�*�{���|��t7WD�ե��A��
���x�"6"�4F�km�� �s�At�����iﬨU	�w��%��$�Ɗ���c_�|S��~.|r��9㘤Tk]�ޒ�&)nc��"I#	j��C4P+�����Z�]�!F�n��'ba���zM�Qz�ti��%�����K%X��X�8���K�x��[:7��S�n����B��
�%�p@���h�c�B�����LR7GG�I�R�nS�KJ��ءUc,�S�7PաK�+m�L��Ӎ0��}.��3�ha{����7�A�����Ar�O�5C����J� ��*ƽ"�d����}�$%G�	�d)�[m�Vۮe���)�F0+�;��#��*�Ϧ��ذq�q��<�$�F+ģ��k6W�F��dA*�m���?����4����5��MbI��h�����s7,�%��������%�9���H�Q���#�ډ�5;�UF�b�}��YUw���g���M��L3��y�X5�&�6yZ������B�Z�/GKΔ^�-c|ID�#�kBp���u�2l����=Q�i�2�j�Q���0��+�b�bH����D�D�j����4T�J�0]�2w�|:5镛͂y������.�#9�ۑN�V�d��#"���/-��w<d#x{x[.8^����oy��e�J������ɹM:�H�Vh����$%MѺc����P����G���Sj�a�� C�������&wT�!��[@����3Ѩ��<vj&�@lP��70!qWL��*E�5��2�B1ObEQ0���>�6���e�cD��q�5�21.�Zx~�0�d�/ӊ�ƶ0D?:�A�3���I]j8[3�{��Dc4�_��v���0�_�� //\1�_�IU�	����S���Nh>*��	�����e&c���k	�f���aX-�Ф,0M$*�Dw-P�fG�Cj��8��
/���m�~N��R���t������U����N(�`�g<�K	�z� �+�S���޿��c{�i���j����L}�U(��2�Nz����E�)� �O2d�4H�TʭM��u	,�_0:�w�t���Hj���x�n����n�C�ݾ?���f�(�VG����{_�����cy�	Xo;/�_̲�}͓$���0�y�+ի��+cl���.;H�%J(�&U�r�zkn��"�]c����=�ޢ���Rw^[v��)B��SW�y�ޠ��t>gx��G�U��=�����X�����|ǧ
�2!�N�,T$r)0�'�SRr��&��dS���Z�=|��Dx S�˷�!��������)��,k����ǿ���9�hE������V�M��Nn^��ߟ���u�)��7���Q`�rq���(/�Y�QLa�V7g�ĝr�c�ABQi��2z�ګJ$���8l8q�:$��¿��Q�=m;09-���_�* ��m����J�'[7��
��4F��a�;Ȑ=w����\	�~�<�>������ˑV�p��W+F,��~�W~,�[�M�n��((���9Ho��\ad�u�l]�?�����n�{�H:I ��& �[~9�����0ȷ�0:pлѨ 2���*�G�G�m�=����� 4yPƐ�AR��#1�%ߌ�ɞ�w���i[���;[(C�y�e�����(�����Cz.�T)╈�\ʠ{�:���S����X
��]��)	a�o�����P-i��Sj�=]'@�)�Z��Ku�ƾ���;�>�JG^j���T��2��_��Ѧ�ǯG��Ȋ�7��k���ؕ35��Ӝ4ozy���a���z�<n�~��6�S��L���9�����0���Q{ߓ؄�fӤ���>�ig����*�u�o;�(����u��j�F.q��m��U�y*&���.��SB-7�5�;�oU��M	t*����24{2���a�O�L(�;'�}�����O�}Qx�C������K�y��19�ا�wg�(Xj�ڴ��(#l��Iœ`I2���=���^��v~ۤ9�SY"�gV���0�؉���Xw�Vh�"�w8�揤�1���ݩ����%�$��]�5�Y�X�Ui��"���?�?6�W*�]|��Z�P�J���|6��*�����3-�{;78�M�0lHT-4+�eq<���v��G>�)�L*��Y�.�(��d�gv���T�E��%I/���D�cn�K'N�2D[m�ɢ�W<����g�)ES�Yg6��Z؜B����ޔI��C�Ӊ�~v�����D�qJ���kU:v S�v�ǘ8�Ϭ�����:?��W��p��:p-L��<����0�j����h	�/5ŗ���Th�U2��,d�7�½��~�;P_����k~��g���E�������8�{���	����T�z�Z��_��Q��΃~�3�t��9��	�W�|�b�V�N�l�;�(������~w�AsN�|F1�Ѷ����OJ��~�0�ݫ��f���S�R���i�r�E�uU���}��FyИB�yÉ�l����J踨wXa�%�x��Q��P��^7��i��L�)N��Sʜ�&D��$���Z�T<������2p&ܯ�ҫ)���֔U	��l䑥W�����	wm���56�MT�.w�-΄H��G����Ԥ?	n$�c���͇���H��{fEK��)6K?r����K���it�7Tk�23�܄��[ne�w�@w�8?��$���+^W����.�kR�30G`l�t�,�'X�|4���13��=��A��Y�"���	���I�'^�M'�{�B.fT�����re�8r$��.�}~���d	퀆f�!�u>�2vj�a�Q_�wI�T;�;�K��'i�ۿ����n�W���Ɉ�
��>�.�V�4�%3gp��#r���Y��}Lކ�r���5�T�r�N��I������m8֩�D��J�2>�{��a�Խ��c�2ʿQ�Vk���-�����K��짚%�
�=��*����8���3�pk�љ���Znj��K�ݐ4��|�Z�Sat��=��ɵ`���������`ƙ����O�(�5AεSU�bY�2k��1d7'5�%b������[�k�ۺ6���х�Y�!iȽ?/����U�Z{������++ߖ6��R�G�!=���D��uW�$�~��בX�ܜJm�e���hF?:��bN�n _���+g�(�5�q�آZӭ=Tc��9�SV�S|�T&���S, ��3h�x�}�3]*�����K!��+�8	��(�L`v��\�B-7���9Y�R$s��#��!;b�np�h��β������=��
D�f��B���ވ������ e�3MT�tcʶu�̠�/�=���,�:�*X<�3[�v��=}8һ��M*������q��;3���E/�ss��R4�E�pө� �k_��cm��Z^��kj�\��z�<��Φ��P�rTKڣ 
�P��l�Ԣ�i��&_����?G����^cY��ڵ[�D=N��TA"S=a�߾`3S?����@+X�@���ꮦ� ��3���1!C���	4q�����B���{3��B�$��rs� "��̽�#��w�J���,�;/,U�+bQ�E�q�-�ofO#4x��z��@&9/��/hV�%Ճ9���0���ݮ�kc�4��������[[0Փ�O��S�
;yw��l:F�𘸊-���������<��D{�)K�o{���o���oj���k����3w[rU4����!_6q�~<�����R�����5��G=`G h�V�3;Ɣ4i��Ь���*�|�
g�S��jPK	��	r[r�I37��Ll@f�����]�8���c�^�>�0>S�]�9&\�Ǯh���p����miz�,����T��urW-��n9���u`S������	[A-��y@m�p��<$�J�܁�yN�~/����f6���r�za$��z��hN^6�G��B�D�A�4��w1j>� }j�@�;8ce��� ����"�88�Y��V2ͥ28]�Nv�wg�O� ��R�R��Q�H�ҩ�i���y+�:b]R�e#�1�����8���d+����y�>"M��*���W�ۙ�q
X�2>�Đ�܁Wе�W��B�*7&�I�Cxe{�n�t@��3L��i�;D�+�Ɣ��*����Pn�s;���^����X�7��Y�0nN�l`#��(0A�Y��DSο��hpu5wՂ'!��!�����{�?Fn�:[�ң��
�ٍw��o��j+{��M���뾈0-�I�є�%:z'F���*�^u�ccf�f!&���� Ld_��Ɛ���3�&S1`Ô���`K���*P����)�,��ٮP`gRg0�SH���pH�7�ϻe��k�>�7<��a6� Q��-�Ҁ sAN�U-�2?��BtOb0�8�qYO;ѫ`n{�X����$:	�Jם��\�R�C'�b�aZDv�f��}i��3�DR��}�O�Wa��D�R�(�N�ޯ?fz]�H~|l]`}���|�Y���A�
��r�R&� ����Sd!3�)�W	VJZ�
h�g�C�>X8I�����9�@9p��p=eH� �z�w�k�7����@f�Cm�s;���'�~R��g(X��=�)7{:[�h��6��\���axU���ġ�����B��r�3�*�����o�xp�ǗC���ˮ^-�ê���}o`���Q�����s'�6���ӽI��j��(��;��F�߁���BHMɜ�(��A���HT�wSL����U�$$�΂����f���z�W:��3L�J<�,����ۈ}�ABՎw�S!��i[���8SGYb�[��acs�]�lBs��j!kd��x4^��~"��������H�/����STT�g7C�i'��	x�ጆ�4&Z}d��ᾟ�U��]��Pl���p8[ ų�'h.����[�=�S��A�8^#5x�R!Q�&I��z��17�I��{�fC-rQ�k�0U�f�31l����cɘ�$[>�*�uCq�%��=���}�ڒ-�e�O2���˅������{��L�|m5�}!�5Z^7(��L񺥂�#5\�G/4s|@����h~'a$|E� �h���jKrp��l__��f��W�N�n�E�e��0�kv�\�7� càj�N����e�����=�O����Gye�����tX+k�D*ca�8�O����Y���]$�$�6�rV��M "�����ԦD���Dtf�Tލti��>3����Z0�bvAF����r�r�i�Տ����UtϦ�%�	�3��j?ZD��q�߿( �F>����'gB����U���{�!a��~�u�4|�����>��;��|w$�2eq6��Ѷ��Ǔ�Ce:V����c��z͡��Ƭc�P�M��+�ǹt��F;��م�[:|�|��|�:��)?�SFG���8����E�a��G¥]�=Һ	˳NJ�.o��R��������+fܜ����=��b�j��*)ٰ�<�m4z�I�6XZ-�,���9Ǹ���H��Ab����fn�U�xy/k�7���f�&�X�Ic�B�yH)Q�}[��������U�����J76-�����t�zu��x��mGI1v�㬢�u�=�@����@{�����C����V��'�����݈�����-m�4X��?5OZ�=ϡp'�����^��ͩtC�Ӳ��L}Ȱ�?d��M�Ib����ʋ��5ÿ=JtMc��&]s��J�`eo�R5p7��|&t�L���J�|��(ȅt����T��d�h�+YW�7�O"�z���=G*!�	J9���8��2���t(4�U]A|��<�7�Uk�Gzy�rPޒA�QE�0��� �惒#\��'�s+>��c����J~�J�y��� 5�p�"��dU��A5R������~7}�9��fY�0����[�z��rc�3��!x��,=��1 ��]x�4B�bX��#�/>|�x���J>�#ͧ�U��Ĺ�K���<�g�����>pzg���'��n/�\���VP��K߃��$~u�.0�s��Y�'<+�(]8�ݦ��0�@#��~��ޭ�T,n�4V�NS���@���F��c?,\��Y�s�M��3}��b��o�X�b�����ڈO{7������Y �;䰁��;ʽ�>nVON��t$���pw�S����@B����u��^�O�����s��!z�U#t�c���Z���hq%C��1_F��kzAސ��wl�YK3�.�1�/��eN�Y{����&p5����L���݋i�d�Y`�#؃x�ߦ��$j)��҅�v�ʫ3>�zI�p�1�J��^���TE�'�*{�'���q��T{�$��4���)�k�n&��� ��fi*�+��ޫc* `{��T���T���X�b1T��	��V�C�=�����2h�?�۴�i1 �o-�	�C9���2�[-��Q��Wf�>��f?I���lPHSI�4\�zoD#���ʔn��+������r8X�>�@��[���a�D�����Ά��Ԧ+���.������Z9K��@x@\��;m��/�0����}���Q��i�N���R��Uy����PS���j�d���H�O��`vE�9��Ny��ՅR�H��x�t�����^)"λ���,nd[0�J#9%����i{{켧�,4f�\?���\�o�!�������,,�U�g5]o��g���9k�N/�Z$??˪�a�c�mb 5���Td�Gݩ��
ο18����̫�w�����`X
;�oꡝ��=��#~�������	�v6V��Lh�m�'YwS/��1�oHQ�-ᣌbj���:��?A��?�ۨ[�D[~(;��+��^ J��t )^5��]Ü6%,�؛����\�bH��=y?���z����#;Z�f���[s���T���%�{�w��uS2C{j��Cr�r� Õ��b9y��Zӈ��>�����G���q�t\�1�=`M]����p���m�^߯hq%���#>5�o/���훅����Tj�ѮH�Щ�δ�䕚�Hd���N�j.4_<��$>��&�T��H�=F?�W>=�~9�;�ZGKB��T�3맕zw5�L�����v�[� { ���;���v��j���O|`�lq"1/@/���ßؚ΁]|�!^��w9�{�"�rŒ0�N9�f����n,Al��@!������? ʝa��!���G%-y
�̏�^���'�(}�O�i	C˾b�>kh�)��	/��������*`�)�Q�r����V�K�Zx�)GUY��S�8j;��X��oo�Ѿ�k+R��3D#'�6��6�k׎������6i��;�U��leG�:(f�!�hu�կ��ō�B+|�J���i�+��e�kK�5*��歡�k��	H�xڷ4=�E^��͝8�9k�>#t��=�Ξ����u&�������C��J�D:��!_m7��io���&4���rO���|���A��2��m�&�a�<�+���_68z���*�P�ߍ�$��C���p�3��ּx�7�ߋ�'(�n��V��o�\( �{�F�
��3X�UP�A����t�P3�Cb �@�C���P��������p�2�Q��+&�rv���c�"U/�<��q����B�&Y���B;�,U ����t�bC>	*ڄ��gr I����'�Ŝ+~���wq�5��w�����[�Ia?.ۿ����s1�)P���i/������0�{�̓=����a����LJS�	������%7�Zɯ�8�q����i?�a:|�	���UZ��W0�a�L�&b��^m?�ma_:f67N�8P���Ǩ�UO,���(�5լ� m�(D��~�Vk���%ͣ�|���"J��c���܉������W>��P�9偭0���Һ|�D�*:M)�|誌�pYG�^S�0�vy���2���3��#�B�R��ƿ��JJ�)<�g�˦��{t$"�j���;�NY*�(��}��Ov����׼^U�S[���:�<��Qjfc��-_�'}v�����#���["(�6ˎe>���� �t Pw^��~�`H�z=��W�.�l���Ėa�yݸv��%�_��K��7zP��Sw����^�mD.��(K��$�qy�L���Zj\a��mg��ڪT�A�&�Vڹz�/�9�v�43��6@��"��\��}*}�uR�s��Z��	�%q�������H
�{���g��� ���g
���>��?���5�ڬ�z���{;�D+k�3� MXc��������}[��j��N�Y�w�(�_�Ѧmz�~9J^NMi�W���
�K���+\/���b�����3�^"t�H�~}������|ۍt`/�7#Z��{�O�/_fV��5�dx�n�}�5�5Ϧ�g4�w�S:�$�a���"����D�zF�s�*��Z�X�Irf%YY��o�Hb�aB�_����A��V���e:�m�p�h}�Q�i�V�<�4[8~5�Wq�![5ba�2z��!��6���=C��.+PY��EdZˌg���_�i2�3(?��ĸ��^��e���&��\ =�� ��:Bv��ɏڌ}�¯i"�sQ�6�WwL|�˯�1��(�ܕ���]���]�v_�`Op"s9�ʤ�2��T~�ɰ��&z���/��#ӄ ���x���L��ִ�ku���3�拓@����tP�yk����No\6�PAG��3rE��yi_�ќ&������8��R4�UZ�����&��YC#�m��֎� ��v�@�s�3X����:�@��UY�F��'xj�f�{��8Y�\s":�R'�J����	!�<�_m��0�[���3����5#����u'��������hk�*U�>v{���;^m��$eq:Y��f�@��9��O�5j��uo`0a�-�~�K1Z���q�[�g�?��Ԟ��<�$��j�����Wyh���s�Dӏ�hX�)W��8K�/;��[�ש�B�=!��^�&� ���j�ǫr�*y��s2�j������n��/����a�����7%vA�|�0�)j0�Ev����^PSc�mv�Q8�ہ���1�E�j��v��n�	
�yE����ߒ��C?��R�wJ�&��ΰ��h|,���`����y�p��t�v�?yb��O�'���{
[��ɕh�摊Uc�J��Q�L�R1v���H�px՛R
���?���˻�G$���u��v��~Wڍ!`�X����:����\"C�ZD��*	��$y~y��'U�"iu��8�o#y��~����^�Y:0�5^O.�C'^���ZI�D���n�2G���l��&��b��aҝ���74c�	��0��<T�K�F�\t�w�$�4�wHn7�3��
���6�{��D*� I�_���1eA'P���~N��9��3*`O�꽊��]�Q�����(w�^ם���^���d�/�q���5�
(h��Cμ9�3�1-�h��ݹ'�	�ƙX��oF�����|��w =o84,�%�"8yvMH�k�sd���]#���e�KB9��F̟{�ȭU���(�AxQ�᧎8�Lϝz7��}B�rrj;�v�M����R6�݀2��t�-�u��H�dz�|��'.6mxgk��S�al`Ǝ���C�J(Y{HKw �Aդ�M�e�iy^��W�t�����q�����9��l#���t��&Nf)��֞���y����5Ɩ�p��+��Wy�d�� b��S#�݃��1�@ItV#�T2�е��y���~}z���[L�lᵧ���!��Ik�۠��> ��<��=[��h:G6�\&'�.;tE\����9!�������5$(�����&�zc���ǝc[���.��]���ZQarf� ���1Ω5��D���q������#��*�szE>S/�2͉t�΀�&2^�y���/����\�`cВ���Q�^j����h�vd��%�x���ǸK��N�pr؁��!���RHs0�<���K�;�l����]wEq��ɪ}�~nv�9@T�]���FԾ��ӷ����5%�MTu� �AtP!�!�cߩFoiY���<?nK�ѯ��e�+5>���AH�B������5���U���:�C!�5�����h�mr �(�*�aJ6]���eZrg�M�C"�$Xj2���
��m�a�"��W��T�5�q΢^�'�J��h[cwwJ�k5�*4m���dq��<���=�*k�m��9S*U�a�+���~P� �쪧�����vg��r�����{��n]�iL�/�\>V�_8��=��u1��_A�]��ҵ&m��eae0�f�Y�z�d��i����1�a����r�w���;G�`�l��4�J�DJ�
��_�XJbl�Ń�^��f:)L�!Ї�1P�n��	K]����L5���� �e�z_��#&~���9|�Fc�zMG��#��(�;�%�0���cγ	}�DEB�߱��'�\�d���� A��c�P��B � k|pb�Ț���m��}.]gP�W�"yoy&��]I�A=�<G�p�������7uA��s&{�a)L����p����N4�eP���]]��|oˢn�X9�P�B���+�~��1ŮR�Ԧ뇑l�JW�_��Ź���Ai�5�5/������<��MQ��S�E�`��	�V����Y%ѽ(-&�H����-ZY}����jd?��Ir?��fK����5a��QMȝ`��Ab\�p>A��!�U�] ob9vA��yz��;s��ل�ͯ���Tv<�d��|:z�Z/j���3�M�R=٭#�W�^g�"�~F�j�a��u���j��.r_�ӫ���V[���4�ov:t���P���d ��s)MWmN�.f~��UZq9t��pOvQA?� ~����-hh�%sd:&Goxu �-��hvZ�<2��a�j&	Θ�L<6��F�fNϼJ�1n��{�� 
F�et���|��������)��_1z*�\�T{#�fK��C߅1|�n�(�w�)���soh~9�;x�V�jB|A�vu�\��vX��& *����l��L�3MM��R�#1k{�����dqM�_����(C�"RE�鼉K���CyZ���ȲC���}qǹ���s�x?V����b2�3�H������Z/�1���w��V�y7�d����`�l`���+Nlor3�(PV�������oۉ�tY`7vR��C2��Z�Y�t�߯� �29J�s��|���0j�"��.��U�
���"�0�|[[\�=���y4`���;ܿ�>tFs-�
8w��<��Y"�C���!�b�B��y��'�^?Ԥ�$EdS��L#�OJY&\"Y�q�gI@8����[֟5G�����G�����6h���δ$�|V&l}��;v��~�)O�֗C�Ns��BZ���cD�Q�`L:f��6>���I�����!,��X��z6��X�1EM���V��b�X�G�М��T݆Sd K���|^B��"f��R�Ѻ��?�1+X�-�eZ}���={��'V��~ϝSM�5���ˣ�M��y1f�)� ��p
L"����d�.��q7�U��6.�k�1�PZGA�y<Z�,P�4 �᪀K�z�������[�h�s�AP���B)��&��ͣ��Y#�S�'F
��,��"[�ax���7�&_����$�rg��H���pW�+���ӣ7ŵ��9�:��th�9�{h<��J ����#�16��؃R�.M����jч�r	~9��<�,���4,�5�4KB�lk�
 ��u�Z��^�C���!3�'ub6�*��Kئ�c�qy��j�\4 pO��)����
��A���&1���~�UB/��ɦ@�S�	g��:�&�s��W]��y�@N`z\z����I��˺��֥�x�3�C%�4�	��$s�����x;L����h�K�q���_ԡ�P�"G���2���y��phs���ن$G��.l=5���c)�Qjw��z�NZ��S~��8N[�s!�ߝ�[m����Pݓ��<G�`��M����<�Dq'���w�a
�M1t	P�V+�7Fov��+��~�82�=�/i��E�ua�����Q�l�g{2�����q�"6Z2r��Q���~�ajE�1��}._Jps¤��xw<���e�PBcg|g��Ϡ���ֲ� �F%�ܦt��*�����C�R�e�Qz��"Y�e&�A�{0�u��
D�FZ���3�}�Q��A��-�#��ʆ�r�n�_ot���cw�܋3���O?>��wh���ežW�橹�,�I��3]��L%r�g�-�X{��������ྈĨwz﹓��U�j��3l6-�p�Y�4ׇmvoڝ�F��,�A�}*0�*������R34�=��|a*�r�:*���Cj�4b�Q��L�>�(�1E����]+!��R���_��Qo$�r�M�^H�Rz����(T6���
�G�eZZ&$�uME�� ����ڲ�ߣ���e6{t�=�f�)�qGE֖̖A��A �c���m���sK�{��Cp�yTr�
U֙�~T�6!ݤʘ`���	�A��셽}+?8���yR���PX�K�dN�����(P����S�y��+
ժyOP L<�V|II��4A/i��*Q��"F����D�϶Y�F��]r*���.pw&ϋ0!ei���<��(��27���g��8�$O�bu��*�������d �Ib-A(?��`nt��6*a����pgZ>�1T�j�\p��r���:rг����a[r�Q��,��`��m�!�F3e>�<n�&�K������3���s�T��0�IL�$a�J��'��L��ߵs:�+Iz��@
���; �&|�����FB�L����m�%��(ړ��!���p�ebw�(�׷/����w��2R�Me��ouԚ��֦����]-g_�+_v�-�= ȕ/����x!� 	�[,c���P�JZ��>,X��&7Fq�AS ^��c�lvF��� b���xf�nS�a�#�Pd� �~KEE���\٘ր���~=��w�c	����7 ����<@q!Ohr-!��M-��=J<�8�RP�4KSg�1F�9~�%�}�ØF��z.2�uh2^���*��xOh�׹$j�hLqo-�H])�c��\���:�7�6�;ݠ*qW��dUnMŻ�1*�̭�u�偢[���Q�� �f��"N���`R��_G.��*�+�g��kO�xzW`�dEF���
�?v���-��Ǔ�ry��H,�����l�,���h�u�p��ظ�J�F����&�6�Mv�o�`y3��೰h_����6�ܖ�g4ǎ��:��N�����X8�����
�z����1���]�3F��%Pb��f{[7|�k�;QJ�y�鬝;�w�t.ׂ�f1M�l�f�1�B?���d�?C�o��oO^��<��H�-&�N��/��Y찍���0�:����y��Xq�C_t��P$�'��\����
���F簛�l�F��W��s?+��O��kR���tz�ƔR)Q�M����PgiNST�m�n�)�~�:>�����&�/'8p<ꀃ1�L��@N��<�4۟4�����3�̎�9����|v�MK�q��6p�����Lc��E�޻Q*��˝�Ҥ�q�vɉQ�Lx<�Kok.�άl����W��=���mf,Vq|��5'�r񮅲ihk�&�[�?dV$H����k�;�������n�%�<��q3�\|1z�o>홌c��\��Ϊ&�՚2ݯW����v�5�����y������;B�U���m�^Ŀϫ�a����>���7V_D����$���u�* ��(Z$��<T'�y\6�CP؅���78y�B��.S;׵�x�����*�.3a˪g�6�M�(9O��6�b��c[#�V��i��@�~�����˪/�Wr}��Vf�\ʀE�4V9P6�×�_�&�wb��vjh!"�=|����P_8�6�6����ރ<Q� <������Ό���Qĥ����i*4����B��w�2Հ� �.�I���z�#��@�0$)Mؚ���~Q"�u�ד(iw:�\��eQZB�%�dBSU�xa����`է4A��Ͳ��C�C�mcW]�o?��VŒ���!�րU����Fg�M���I�e���X)b�=A����
 )����`�Bh3nJ�������Dk�_z	(ΪiDs�f-��&�����H-�/lW�C���4y!}^��gry�#;i
�)� uk�M�5M������C���K*)���Nv�D�pq���� ����H=t�ڀ�U��[�L�4q�q�)�F�P���Q. �J���0,n�g�V	�x�����]a{*��.�KaB�\�}�p���&�ct1!W5/Y�=�癈._������2�͙3�:E�����w�� 0
%��8�A������3�ś��|Q���_V�d-�뾚��B��]�9���Z��H��[m�;���f����G׍���l�^wׄ�N�%��:K��� �d�'��5�cj|���9����u	T�9˯9_9Q��3ᔑ2vL.�4d����R3i�`B��U��@sj+��A�e��rJ�;�Y��i��l�"��B*�Mq|�LdY8��'�`�{�}n�m�X����m���@$w�w���~�IƦsh��_��&���7q���ǲN�캋_E" �i�^j���F�u5�[P���,c [MOQS۾dR�	��j�������V�[$�;�WES!i_�!�u����~6�2l���;�"lʞL?���#�k�ئ =D�$9Z�i���o��C ��ȸ�U"G|}���W.3��N��U	��];�z�k�Tt3�^@�`��U4�X�]:���@�D�W=D����\,>�ܔ��ߘ�r��9e!$��@�]���	��+^ƾ���]dC1���A��j��$P,�۳T'�KyP���2�G$ړ|��|":�{�)&�j�Xo0�Qz�ނo��>�m�����"#����7�\RP�!�K��N����S7Y̥>���m򺾗�` ��dV�2<	G�� $����~�K9��(%����Ac��S����ă����F�Py� _��7м��;��[I�Nl0�T����SRmB3w�?n[9�д/�8R07l����>���K$lF���o�S�E$�xX|��*$������8s�F�+B���ߝ�*��#��-D^��q����4�8E��+�w���w�Ќ�����;�H�q;n�mǏk7:�JP���m#N�K�lvR1�YZu���P���K��q��i&����ږ�A�ѻ'\-f�E��eO��*�+{�����#�<*[_�2�u�;KB�tS�i9�b����|�#8�>9O�l�C��鳍
�(u���]�I3�?��7H`y��v
$� l�;��4�Y)�!��_�~�J�P*ϋ>;�2_`D�&�Ԕ�Ӧzh��_
�>�?y�F�9��������U�r>}�?���q�'d�1"��? Uޯ�BYPk���暊��yf�{N�,���!��N�}~"?��7�Yh�tP{�\t?��Ii���gϯ	���pr����S�azF &ׁ�+6�~�͡8��Y8hsb�\�sSb�l"�ĥ�� ZNA҃��8da�*����|w�v<��o���]���Hl��V�jQ��B�zv�:��?0ѿcc�1��0A3�	�C��������Q�X�w��|ʂ�;�Ó[��x�ɮ�>͇����b�=�m!͠x�����/�:�URD%]�є_>�&f����K�D8d�]1�~\�}�G�4A? �ԧO1j���ï�-�r^���?�MZ��q~4�,|�)*wR7_��R! ʴ��@���.��!S�`E���-��n��'��8��j�lK5Ѽ��Q+1��?r�A[r�5Q��G�N���@^��c�i0�S?���2�T9;r⿴�N�m$���F�C�BXGz�򆺮ّ����u]<��p�Ω�تM����`�-F���3g���-~�ƶHB{�]��UI)Le���66�[#,�Z�8�=�G���XCD%��9-��蜟 �LVrL�\���&�����j8TAЖ���S9ﳑ~L�䗒We[�{x���*��h���-_]k�@_9� �`.s�����cIg��2��@3Q������iqOT����߷���I��Th\����=G���5@��ǝ=�-�M��IZ�Li�w�)��(�oG(����X�Q���[4�����J(Ҋ���X�*��>�.���Ê��}"ɡ��\�p┳���zӪ�<�*�Ju�ϣ���bpO���S�^���R���Ԝ�ś�p��ke���?�E��	�?kG����e+��g�<ЂM]���$ر}]��C'	0��:�>�/4�-��m��E�����w��K�?����W� ��x�Bg�����_a�Q]��Tژ�->�,>w��Ud�����Q�f��f���:��wR�)`��p������ex�F�C9%�0�D��
�Ӏj�Qv�����9
�k��cotג�x3�kZ�4���?�R�%L@��~�Z^���5�LD��ՄН�l��G�\SR3�>��X�7ǫd�4��������^&��i�mg��zFI9��mm�]Э�O��m$1���ʍ��^:tw�0�YּX�"�8��x�68���EL���0f\�����.�'"y�G�o]+J�Wc k����"��a��$�}�����8��\����4ڋ�U�pɛf�$��G^�z��Cj[���7
s|UVK�89g�y�f�)a�}�\���e�'4��|�Xo�ƽ{���DC�9��W�ы12���/ބ�x�g��j�Qt� "�N	��ƣA��i���\V9��� JϹHV!�ֳ�ָ�#Jc�P�d9"�*D�"�2t�H:��h;�`F��,�s/��xI��������
 !a��G�g�S �<#���b=�L��ޜR-G5w۳ϫ,�{(L�o�r���0� F�
fuW��mlw!����13r�h]�z1���<9�e%���-q
%��7@?�i� �ot���g���M����ŢNR��>Lum��?Ԩ��Mz�/TL	�i�*l5�P�煬8<@�5�0����7����%J�īY��8���݁G?9��@�I�8���1���͞�����K8N|w�G��Q�ڞ���hB�1��aCI��*�Q;seoFl�d륜�j­�N�f�@lS�	�aK����O�[">N@b'%�u�bY�jX����r�1|��|Hp�-� ��x�ͅ�a�`�l5��|O�1k(�c]�)!::���!>�v�U�Ԡ�E��4>`
x��kf�Y]<_p\���	��)�f�������%�W�t8^LU���z�A������(K�|b�4�%gaʆ�����N����0�B����<��<rL�<Z�d�&'P�� ��v�� h�yc���@�vb:���ie�y�f�ӽ��q/�C^bnua����q���.W2xs�E��T��J�x�ᝏ�C�$c�>�D���Z`(�$�-� m^^o����>��_�[�F�T5|@Z�ט3&��q2Y����좢^��?J��6/�fմ9+42� q&����g��s����m�'�]�`����C{�FE���C����:FlgD[H	�����k#o<�R?�������E��r���­�e�/"c �1�.j�pF�C�f����T�A�|�d4����C���og�Uі�C�)�!��&G)G�$'�C���b�	C1���S�Bh�8��� �\��N�[���U��`���]�"`��4�	���VO�M�/+MA'��@D� f�)QiO��LLP��M1��� ��T[�JZ�՝��쏆��{�jd�t�p0�8��*4��B��s�3<�Z����e��]����S�G����Zm���n�P ��g��7���֝d�y����cD�*�8���؀_˴jo��FB~h06�nL< Ek-/��S���~z1/���к���������w4����EEe�yO�y�łoɂJ�g�j}r�H3`ܬ"���xۜ��&�̙�v��ԙ\���Qo�����ߏ7�JӜ��Z�>.I@��TJ�\���o �|@�ǒ��6Ka÷tJ�@T��"���s	��Y����aƇ��hH
��Q�-5/�&�]��̲�udh���pm\ꥠ�ߥN�I��l_k����Q���X�n�����y&
qsK#�)��B{{�Z��0��i�4�ܫ�� '�v��>s������N������c�)��Ѩb�V!8j��c#��559��J���uS��"�yZϻ5s�Xܘ�� u��4C#�N�=�X�]��]����\��Rxp&z�˳�g$�\�DC*'T�4�g�>#a �-�0��3��0|f�����=���G=e�ru�Ӄ�]W��U�	�^iB��j�i<���r��ޣ���rRe�[���]�T2�/sːfܘ��v�@[���6���lZe�tx�9�MT���U��+z�{u�67PM]K^pDм�Ƭ�x,���_[|>���H�7�=]-�NA�sT�V~��p,a�}8�J������'Qpl�^sa���^���-�-�AS�Q���ӣƚ�<�l�F�r;C���S�*�p��ْu����$�υ�Qf��Sѣ���hh�T�"�3N5����6���G#��)%!�/��?b"����
�v�:�^0ڡ���F�Ȩ�q�`��&�����������F���mN�J��
ܮ�T�웤�"�i��Ǖ���9	v�dBH	�c��_%oc�N玩�L����m���9��K��}�EpQHF����x�ؒ�F[���K�Q�]5���ʓ����g���Ʃ,.��c�.{iK�~�/3�d�Zn̕�d��o+��\b�d�Ҩݤjh|+{F��f�n��h�s1��Օ�����B݂�iF ��!U��e-�#�S~I��U�Q(	
�8 ��~FM)��rz�y4���drzT!nW--��.;��K0,���1��6+���4pP�`r�`8_L:�k������#��]��K{���'B�IW����J��=|�M��,ڣ�YA�}|��mޜ��&��2����%,�i����<����J>8�����m��/�-�,x���Qa���a�\[� �2N�#?�e
�!�f�S���+)(�z�h��=�}�����nյ�wCD���؁Å�`[��MQy*W ��ǃ$��6)�Τt Z%��⧌�!5�d�+�$z���OD4��6�y�� V��y�@
�W �3��:�MW
�|6��~�;i;������8g����~z�X�����U�܋3��FQiH|K�ܱ��Vq��Ђ����\�Y�52��[�PsA�y�֚+�	���7C��T���s��U;�e��U��%�;=���Q��d5�5�Z���������vJo�X?�^Q(u�Y��O�M�z�k�S�BsNQa��̕���w���-���N�;�"6�^g��De=~����H442�Q˯Z>���EJ�'� 4��*��"�n�4�1�8X�ꭨ�̽#=/vyW��I	���M9�~��X0$�~Њ��ؔ3��s��
�p�"��6up+.��:���9t��c(�B��[���y�I��"��DNB�R�JVj�����g��y�r�8P��U��̀�1���#�2茴��:*��7.�_B�{?Q}f���P}����YE4���j���jUd���[uoCHp5Ӡ��dg�"a�Im�Ny$?������< y��~�æ{J1���2�2);M:��-���n��\�����D%��Ƭ}` Z�	��P�M�oƓ����i�\��jT�p/ԧ��
 r� �y��mNwa�t'z�\u6\�lJ;�n%bNT��`��v�0�t^1a�:׻E�F�	�����azO�g�%��?�Eɑ1''��u��B4��� &߷忳������@!�y�\�\����K�3�m;��}����`��S|Bӷ1cry��S�������������iȹ���x�w��W��xR[�,xq�4\>�#>������(2c=lI��!��}ic������U�B��yt_��%4��N�<?,�
��@C� 2}��_�#'�mJ�{�dREnI
�[�<[p�����k��M��P���v���j�2�|"QJ	a�@�c �z��,�!���W� -0��p#���U��n�an�s�'%��FQ|N�����?�?�`�<["�дDT�(\���Y���?n��MD�8o�wq� ��MU*�0��_��g��8�*�*�"*]d��S�>I���r�Z�-�<�nL���L1.�33���_��}�"��u�	.V����gW/��m
?�f;W�@��HX��)p���1f9K�,��n��e���\��?ʚ]z"�E��]�<~ �� �e�ei�<���&��1�oz膕�(�R,oq�	�D�� X���"���K<Q�5)u|�w��\���E�9���������9����+�^2�~	g�p���� QZ�|� p��L8��W�X�G����ʤW��ƛ�3�+!�s�\mщ�����p��)�"dQA@������]E_Ҭ��&��f�ms��tw8	
�%~!vҋ�k�!�a�??ͱ��)4̈́
�X�U������2'�Z]�۰G����ҽ��.� ���cz��	!믗���%���9��7ɵ�Q����% E��Zd�ek����?�	�������X���c*�ǟ(�j�7��D+�W��ye;�^�{���d8�/�P�](/V�27�j�����<@ET���������S�m����w���\�TDJ����$F6�.�8�L�� T�ˊ� P^�n�V�*�j�d���`��8��9Uב� �T�p�^���w��O�\�	���>�Mi<F��1�i�Af���΄,L���&>3�
��h������,Ls`�
FE��B(c�_7sVǺ�1=ǰk��Wp��s3<�c�shqM���Uu����	z}�u�`e�umt��>�*[�;�>��_%Oyp�q;�D6���i!"4��?cL�8b
 Rx��G���Z��[o�����6<� ��K��Q��n�:��M���������R�CX�,�k��z.�4@�KL?^b,Iv\�)=��[�D.�x�|>�S ��� �A�ҿ��D�J8\���:A�+�{����P�>�Ǳ��c��@�O@CU䵢��G���_�����N�U�=hsI�mOMwI|R�%u�7!�;N:/�߲j�&
�bm��]C=����ϸ��ltJ��\��~ԩ�$iO|�0j�2��qA<��L"S�q�-nw�y���V��˨�x`��-o;�|9y4`Bt[y�TFC�J�k#/_M�/���7Y#
�qM|���EFF�ѝg^x���J�ػ��[20�l�T�޺,�2Mb��'a~ �ź�ic�m1*%�:��+`�qc�����ǭ�gi��0����^�����g�C���'��h�	�I�-a�Y����<�yD�h#���A3�2"�8>&ڶ�h���j�]�K�{�{�#���5�׀�G��9�C��x�yco=�%�\rI:�-@J�D�`6l�i�S+�kX9��@[�/<k6%��ş0y%,Ǜn���@ ����#˞B����vדB��G%��p��]��x�����U��Ɋ��+�q�EK���̧�+,���礪�
��E�5GC��o2��&�RzqBH�Y��WY���N�2�
%�q�w5P�Mh�VbY���/�ԏ礓I��$�
d�{fY��I"2lzφ+�ȎBZ���	D��ǏP@��H>U�i�9b��dd��f�S��g:P��R�O�qA��g���!�jg��������IĲ���H�B�������G�/���"���P2f�%DQ�<����`�Aq'���FA]t-5�Q��� .�_ȿ�6KC^��p��ݙOv�'��V~ɼ�{x�O���_����b��B��\�J�5K�9�k�Y]��[D;��Z���T{;�ѷ�����.)�8f�ݕ��0�
��Ҟ�lp�OJ���>��0�:霿��
R��n?��͞e�t*�M#���
9G��r������4� �Ʋ�*�?�JS����	'��� 3�����½��	���ԧt���Y�	�"�����{�ӁH�y7ua�nL���^*`(B"�t��M(˅y�G�ڙ�ǽ6��Q�]������e���(U'P	�e����><�Ԗ.�0�ئ�h�P_ Z:/C4ja|"DM����/34T
���\�ʥ�7�_i�:k4��'Ǽ�$N�47��yl�瞰���a�����7�
 o%��"���v+p28e5;�I�l�Ȭ���R������"ά$ch�6��e{GyPYxk0Wx�'�">���s9�)R��m�0TѼ���/k��ӊY��(U�,���Ph�d/G���ҳ8;W#1��ўH+����@���ͳĞ���6� �y̠r�#��,7M0�U��������nT��n=�h�<������^̟/\)��K8ʯ8��_� yQ�)a�s�U��:����Bmq��Ν��8�IW^+.��������S���"������2֩��LWoi�����dD��R�{����#���y�E��c FdB�9�x���=V�c���f@ �FM��c�|}��A�|_#-#��N(&�N=4�Ϛ@�o���y$�����,�G鱁8��Յ��[��V��4�Bef� 4_ ��b��O�<�I�W�#��M�ENV�w��B�g��@���G�`��ڢ�G*���q/)��Y�Ҕڨ�?�m;�<w�{bGL#\0/�����\ε������0r�_����cJfx@��ȐX፝d���&,h؆�ş�,�����4��-G����i��:�Ul�J�!���64$�i�A(��=GȎrIA�������,K�)i��LD�Z�}f4���:�E�K�)��	��ݽj�$yF��^��<v�R�H�R;��4���?p�Zt/޻HB�l)k5)�צ����X�H�@��g�v$�&x�������M�,1[�_,��]85Yg|4E�SL�n%�7��.[�dn�\����� ��'7�����|�ys��JӌA[#��� ���[nY�0�T)a�a|ə����<����MA��܋�{�����L(.��e&����T���Mu��k�G��5�0�����"��}�r2v�H��Y���81���Il��
��K�E��ޅ|eO�����iJ� V�h�Y�t�C+{Ii��7-������$���WIc	<�dS�c�=��F^qP~1�,rdtN�M4� �'�8ʡ)�p�1�0�&�zӸ�	�Ra��s�`EbZmo\Vā���U�R��)�R���D�T.΢�JqU�OV�f�1�-˂���6�a�M�+f�f���V<e���K�G������<�!/v<�}�b����Dwc��ٸ:f��8�l�x��yt+�����Üɹ+iq�C��6�,w/B4�1����Àa�=����6�3���sc�2y�UMа���B�d�������t�y ���4z�̭9��5C5�Ʈ6Ϗڥ������Y��D������.��.�)�u��~�y�D��v���ތ7�l��t��Xd8�F��ڳ�����8q�����l��6����m|$ی#`f)�2����D��{qN�Ϲ>�vb:?|r�y+b��Y۳�Orl�U�y=��j.H7�v��]��Q�L��L/[d
ݣ-9��b=����
��L�b���	l �~Vuh�P��� �1�> aJHqoN���tCktŽ$��^�r�a���'���\�_�i>F���_�}^���oه�/�l%�Q��y����_�~��!>��=�'8�f�!�Ao�&t����F0��.�O	T�'�l���4���طA������OGpQ'��+�����x�^�~��u����[�yl6����+I���NOM�W@�4�ͯ�܏�j��U�����'<*O�IZ���YƼԔ�ג����6�;I��0Q
��Vc�ۂ\�L!�ΊGAl򷱇����ę�RE�8�l6�c%� �zf'���#
����ea��֊e��6￐���|�������EDm�:EE�����s��,�[��愸>!r���P�/3K:��7 D�9ě��k-PH����<��s6D��I�,�鈝��D��
�+,�@I&L�u���W�0@VV�l�\p�®d�?�g�m)�p.��`��;�y[.��8ne�<�j�HHa�W�# su��p��~[��P���MGJ���������5�w�=�X)�6�n�k���[��3�%���N���]{E��f%P��u�6���d�5��R�<��"��>�j�r�!@��6"���оf�<k���>^�4_!�bT�=�Մ]��?�.d�UP�:�@W���v�X�]Z��U�̥�;A�	���ie�c~bd��fZ��S�[�L>	{�cQZ��/���!�b�KML�*���[�n`UdlIT*6L,,����nl|Hk�	=u���d�D�|D&�i>�!����I�Dx�˗�?�����cy���'��>]���#�ob��ǴL��� �[R������">���L-�ee?�v}��E|64��a��L>�]�!�=�_^	p:����u���<��<˱���B�s��"�.�#4�0!�����fY� 5Ԑ��#��BR-��L���Q<'k#/��S��̝��R�H|��V�]_����2恰9R�2|��Z���J �{9Nqh��!CF���k넄�B�����C��ă�! 'c��wv�s�b��&�^8��G�LV�+���6�(�oi�����2j�����1�#���:�ZOz�D8 w2�CL�phP���y� r_���Cŏ�yh��2�O�
�!��� �1��s-4����_^ߐ~�E*��d��5g}.R�i��E���Z�y�B�D�ң:�o�"t����nzr��)��q��Gx�Kc�N1���q�x~��]�.�~|ʼ��o� daj�8�M6m�,<د�i�XWAڷ0��J,��Өr�t�)����.��yk���1��P�6ǗG�/?�]�}LH�X�'W���*dz��lY�-mK�n6�m$+�9Z-K�r����$��$~ ;;tvw�r}�C���08�</Pu�[\��6���M����}y�s��Y�/����h�����f�n ��5𔣂9��e�[����9��?Z��K�j�v��&��R��5z
�逰<�|�$]͖2����4��$jBd��2� ��,�z]����&� �|����D���$,�?v���=-^��Ca��d�W�uvCrW�>dY��{7�-|P4ŢNG�/i������x�Ӕ�js�����Xk����.��g�T��bBGa��}Tj�f�&Bx)�Α�&a��ۥ\Shq�o �9��f�lUp1��j��#/x��T°i�@�$�f%�y�6U���by�~
�u]:����R%2j���ؚ|��V�]ư�0��Aw���]����s�Q�?Q=��\�~�_��YY���2$�@0=nl-��$�lY�R�`�W(˦�I��,8�D�ׁ̪��w����m2���e�qC4S<�_3�a��}�5�\�xɟ������B��~LZ�52���f2�����s���`'�������^��<gOc�X1��*Vm��+1!~�O�E<���=�۸ ���3b��0ZJ��y����w�P&�LзrEm�?���+��.P��vܙ���M3y
_�杞�p�}���kK��n �h6'��_��;�l6��da��!� &�:�gM�#cҬ�U*t߱�������Ϲ�C=P���͞�b}Ͳ�S䶍�k��ׁ�j��Q�������`0��J1F���B#�~�����Dʦ�R��V�4-}	�>NA�ZM�b�JdX�;/<���Ȉ�{Dۼ#����WxE1��c���Z�'����@Mz����fq:b��'��0�s~��V��7����2�&oN	��SP�! �94.m˄�|�.=�N���1L��G����]s |��Uw�<yO*Vnn�L!+��̻�v��}1���i�ú�7mOӚs�~%C��k�u���0���k܃�^���оk
H����[��{#e3��e��S�:X�[���
�d��i�9~��涉ֻ����vΗ��)<O��7�(��c��e`82�jb�ۢ8ԇ^�iPk����R�F�B��)T�#��.�f*�*��j}L�������Fu�9��COi/�vƛ�!�?����#��\�Kr:.z��J͛��-t�-̏$��-dG����:#�Uz��H��8AIU5 ��u�执u%O d� W�N�M��H�����S�zFn�/� �*7���F_Du�lV~#����$#C�����߲���"��g��w�=�4M�P2��s괧D�c�0,xՋ!���t���e�86�Pf��G1��$���&�/�a@����Z�Z����mF��e�u�Ϋ�2�:�ϰ�S������ء�"�I|w󓉧�C<V/�����dhU�����Q	����U�>�=WQ������SX�Ɵ��qt��Du��� �Ǧ���D�_���D��x��9Ti�����%��U��a�;=���C(��C��*ы #��nq���o�Θ�%=�7h_3f�0�J�����>�g�{N��(f�~�H`pn*��t�ؔl���܏��U�K�iq����	L��3&�~�%R��S;G��G�d�q*)�z�!�E�l�Z�yz��-
�^&$�:p�fH����X%����%�f\����]
����kj�1��;t�?�]~��W�`'���f�;$ڗd���i�6ӓ�:��4���$������i�jE+#��"��;�ę�����.
⍗�b��A �ʌ���.c�Vh	�鋞ͣ��N
���(?B�إ�S1EV��Y��ү}�I��T����z"č��7��z^����\��"��i�N�<�����~�Cw�ئ�x�p�ࢱ����{w�TaRW�-�N�����;��Ԯ�Y�_	���jg���9�xRf�9���.Rn��'"=��l��̐�@�oj���$�i�Njn��v�1s{�I�Vh�C�p�+bu�uZ��2��d�s���u��2,�9��˛a��H���%�U�Ls�����N+��9cT#� D�(��B�$�Z�9 ��Mٚ5�=�Rb﵎"����3-gl�5<�Gk��9!K��x�%��iq�q����L���>��^w��J�b<�c����ư���+v4�h�N�pZrV�E�� �d��5��(ctY�n�A�x>�p?)��ISY�H�5^T)�*�M�1�u(��L{EoA�����!p>8��;m�8a��ʕ�]!A	
�&r��lf���ڪ��Z�~��ZH�wX��̷F�*.�3l����
8���j�-���R���15�s��k�+��*��j{a�,�� G�II���!D7�DO�4j+o]�H��я�;Z�wh��cu�
4?R�DE6
��#�cyf5�po ٩�(������l������7�Y� I͘"�h��l�� 깪Þ���V�z�ϴjsc��̇���c���若���/K�w����$JJ]��&�+5���d
5˹d���M����Yh�K�dG���|���[0�	�|Hz_o�04ߚ��#y&Ku��u�`t�]�V�gN7���e,�}c[��χ�A�aTF�p���(7���8[�/t�eU�+��y�f��%���<�o�6X�l��B��Z�� PI �.���&�B\���SaM�֝|� 00A%�ȣ�vd�U�r���	���web�}H@�s;��8Sp({���i*���L <h����é��n�Yx��Kk�Pۃ���T���̞@��@:$С�K�p�xvse��4a��X����L�FwѤ�o�b/��#�eH�O��䎻�g�@���j�s��@!r[g��#�����^z�Wm�\�,]p+�B����&�X6}�%ْ�TU���Ӿ?�a��H���"�U��	�,h��_�r�1�$��M9�-��l},����T�Y����AQ?VӆM�˖Z����kMC)�cD,�|^&��S|e �zw���φ��S�D� ������qarw=K+\� ���)��(���!�%;�=�e�H��q��`H�{����V;���S$��ƣ`'҂��duM@��[ͽm��U��{Ѿ>�O�×��Ϟ�C��z���TZ���>��u�Y������"�����u�=�Wh����h�ۜ��6�Sw3\Gd�T�l��]�{������O��I�F�v�%Ȃ݋0�-%��p���2j��4bm�����+���V�1)0�q I��.*�~�K�s(��>棺�kLظ&q([󠷕'����=O�^��Ie �0Ö�+�$҆���&T>��o��:��b�ޙ)X�:��'�\H�h��s	�e4}�VG���� 7m���oq�*���?����W��Jc6�v��:>_�u��kb�9"���-%yrqZ�$8:I�n��+� ,#���mP�M^Q�;���za3�=x�e�RV���e�n��䡉y�%T(Z2HLjq`���ם!A)���D�t8��"���ڵ٨�*Ť�P�f>�b����
JV�:RR��e*+����d�k�UhX��zR�ȇ�H�<2
 e_qi�.6��7b �W��N���^������ �ٟu���h}��פ���R$��� �vΕr�o��t2�% �ɜ
45Dh��B˔ ���yg;2̪��y`O�Z8�"���@K�Y��c@4�c=g�5� `����-.�Q?�ź��EN�/��D!�_�8t�x�������9�J
�"j)ft��-_���,ž{�z��%��D�y��e�-���{��)+�v�u�xQ_� )�[�"�LQ�8}��u7����C�~�����ko&
MH�J]����;�l7�����6��^[�Jz>��`ק�xr*ܛ��,�L�'��Gdɏ�UlP���.A��R�TP';x{P�sծ�LE|+~�_�����c��X[u!��4�'�Ī���1.,�9�k�ľ�������<!_�	�@"`�A"$�;A}	xO��_�0n�����o�0��5&�e��/URKT�Y�~;����Yݢ�ל�ص��j�>�"WD*��~��a��<�:%<}�R�KU	.E�t _4��ktB��3�ek,��@&��~���+���f����k����Z�>I�:��ܸ3��!�=9��f%���K<K�jT���U����+T�����7~��	�5!u
۶�]:>\��57��R���;�ׅ"ZCJ��s!Y�{����.��ޮ�'��2ueo�f���W��x�M�ޫ{�� �&2CI�?�}��[rTo4�EjFy���tZy��D�Y�ć��A[�������q���S�*���pj[��ݝN���q�����S�b��lJ��k��J��{HKh�n�J�������������j��,��:�vEC/�h^�d]��w��I����vIb��^+��Vi����u$AVj�	�"��9�������+�q/��<��PI
>�D���538^���"�h4�0�$~��c�+�<ip}�v�E���Gc�f�
���ES�/YH�M<@����o0�}Q�?H�0z`����f|T)"#�w�bG7C�����,�r�W�L^B�y�b��b��g�d��6u�%7B����7o *��q�D!� ���%��V�\��/�]�*�WFn�3Yl!mx���6���d���`ȿ�a���|���a�!X���bs�����of@�qB�4ҷ@TU龘�W��������8�*p���)�/��b+��߁�2�~�Y?���*���WYo��kE�&q�d��)�8n�&�qi���^�˃q0ͦ�ƏHB�8�1����Io������:>K*��*4�;�EG
�r�%�'�Ayd�A�,"���@k]M��xڴ�����N���h����	�y��Q�V�}����Z"&��Gu%�@Q�'x���Z<(y�	}��T�U�*��^s���o����7�"��R�Of�&�-�G��;t�S�OZ����D.����}m��!U����K�Y6m�\������'c۞�٧:A���g���k�`����E���F1*[?���eo�[�J��ҾQ	f���ϣƁ��� h�%��$gX�p���7��'!�'5*$0䏇FϯS�o�y^��3?���ti��{{�D�Jq�xR��T�[�Y�m�,z?0���;JO�k4�S6q��4�yx��w�~"�~��M�~����W�e%���'���B�0���ݻ�^7o�2��-�T�v�]�F���a�Zj�'���T�F��V)�}{s*��X�` {$��aO��H���?� �^Vk��Q����\��-FD���|�|G�_�d{��W�s�D�d>�P�(��ŉN����(�_�x!~�v����f������E%n.�����-އ�� 4��XtB�>Iw^[�e����7���l�)�bZ*�I!D�)��f ���rA����y+ѣE�Dʚ�~s!Ct���΁�gY��(�����_u�\\�rNG��x��d�l�2f�wz;?^�� �a��z�?`D:wƹ�_�Նf�	��ۿx"��o�s������W!��fԭ-u�j��R��g*|%߰UF���&o;T��s�k�zL�ӵ������xc�0q�J75��'rp��d��T 8G%��A��kb 81���4�v�.��R�B�"."�fU��vU�n��0"|��܂PBm?x�@b��_���t}&�w�s9i�^��szphj�7�C�����Z�s�"�q����:6t@�*� �U�!d���[���km�r:�|��KԿ:�˧����'�AG�4h�g�Au��
n�Kr)�2�Pn�Of/�HG��x����"�	�Ĕ�~^4��`��T�2/jYҤ�o�Dƶ�ݣ�xp�y��-b�ZT՘�)df��~�>�W֞��'Ⱦ)u`2��iΛ��n7��el{WIZT��dF����v��+���߶��z޼��D�B�2g&O5���'���ID�-^������f���ǆ�C>Oׂu�8y:�� >�C9�֊�9[�:
��Pc�+�� ��&�Z%S�'�F�/{���ö��p�
�]C�3���i싆�A� �G�D+��X�]4E�a0�.Xܢy��J�fn�%;����ܿ��屮)�ZxڲS��DAA+����/̋3�L�"���0�#��|�ow�@�8�a=x>�����)2,�K�ژD���4���,��z�O]XW2o-J��㺖w�S�'��������#Yy���E�#��eM�[S�9��8��8�L(�u2��*z۷+�p�9[�=���Ze��Iт��I��@ ���LB�	���1�녯(�ی�/d�R�`
�*��?�:�N���Asl�=�W��ƛ����Ny�d�W��=`�4��~ I��p���RP����<���5|�-,D~�3�8 M(0H�n@��/H�25��T��0q�3U�^/�	R�uI�a#��>l��b���{�4��	W�%P��~T�p=vm��U�8݊��s��_N��2����4�43n�0���e��`ix�~���QV�@9~�6�!��� �^��k?Y�u0�h��i����EeKGA�0�l<i�}���=ӻf<\D�Ϙ��f�ևŏ�f�����o�M��!��b�Y��W��^�S¿'3aā^w�����[t��M�N��K0j5�����g�%��0d�j�l�z~���ޡ_�x��8�,�IqI	e��Y����FXa)�.A1�{�2������J6sI}��eO�m��R'�?�FCbP-�]�K g���˨t�?~j�gf��J�^B�S�0B�;�dRU}@�h�U�0GY�On���ǳ�d��06������VQ�!G2D�G�!��i�#U�35"F-���>���h���>��'!�Ԍ/���f���VV�
��Su���4mN����׉ei�c����������M�$�DScqH�x�����IӭW�>މe��>��v)]]6�̫�(X�&ɈԲ�1ی��k#�_W����o�н���>�}�
�P�����~��M���B�4ЅXH�$���k�X�ר�:sD�\h�D�	@��U��%Z�}�ۄ�C��#;�*�a����nRxw��/J�UDL��5�(΂\D.���4!,ȸr�����l&�d �GU� J�6�����|��ye��h�mփ�S�Q亮�!.�tqdP�B����f���-Zypp�����9��@N��%Վ�ޓ�3��,�J;���)�>}s�EF9�aلv���'ݐ��(o׏��lS��V�$�@Gf-�݉���P�_Gv�栞�L4��y7���$5�k�!O������9�Z
�o��Oq\Co��ߊ���W����_��k��o�ߗ�#����
���qZ.��؟Q9��3�H{r{pEz��x#5�����X�����:�X|�g��I"�wUf|�6i�S&�����9�!�?��l����_�ϵ<00��4^�8àL��I5x�ЎJK��?�?߯��7KHScGL���Z��W[M��T��2v�M�#���^�4�}��{��ij^%4բu�1��;���/�V��Ǉ�U��Ԯ>�e,�v�#3�a�L��#�Σ�ā�U)p��؇��Օ��ּ����G6�[P��Y�c6�C�7N1�Q�MM���E������kώp�s���+vI�
���敵R�D��^:ߝt�80��Q�i���u4��A$��mU�"�U�������\�F	�K��;��3��D?�@o��]�V3G���3[u���_[�1��C}��������v.LW �ѾϚ�+`�z;�
ש������4��k�WP����2��Dbw
ַs�߬����}�f�t���%.�ՉԴn���Qi���$���CH?�D�)W���Nu�� �Rr�������W0�+�/��s�Q�}�~����C�nɉ�c�Y�۟�p<lO�$}�H6�>�q1�Z���.�6��[S���N�T�N��+���~�țd��s4�X9�L�
J;F�Ԩ���bu���l F�Q�$��9�+�)\a���YBL=�v��SzD�$C��z�F���>@��5�~V(̪�pέyI"��}������"��0�3�:b��M�Nwا6V��v�E�I��6���>�̂���,�>��h�~qa���_��J����\0}�`���ϳ<c��[�L�-��nίyQ�����Ӏam��c~�jԼy15=���W�r�">�M��>��#���b���[ 9:SD�N�a86'��)|>��������p(n ��-4F���l���Ki �\a�MVA��I�z�A�����eU$Z�Ic,���u�Ђd��)�X3��䂠(/�2����k�[ �'`�6>[Y��84`{�=�wQ����0sg�TUc��� j�ߩ�=�(����g�T���8��I-ɱi�~n�����[F9�M�k�I�㞂�����U�����㥘�J��!d��8	_�n�� �8���QOc9-���h���CE]�Z�<��*�^��O>�K��'�y���ꊆ{4m���ۄl
A�*�N��wRZ���l�zNRoA�O�+4��(�h'�D�|w"T��� %�s���m|�C��˗����F�<p<���led���Пo�Ɛ��%�aa�\q&KT�I.����q�8-ب8��X?=T]�
`�]el�� �F�uo���?�e��<Yt2y�s�*���R�/�|N�ؐdz�j���8���i��b�J�Q�{��z �����i��������y(rJ�:���ⅵ8��Ɇ!|�ٔl���$F��9�\�L�͹y��ĝ�J}y��̇uu��(������z���u���hD���f_�oy��F���A^Y	c�Q9l�v���K��ך���RS��v�p8�ұ~������}?��F90�d����E�h�ٝ���%�W%��� J��XwPHPmk
]j��i�`��Wz�M�EŏΡ�';���/���X�c���ޢxf �7�Ҷ�MZ/�O��G�^��-K�ђs�dk�t�1
�UKxF���s�߲�/}��V&t�ufSd#�9�3����bIW�/!���i�}mhYl��@i�T������������3  -�ߌCϴ?xr
T��Gߪ���5E�鄢Fj����Ɛ%����%��۴rkU~ 5�v"��y��jVOz�����8��`��*�R���R�C���b?��L^:�j���+5F��9��z��ws����7�<���J�}/앺�I�L�g�/��XF��b�hI<�1���5��}h3K���u;��:��a�|�zγr�'0���8���&#��Ne3s�kػZ����eۗ���[��iW�H�p���Ja����Ǔ�ǫ m��Vrthf[�H�@Ͷ�W��Rϑtn�E����#���M{��.)�����/�u�JQ� 6!���[�8�~��S��/��h�x�?��֠J�{���uF=�(r�pA�� 
�K�tc�mz҇n���4�r�VA �_���G}2�-�ʥ#��}�*h���a#�_�,
��B���\���̉��ֈ�����X]�=Dؕ���
��ie�h{@���F�����P� FS��F�����`
��g�bQ��+^P�&�z�vm<�J����䘄VKM	�T��c*#��c���p�`���!-�>۠�=�P)R9%�eq̄O��F�+,�-�k.����ڷw}�wغ�����`�w��Zc-NM�~U��R���lyhlX O�cw�|~�:d�_p�ƌ`J*kt��ˑL�>���t����
��s^ ��KKr�5Y��V��ƍ�*�g�.���R�۴FES����ߵ����Tͳ%���������h`�P��TE�V9��5���)�hμ!�ԍ����̪��vV��w���Q�?$a�y�_�lf�bn�Ū>/W׺Zl�U�|a���l\݂�g�G���ԗ�Ca��j����
UOA��E��]��^`h���e ��l��q�2}�]�0��L<e����5[AA����P�c��QYF�i��[f�#�~�Sja�]z�K~xY8�J��o5�(��a"F�u��3����ݐ/�^���=�����~���N�8����#_-���bTI��@�}4�@ȔH��` ����h$l�\������K'�wL���Ɔ1�S���T\�
\�I���M!��Ѿo�t2�~Ǉ�*@|��"V^Ւ�:~+�g��$q��V�[�I���=hK��&TL�D&�RQ����<�V�au}ɶt��"�������-Ųk��K���x���y6%��B�z��mbD[uH�avwd�o��*ז�&�(�7�%�gH���U�'H�=���B��L��O2|pr�?�x�/At5������.��z�8=N7R��t�.�A�n֞�c�{�-,���o�b��Q!��Ho`�p���ǈ]J�J䓈1�b��_����>�63�9uͲ.���)Dؒ�g�1Q5���6O����	���Ũ|�׎����׋��w߲�eȝ	I�Nk�n����Dr?>
.��Mħ�u�P�3��U�h��YX�2nj�h�� (g���g�x v����?}��C=����e@�Z:齹7�����H��¸���/Ӄ�a�;#Q	+*��ˎ2��|s59�)Q!|UE��j�:��������������J�x1hO8n�`|�š�������?�t�P+� ����M�db�nM��P*���ka��洵����چ>$��L/£]�t3dՄ��m­��( �������>?���i�i�P�CIH��h.�v�x�����B}N��0���Ŗr@?:#�j�q��83܏�iR� �bi0x;8҉*ݎ��K
�V:�-^���u��|6Ϥc2�*n����v�"Z�@ү���0����j�X���ĺ�a0��J-5�h��oy�q�(�[<E����5�%C��k�"-�gYew�d�[��;�	�����io:����	M��a�`��X��m(:x�b$���Ϫ��.�8�4鈕b�^$��s;Ӳ��o�*?Ps��KQ�j�Qg�Y/�1�P�R�ڧ���)t�^���hMx������J��ho�)f��ZK�0*:k�p;�ٜ��K�g����?y�m{��֬�14�#%  �9D�VH����2W����=2��ǂ(��*1���!l��(g�#��kDt�)(�a�-_:���V�\SH��
� ; �E�z�8����1�O��AP�jN�v}��s�~���	�S�N�F��396"u������f��7�[*d��O�U�)�n��QV�ޤ�|k�����p�5u���8�����J�c��� ���dW�����V��~���� n� KW�xLe�h8�L��gOOE���ZIZ$����^2���L3^]=Ndhw�lT�^�����e����/*�X�#�1�P�t6��OأT���5���m��<ڑ�$a����wP��&D+�[[0�U�Q����B%V����iGp�ߦ���t�����N?�H�Uw�(<#���=$#�����+�[�M�������8]\�=m0�"'�K�,',�����j���t�������d�:ş������g���C�D\;_��g�j�����Y��N���R���1E��&1~-h�.��ZE6��[�
@�Z���5�LAx�$ģ���r^�(��4��1[36�	����k��������څ�-8;�+�]��,�q���@�ޭ9{�%éc_;%��1g�'�P࡟�0��iw�Z2�,l�>�aCa̧` <;'�J���d��_;E^߇:�"��`C��r��_3���<M�:�S����X�M�:>#y�4͑I_�['n�u@�SGs�o���q����=C����W6�_7�]8/�rE�2&r~$
6A5(iгZuq�`V��ьI
��6Fa42���N�G>��xJ��ǬE?�e����L���#�e�)nd����̲�G��� ���t��� �o�0�x~8I�6�C;Hk]��v��(��AV����@�Thj���w�2�!�{��ߒ^�Oo�[iYq)xjt�e���I�5m�9b�8���;���vj!.��?���k��}ڄ�&,���#xhP�P<ÞAb�/̬m���u)u�����T5�E\����\�S���␂�š{�l%�Zܚ+��s��v?K�NY���	^(=u�p>,�.���&i�R��jp&����>�����Ǆ���T+ږ"J۵�f9�h�u�!��o����M<����1R�]��m�s;fV��d�JAc�!kO�,x���d
}RT�^͠93��Zj� CD�گQh���4��J�;�������K6P��Yq�2�W����^-1��ưӣ(�8���S�,�8��8l�t���3U�J���P�B�^��������iA��.&�
f��,�v�;�l�M��m ��0�W��؊��R26���8/��#����K|}r����2:$�L`C�o�kU�~�j ��/;�zO��`��U,8�t�-�\�S��^��q&�]ǜ&�L�Ev��|{KyBV�{0�Pxk/��	Yr���z+#.��\p�o�`�u~J��Ǩ��B��٧��}�j�'�Yr�k�n��e��V��vDk{FmY���Y:Ze���\OzK��eo3>��t���:����.1$���%�ڢ�� � q䌈U��D�´ky�jx%�fel����-�AfƎ�)�]�o��Ѹ`;	�v�hF!���*�t���=\9V[6�=̏r?�s-��:��x1+oyS~SO�^˯o���p�2��` �/���:^���WU��c�z2���]Pun&���%���?5�$�'�^��O��Z[' ���Ґ��;ξ��$T�5!j�e��A�=�����ϳEv����;�rps�� 0H�[ؔtZVg�o���1jۆ��iv,AK��(��r{wNW)�h����N�|��P5�=��J�>D�������(Q�
��P�'���D��i�&��	)��
B��$����э�e�`^�>�aG�=���-#�"�d��e ]G���t��)���j1@���VR9C�]�3l8C^���w�q���� �w�,���E�(^"���-m���<��W��}]���<���=�a1�<_;@i�b0p�
G� F^$'�7��I�O��I���T���s?��&'1����f$?ԏ؁*�9�9�{4��a�-ن94<7ۼ��H�(w�H��˥��;��B.)���?���>w�( �M�I���Df)h�_�V�u_���{^��.S��.\�S{5hX��|�J���m��������?՚A{�p�F��[�T�*���FV'�4eѢ��	� xߢ]V�e�6��Y�5&͹
k�,�r,���B�~��ԊC������XhTɻ���hi��+�����n>-�P��!�y,y:��Ѐ�B� CS:E����P���(��ĞmowY��w}ړ �wP� .�/�"���Q����1h|\���#.��p�V��l&��Hk�ÓW��M��3�@Ȗ�۞�+��}�[� �WT�����.K ���(���K�Q�!�۱�	v�K�ƉbW�Wȗ�K��f�7m8>�h�VG��vqvEyu��%]�@	Z���=��d_�qz��V���-S�Wu8W@<��(t��&uA͇�kXsM_�o%
Pm��b�t�=~d�c�dY���.��Ϛ����{�I�x�C?2�p�]�}�B�,[cs\Lq�E��y���_"֞�9��G%��Fӄ��r���X�� ��r��:%,uҢ���$�Xmݩ���bxGv=���m��,����$�T��3=$��^xc���#�x�O-�!��U?��l���)݁���V���w�]�At#kL�`��S��Ƃ�ԣ�V������J���B��
�hiɫ�#P'�����7�f�˶�a�G��m��d����%�����#��Q6ӧH) ��_ʮ�ؔ�(󔧰��Pe4����.��E���������g �C�L�_�z6ϱ�����*]����O���!s}Γ�w�7��y��Po��B����Cq,��7��r9��G36�-8Z�࣒D)|�5���-��X��J�P��$�?�&�qv�F�D��A��B~�X��.��T;��I�rw��Cd�\��� ����b���"9�K7���@������耕\%�w�zq��*��ŝ;h**2c>P��VZ>-g�6�lv�I��,:[fr����>!gP�T��@�+�u�#�mG���Z�c��#�!.{��� G����/�.�-�S�1�����>��c��B'���Q!�®C��a���>E�����D�z�e��L??,^����l�7�p;Sm� t{K��7��6���e�ȭ��(?��QY2^�C,n6���.��t�-��4���m�]�� T.�2��|�BG�4��A�L�f��{�)f^,��
Nt:_lH��U����Gy+X>���Tt�h����I����.C���Dp��_�AYr׮��n>�|ٹ�v=l�~�c�E������� ' �d/=�ߺn fQK!C�Z�,�6  �i���;�@)�y������&�=�y&K��ߘ��(W����~��i(��#�7�	 �g�g�J&@�e����-�JG����L9�c8+I�!}J8�ZI�� �[�O'x�X��aO�B�{��#T�1.96�t��^ Ώ��O.*�M6�j,l�cp���JI�	,Mx�@vP��!�����B�U�k�6m�j��5L~4�,��m���M�v~k�j_�1rhm�u����һ����˺�
��7��M8[*�GJ0D�j�Y�L������z)܇pW�dXx}p8�﷊��@<PM���=��A'%K	v�%�������H��������lq�7�lW�ǔ�?�RD�j��2�-��WI��#*�.�6�f�p"�?��;;o(͑��GQ���%������p��5�7]��}EU��#��)��n/n5�}EZ��o���O�9��e�`�$�E����%��Ã�Ś��Y[]"�+o~>�@���j�b>�;���uXy��s�d��d��s����ư�T��J=ߠXL����r����U����Jg�~��7���qO�X��OM;n"#�:3Q!�Dؿ~��)}~k��3~#��F����B`e7�7�F���>�Q�`5�%xx��Q6�mJ�2�yҫ��A�~�C�)pޕL�spIo��݅]��S(��	�|Dfd{mh���T�{��;OP;]�:����&��*R'`��3��;�K���=�Ţ��(��D�zj0�r��'�5����-�=�MFg�IE?h�N\t����n���k,�'�����l��Xga�PkP�F�R<�~��4�X��#D���EX�Cϕ9��Ti��z�7��*B��Gcb��椻R��B�>la����0I!S�v<�/&$vl	�[j� �f����mg���ׂ�vn��t�uUUܤ�����@y��lF�#	��a:P��.܏4!sJ��)�]ǖ�L��Z�����u��~v/�}����A��:`�65�bӏ�j"u��,���%��Ͼ���"����PI~'Ù�u�L��SGAd:��Ӈ��ۆ�9Ҡ����\��d�(�+b�ar��o6e��?��c�Z����1š=���Q�:zT�-�Vm������YP�#$�ܖuS�	zY���6�	���ت��y���0�X����L�	�w?o~��V_o��"�a��k�o�گ���=$���t��&TR:�)y;���EF���:?K�G����7�:x�b�y�S��_;�u!蛲�YA���f��DU�jC��WL���׃ۿ���]���a��>aPi�WK���`�E�����������R^�&_�Z'���$+ّ���*��6��m;�l��__~L��B����!��1|fKj�7p�=s B�j�z�Uq����(0\ �9��.M6fΏ���m�v�a?� �'�����y�lE3%��5Ի��nm9C7�.����n�6��������z�3*�۲d*�9=���>�:��"��@��<�8��UE^����A��盝��u c��_}�����Ĕ�:��ɕC���3�t�~�9�Ly ������x.! "��6�ս}��'�� �����h�ot��ffEt��qTY}�9�W����]C���K��ODzGpư���z-̋��pg�m癨�j� �G���ʢ�`��V�=>f[X����an Q�|���7���.-���:d���s�&��_q���������q!9�r>x���&Btz]�R�b��<2.o��]��V��Z�x�R�e
!z^���ʗ�pqa'E�E�9�B������Ņ<5±��3.&&h�]���#�sK�e���cN��ҹ�������v��;Ǌ�6�
�ƼZ0�A�U�3x�s���E�[c!~8�=cpa�e�3&A�| �ӌA���v��^��um���|7�2c�֎C�n��h��um��O:��s��[Z��Q*a�����I�t(.�@����=�>��b|���.�B��q����o�@�_~� L_­�F���n�^{�ۧ M��'?�M��֫�PdǓا�^A%�}�|[�6�	_���?�V9WՁܘ�!���QZ{��'m����&-F9c6��J�J��qbyT��\�j�?i"����kFu����'���a�6=��%t��KO��&�e���QĻx@,n�[�t膛k1}|��8CQ��C�4IB�$�o�mWe��Y
�~�PQ���f��7ǩ��+��j��y�kuGv��b��N�I���s	-�}��07,�UW�m+ܚ��I�/��j�$�g7��MǢg�*t�
�����R
�A��1���s�c�WPK�9lS�/��Uj� �N�YB��f�_���l���<����GC`S�)� ��/X���1�}�p�LeǢ��(S�L���c�Tv��8"��&fm ��)M�:Ex7�t�u={~5�g�,ګH�I�@Mf׌ICi|0�E ���Ÿ`U���An)���5
��ˮ}�cC������(���bh��fd!�Vy%��K�Z�fd��G�.�n�F5#��e�x���]�Z��Ͳ����V2$�:�}.��@��1"a�W��;��𧹵�V�i��O��; ��ڭ�X.��5v릮�0�X��dB������<5X@# ��q"b_xY�8uuЃ�(U�����n[su��84�R�_�+U��)2}��*�5.�d�d�-Co��.gl^a��jH��f����٫��[�`l�ͪ�#O�N{�;C�H��57�~G-�����Y����+4yzےe�ٞ�,�U���-kB�V����u��W�gr>����)����,n�����h@?��pkf��0���YѮo� K�w��>$�A���6�b㇌}P� g�&g)y{	&u����:����V��{U�w�b�X��"�j��K�K�]/@ݔ��#[Yf��,�횘��}�\�ꇁT8��X��C�!���������I~��}24���9X�o5Œ�d#(�&d郮�:,1xI���һ�:�ȋ��?S�w9���dȳ����W�b����R��ql_�JT����|��O�U�)������y	�k�'���)���ZB��i��>����.D�CWa٬쳏�N�~+w�e�J)/7��[����b���\Rx�R�Ф�D��%�N��_/
m�3!�9�r�u}�P���0�!-�ۖ	�l�*Q�u'��.NΊ/�˔�2�q��F�^��8Ƿyb$�[Q�|��e����C	n �����RӨ�M}�4f��r��ŀ�i>d��I*$�?�6�Ga��\�U����i��Jɍ��r�X#V�̢�j�G��� @���C,FTo�����X"��9�WB�E(��E�45@H#�ց��d҈��-	I4��b"S��(	� ��q(�$���p+�5�&�5�|?�y����Q�z�5~� 8Q�E+�ADF�|��D����
z��^��N)��'3� ����d`�eM]+�*��2GTŗ2�#X�R��~��3�B��)|��Ξ���N�S������-�Tx�X-3��jsS��n��X6gN~3]���%�
��[���4���6gZ�(�lR���dy�1g<�JCA:���E�O�4j�-�fs1o��'��ap�Y����]�"��y�˿ĵ/ڏJ&�:����Fkԭ!�tr;=P[s`V�j�e5�L��JM��U{ߠ6No�����������#pO&a:�/W@G�4� B4f��QI�V6���� �j�<E��c���D��9�:��o2�Z��F-��V`�pO��˜��ζ��?�.���п��Dj.5w�����̎�Te&A���Ǣ/Y� ���p1d�W/�){ -����q�� �p;b�V�y�,��?�c����B9��T�{��&��K��Ԥgc�sHa�%�;@��>De=�Ib�}j�o������h6��C�>n���ݒrD�5R��}���w���-�vqH��,���
��Oʺ"&F=~~�~�ā�5����kYD>���] �cx� �����SFn!�.9�2��F~h+��mߪ	������b	�}b���䲥�*���)�&����N;�_9���\#򗮟��K>�Wٮ�a�=�on�Vbp���v�
�h�u��Ӧ�ѹ5O���)���/��s���>/���y����ڕ�T�x[?�s�>��ts���l�r땳�3���Q*��\&k���Ȇ��cTm90����s�yx��'2nl���^6ѷɲ��={�p���GC�/|��O�3y��n&@s�,:�i]2���|�>'�g�`�M�;�s��
K����2O�3�.!�g�z����;��oBGy�V���ܭ� ~>�����Z�)m��(���V@��v�@���5�7V$��d�-g\j�)�%L엫k��m~�^C$�@�g��b;����Td��*�'����^ni��~N��c�zpr�����tV�(�X����k����%��a Ud���]!u�@p�krnK"*��8��^�2��ΜQ+��S�m�7���{�)��LF��@�v^�Kz��F�J��gb��:t�����Eݹ[���#bt��!a���;VQJ;��D4�)_�xURw����sƢ�D�ڱ^�bf?�	��_��RX��șA���.|�fMQi\2�r�H�B�~�}elO��ʇ�7�P�����Ð�rY�#�]4���={�%+�������n6���WO"��(I��c��g#���m�Z.�kt>�p�Z"���=��`���l���u�G���k�ų#�va�X-�a���vU�Ǭ�-}G4'��/�; �s��6�w~T�Z���['�=g�1�YK%�������>����AՅ�*�{3R��Ὂ���%�2��!��{^v�b�{���a7
6�Jwy�JX�_2ep@)[�D����\�ޒ(,�~��_�b����q/W��m��H5��Q�s�NFpKʕ������5�ܙ�3;�U�/���F\ῙD=���6�12��D��ʣ�p��c�̋�ݞ�����s�=K\�׹
�D���Z!͖|�.�5O�|3_v���g4٘Y,���~�!\1��;�a?�QB�w�8��D��Ys�֌eY�,&��qI_�vA�>�Y��snE�����OK��4Nd��䚸�����̘R?:ܠ3Z&�\}�����K�"%@W��v��a}̙y����WB�#[پ�f�W��c�(�
<I˸7�0'��N%��B��w!�R���D��/���U���nn�<ɢ��P�*}�&�ϰz��K=���B˅��R�y��L|_��\
j�ی��|�����g��@��f�M��"7t��^���&��s%���;���A2���n}B��������d�i
��e�O<�0ݽ�4�>��I�����H�Ld�/�Z����PJ��5�H%'>R�	�OPTz'�P����9$^�	�!�
`>�Z8㽃�P%������T��P�=�d��k2��&`(�����W0��<Fgu��\(?�)��!؊"�klڞ<�F!��7ԃٺ�����B��U�`�H�&}�G�0�"�o���x$|�1�F����5@�B�F;lH�,����J7QQs��� �����o��M����˛��2Z_�P3�D3���� R�|�De����
�����96H0@5Y�������|)Ή�e(�E ��?�!	�P�L�@�ĨTbh!�7�A(<:���&ٓ��ɣ$x�J�.c���'�#Y�˘Nо��ZT�����\_5;��Ip�#]�M3-Y�v�Ӯ��Fk�AO�@A�N�Wѳ�/�tG�N<����+p�O��$/>c��(���EI����1���[�k!"���	�xwe��PUu��Ӿ[xJXWA!��T�lz�����ɽ�|���"��2y_����@�}��������A7�Aj����}\���N�0�a0��M@����}v�^f��8��`ߨ�y*6�m��g�j��oqa}|�w}�'��17��U��X;�L/'��	��a��A'"9hþu_P�+��ֽ�>�;��x���E���~S�� 7�T���ዘʍ>���9�g�> r]�_UX̑�qT���nB�@�,�WPf��u;�R��&�U*�5ꚻ��LUP�H-Re_#���g�����p��
^b���w�Gd�xmɟ��G]�Ex�񞮨m_J�"+xq���&_�7�G���|ل�O�ʤ������5A,	�di��B��f�W+	~��#�t�Ӯ�UC_2x�\K|9m���7��n�v3V�n��\o�,waҵ�'���2�}���1;#��h�`5�����N#!9�SȾ��}i"����{��e���/c�dC&2j�"�ݩ�i��"��R�"��N�vqb;�����	�����O"��rN.!��^'Çd��d Zó��R���S�ʐ��-�GO�Z�_{V$�$�-H{��!��D�&��Eks�y�}�sy֏!��ڮ=�H-�107�e��_%~��R�ʮc
�WJ/��1ѭ\�|��]㻥Ǿ��~&���ޒ(��엟\d7 /{9"�cY��c�o���Og�m��u��Q�VL13��*�����~>�1:�c(m�j[��54�e�/ A�����.;��H��O˃�ߑ�I��a�m��g��F�B��ϕ��3��՛���Q\����,ڒ5<w�K�D�K�����>5#�
Y�U�����z��n�Q�+�"�Ү�d`�+��]5�6�q�H�O��u�ǖ%�G�͟xd�4g�H�.��]]��
e��	O���UCe���(���ҹ*�p<�YnbQ�����t��&��V�_�Yt8����n)����jg�˵�%��}Q)�jg4����͛Ձr��ћ
F�*����sQ>XI���m��xsCU�c��A'C^O1�s�^5-9y�5�ꬖ��[6aP���64�i��>���:(9��y!�Q�`J���� /7w�D1�o,r�����'�� G��a�@@�XQ�mq_��gΟ�)��H�M��Ȇ~F|�֞��c�^r?�1k¤�\�*�=��:�{�q��V|��Z:.�uW['�箳�
�Xk,W���i����7Q��8�byc���vP��I��52Nk�I���L�G0�\��~��@ E��SD�U
^l�9��T܄B��.1���3�&��o�R����Yn.�Ł8`�����L����NpG�R�0�LC��!k}6���*����ΛEm���O��ZB�<de��7Z}���g1eXn"0�t�e�!� a����B	IG�k��K7��H�&>���'���Y�2F%�WE�԰�89q�ܮE�}�/�Bn�|��q�fú� ��p
*���Z��3��G׊��3#���܀-��
Wm��=���)7B����!+	��Q!�R��V+R'��O�OYV@(�fW,̶۾���s�5a�ԍ��*���������bg�'9~��S��o�����0e���k5�^�,r{�tF��	&��/���Z���U2KW�v��_�^�Θ5 ���b��ˍ�$`�T�
u�� %W����a�m������A��wVT�
?Y���O��$�aGkg�eП�۾����P�5g�15��X�!�8�p�a{�+A}����K�0Qz �(ҷ4���"�f�S<}*C�}X���g��r��w�F���/ͩ@�}K\��x�퍈� �*~M���ڊ�p�`��	O~�.T�2YC��S^��Ov��<\EXH\SZRt3SC��g��1X�˽��E�*�t?t��?�����F��	����=&��#���6�ԙ͈A0-KXWQ^���)F�Hc��߶U��f#��8�����w�*4�%}3z��Ս껑]�����R�K����"�+�"P��y��}�~B���AKi֙$x�%�1B��B�	qec7I�윓b��Ǧ��|/�D�6C=rm���m�ĒP����=��#��A(z&�Ћ�;��*&e/\V Dŕ��1r�k�\���1�־i�_&h��L�8���Sl�F��Nѐ�`����:������Y��`J ��n�m�Q1YѾ��F�����\��l9�[	�Oy�O�ߍ��T�&@�T�Բ2ͮ{CD�ȟM��e�#�x�ek)�d��gyKۚ\�m�1�k��XN�C%'�� ���1�^�m�C),&���H3_C,l��%O�'?�`�\�r����I�6E�S�������9X��Q�9N�ι`-�� �g�` �o���?8f7�`��zY�z�"�.n���(����s�,���S�j�`e�7��^�v��s�c������[{�i��Q����뻖v�a�V��OX�fpdʇ�Pa��rF���{B<3<l�Zr9re��'`"7�sڼ�A��	JY>AÊS���2�rM�oP��c��:`H���y���iw����٫�����1�����>��ͻW�`([]��򶒐T���-�#�%փu4'�ֶ���4ٙld��������?v��S�i���~G����qWnw�o����3t�ǎ�R�b�~ku�QFBv3��h�}?�m�2��C*O�eF��8�[Rj0����.�P�9�Y*[B�8��K�f-���/��k�_�5�rCbA��h�}E����V41��[4!ã���X4�A��q�Z�k$���Ϗ*�
�/��"(�$���������Qx�mM�9#dО��F�rC8��-.A�o�A9���rrH��eR�7X�;ld��1Ei!���:����Gg�w�o'��p��Mh�
���3�X���8Lg�$�m�c�-��'�NմO��#�Z�7<
[f���K2���H?fP�_{�=�Ea�k�����9_����5��������n��]c�`۞l�s��T�������7}�4r��Pk�J�:*������!8�H��FXQ0iE�@����3�](,����Ϳ(Ļ����bG"Sr[��oqݶ����<�[�꒑s9�z�`�Mm�i����Xm���K���u@զ�pY#�����?X���#
�(wߣ�A���'�?�43UD�c+4J�� �]��U��p.�`�З2��P��~ yٚ�d@̗��]�$�"�	_�wp�w#'dpb��Q�eu�yxa�ߞdZ�=�P���� �e�D.���+�l��SL�e~�2�|*��������<ꞏ�Y��p*�W�׌ei��~���c6z(�vOJw�1�k$��HqW���L=7�n�̌+�fM�CeK�,ltR�fڳ��B��{���Xm���ǯފM���#dLO,�&@�F�V��5�v�hn!3�L�z�9�C�`�ѩⓎ&��L�s����>c�l芄�
ҊV_����N�N��q*�Es�N��-�m=�-��K":}N3f/r��N��~ܶpA0��J�8����^7�'Cէ�\��g���	�f�[�Ҙ������F�)��&Hl/�nb��m1����>$�.��I�����[I���S���fЬUC
h:��1яI5���9߼�"�l}����n.���U�G�����{\�����	��t��ܶ6"�����dٍ�R����]�p��z5V���-5���<�A��'�!���ulf2��YV,j:_��4*=H���i/T�ZN����8���-TY���*f��K �6�(�S�tG{hH�(�\p�n��;������˓����g�U�,���2��?�:�Fӽ�5����y�Rx��'�b�#8(#ԭ� �X�>�"%)?����y�=��Fėn�A�u��[�n��Jy�3Z�����U�6�_�4���w��(� �RL-Lvx����{)��7j�VEC	4ON>�*���J�,�?�E"b�ߚ��xsL1+r��!��:�ȘA!%���aR�׀������8����tm�]�0L��cO?Q֙	y����p�c?��2�/����r&L[�0TA^��ؚd�����������6���D�feWwc�CO���^F/���;F(,�,�v�Wk��)�>ǒID�O������P
�}D����[�Ma?jB��e��.s5O�f[��Gh��K��(�%x�d1��)S�b��d���;��jt��9�Fo�5��{-�ه"^'hdS�,=I�
-��|�I��-�X4 ө�h@���F��1�U�+���>�I��{�t�Z���`�y��Z_��_v	�bU$!j�R�9��GI�������,J�ɕ0��>�n�%�ɝ�V^���Z��⣸��y������V�fx5�D"�@`h��#��dN���F��4N�����+���u:��{�qE���׵E;bX* X5��`�C]jᕔb~Qe�02����D0����ϧ�����DM��ie��:�9SZf�G��B����%�@0���|2x�%�p���m��s�)I�y��B`*�OH��%�^,X6"m�����ٮW#��zۯPsR���x��y��nt #В����^����}r��f��μ�!K�q �����|��P�b��:eSj~A<b)���DJ^������hυ�Ǽq���(9�ف������؟�υ�Y$t�9��pf/es�'C�pN�4�� ��$�GN� r��r�>�K���Y���Iҋ�&�{[N��L�Ks�Y��$5����	X�C�p)+��CWF�.���+S���2�]�ߚ�~f�Ҩ��N�!�a���/�Q��$�R;�:|�F���(2v�\e%�u�3 Ɠv��葮"v��i�B�ݒ?HG�u0m-�-n� V��6gF,�!�A|��9�ȃr�%�[z���l4��,2�Qx�@ƎcӖ���J7G(wz g[+O�E��+�=b�p��������q�.�5R�VIȖ軅� ��R7�� �*4���\�R@f�:����r������Gj��9��]��,��pC\񛿝�nAi�������,;�U�m�B�[��0Wh(�3�ɺw��P��j@bYY}�#Jp�
�� c�E�e�R>r�QbA�N��Ց���\g��������[{�A���&vo�f'��ǥ,�V�tV2��#RT�H��\V*�N��r��tH�"��;[���]5\F��r����������t o~����Ψ>�f*��2�bc�V�{�֩��~,�!���W=��	���!֘)�ۨ���~�n"�7{��O��;8���咕�٭�*�L��]�&t�l������Έ��n�;⤗y:��Hk\��W�7�^b�!��%�*����=������)tl�Sz�(-��[	��ؖ�l^�19���.˼�l���~^�͒��I�\x�Ѽhb\|���%�博X�B>cQJ�LhH�3���w�%�BU%UN�\0��ij��͹r6��%�#���M�'�!?{�>ѳu�j$����*'�a*�<6�c���*������kjU��Wh���/��#>��Ga��r�u)k�㌎a��0��m�<i<j[_sX�d/�O��b��5��ݰ�v}i�HT�8��P�O���-J�ۇ�l�d�'�;��utF�c�(�R[K����M5��{E��gƳ:Ti�I΄�9Mg35/͸��%l�ږvN�C�Vپ�%�a2Z>�X��K���V|���
flI�J�0D��*iNږ:�w���_��"�s�5��V�����p꒪�,�=��@��4�kf������lc����ӄ��` ^d�vڔ��8�'A���j����Z/���=���{��W��i��]���o�����x�Q��N����`;�&&����+h��0`�t����p�.q�ވ�|�����{���(L�뤡��ݍ����kN��?Dx٩%�����:�7ý(^��u8�WM�B�1���G.S��?���Cei_f?53�6��j�ʥ����>�KF�bw+I\y�4�u���1vԉ�Q���6���O{��}�Htc���V�W�&L����`7r�ؔz��%>�:Q��'���N���e�$�~6ķJE�1ڨ�ty��P�v��˞R�ڎ$����2� 9��9o�'��bçZ���+���D����˝..S�4ߐ]`Ngo���w�e�+o�l����W�4����Z�@dX̛��£O�� ��Q���B�2��6�:����7ز�k	]�>t,����ĎaY��≙u�V�?�[�"u�����:G�+��z�ttk�y�ZX��G|���?�]��O�Y�~A����?��@������:CL����7��J}!b�z� %�!�) ��h��X��`�v_�d����|A'Am�)�Y%���b�=�v-��"��7<lv���@� ݕ�����C��\U�����G�0ꀒ6��S�����?���GC׈�с�A�ZQ��F(SQ�}Οfr턶=a�P�q�x�;=�"�ɸ�(����f�i��Ow}Ӂ`w����@X��6M���
����dA���jB��[/ʅ��e���'7�͛��ֵ�P�/nZ�5�@�z�Y[;��oU���?�ק�� ϳ�'�p	#8pQ��FZ?Q�
���YS9Q?�=t^Yt�����ϝR�m�M�9!�e��o�[I6�Qr�V�� Ha�����3��Z"���%RV�UHB�o���\[��TN{4�%�����#��*�5���q���|�ۓ�yf��G�YZ�jK[���'ۉ넹��b�� �o}��9�8)$Ov�y���AA�߆"��ڢ���#�ho�	zގ����!*���G�.��Q��q�:�����5�p ��(����R:f��Uj$����L[,���C�P�ES`�+��B��מn��`h���C��pq��ww�B��"-yi�.7���O@�K��rfr]���ޗ��'��P�xa̮t7b��(F�(y�䎠Y)��.4�΄^�m�|�yat�Q��*a�P�����D���Y����A�S�.��ŋnހ�u�;d��.��n��L��#j���$��]B�7О���s���W/:P5'6��@C{���]`��M+���*G�f�Mo�*1d�C�h'�yG�����j� �kTj��.��D"�!��a��fNӣx�����|�f�)^2uU�����6�5���@�� �m�'�ˉ���B�]�ַ&�+O����N�v�t;�0�q�C���N��8�Ы'�����N&eJ�Y��н:�N��t��Z��\�n�@wD�O��:9(�W��d������H��3��1���x17M��^S�82�>x�㣗��c%Q��]?����G�n��"ƞ,�
��3��s��Ju�-V������A��ZJo6�}���!���lhs��i������Vu Ob��J}\$��p嫩롔��P���������ĥ���^���ZvJ)T*��&pj�)m���h� �QV���L-�#
+�����*���ҌS�y�I6�V~X'B8���6ۼ4u�nTTHjy\i���i�U۹Zx���P��ش�u^u�Ñ�5��k&2�Tۗg�LuV�5���/C���/��wc$�?�6mHh��ύY/O)<�����^�!�!ۅ��0u�;����M��Qǯ��n�14�7���`���f���A
Х������R���Un܉���h�Ø����<3�D�p\������:l'��
�͵6{�ر�c=N�1�X��]�nzc��.{}�㑛�[`�Gw�2�rM��u��n�ü��Va��h�7�LwY��ęs�&�E9]���t%T�0�G~&§w�?=VY9��?�>�iV4.�p2�g2�Q9�����ɃK,dÉ���vfUn?��85������5c��_* �_"��,��K�\D�@���o��$�i?��	8��)����o�_c� r ���?Y��KN��*؍�=��!�z�	^w�dW9G��|�ӭ�^�GQ�B�NCj�U��%�Kr�lp�Stb�"�����v/�e���rn �����	rmA-���`��7*Oh)xU�j��-���C���}��I�n���1�� ���ηy�nB��* ��˵ķ��Q�ۃD��ĀA!����?BN�B��/w�*�n'���|E�@������cO���vK�\Ξ.̎Y�z�ػ��n��3�?��
}J�Q�8St�.W�����W���"\�k�O�a�O�|�� �	�u3��t����� �cƨB�L�i2���i�����|Y"�QS�c�{�Gj }*��Z��u�o����I�(~�F��y�����*UwCփ�9x"3�d�P����)6�噏Á��&e���Ho�f�f؋�3��'����k��͋	�7�!Rs�1������q)�h��k���X� ������\��B���D�}\F
�7�+�p����ם?JKh6b�E/�~-k��U�VH�]�ɱ�>4ˬ�8��mj�nF~N����i93��5�'a�c���gCU����M��,�c�tw`��ІZ���鴚�-���E�_��su�t�jɏ�h�6�s�F;����4MBILmg��qZ0��,�Qi����T��I�O��b}�CT�� ,��^�t >V����h��׆r��5o�7�|�v�;�G�`���>W���EX�N�0�|�Į�	@9�f�Q���iUe'� i��X�K��&U�_�̸�$U�CY�BX��B�N��;�Xgҫ�X4NzWoœd�YZWm���9Lg��V�b�pX��IEfҸF@}��KV]�i�7�"�{���#�ncT�$���]���L,˹X��p�9���u]��n�yZjTϊ(Q�/!�@�f��_5V2�K~��+�oC˴�Ξӄ=G�}�Z-���Z۷"�qt�Nr���l�w��i`쿜�왌`�\��ö��w�Ԟ�y-��0U�o:�0jJ���Vf�"��u���ٴ��/��>�M|duP�#�}y�C͘ꈆ�8`5�7Q)����tw�N�����N%��S�Vm�u�]_�����L��)��%�,���I����(��gc[�)P\��:���!.o�{�n�����Z�g�%�]x{F07�lrk�E�Z_|��ۄKӮ3���C�uN���<�K��J��'����8pϪ@���/�` W�y�d!Ǆ�)�0�e���W5����(�M��댹��e��^�OS�x���]/����)"~np�F� ��y$Ih�D����)U����{�����O8jRU����5���O����e&��X���T����2n�����U��Z:�,�*���5e�C���i��~�����s���y��'	�V��`�F�/|T:Gq�Dw��� �u�"��Q�'�1��F�]*-p�r�0�k�6qdôFe-3:���*Eg�i���gn�J	��	�dj��u-�N�k�����p$����P�`9�#w�ol�-���*�0�)�F���L� ��6:o�5R�ͼj�J���Uv+��z}jP��?�=��d�F9��"ЇS��zB�-�e��kH���Ĥ�٫S���1���D�ϼ�Z
5��bS(-u
S���_b��L��K�j��<clۜ�x���hy�P���7z;��E���p�Ha��3�Fxo$ �`�R.���2��y�.?М�j��V~F�X�g!)��Z1������_}�FDФ"�~�� ��1LlL�ژc�Y�@��8by�2���{y{��89K̰z���ľX\Pg��$I�U����s�tXY��%l|���D��M��#�@*7n�p�E-��	l]	P��4���K*%5�k\f�󖳆�ab`��dǀ��
��l{�k��)r�~�Ks����`P�����Dvp�NvD��q�ZR�j��q�g��R�L?�D=f�SW�r��N��/����A�?�jԬ'�w��A���l�����$��`�={FZ����k����T�~������* ��u���pe�{+���y&Ý��ɘH�CH��= ��GX�^�l@�W �ѯ�+�8���PO� ��ml���^��įԑ�:����g4���;hO���?�P��~ig��<6����|��������f�U�1��`J�%��������`��R��)#!�i?�E� 8�*G�d��|��)B��H���Wr�k�"�`�E�eA �؀UQ�|�	U���j���"�p��T��>�����<R	A�~u��n���1|&�Q]n���k�޼�/m��܄6��U���>7�BZ@z�ȶV��`�c����ހ��H�ll�n����VϮ�9)(���	���tR?m�'�E�O"y��A��0�2�F�����SM��F���xc`�u��3�t�G��s�ޡ��vC^me��w��vaJ*|8y]ES�_+na!�<F4;Z]�ݒ�i3<d
�)&��Nkx�s P�;Aꮵ|Ǌ��]�2��I4�8���b����'�g6��^�M�(J���u����������M�����,����7�&��Vʎ�������AhX�j&�n�عM�鿚=�D{�L2���O�����K��
o6
��x�j�5�W������Ņ�G�L�&dy^�Ȫf���ח����A�L��*j�M�ݝu2SB��C�E묅V�o���S��G,�ɻ�st��˘Z����xtը�m�����|k��r��/Pt���S(�p])`1�b�ܤZBP������!�k����%�@�nB��u~k\�W�M��T7����.��;d� l��
S��E*x���j���/����3t�牆�bW3|�ϪE��`B��w�H�o�2Œ6��w��ka���h���C�d3�~�/�� �M���<� ꙰r�zdt�rY��_$�F��G�L%���t����WM:y��E)zqmê�L͎8)13��乓��|>l��Y�R�e��9��Ȁ�����'�,����.�2�1����7�p�6k%w�	@/���@Z��x\�ù�w�P�H,T+��u�?����o$q����h�=��HuL���1VA6�~�v�d�gH��Ցg��G2�Pfd�0���a�[�����l����d+;�g0���L��$�b.�^�82ò�g������� S+�lQ��K&M�T��#�^r䛀��3/�~j��Ż)*c�+�&�ڇ���[�$�����+lY/�~<�o���Qw�
��P"3�$�Z;x;����4�.���Id�םqP�v�xdL3%O^l$$��=��Ku�ϋ��n��CG�)ƲT�D��̕"0���t�ڔ��:��	��{��"qA��K@^�4i���h��g��	o�;GK�'�����Z��8���ĥm�}�Y��b�˵��߭avj�=��2>�)�ʙ@,![l[�'B���_��ҋJʬ�#Pq�d�]���(�:ր���HSš$���O@�ڽ��0�o{/j���x6Ei�� ��8!�)M�Ƕ!��.�ǣ:]o��ތ8��$���r%�>%אH�S�����!ƾy�S�B�6����x�{�Լ}��K�{�ޱ��Re\�+V�0Љ�V��;�;G��K�W���JE� J_pS�Y�����
|��5��!�=!v�����H�����&I�u���[��.}�d��zb)U�Q`����r��E�.���b`�&��\�ѠKb*�����L'�+�&O95����D���N��j/���Uwף�{?�΄'�R���u7Tl>)l2 9R1��!)��Ͳ-h�d��E� GָQ+����%���.5��IB�c�gfΠ5h;����� ���c�*�ۏ~�m�y:��F�u�c+�(נ��I�	��s�����Ȫ)rl�[7q���܃�w�Q�g�Uw�YI!4&�� �:�8�1���R'd'fPV��h�7�q����B.�fT�W����!2�;����o�1s�֌A�����P���\p�����d	Sl#��2�^ ���KbܝТk��	n�
|K���'�G���(�J�؂Y��`�j��6�p�+�=�S'��s�2y��pRcA���X�=�X��� z��#���kND�c&�@�����,F�Iu����=@��c�2���?�r�s^��u�M:�7(�����̨��XUY�W�nq?|Y=��`]ދg2����g�����;s��;��a���CH���#-���&���A�r4�Ais�nyF�C8�=$8;������/������Ig��I@C9�bY��m��r�[�l�u���<rW�g�U����x�ԡ�I^k9H�k2G��DJn[�Q9���@` D娍('�㑨u���l���;=>�e$�Z�0~�O����(�G,jpԱ�/�����W���s��q�C�տ8g6���z<g3��x��h��d�����,,��/9�=��V�a{��9_�s��!��*L��s�A)��`��y���w"R�/�砦��%��:#�&�b �*�~q�۫8ѿ������������>j7�pt��>4|�ih��A�����̌�x���z���φlZ�h�1�#1鉣�C�Յ��n������HsK���CS�`��r���J����D�8�VaY�Io��R^�a����M����g�q��v��S�Έ(�#�q��(2b;��NQ_{�V�_�c�B
b�}v�9$�/���%!t�KQr.���P_�e�>�Q�X<�1*����Stz����Z�V7�?�;M��YJ����W��U:�5�g2�d*��ȬY,�e��}���M����D�X7B+���{�B�Y�ӑ�2+W4�v��}��QV���Yc���=���U��w��l�^��Q�k��D��4��__�Nt�&��b�\�����8�N�� i��D.��#;���0��Ro,sv#���S�h�c�wD��2Yv�ׯp�o�\�흞�Ma̘�1������xm�������ԳcS���zO
����6��_*����.�e������X]UΗ_Ȯғ9.���W	�Kh�{���z�$k���&����,�	`%Nx��@f�����Q�G�hr��4�C�L�oy)�	�Ӆ�������_s2�x�e �_;_���|7����Z�&Uo��_�s����P�W�� y)<�-����%H�h�H���ILE�GP/wE�/׆wO~�en�R�ǨQ�c�Ԍq�^z�vK�b�8Y��?
��*Dwb[n�5�C%,��_n����]�>�I�0��Ք�w�u��М��'�!�X1~�G���ﺌ8ה�♫@��T�2���B��pY9�?��Q}�f�ˊ�.Й�$`45�enJ�̊�Yl��R��Z���NA����!x��&߯3�_���]���М���af�:��#��gxn��d� ��������×��!VI�cf��]�b�ۯ�s�y0�gN��������`�Y�� $yV�(��I�h�Y6k6\��>�\����t�"�^��2�̵iE��߳y�ʡ�[��fN��h��A\��guzE�~���ub�i��	s:�F�� ���m����-��U'�$�[C7�@�io�FQFZ����Co@7E��>^$m/B�ڥ����a�@�:����$����������p��kL72�D���y���Ho�ܴ[W�:���ɷ6���nK����bvR��L�MЁ�wD�/K���y�3�[T�\�v��ppF9�6C�F�)�1��t�6=���r.?���B�����r��q���$vP�ލ�ng�x]M�q(]��NZ9�]/��4�|�UF����@ S��H��A�|��`�`6^�n}� `�f�]}L`R�5E�c�34y���_�z@Rw�k�n)����w?+q���-U�D�9���r��V �Ag�&3�h���gn�&�PfL�ܠ�L�+���G��f+��~�YU��X����<�z;�}?�px٧ -I� &8�!��R���H� tm��V�rB|�K�����,1^�����*�'�(:�����S앨����6eS�v��{�t�T^o)2�E���8�����^���5$�V_c�s��dc��0|��>�W�ȵ/j���8�ܬz���M�.�#9�̲�cn)�t��9of�,���@����;��g-���1O��zh�J=���(�d��G�'p�+��bSX$�-	*h�g�CB+!3q�ά(;���	to�
*�;7?�q<��Bl�SN�o(1��Pl��YH�}䚨�
�Pu����j&��ۖm4Q��H����_`�r� P0�B)�H\���;/�	9 r�i�9��q�-�wR#[,R���"�ZG���C���Ps��JduU�*�߾��n��_9m+��)�9��3���S���I+ೠH�/Ԡ��ۓ�egO�����	h�xe��#L�sh�k�����O�6L�kU�Jg�$�����>|��E�r��NL73��<����w}�ͲE� ��iH��.�͕,�z�m�"�]~�8EX4i_�����G�jP�K�r��&�`irJpż�(���n�>���DV}�
]�wv(�n"٤�*c���k/�L-����E'7�n,��Jۍ��r�J�d���8��I��.���a�Z�0�QR��'Wg���L_�*-�9�phs�N������>~P�{u�݊���� �_[g.���_l���!C��'���Έ�sp'듬�~I�.�DW�:s�Ww�A�AGe����\�X�b}9�*�T�����.���������r_>S#)޾����-��:���ޜU�X3kDM2�-WV"��㹝������P����_`��ܒϺ5�#�Q��@制�1� me�5��4����E}K��R��}���>U;��!!��_u]�Bo�N����8�'�S�p�:��t�|���4^�A��{�������u�B5�Ѫ�n�-�?�=�:�O�;������.���cF;"~�_����ʎ~0���B�|�%����S�/R�������F1Y5�J ������,*�%���o A�Zʃ#2�IT>6��� r��q��b˒-C彲��ز@�G�Ք�x���Y"������Z�>Fl^kF�{�/F[�o���U��i�^� 48E]��~^HV�3�W�I/>?�#Y���K�u�	u�z������aQ�4x�yOXL˖,� ��AuO�TCB��B�Τ#E�`�h�TY'`�Z�r9��#W7�X�-����ψ3ܱ���Q��vG�eޜ	�~2ᓊ������W��N@#<M��ς@"�v����1���I��x[�Q��1��3���rg��@=\�G���.`���
վv��JT��K�R`�;k��P71��o���©�����a.'�W�)Q��%#��S�����[&�$5^c��f��-v��]��T[w i��ӮNp�e�|y;�_,�OG��'-�o5ν��5/r@8ji���(l�\�;���A��b�=8��YĞ��鹦0>�y]���[�E���:�w:�6����1X��~�+�0h�v-��i��䞿'|E�sW�㡊G����@�@�����x��%���(���Z��(�̾���5/2�����t�Y��L����))5��5�]��5��y���3��Rxm+o��NI �n��7�8�;�ϓ��G��!D���އ�>��g������Ƅ���9B�/���f<K�):�/��~ub�g �|ju��B�^�"����f����~�>f�7.��븮���`FLH'8�E8���E�9EIB�V���C������	4��r�V�_0�~l���܏{,��F�%�E�ވ��ԍ�W�,'	\�z��t�p��c�ۮ�\�ޚ�`��*�-�t��P���c�����մ/�L1�ā�K7a�1��ݗPq�{ *G�N�'�^:����!o�x�����]���m~; ?�i����[�Z��soW��Ƙ{8z3��B��'p�p���-�R�.�7ӷ�Pʵ�� 贃��!����O�	�\b�<��p���3[3��܍X�b��a~S�b�~����@���z�W��/�:�W5n��)�syي$�*IKkO��=W�j���S�Yl���c�V�J1wCr�"�z��K?{���0��}G�]tUj�����ƴO�����7K̟v��4���L���AS��P�R�|����#!)�{u�=0�3���a�)g�Y�0���l&b�7u���I3�&ǖ�k��� YE
c����PѽW�M��� �vA)��\Z�Pz�W!�����f��c�G����h,.+��p���U��t�EU��mJA�}�"i���䘎�o\B�;�,��@]��ex;&�{�'t�uB
����\G���8�Ld��<��$@���m��:R��8�e�P�������YƬ��Og�~Y5c�,	,}��}�!j�V��DO���1s�T�~�~\w��T�QɁ�nFh �,u�M��N��l;D) P.z��8d2:�k���MUql_K���0}�]-�qT�(�<+J�ɿj���T�/vǄF�#�NQw�u`ӧZ���m�X��XG��F
5�;����b]
�tH�j��@\�0_����$�[>E� �Ph�3H�å������jg=kx���*�%�m|���w���þ\)Ε`�(��S){?~^~C����6~]ې��$|�ZlL$���R��~�Mc<7p4謾�ͯ^K��Y��pY��#���!�(Q�t���y/k���Q4N+�N]ʸ%8�����2{��j"��}+�R���6�#�(����C"�v���k�ft3�j寫�f�B���^<1���'h�:�7�s�{���;
��`��A[�Ff�*̀n��5�V!:�
$hW������q��_���C�gg��F���:L6Ǵ֓��/�F�ʇ���ݰ��X�X����j�dxmQƊ�tՂ�i�1k5�[6�3n#���*��n?�:�L�\�(ԫ���E�{y%W��x,���Zip;MA�	h���/���hWQ
}�5`�%���1�
��U�KY���$w5��W��������N� � �7@��ϻb�B1���fF Ͽ�ml�Og�����sO�<Y~�����5���+&����æ7p�C�kr����n�Ӵ[�̯�=_w7!�H3�l_�k-�b����p�*@֘�!1>Vb�֗�b���8��G⢊̜�ۃ��&���ܼ
���YC���KP��W~:L�!.o���/Q�>WC�d�qC}׻x��Ҳ�����Ʒ�T�c aSY�~����>�Skgb����C3t��#�9��!���tz�%y0�PI3�l�z"�b�fE���bA�`8BT���+]$�3�_�l����}�ӛ��eN��Y^Z��:�� �]�ԥ��}��H2�qLf��[�	�u�`���S��2p8�1p���!�x�!��J�86�������v�d2��Ŷ�y�r�̾O�52!�AZE�$E�IG��n��`۽=}���b���(_ش�\� 2C�U�nO;d��021�U�;�~��7n67@�^���gi����@+�3��2N%�.(>��K�Cx���#u���Q�����Ę�d�K�Ƌ���	ɂ��L�{Ǟ��JS^��r�"[�h�K�9��,-�����S�o~��]� �t?4&��w��iX�Ħ�#��r g@��U��j���������gL|k���bJٮ���A��W�ο��Rg>̯�_V%R��0��'�����ɼ�ڑY�e��T��u q��o�®=e�q7�3��98��v��}�T��	�Hn��P���%�'V���R��Y����O�[E���u��t~�{l/��;�0�ឧ���<�+e!i41��������� ��ۏ�ؒ�C����J�bu
$�?3�P6�ط1L�����e��A@�˙��[�B�f�*�1�M��$L⪌���z�K�K�6���Z@�a���)�ՁА�aA�������k'��~��"*ٖ�]	k\��9Z�yW#�K��=��˅��"����zս�<ٜ�T�I0���l�8/u�I_�W�K6�
��/R��r�ʽ��h��{Z�5훘ۍ�qPn$���h�p��C��XB9�|c��d�^r��uR&�V�j����٤�^�1M/��kէ��VSD��/�'���2��ő��oMP�*T��/S�6��@��['����r�~�����Y�xa[$�ǔBM��.��Z9��=0�cg y`l�L�G������p�I{WO^�eQk����k�!�h��4{���6�'�G���/`��z�؊�&md� �퇔;_�G�|-�}�	.�D���hof����`���.�]�&�m�ԒL�J 9-gꑲ\�J;}ڝh�	(�+(D.=�?0�>怯M��6�70���!	� ���<�N�� %�����o¯�ǿ~l�{E��>g1�Ӑ�>���^u�W�-��q{=�1�qvZĽ�܇1Ą�~(�g�J��T^,{J�L��e�CUm��S=�ץ��r�'�_A�����і~����O��{���2��йh��y�+Dl��x�����%�)#,c7+��/W�a�,����&l�Ok,E�i���\� ���9y��&a'S_/���,+x�=(����ڕ���Z4�ޱO���fɊ��O��v�Y���eSW���0]T ��Cd~!-ro]N��"��*Y���e~ȗ/���|���:˵WZO�pߵ$\^xj�@����}۷8
>��s  ��M�8�e��k��n�C�O}y(n���˸֙��]��E)�h0�������ǔ�8�nmL��|ʪd�y�hn�濋�A�����+�v#7�S7�.]�{�b�����A�Ǫ�n��S���`�	�/�^t8��ܰ��=%M�W
�(�[�Ìa�x�1�4�����۶AY6Ȭ����S�7t�NK�_��E�������1���V	|:����-r�O�hRH��c`}x2(��9�z�=�>h�E%a�x
��H�(H��Ѻ��!-��gh�_N>5)'F�h�/��"�D�H�#A�>��i��14�
��{���Is��x���N���(9�K�
5Ƥ��ۗ�	�����L-���p�a����A��k� ���]�9]�\��O�߰�&�M�,��-�BĤ^i.XG����&����Y��e9Z�s�+���=�u?���'��,��8�f��n���=����iZ�^q}�.ȑۇ��y��
R]����sQ�%�{�z_͘�T�O5/���2I���5վ���&N���6�m ��e\o�C"��˫-�p�Ĩbd��N;��8o�e��f���x��V��dsA���{PK?/�	(�u��K��V�+����`�/G�G�4e�[��k�94�q!>Tb�	���V��5�*�1�����
{h���/���]�K�
�F��.u�x�e�f�G�y�X�v�`:-K�o�mN���޵o��b3[� �Pk^�w:�lؚ�}���EԮ#]Y�������n���!�M N����WL�(]�g�ꋭ���F�w3v\·�4;���=��	�{\<Z�*,^�M��#R)���S�X�'Qq���[}do��\�ة[�sr��؋� ;M�E�~��Rzx�@j;DV�[i�m��,K�/��m�t�ߙ��Ϥ�Dw����lBt�&?��V��Yj`�Ψ��2��:ϲ���������NY���cު!��[i��#)�K��Ä�I"ת��Ö�>J���S5Ơ�ݱ�{�G�z���HL9�X�	��ݩ$��M6�C�=~�L1V���8���ɒ�8ǭ	7P����u�E�.�%Cu|	���K߇�;��@)�����'��>�Q�or�!foߥ�'��OХ����o��T9�����4�p�Ҵ'�;�6�"_��{w珚�I3tɇ=i[���f�<�u�B���)ŝJ_�Q�>)Xē$�j�B�i	�VxW�yh���Ft�KOu所���i��?+��� �fܪt�����h�l��Ķ�JJ�_y�7q�s�{��B��d���LP�qs���UՅ�$%.�Ms��f�2W�`p�\���@��CP6E�f�|p��}��7A:{i��m�$�:�n�5+�M�H���sFcrc�8����|�fVf�\YL���lP��(�
�|-��IN:��]{t���̞�T�rE�a��������ߤ�xB
���M*�����`Űq�=�a^��+����H������^�P�:#Cr���$TmYwFƝj4� ���}`h�\�c�f>�j��US�T�����	S����:9�RF�L�6�v�M�+�1}��aS�ճB�f֘��O\QS��L�z��6ѹ�k�*H���"K7�����>�C��X2�5�}���{ʨ����g�G��4�И��ݘ��Q��(��K��P�7�x'�q�m�>Ő7�A-����iӰ�L���C.Vv��r6�a��Q���4>�I�
�h¾�E�\�Ӧ؊A�Ф��¬���xd�ŋl�3v@w�v1x'@Awz�]�D���@�6����~{�������N�n{�Bt,�q��uήe���ō�Iץ4�-F&�B�0d,�_p7���3���+טʳ�J�L��{z
�%,���N�;R?@s�z�lEm���4U�43bHW�Y��>(�e�sW!L*^��^+ u4�>�g&�Ĥ�d�"�垼`�5�}�⣻KZ����TE8�Y�J�B��u����I�@
ܨc�yׯ��mp�� ,��mƾ��ֲi4��y :/4�·/�q[Xq�Q]���C.��t �$�PN���ձ(�P_h?��^�)c>�� ���G�G
Dd���)$�^��JG����O�,Igr�/��zw���2	`��d�v�w�ރK��{�G;���4?�k�*$�g&V[p�	�_~��c.���>���8p!߼h����|�������۽(����r(]�%�h��/(��AHR�������*= ����g�Z2���� �>T��V���U���qJ$2���'�����N���cw����G��4^\RF��f�!Y6?;9M�0�	�.��v�OHq�*M.�֠�Ǒ]����k��+�z�֪buyϊ$��
?%g�+�-�*=�&������u���r���*�T�Y��&)�G��<kX�*uӾ�_cE`B�
2fJXC��W���5�׾�1b�ʏ����4X�o\��5 ��R QCO��uC|�@��R+q3Y���/h�������m�c�-�������m�!@�h&���l�����U^�M��ȏ�:gPW'a��.�Α�7Q�"��f'�2����9�{ǙF���'4�.�����7y�uZ+�!&��Ţ`f�s啀H ��f�Ŋٟ�k(�?�2�rӻ��t�r�gp���.xo��g�맫(�$��u
ɌҌ��:��h�D�HP���5����h�=	�S]�gnV�#�����z3�fp��q�`"f��SL�|�穙�Gc������Z���\0�A���r�v��1`��##u�U��gK"���H�ٮ}��ȧг��t�Gm�̍8&�i_F$Q�������'Ǭ��!�o��s\p߾�\�?C�Rd����Di�J�]��͔(2�6d��t�J��!�����[�(�Jy����x��}�Ō��29C�՗v����]��{�1�E�I�N�X�)EV�;uF�Jp�&b����K[7vvxפ�C1�Zr�JJI�ǜ^閂1A�B��ZR�kFZ�B�p	��k���h��+��1�ޏ�#�Y�y�^_٤���5�+'���Χ���ʞҤ����Y��喽�o��r����FF��Fu#�9���0���<���flQAM�N�w��s��LxLP��9�$����ӎ
�]�|��H���p�eE������p5H���n�e�	?��M%����n���ϊi�է\+�Fx������gV�(����~य़)L���J�O)��zb���M������GQ���¸���va��.��%C9)�̳��=��!:�0��Ǯ�i`�U�T"� �]�������.�ڥ:q��Jl�d����\2l���@��o����潫�PpG_So��=۳�)ġ�ux���1���"H4XF� e�p��d-6��{=7b��kB�X�f�>u�{��K
dYC��q�@Hga�K%#ܲ�/;�yY������}F����ǿ�NA��3��}�l*�q�$2��;�R}cR�Z7ɠ�NjSZ(�[��Yw���Q�e��w<k��h>k�1��\��&]`z��'f?���S��V�CW����Q 
 i�3��N� �5?}s���ƈ�.)9ħ�|0Gk��P)d�9���E�~���B�U��AU��r�,KP�#�,~"�F�&�=�Y��� 5
�M�4g[QkIŶbS/���ٰ����%խ����^�����3���c 0!:�]MY���"pe� ,��"i�}~��R5�8�f'<�]�2�]����W<�� )v�uי��`���ԗ�E�RYj�!��ۗ�l7~�tE{3\%�����oGxn���Y����W��7h��|���ᚨS0��Y0A�ɘ�1���U�mt��2K���HH�<c��p���Gb������������33,�@=k<F��y�H@`�R��V�0lC�x�������
s����C#+���t��;�*J�i2�oC���3�z$�~�i�%��E��>�I>Um��ʙ.#ѱ�A�0��疦����j��d�����.O���A4O-��M�eD�n��Z0�ѯ�{��M�a���v˪oj�x$���Kb,�%Y+�#����l�?iI��uo� �atN���Ua�D�n˪=��QSX�;��{��~��$i2�2)��4Ŷ�<�U�>�y1��>�#��jH4��k��dV���09�`�p�!s1|U*���xs�ZE=ӟޘ���	��
#8g��t�@������+|�}:i2�J������k��+Cg�$��"@�!�!�}��&
�C9%a�c��O�5���LB1y&�ik��Avi�؂���8Y��^��}P�-�+Nl�����N����9ytbp䨞�eO��c�������ʻ�v$�KJ�M�?<������z���� _��>�� �;.#7K~.�}O�,Ɍi(�˚ i���ݩzN-b����k"2�[���ȗu�Y���s�D=�	�>rV�J&,wx*b�lx�I�>���1�G`��N��)L����O�m���/2�&��S���/6��4��O>\�XnO�S�/���><nn�j�Rf4jN>�� �fM4�cͅ;Y��"�A7�'�¤��8O/��;�J�V���3Lƹ.��'7a*�q[jC�(��}fG���ђ�z{p^v!�k��wU�������:펆�/A�!4�a�i�!;*�)�j�-%��~
�J�À���'L3��I���Y�xl���� ��>��,�i%�Ԍ�)���y���7 Z�+��4&�r�Ē�����ԟm��o���~�(�om�����Ն�9Pt���q �ͱ���)�L�\T�� r�	�b�Ψ`D�[��GO���Լn=�i��F:Mh��r��
����E\��i0:�!rzP��םA��N����w��o��Pm���K�2چɨ9%M�p�p���5���XV��VW�Z�LQA`HjW��o��؝���	�|؞�J���UBf� �����A	��e�H�-�f\�w�����Ri��S9�����0��8�={ק��1`%��(��c:�ymI}>OH۲/��l1q�����篍�l�O�ɟU��E�*rM:z_	GZ?t�O��w��i�R�Y^�#Z�Y&�^�,��Q���:\�?�)�� 0�pj)�"P^��\���TV��OI�����M�57�D�i�Gh�`%����(�Ł����4��Q��&����F��� ����'D_�og換��n�k����Yt1\*<�6����2 4~ M�Ju�j�G} ��Z�6�RW���1!O/ǉ���{� ����.���L��Xm�J���Pu�|[�5�o�v��v���*i�s�@�"y�O>������E���A���������i�	�+���??^»z$>.�@E��aQ���@��A��Z+�2���&@���&�]���?�u/i4]t�獞]~�ѓ~�'D(f��b��(��/��G�W�c��{hh��.�]ϋ�f��㝰��Tj�
ֽ8�5��Y��D����s$-X��ɶ̊O1ҘBL�@�``��1�r�"%����ꓕ|E�&_�?P��<�n���t������8 e@"�h��>>�0Mh?%� !��(D#+֩	c$�ė(�=i���	�(��Ҩ9 X╓�|�.��Yt1��r�1)>���{���g������v��79`��ϊ���<!2~c�5o�nl�,�Bg��%L*�6
L�F�'MTb!����π+U6-Y�OՑ��#�WM9p����V˘(�P̔D���Q���Z�e���"�R���|X�K6�1�yˣ}�,��h��g҉�%�J�1N}U+���rϐ�����d�jJ8 6��l�N8��=�t)�Ԟ��K�2Y������c��[���V�5jNr��.)�Z�6�Я�iҪ&^����Ş��09�;�4�ć	�i3�������6�V��K�Ù�)X�`��<���F�2��DS�Rf�!#�c��g
!�|a�^ :��L��z�޴`�e�w�}� �;��Df��k�-������K�w�D���UmZ��F����W��<�s�j\I���#g.4�Q���t	W.t��:�\�s7��%5� ��L�Y*MTo�/�Zi5��u�oc�����S�!?��g�'�x��m̵��4��6�
��mJ�����|O�(O�H�"]��*��.����kY,~H\���z�� M��ݰG'��g.,�VCx�E���7FfXN���-P����Z2���m�Z)�t���.�/��/�zn�7ϜK��:�E��L�$ �;5�����=>�F?�J^��9��o�J5��$��OE��؀?R�/s������9��6�����bᲰ�H��A*ռL{�)ͩ���`�P��*i1�:!�,1��{aj0���Q��Tv1�J1S��zF3[�xpV����xf��JW(/)Z��izʋ�x���R�<ۀ�t,����S��1VΕ#�u��Խ{J0��Z�x���h�$ܥQa'���@��ǚ:[靎طK�]b[x���a< �?���*����s�oFu��U��2�ښf�&Ĳ�+�oϪ��yD8ƣt�֖hY�Lx�J�T3j�Y��&Ƅj����ٓm�	�㪢9*���>��e�*7]�Ӳ�E����ջH���w����>^�u �W�!�ji{}_Y/��'{�SY���
�M-���!�o7|+�	$�$H�,ߛjv����b�{�,=�O0��#��;�K	��A�S���hF�II||�AT"�!N8.1���c��*�S��#��DbS��b�*R�{��l����P��6����k�~�p ���\�G�E;j�{ZB2g	�v�ڑ�D����wg��ր�X����w��}���m�0̴��u���R#��3���H��
M�����a!]��KM�.JU�V���<ݙݳƸ{E�R*ԣ.O?��a �ҚT�,+Z"6P����"U|a0�H��k�[�O�2���O�P����-��(utm���A�Y0k��,xj�u
�Rtv�^���b���w8,\��8�і �ֻ�G�	#럾|j�Oɩڶ�ꔞ�f�}bV,�	�[1B%EA��_�^�%���-�1��h8#��p���iu�v�8A��#\sKT$G��D�l�{�|��lg���2[�ဇF�FC�~�}m��{2�]?��_u��:6�wtBOo(�Mk��iȸΰ��2a9�������2�˧2��V����� U��;��S=��<��kş���#;�}�&������x�]���!+�����������ԭ^
��M80��`nYI�/����z8Fѿ͖s/3�詞#���0Z��Mb�אfP�y"4
*G�WUc��-��8�HMk	�e�,�FlH�V9r���՜P��1�B�������j�������E5�#H�%>֎	��B$��t�l�Y����t[gq���"��:��d�7g�4r���!3�~��)[��Q�r�)9
���ur��)��Q?9M	�xT���{d�rE�u��Q=
ߙⷴC�%�E2̢��>>�x����^���ڨ) ^ޮT�n]s֡�i]D oc�H�z%�y���ik�[=�����~
���9m�!��~���O.�vb�z	b����p��`���/ ��띯�̊�6��Z���r��ja��.��{�hMB�V|�.c]9G1�ܴ������զy�7~T�u��	ZU��aX889b�)�lh_�~}��_�H�舽^�i�xI�.�����yu�k�;�C�~���M�ˎw��5���8\C��r@��W "��K˕^�v�B�
��Tq@NR�;�`{;�:��2����e`X�d2�/�4�Ȳ�aJ�u88�e�#��C��)(�O�4�Op,�����K���rvӍ� M�t]@F۟BZF���Kꢱ	�� ���ʊ���w-�-q��?S��#�ǫǸia�,�\p�Z�9�� �ɣ�|���'��ϔg���ܿ�O��(ݠ������#��[D��R�f�|u��y�z��#@0���a#o���3��&gJ��l�8�z$�=�3���E�]��O�d��m���*���'�%^�������O/!�꨷�cow?H�&U'7!Ƶ�n4Ju��yi2h�j!����бv����d.��C�5�'�'.ԩ�R��\P��縋̮��dB�yJ3U�W/�1des�N���,bx��_%����d�|���%!�Mb���S �eH�x=$N#ϳ*|��gY��Bձ�60L��x�r�X�~�W���������8�漿����C%��6F!���,�@���D��iF�`l1��K�`�:	���E5��e%�@I!�K��h�>a��D�]�����7T�I���m�hhbV����թ�x�e�O�r�W+��*�dp|l< ���ݻ��j*��cQ	���Q��c#e�,6�G���M9#|յ����*��jS����E� ��4��E���j5��>�Y�</�:Ȇ?�$�p$/��+������ i��7�N
��G��	r�d��5,5�{�/$��I�00%�q�a��Y�P�C�3�kj�0#s�պۏ༷~��9�u���O��F��lˡDY`��6���u�����e��O���w%�Y�:�5���J�x�M��JTIr�9)�������MfN ����F(�"(��;N��Z������9�~ܧ3��x�����3	������vӛ|x/��/{�'Bh�o�W�G.�bh�U����p�j#F�o����� _k� �*	���f���ހն?(o�p;�cĘI'��+�M����7����E�Jk�ٟ���fJ�/�N��vX��nMB��8�E�����a�d���)9YwA������r�k�J�giU�qu)���#�dAd��.)�8��g'��4=S�� ��2���.3~��&c�����b�	�@��D�����������)��G=��	�;	��.�A�g#����6�4X.�knnJx����l)��<�D�:�-���ð�X�C���D=d	�ƀ~w�D7YR��&�D$ͤ.���u�U�Z��9&2WDʈ���X��:L/��?�d�¡̡���c���r�}�C0l�|<01�dx�b�H�_P ��l�FX��Xt���%{�S����
`��[�*S�ިH|�kV�C��C�QX���?8,��0�*f�nHf�T4/�4�l��%�1�������
J*��3|t����Fq���]%��.��31��H�,�.��Tff;fs����)��n�<� ���pO���������D<��Q-5��˜ЃRf�$Wb$g
tf���%t�l[	�x�c�HtZ����s�Ӭ�n��k����W�>o��1�C�r�K��pgt�8s��>��3"y<Ӟ��kv(u��a!�9����>�)U������J�_�gt���*���3{n�t2�r�h�������`x6��$A�T$5!�vs�Y���n�yqᑾD� �3<�	m�q�y��88���4��ˋz)��ŕ�ZX(��h�f.1�<-���n0\���'H��r��
o/#�o')��e+��l�.��Q���6�NS���+Q�1-Ҝ�b��yTH&
�#���)]���\�	M��EwsM�d���[S*���W��7N�0��9h!���?��{YͯbK��Q�������#X�������jr{��-�qX;���N�����VE���[W��u�H�]��$�y� mĉ�Q{n�vӞ_�%�� r �IQo3 �������$3�K6T�(<%h�l��"|^|U��ǰ�y�]6	ݤ^"�!�k�����38���BH�	�w�A׽a)$�����+��(��3Ï�oh����M�ޫ�#-M����N㴂�ő�Sqixޔ1�B�V[�bn����۩_���Ǹ���:`�w�xdtW��/���}ŗ�(C������`��V�����#2AND�7�x]���Za0�4�Ld�ӭ��N5���R�c�N�G~ �b;}ţ`2�J	*�ő.�& ��I'�{��s}@�8��-��U=/9+"%'7�{���/% �Q,3���� ��O�t��ĐTnu����]�J�rvc�~� =��.��G�lݏ]'*u��4�e����q�ԘN�Mh��ݱry;��Z����U0Sc� �|Q!/܈b�u�>�5������b1\A�%��z`;���mcy����?@�@��9�L�n8�ϛ��OfP��kf)k=�$�³3��1#�~��v���u}GB#B�i$C>=I`����L�V�� �0�n
�*?_�{^hU��LY���vo|4�� tZ�H�=c�冾�v^��:v[�J�Md����naX�>�s����'CU��m�鶤RuO��4F�<�d>�����h�&�o���K޿�pe������tR%��kc�.���x��}�$��{��Q2̧-]����ou�y#��:�C0�松 ����kC�u���0H�~���hd�.6�5���(�Z�u����dJ���&[ !s; k�u��h��XvmL�r��^ʇ��� �1��.=�%e��?d�@��\6��SO��KA�Y�u�Ps�&0�ve��}N��FC�o핡�ؼ^�,�֘���	�e�; �lѫ"�zᡰt�}�'+���RgDl��5]�k�@�r�K�.!Sg��ux�g���O=����E�	1ιׁk��_��I���RCx��B8�.`yw)�"��8��ͬUI+_ɒ-`�14q�jk���A �BJ�s�>3���nR�MŝM��&��md�7ҫ�Ew��pL2�gw���^d����r_�������xj�>��b3�~
/���D��1��a�ĎQW���z�Bo<�(g����_0�(@j0�zG�)Z"+�پ����9��ꪖh�da��{���R� ��z$c�ĐB��Ds9��xm�ń����{@�3/Z��:���P1l��Q�*�[m_4۷'nt`11K���	��T.����z��1���4G���|����fU�M尷'Q.���\\�v�o�'���w>���(�+�fWi����[�%Z������Ot�ܸc��|�l�ȇV��$}t�$Pj���x|������
 ڽl��K��yL���[��������=�v!n��h����[β��C����x�\��!��eX��o151������fͻ���Shl���u������X���(.��cg_#�Z��5��\�;�{$KUx������n��޸�eJ������#����?�� E�<�K�PW�^�

=67OE�7��gR��f6�YA�$]N��y'�S~�@I�p��n%D�@,��o9�C`R��J=�ot,'M�ݍ�(f���?�~C�,�H�����VWJ�bj����]���&�o躉)����-׆WdF�i�T��	s�0����wC���=�,���v���~�'Vf)��-'s������Qb�
l.,;-
�-���T<�)�B,:���e���%��b�́j��JO%�|_����8���x�)ѹ�������%�t�I�y�%�d�v�	�a4�>��*�w�m	�9�t�dH�(��qP	��M�����/`��ۡ�������t9X�����yp)~�
�f뻀W�?���e���]���d���������@a�y
x�����r�;�&f7��O��Z#��m��yի[[�&p8VR��誉`˸L_�i�o\���M"2�O��:��3��*�T�N����~ÆG�Dv���G�гH}�E2'�����P���$�������(��O�� ι�d#�;�} ��Z��v�"��j6����'q+^�.%b󱿜��K>R��A�e0�J����M��˟��БozZ{6#>lؘ����/ʜG�����u�B�����D߳�O�>c�ּ���'ZM��{g�aSj�_�Um�_S�i����߭<����O��HKZ(3����7/��#fk�!D1�BK����39܆1\�,�f@�fy ��7G��|���~�;0���c�����li����%�$��h ~Ø��#�)���f+���kcG��[�SV��bF	��F!�
��
t���pܾ����,UC�Y�Ve���|��21r;n/�PR��'��1����Bk���X��RQ����^�c u��f�	h�S��+�#��җ(�6fe�/9��N>^�����i2�C�>"���`AcG��s�A�tv��φ�W@�	@nD�I�D=���hjH��m�v�ZP��ă1O�U6��O(f�w���+�me�0 [~��.v�(Árb<�ʶo�U����e�
�'��x'�	�t)2���B�7�w��6���{�^p4�.�� �+�U~#��*eW����M�0됏yJܵ��糄|F%䌳�B����M�Y(5'�U���{L�W�N�ǽM����a�ߞ�h�{�v��v��eǆ��0(�V Wf�(ű�)�A��Uo��Hц�
�\7.�I[YU!�19$� ZE��NwI����7�1b�m����<�#b9\���tG|-��ρ��	(k��?3�W!m�RG��K�Gj����#�/�!����b�y)Y$¸�dWd.o��A�'��qَs}�����l�f�ͱ1E9�K^>���A7m/�iGw�������&#��{_zb�D`�������`��B>�QU�L%� ?��7�>:��n��k@�g��R�Vʚ���/#g�o_�-����l��X\��Au����������2Oo��7�w�A�F�Ztv 0욣8�CG��^� ��y���C���Q��m'�_�7��B�l����Ss���v�`X�]�!3��6N�������*65���~�`"���ڣ7ji�E�{��w�gF��[�����仨u���������1;���!���
�jݗ�]�!���_$n�w� �����@�ޛ����-p��H)�y��\�׫!ԛ#=�'��=�5H�	(���y������SX|5�s`4 ����jW��:f��;,�A ��"�뽉�cG6 ��`Q7�qt�c3��S�SDx������OwF�n�0�\�:7AѢ+9�����0�c{�	:X�j��a�������`�z�	�C��)b��
�#ë���Gk{}�<�DH{�|�����	=�gw�`ut}��'돝��d�Sat�cMJ��:ů���*�*��֨�!��,�/���Ӹ��'2E��q~
��
Շ�(D	J9V��.�-ԫ��d맚���L���i��(|�T�O���ھ�K"Y�ٷXÓ	[^�i6
ق�v�N�5 �b���}��?}�8$oZ��*5��b#rRÿ(�1�� �2?9|��A5��I���l����?���ت�M���L}�9�ˁ�b$�� �C8����22����d�V�7�Js�A�&��?�ɑ���~֋���+�{��O��֢��樹�
\�:��N�XI�k��b]�{�{g27��b��D�=s&�c0���gR/%ɖa�}�CE��6*Wx�֏�D����e|��Qf�6���)��P^�J�)Y���{�v���J���^��J�@TG�����NL���T>ӛݧ�W�9\Ø����F�3�P�a���F<u�K`���!D�#�%������,�Nka�"��!)*�������~�6v(���1�3T.����]��l)���ƍ�}�LiH�"�Ҷ cM{�.��*��91����l���.�}�Y8��P��Ωk�i��ȃ"&@@`�&-���:A��'~ܘU���PuG�髆�Y��<��Q�?�3�7�%��@�SI�v��ꑜ�1�
��!���w���/���,:�;��"���"*O/� dJf������##��=�'�3l;�Y8l,z��/�5>4��Ѭ����m�}�������^l5�\�����	~�A �ܕؽwR�'7j��?��-���>$"TC[�\�G������@J�a4-H-���X�D$��l;O{�BD��Fƕ@)k�JSD��ܫ�����>;���o�Qp3)�"4�]����0�O�[������D�nJrD��h���WD�3�c<@z����E=cq���PK�9���Lҗd��e�ӭ��3��V�
��J[��ܒ�1i1]H��ˀ-����3�TlK��j�J�נO�ij`�r��P����9y��7YK�OO�Ҧ�����\��'�#��������%����"0}�^�ϯG���k��˒0�f�U��N���ɯ_8O#���`̼.���M`�������-Ѹ�KkV���EJ#��)2�x��x߳�V)S����)��Z���3�`nTt�d1/@��&��뢐�����͢��.��\2G�,�CN�X��t^��!TQNӹ�/��Y��@M�~�[e�QQ������%�߆zFEf�8��D�j�3���OS{�b��Mj�?�
G�ja�Ӕ�~B����1��`�;f��>I�#y�=��Ҿ�鑴Ҷsg�:z� r��[�@e��m�G�I��h�b����3y+�3��H���k��ڻ6�Ϗ��wi��	č֨zo��x��W�Hj�Ha��B	`C� o-=A�W��U���ZRo"&㕜�[z��'�әQ�s{���z����u���z��R�қ��(�hi�*�-I�w=)��B�VC�>z��8aL7��\��tZ��]��B�d�W'X!��tb(ҩϡ���V	"+DU�-��ReơM���eDOoڕ[d5r����:1_S�������F�%h}>�^���"N.�_����u�;����h ?����|����5Z�鏶�/�nWz��kڱ/r926�H�C�NKz�M�s��ؕI�i8Oּ�׽`!1Q�=%I�9`͵/�M�u'XE�e��a\JPm7gJF��6��H%��<�D���;ݵu�Ѽ��Ά�5h�o�,�����RW�	�G�Wt)�sj�-������a��/��X�P�{��P1։�>�%8�<�lz�{GwpS��g�ɡ�҈�eu�LQ�ӽ���H�g���*I��u��O"Tʷx�H�M���Y�5��a����6�=qp�tZ�˷�~룏`M7��˛#��K�w�5}��C�n2A*,<5c<j���[d
�F	Y��&�w�x�,�틓��P*!�0_I��g�v^Ioz�K�e�.6����dA�d3K��/�u�H�r&P���agêU?�v��".�0k�H�(cnR�_�B9}�F��g�p�,�=@��'�)A?�:����@�+���r�̎��|_1<����딏�x�(�K�]OWD"�Y�N�G�0�פ�"�m���S"�E;�m��ؽ�}N1hw��|� ! ��s���/݆9*�����䑽^��D����1���(���ǫ����x�I>MK�UAin��қ�$�ޥx�������G�c����;ȓx1κKhA�%.��qw��$t��+1^�:R���*�_6.����̪����~��X\ �ky?�w�G��8K}H�	Ü&�X�k"B>�ʖ(n����h�8�=E4��sy|��w\�W���w�k�p�����4�	�A)�cu�hk�|nG
0�����w���v羵��s�� Bm���m	��v�.U#{>&�jy�PJ�:�t�/�����.�f8Y>��4�}����.����ww`�k;�����JQ��t��<,�x���{(L���L�9��<�A��w����5:��F�b�%glI�4�t�Y��~-ޏ������eL;J�����ڷ��a����tTY/��`-��<�R�W�8������u���r��£��D��z-D�@�y����U�5Z�P��T�u�����WL�VF���ad�e�O��pF�+��xm�}�3y0Nl�j������b�RǷ�5(г�^@� ���VW��R
�.�,y����8m�����I�?*tz<NhL��qf�8eO}%)2��A��:�Ci]u������ȫ� r�$Kkr���E��l����k�J��\d��e�k	���{i�����!ݫ����U�y(S�&ԀB��+(\��َ�_���g����Q�a~�S��⽬�x5"�|&�y�&d�T�ot��	(��O���v��0~���N��]%F]�5��:?g!���\�� 2��)lP�Z��
���x�����8q�.qd��~��f�I��� ��29��B��?y��s�ic��ߤAw� \��pU��7��ˑ(.�^������\����KS��S�K��We�D�f����n���x���x`m�wv��Bk���So�(����D��� ��I�ep}+�Ir�(C�)��.�� ����xM"1��ю���6��wb��vؒ��9B4�O(o��E���ͧ�,�ޔ� �Jp�ȳp��{�9�(�c��_�������_�V�XB-�#�:��E� �)T�FU{H�\�3	W깄�H�g�:�eT��{��`b�i���i?q(}�����X�̊��2'U
*�k����Ra��'�V�~,Yu୦N��r�q���욙򔯩����[:,�)&����}����4J�H������s�E�" �4��m�A��?��pf��*�QF@gZlW�B\�|}���ܪ'O�Zu�X�,O�@�oa�w<&8�������=�'�fa@�-�t>��i��bb/�`����%Y�K��$#�d�����CUs�r��J"�i�0���5�ކB&��ޑ���tLi�EŠ��t�S���H�v*�~/�DG>�V:�$�N�Ua	�_���<�6�˶�d�F�ѓO�]�l�~a�t^�NM�=;�><T�w�v�ۤ%X!7q�ݹ3]��.GZ���O�:
Js��Pc�Jܦ�$]Y�4T������{�6r�h�~<�A�Q��5�'UH��T�C>)>�q���(w��~���
�����`��k�ƸT�{��pa;%��;�:2��М6����s]������N������M���Cj5HԌu��6���mJ	b�-F6�Z`d�x.���������~�:W�ke0�A��&���*?��g5f�Zv:�%�OY�Z�i���p�u�L)�����p%½N�N�r�.�����f�L�݃F���&�T�x�E�o��,��*C�N{,!q�j�P	emA��6'ɹnN�L��^����l�[Rt��m�ڔњ�����c�Ȁ,�#޳�W�gr����b�qMlZ+�DU4SO�\���
�\�}�Fܦ%{�~G��+!�!f�q~�E��^�vYc�dL~�Mq����1$�V�-��ӆ6ə�@[f�;�~S�^��9ZO]�Q�/��\���	���6H�����x�e�;�@ʥ��H����} �''
��Z�ߢ�+�h���e�kQCQ�M��k{t����C�x�Gw�
�t����-���ʪ�<-TS��k�D���ۚ�P�2͐Ќ�P��1�Kg"$$[�P_om�]��+���Hsx����������x\,��յ��'�����������f4,Sމ��u���0�<䫝P�<����t�����s��u�9p�_�O���b' R;���7 ����T��n�F�wH_MnY����'\����e,a�֎p�6v�(��s��N=� wz���� [A4��4j�ə�Sp�ݠ���[!� �=�R���Ưl?�.��5l0�ώ��j�5N}8�I�1��W+�C )�[�14�����xOT=�ēX�������v���U�Q�M��> ���7�n�O��z�B9��q���W��Կڴ���K����r���� a�QđMLt��.�[[LS�a���D�L����,>%N���F#$Q3ٰ�Qn��|�!�3)����A�0w��:[�\XBa����`�H\�բ���C�_�s=�z-��S�#U��`��O	!��,���Ƙ�f�84���(�nݗ�� ����j�e��������9t��ȧgvS�_b��e	1M��k��W�V�44��qLK�gt����?>
fv	Siz�u6���"��޷�h��-��%��}>7�&l4G�u���b
C���n�0Vz��������䵲�������+��9����*t>ON�nάj�M_Ip9�%|ިP�"�L�}�v1�����]`��p�^P�
�Y��� o�D��j��U���A�q�L�g�^�k��_���eԏ��z�"#��12�mr�J� \����Y&?��4���5�5��ٻGl���j�T�;�]`�T��yqWv}��1��QS������8g���2M��f]����t��'PE���ְ��첗UZ-00�_f����nvq��q���#9� ������+�<�Ȧ�\��hL�E�� 1z�G6c��7�!���O����˙Pp��f��b}!�p��D�'����$��_ܐ^߄pk3�{q���¤4K0���X��������eݶA���=]2Z��~�-1�c�;�,t�l"������rL�&q�Џ��WȆ�Cm)���N�
�%��d/�'��#�s��b$4VkC
��i�(ג�]�t���tݞѮ����1Ih� Q��>�61l�����y!�E:�vGcn����r1a�b��u?-dt��܅{=uӱT����B�q(}\��q� ��2<ߢy���KGW�!�2�����K�Ą�� ��Kk�X�F�V�|��&�����9� >�z�I1�٪�	� �]�^+t#p���֣wG\�am޳��󪽻��tS�)7�Q��r`oW��%��,�mT��}�k4���G�#��]��̵J-�(��+�����n'��`HV�>
PDƍ�D�q5�d�0�LN�s�d)�$%��$�����(�`�=�S^hنl�ڤ����k]�-�5~��"&{qY��8=��"���W���poi�p�8��Hlis��*�����'�n?gu��8A"�]�'a�^<\^{ �c�-�"�IK�*=�F����4�CB�\���5��1v�/X'�p�b���v~b
 pm��X��KJ��oԶ��Dlu��خd�s*a�_C����˳�͈m�l�.�ĥ�F�}�E��-.4U�6�av�Wh�v�'Y1Yë���8���C�;!Gu�Q��;�+a���X�E������V��s��ǯ��8�xS���U�@�9ԺbE�� "�8��-������|N1�P�t�X���e[���{=�l�u|���/� T�( J�	�����-�t�h��T�p�q%n$�c��m%��\ZǊ9<�o7��Qn�i�w���X5�*��7�Ҳ�a(��mxl�~��J�n�A�3�Y�{�.y��҉p�+��J���t�nF�ZBP��w�#��PXZ�A;���Q�'L�N�Ʒ�؆�w���6}d�	��y�(b��ȡe ���fɧ�F�`�q�q�`�N��H�U�eN�}�ߠ7���_zEMJ[E��Z۲�[P�Qa�Aa��L5ӛN3�lvt�Q�_��QU�<X���/��[LLh6l}��+"�L��14��� ��zz�W\�<z3�� ֻ�l�-1"���]���u�>쒒\�:[��;c���'&g�T��X��47�E�;Q��ɋu�ƞQVI�XY7;�l���)(����^ڝ?>P�Rt,��{m�Lq�^�{�(�#d���ȅaٲz�u��/30��`�*�u1�qd��Kt�%���t���z��P�z�p�8��Y��6����Jpn������S���:����h2IK�;��,��C�R����#YϭU@Dm��P��'���L���ʫ����o+V\���>�%F��
�3�.R_hx>
9'��0�0����y/����q*b%(���²���ڍ
�FB;K��F����#���w/��p����I�ѻU<��"�%"G�$`����.�,shw���[�>s�{�M�$hݮ��0*������5|y8r=�
���e��ظp+,o�qu����[�x�ҡ�����j�1ۖeSq�E�1՗`�m,��c�;�, .�-�9�
V��f�3��s��A�zo����^B. 򹥭���ZZC 8�qf�רI�U�� ����5�/;A}4y�*��AU6�0��� &զuYUh�,Č��h�����UC^Q3W�j��Ӡ@�3�I��AY���	������3X�=�؟Y���1Sm�v����1l��*>q�HE�F~Y�C�NT�7@�)�7w� oy�e�v�w∋ 1��5e��uV�S���y�S��"�a���Ø�o�zV|Gh.��w0�e�*+^�^�#�xiE��3��#1r���J�]���T�����o�{~���4���@�{ا�Õ�C� �l�  gf���bm����O�ƣ^#L-gЪ�eeXA����h��O��\��2~ ��(b��3���`J�� β:D���e��� ���ΫB���Ó�Za��8!.te�S�	�起V�͊�%���3j�F�~�zƵ�~�z)r��*��`|�^��ͷi�4%�
s�X�J=�l�׵D�_�Am���=��]6?�.z��B���zI��\�OߝS��[���TKlS��4B�R���<�(�s�=,T"ؘ�g=� ��h��q��}����S��ݺʟ5�s���T
�9tރ��������f}��J�]�6���&��k,���F�(H�P�0>3�gSJ�j�ݷ=/���
���6b�g�:`���b��J��)',���_��]�z�����D�O��r��veKץ�-��19�0�����<:�6�.�IC����������-�:�Q����d�{K���0�R�}�PkF��*�)�L��\.��J��cVe���I�c?�@k����>�HI[E����*��X�Աr��vx������B����ԫ8�U��]�3��J���ܓ/*�?!8ƫ��0��"wx��`=�^fea���u���=[`���k(o�2�&J8�_6�-'<���)XxKO���w2�-���Sd�)�Lޱ�^^��u�j�Y�a����r�Cr]Pj0u����%NG		J�5�7��D0�ʩkvU�� `U#�3�0���X���l���
FbC�vP%I��G���z��n�H��� �kѴrىg)�_H�A���}��Zv�?��P�傩e�/���ˇ��70�@��A����/���D@,� ���Y��/��P�Ċ)􀄈�����T�[%o��!��cθ�W�/_��O��)�ئ�^(�?��q����Z?-L��rؽ��Z��j��d�@����c�+�#�Íe#'�q��5w�qJ��%ᢦ<�Q����s~*�%�d�^gs���o��هa!�B�Q��3��б{�2#`��N���	��v��ݛ�L�[-�Ǉ,pW��<½���w�7o��������%�������jL��l5�������b%��7�Ҿ�H���P
!0@�4Lw�8�#��|���з}/%{l����ZL���/*͢�&ב�24��z �o����jַ?��iUB�fF��/�T����ڻ�|��u�b��M���vA�$q�+�g�u�P��}�كנ-������sU��ߋ��.�U�Ň��̬v! uڛp�A z�L�G1�n�(R�Ċ6��F_f-�:��ӣ)uCeQ$��P@�%��X*�t����u�O�;I��j�S�)6���}R8'�������W-f���q�2�C���1�o�>@��ږ鮯��}����u���,>΂O����^R<�q�5�t1(/<i1Q�}q�nз. ��b���vU��H��q��[��d��q60䒆�F)�%*��(�G��L��х����O�8��X�c? &43@��(��.V�:G�3�YZ��"����sڴu���]J줃s����1Or8!�5�o*�F�Uy\�=�)�!R�m�6|na~���i�f�Y��^�7b���Fg��箁!�����h�=��7;��b˩�S�@ 1NwD�a @�������JPH��ۇ�+eړ���U8�����2GĴA�:���?L[DG�is�䍊���4a�hD�_Ѐ�>�e�>��:�kʍ�m��Q�����K�	��f6*W����������tH��X�G^�����-��xOV�{T���X��l}���5�}o��	������J|M����jd/>C�J���H��O���4CI%d9�X�#��W����+B�{��m���b���]�q�%^y���E
g�0E:ő�U�́7��V�P�-�ǎ���ʨ����I�[F*3�v܅7��U[�[���-����o�l��?<�t���|�7?��y�_�
i��
�L(_ot�6���>'F\{�ó�:�=*��J��U�v̒������V��L �+ @0	��3��&Ҝ��e�4nB��g�&�x�O!)��@��o��MX�9~-r̼�^�g��v}n|�f����}^-%��"DV[w��g��97�>%f�ӳr�-��Xh_-07ND�B߇m���������"_xIi��j0��M\��q�::E���^��F�9�I<Y���o���KTa3Q둶�;�io����k4� ��c�-�����2� ���������/��y�U��)��������r�Ue9���X��+(�iq�QGA49�����&��v{Џ�c>�+�t�_q%l���E�u�(]j������->*j:I����϶��cE!6��Iӭ�<՗[҇�M78Ood־�kw!�eP=79�<�zsn�ΝC�h��Xp֐k{(��_����Ai����ͱ�,y�Ė�eF&Y�UE :.Asq���Q'�?����-��|�L���b/H�܌��i��#{��'�R�il���*'���z���PisB߯�P<u�y���=��pj�S����4�n�������ٿ2�����*�.��f��m��i�I��m/~LM`C%BWŨs]�~��_�`:-�fl��Pu��w��DL�;I��Ka����_t|�v�pȕ��+丂l��[�y� �R()2�l�c��=�M\��V�=ӼCfP`��O)&X� ,.j����b��i��1K�[n�7�VC_;���yMX'�_@�qsZ0v��`tK�:���(�2V@C-L���r�FK+U�]�D�� �����k���8�4�Ӡ0U*�{V,��L6�m���fƲ��%�֟�E��r��x�ZĆ�z{�'|���N��ڼgzc�n��֬d ���1�k\bzL����~ޗ)k���6�*��6 G嵑�D_�fs{�TZC��� ���>-�	�����g	5Z.:ˠ>�6{�g3o�H�^9ж�ϴ�W�ՋI:�,�P|S�k�֗��Yd��(ߨ����
�w߳X\�KL�)�"���)���&��7�@�rFs�-����65�ٙ�ok/w�}���i��8݈���_�9�Z����?^�˙	Љm������'� ei���U7�R�����ߏ�%Q�T�r3��5��SL���������skh.�ޕ�i��k�F"�ϿkLF�;)P�Em��W||{c��
�jyyQ���p��S�3q:'��{�<���n�%�fl!z���Q=�XZ��IY��Zj4��fr���a ���r0}�MV���׊���m_Β���`��z\���N"O*{����E�t�Q��tR:ls�����so�B�( ���V�%�y��@��E��AR�umn#����a#)�U2�F�y�����%�~�eV[�#ٲId�6c[�5U�4JZǖ����9a,����A9����X����G����֍X l�����~0�f�Na)RQ�FL!闖�]�S¢},�`��A0��1+s֠�B�l*�;	"�"
���[C댆-^�fM��xkWmBnSxD5��� m%��:��[l /Gj��+B�t��]���#4��
t�&[�ǧͣ�6�c}�g9�$��|��7�iɷ\�u��=�hf'�B�p$mxEԳ��;aN�U�c�X�����Q��fE��4hr��8�C:gm����� ��<�hd�j����M�(9c�1t鬑�r�q"���Q9� �s>]X����q�]U��x�-�k���گ�|�'�z�߲r�rX5)6`b)�Y�?1t�O�fS`������Gc��C�cr���Y� ��>���;
��ĵ�yxJ�Vc�3��Pj*xL���y'����ȑA�������$��C%�e�(9�YY��xW������PS��Cc�\��۹�wu��$���ZC�k%�+����fTq�K�F�S�n�ך�!�C�8&$�wMB���߉Rr(^U���7e������U�X�ń��2(�J�����%�3_8��VzK�7�Nt:P2Fɺ�H�_(�<�*_�B�	���>A�t�7:3W���S��x��O�',�^vf�$DM>*�%��.y���f��$�n4n��o�|.�RoEckz�8�M�T�Ea<�< sq$/�� {��@�����0<��H��XNoj�-���U�`��2�Ē�#� �^P�J��!�
!�h���g�B��&c{�}л�WHr��3[���7)F�P���֜2bD��Mj����Y���O����|�K�i�1��v����e��L��D�� ��y�Z�f�D^��q+�$�������↹��H���/*�<���L�WE�����Sw_;��heU\_������H�z�OE+��|�E�*��ܵ ���#N����{V�QWC���Du+ݚ)�#�$�l�:4��1�s��$�A���ŭ�0m��K,q�6��8��I�Є�N�NŪ���������0pT����8���`H&��q��ֶ8��|��	2`m	U�R�|�:%@����w7DuY��( y�W���P53e^��D)h5��wy4QWA�`ݞ��
��oB,�=��gj�0�Ȳ
�E1�(�È�G3ܷ�,!@�,��Y&��OF��ew$�7�@���~"yR��_����&e�zjc��p$�+��v| ���wE��u�)�3>�p86KQ(���dh��Kr;�;5�Ǵ:�GC�iT]U�&Q�Ԛ!LܗB?��ؽ�uE���)a�z������]��[	��C�X�H�5�ތ����T#?-.���lD�����B��ޒɷA����q9Ȥ���8���wbS�}�V��ƣ�	�� ��Tg�b'$�h���Љ�%u\�`�̀f9����a�`�J|d���5O巛e�O��y�2�'���\�.E`Q�#��Z%I=�fP���_sE=�����m���ȰڜE��K޷ȫ�f�4ʰ-�~H�_�e���W�k�;/���X+>��"��@��~�6�A��[���,��l���)��|���~͂>�z�F�8���|t;$�s�=�Ƴ�'��I��:�;FB0Er>�k��~��P�GZ��gl�QM$A+� ���3�F�'H$�%��[5���)ߨ���2h&���O7"�اž,��SU�������*�k�@`����01�pFK���o�-�T!*�����-��Q�uu���1Wj�U�Ƒǜ��򇿓.�5���.-�@�5��Ǝ%���T�q8A���z�]H�6��WÐQw��
ʯ{����X�%������R���R!��e�}7ޓ��1F��$�a�1ǅ���Bb�V��r��-H��і�C	fbA^��&2B_��-��)��䇦��#x��G�?���߲H7FCla�-�,ŗ�ϕ������t��Y�&c]L�d<gSk3n�7d98#�s�8k0\8QQ�M�Q�bG��S]�}�&��9��+�����{*����W����מ_��We�GWՈ�=�}%)v�-�esc�l0��f3D50���x� ��7 ��-���C<��)c�V�'�&�����]���0*Ў��̓�U��tR� ��iq�����
��S\(�)i��ٹ����ؼ��ed!@~+N��4�*[%jVѩE^*��耲�ަ�w��N�m�]����T�.f��v%��^�����6 x������._�4HQ�����G�:O�B�`�N��x	�8Ⱥ�i�JW#��ɻ��5��V��D��&9? 7�;��<��Xn�}���_zD�2�B⺤I��J5��u\�)nћ%��U���n9��ԻcwL�-��J(��'ĔTv�yΎ$�<+�-��W�	���S]��u��t���R�3|��{�#Q����_��:N��ۇ�&$p����;���釶=�?��X�+�L4�k7pާ`é����e�R�����9lK4��ot�4v�OXs�]5JZ.����)k��ʹ������=͘rR�;����@�.�q���m�N#��M�p�ېu<9�!��7.Eo�i��p}�5����퇦/�\d|�=�����8<��H�	i��*orud-�p�����l�u�i��
������F�0%Z�ݧ��V��ܛ��J#k�9�"���um<vdE�Ӻ�0ߴ^x�t�z��z�ݰ���u?��-6)@�|��&�K8%�ɲ�ɛ��c|6)<��L��E�/����%h۬�b�#�o����-��./�Dz���SY�ߔ ot�Q����q���h��G*�HC\rg�9O<4� #��o�B����a����o�VI]$����)��M�7�$�O���ƨ3��俒}B!�M+�R��L�����J\�K����&^&��F�)�'G1��ѡ�[��"ò���:e��w^����`)��Ŗq����~L�,)����%QUnoF�B��c��J�*p7�m�V��Ab�7�p�\Kؤ��>���d�2�M���M��������48��:Sw.�Z��ZӉ���)�B3��V8���9�%�o�R��[7ԕ.
3X��Ϣ�̵�qg.j�)L��� ���։R�so�%`��a��Jm[b3[��V�����\U�r�1|k�;7��o�Gn��,��6c�p��o��J�m��IW؆~��� ��D���܎,���D4��k3��p ��B[�RJ�������>ka�疌�"��|j*L���JAAY!�n�9��"ཱSJl�$�c.��G2��Pʀ�b()�@�'�컁�-�!����(����O���R��,?��\�8�:v�H��(2�I����y0>[�����6b�+�Ej��d/W"_\<�6.�v����)>j"�d���a,n�{��}f��1��n������䈮j���/�V�U3$���;�h W�.}�!�0��]d)�+��Y_��TiNo"o���y�� �z/`�^��m�U����;�i��I�W_�Y���6�z�U.)X^��d�c�hH�n;��¨�f���d��!�RRL|�ix���v
����(�+�w���7��
1-/�^z�m�Oظ���t��V2aM�%Q�uڃ�p5�J�W�]$Os#G-�>���I�d��T�/JV�Ƃ�B�B��L�����-Y��<�w?I�5��5 C�v����̙��� y 8?�<f߈����#T���^��.�>T����*�};P�pŊ#���_ ��s������G	A�{�Z5��R �6�Qw�A�{+,�����{�D"?*��݋+	5�>(Yl翁/K��~F���x:�گKzx��]�~ng)�1��-|����T�UrdM���K3Z���\t�h���[(�qY��]��A:ɴٔ���������n�d�"Tb�F'�D��s���J@^,�@�!����%҇L7��c$1���g�*+�`�Jm�G����'6����b�6�e���#CZ?CN�Uh��K�,�VTY����K<�����*�}\2S��:�y�O���#	1?�ig"���U�g��@��FM.q@��d�e����"�����
����E��X�tz[GaW�Ѕa�X|%	����]���}~��AV����Aշb�j�W ���5�}&�c���[e�#-<rx�/JUŝ��m�m��\*��"���e�8�U�����D��criʷ��/baxW��͊Tw@�x�=B�a	�?��Z�@��b�^�	��#���4 �zz��3�����~�i�	�"��$�V��'����`d�F�f�xZ�HF�.���Hn�_�?��3��	,z���ǎm�~��f �Y�2.J[��|[��q��-(��c��2�%H�fd*�]����÷����iK���ֆ@A.�W|n�ky$���&E��\���}�Q\H�F 7%DH?��^�@���H�9,$�|S�F4�`}�S�9h:5 '�bP�Å��wT$�<�eC'kA�T
�J0�&���<:@�7�;s���#�Cک�(l��$ �*�����'s��OTJ/��𾑛d�����qx�N��� t�l|G3���j����I�c���3b���3�.4�ki�U�C@�@M�?��5�2�%.�,�g��V-����MΌl�5#2�.��T��*���m�Sɘ��$�<IX�B�e�B *"�����-���Y�
m���(�N���/~!��R�h��(7�_\V;��'�2R�����N��Pa3y/����@��/lgӲ�`���x0����gƮc|ўЇ�#��`����<;Y\Q~�t!���Fm;�(��"(�BG>�[T�+��ŌD80���������ǽ�gi�����$����S
]Xp5�	��O���=R�����X�~+O8�����
��ߏ5�^����aJ���Z�{�mIC��<�J�R.��$����W>���c[bJ����B�<S'J��t�B���LlPIYD:����O^^�MG�8ዟ�����ܤwg{�?3����F���d������0����cD۫�&X�ݔq �nK`+뻀	�Qf���Sfu��Lc���N�����`��5_<�9`��L��b7=��K9���+[Y��s�F��i�\��;�W��_d3)�I�\�̆����|��!^Cr��>�K��F��چы?f�b"L�X��t#���-�"���-oJ�Y��Z���ߑ��ʏ_	L(
jF�bN�!�~I�o9��GL��Y�\�����p�"��z!'��!��:��m[0�eXG/y��p��a1D9��e�IH���'B�ͨ��`-�`��8`�8/�23�q;���8�ச�I�WL�;�
��E���0�q.!�#�A�����lcN�VR�F�#�=8{������1��u��[��:l�i���Ź�B�jY��n�|<A��L3�o�����e��'<��m�h�� ���^�Juo��2)�K|��铜��f�p�g%�Դң�-�2����!���{n����z?o��y��ϐ%�������<g�A�������+>�Ø���Z#7�u�R����?�N�O+ �l��� W�e�4��"C���r{�lkP��$�*�������oȫ/~��26`áPn��`�rK�p��"��|��)tt�*_�殍5*=|._�аw��ώ���˻�qu��{��u��e���Y�ۗ��}�H�~��6x��i�����c�rS�/y��o�:��%�D�>���x#��l¥2���\�k�`��j�F�����@J�`-�a�[�������L�ʻ�b�JDπeh�7P̘7�pq~3S�l�=^љ�/h��*B�ͻ���o\����"�ej�w�O��P�^�� �����M��IպTZM��R��G���V?�v2���o,+v>��g�op���ȬV�d�꩷����gF`!*����AW�ȇ/�ʻ#S?��M��_�ߞ�)\mΆ�(W��5ؠ�=\��$'K�#*v�d<�������G�j�C6��/)\��A�w�]�yD���(�)&�����)>Ԕ�u��vm�R�b�����&,�Ko��2�(B?�.7i bjA����� ](p2�D8-~�����y�]SP�g�@��1�^#�_�2Ñ�&��X)���5o;f�t�ù��?k����C��n�>$�9 �}6����(1j�<ڪi"Ց��?=��o�h�/���5Og �)��mP4f�vC�lj�������Ç�k�ȕ�"�TNA����K^��&c���:�<��!������s|�z�fvn�DNO׎"W�\�0�A�������_z$�Z���Æ�{L�SO"��0��H9�}�X���߮����ERK{C5po��T��v��~K���V�����?�ړ�O���a9����	����[w����ǯWY5IY�z����딻�͗J�.H3�{�!���:��0ݙ�0��*I� �S%�K�떁)��`_̔G��|�C�?�n�%��ՂO���.��R��q��|-��ua~�H1#�=cS=7#:��-:""/��a_J��m��kOl(;���\�:��:�}ػ�%��ɓ��1I���4Xv�B�}�]��f��]|��HpEa����Q��$��ڑY��3@�O
�v�eN:��ؤ�/r��2ܲE<���NI��;�hL�j �)�g����"w���,�3�j�d��Y�$#NP��F��������]>�.M��Bۯ��$��(6�����2Մ�0
y�����['r�||`����t�U$�y�¤��5w��"Ek��������+��_58t�U��\��6��O�(8`P],}x_l�~��㓲n�'���-�1~��5{��>��+��𐮂ޕ�k�cB��� ���q��(���-o[FB��wE��I��~%x�� 	ɁJ��Ş��lYLrQu�AY�ܶ�L�d��0�#�&ѧD����O��i#�a�M;���:�P�mG������	�R/�<&G��9o�zpŏÄsdk*����Ȭ\�*����zW����I�Ao��1,&*�;~%l�>d/�p�uLm�u$��`l���I+r,�����@�g���.xO�K�݇.���$�D�����X�Ӹ���1i�|#��[�!�}�L�ģ�.�~��1)/f�E�E��#��=�e���S�'i���&5ڄN�B�����v�߃n���Q]p?ʹ��fw*9�o�ݲ��3}��SN�\��!����*T�5@䛟!�n���L'� � �_�׬�;�61v7�h	�V��M'٧�@����L��)�o7k~.�e� *[��x�O��S��`j���!rw8����oͥQ�k��o.�9�N���.nm"�~��&Χ�N!D ���h��;M��,W)K� ��2�֊L��ԦV��C� hC�i�7Y��2u������O�md!�d��qҪH�Է������%�6f|l����j�tք��u�.Kh���s���3�t������o��@�	��R�P����@�n�ĤwCUɡm�/JV	P����Ƥ�&g��-��͈����=�Д[}�hla�wq�wWc0mi����
C����XU��-�i���f��˄��,5�CVId�~Y���c �l�_�����87��ݶW�z�����a9����@@�ޝLjN ���/l|-g�j�,�	:CQ�JL�r����p	~�#�,�\��tY���Fk�D�A���2ٴ�����O�8rZ�܋T¢kp,&��4/ i�Ɋ��"��s䙃�G�h� 2�>��Ą�xY���pf��`�sȗ�j	�2n-�x\Sg�Ea�7$�r1��V�:����q��$�����w*8W�W�u��yOO��%R7��K���z��qϔ~_���"pc�e�bO��~M���050c��GW���E��`N�VuN��d�1��	r��`I u���<>)��kb~-�������F�Q��p���<b�n!��IC,"0�v�s1`y�%9_�H��k��ЌyڕD�B��I���b@�0&�k�m!=��6Z�"�)SE-:yC��'�`� B ����Yx�.�!�lu�r�)�j��C���*�����������@҅v*d��ծ�&#�Gt�-Ȑ6{�kF�#��=f���m���c�F�|B�8;��cW=ј�ꑂ`���@�(�������v2a�#V}�Z�L@1	р}�\�)���������H-?�{A���ip~w85�?��\��n����у3V� ދ� ��K��9H9^��J�E�ݛ^$+M�T�iW�F�$g�"4��C���ɸ$P{���CzC�OM1>�/���>DT�ҫoK���w�O�΍���	(�EM<�A����E�a�Y	���ً\y}�bK���vt-�,3^��an�IZ���{GD���<�rq�j<#P+��J��$�ʫ�=��iN�>oR�d;\�5�3�	��U��૲��� q[/�,���oL��GP*���}���I�<��z+�%��X�
V}?�d��=9f~
�����V�
�G�랼�)���py������B+�9x�pj#���T�;_�q���9�8�C2���ֈV�%�e٩ Q̟�]�/F���G�����q�[����/�R�@�ZJ�Q��pA��Z�apD=���y^�ྈ�����,��3����7����+�n��=���:DJ3��݁cĒa�˼D�����3���Uh�)@�0܈��yta�<݄�f3��o@h@���p�q��r��o3��L&��y>�E!r=Jx�Mfv�8����:B�K��O:���!C~4g2�`�K�xN��S�3C~��	�@��V��ynl�Ӵ�0��7崦�Z��?�*\ �I2ި/pM�+��?;�����H{<��h��_�M[X�V�@&���V�f��Z,�o[��9�d�x�����y��x��ٽ~�
v��q�ʯ��k��<T������zc�N)��T�l�":�/��>}]�M͓y�hU��ʢ�^K���2�è��l����ܪIH�8!�����|@�v�r���)���y�p.�K��h�;�)*u!(��8b�ɹt�G�,�5��+���#��Ώ}Do��).IGRQE��Plj�e8�A��Η����/˸�h�Z넆(�aX>-��X�\j�}LF����^DIӼ/ѢK� ?!����H}Nh�>�i(�s+T8.����H�k�J�ӡzZŜG�=Z,�+�K+z������?��sZ�#[E�̗�-�#��n!k�n�t�c1h]w2�b
�iu*h�HX8�td$E�^��	��#��ʼFoy7�8H��Jn�̜��R�GmA,͓R�y|����(���CЛ]���
��)�V��ҼϽ! ��5ņw�@�4�]����<��?
����U��N�(��)T�M�B��� #����ǝ�`|�	���e2|����
����d�5)B3�����wˠk+ơ)���"f�']Fl�<��T�
�d_�W6ڣ���6��$��Z
b�Z���:Ty��F�������V�ފn�t���K��QAkf�x^c�)+�h^���܃�G���_pіci����[/�t=����;!�&/:�Hmd����#2#��R�4I��Y�C�Y#��#�[��A�#��+�ED�w��u���F�8���筽,�Wϗ����q�}w+駐��)���^��\������T���˫��S.|3̰����V��C�;�����f��(��W���� �D�n@���˭8}�-�?c'�_jZ"���µثTݜ6��? >���-�t�^5�`����p�(�974�=%�N`�K'ΑA�P���>�E�B&8\�>3pJKyg���C����3��}���l,�X[&n�g�-d���0d$�
E��Oғ���=j,<��;�=��~�%���d�>1���c�U��B����r�N�������aRۇ]Ocv��w�}�[�]F�Y2��Ɠ9L�po�V�e�J��Jf��};],`M�(��v�*/�0V!.r!� �Ki9d�\k���������A�*�L4��H�WPD¼��j�B�2Уfi W�bIN��uم/�ݫ�&�d�e5"��JdT^�5��I�/39~ŗ�0�Ͼ��"Z��ղ�M�p��������{��+9�χC��_\2���P�� Ͼ�[�M����~����F�P�h�â��������{�ކ6�a��\�_������:��s$E)����O���S#�1�|VfMz�|���N�Fsŋ��܏���p��Q��E1PǗ\�$|Qn��Oi0]�j��G��P�8E'��ݹn����	e�T|�������� 7gAM}���%[���/NQ�͏D=��w�.zcCCַtnt,tD��z���-�F% �sH��D��tY�+>���THr�M�بs����궲ɏ�u*�v��$��z�DJVy���hy�%��$���\y�[X�J��n�½q�;&Z;����x�XF	N}��%�L3H��S�J���1���-h%kxx�ޤ�����U.�7^��a]ڈ�h��c������Bg�Gf��=qt����QSe,�nrN7�׏�e�(�"� oC���ߞ���~�	��!�p�l�u7�uk8gk����c}�S�s�x ���w�YcX��E��W��PӶ[���3̇���"�?��Hs�@E����u�d�*����&�8>(��|�9�D�)�O=kb�L��❩�S^�r���2%N�ZD�AhG��M��(z?)��Q�D%-����#��<��J9�X2���Z'.��|�_��P-���X����� �Up�>���D	o�8��ez;��7_+%��q7�΋�B<��F)�^q�V�	�&�M8����ߥdl�s�	Q�?5xL�Bq��w��L�fƒ���Nw�Gl�����"�Gҥ�c{f�A�y�XyeH�0�~-?�aNE�j�3Ϫ�`�'oCO�}+Vx�_-�fN��V0��0:�0��x?���Ʋ"lt"��iE�~gVH���MEB�2���*�k0��/��-�j'#�g�Ƌ8��t�|ѩ�c��(���O��,-��4& ʹ��i'�u�J�1�fy��J�F���ڽALj�0#�(���f��Y����3N�֚��tѩҞ��>���L���┈u�a���4�����9����0%��� c�m����Fˤi�eCE�Ĵh��q���R�g^i⿍���x��`Ir�tA�<�p*D_F~9�S��,�x�@%c�Kӄ�^:<�[4`�]�2ra�o����T���5$��?2o�2��4�O��W�H E!k�C��U�ˣ��r�������u	6m����G��O}�P�hc���v 1��a]�ߍ�X��3�]��=�A�ȇ-Z@������)�8��A��XE�qM4�gb���A|��F�ڷ��ί�S��Yu�z��k##�b�Wy)�9��ܣC]��k�y[/O��:"4�wn�jRo��-�b����:���_��u�o�*�|ggiC��w��)�\9��ڮ��!���b����>����tUK����jq��~��`�nu=�