��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\����q�?��e�I8�b�Ǽ$��"����ׯ1�V0�����#��+�3�Xh�X��ȳ�k���(d�gƀ$��ǯ���'��+��,ھ��+���\�5أ�7VE��4�6��æ���IX��U�o�/�lH�f��Y�J�➍z06b�Fee>X����)��]lG����gvRtF/n�z�Y�4 �ư2zuQƤW'�*ֻ�d
g�nd�/�h3&x0�B4Ƿ`Tc��o��R ��;���B5��x��p����n���Q��U����bo� `�|���sb6C@n=��me�KN~Ҍq�e(�䬡�Q�����{v���z]J� g
[���c���e�վv�s�v_g&VAT�0
%"�p�D�~KVӻ=�,H�B_�Z��x��b0������/���8eF�6�n���D�*k_��3/@��D@����dp�ʻ?O:�i�PZᖏ�$fu0��&���,[����0�V`B~�ѸM.PE�mq�^�{����[b��=���#U�[�fLv�����"�1�EE퉆�g����^{�H��	1�ET�Y�� ǳTeg�Z{�l�:&_�#,��.�ߟ��Z,�m��=Qj(dШ��o��`BZ 1:Y�T5�١0�9�P��!�q����,ǐЎ+����3�&h�2r�wP�͠w��S5*���`- A�vSD�d4U>ݘ+�z� {vb��W��y,���R����֫�������6�'XG�H�ÛC�����dȻLV$MLr�N\��5ND
*Ux^�Nn͝���ę,��y�BG˕7xk�7��LR�c�ږwk,i�@�;����ǓT�fP��	T�"�ꉓ��? I�ҍ�\�׺D�X$��X�ʵZ���H���m�4XJ�x��c��6x����-��2���FC.��-=n~_ѐ��Z�"`�]��[gh'�1��U��s�a�f"}�+�%�h��m2j5�kp=<̼�v�;�vUȁQ5�C��UyP�
g��?R5�:�O�i}�b,�Oʹ�CkW���p�h��V��R�2���P�Gc�o[�]3ӣ_�K�2�m?�_2�<��Ō2xu�9{���db�
#���zfշ�^�T��O���$��~1�.�� ��i�{���0��HJ���o�ű�����'�^�hכِXiϾ+��F�!����[�Co��q�P�i%�������c/0C�m�x}�ɟ�nà�G{�<�f��ϼ��P���&��WP�ѧ��Q��M�A����G+�o�~��	TK�c�j�+Dy������f]Y��tR��r#>�]�ڰ�`/7��c�L��	|��L�z��kv����q���v��Q[Msn��2�A{N��/���׃.��` ��ʳ,Z�ڇi�D�N��=z�
�$
 �g3k1{<Eฏu�G��p���:L����G>�1��!Z���j�拊��e:�B�Z�Um�YP�r'K+����O�OxJj�Dg��QM<�nCyN�>��S>]�t}߸�e1�����!���~ȕe�Nq�4�2hy��N���.����v���|ށ�/uDB��û>��z�%rly�$��G{:��$`�jLZ��}z�E�?�I��C z��7X~ю�/�yd��B��d���L��}>�&4��O8ua��k�~K	r�>�ԧ���=]'��l��^��r3�Lމ]g85�/o�=�%"�t�g�����΁� &z��-�W*[0X$]���N}귭�:&���"RM��ڷ�6?-���3saH�p:ӵvǚ@nA"o[?^�����U(�*`|H��ld�y5�!"T�%����Ưg���LS"HK�^_r�e7�3	�������}�|����k�Q��w�"ɗ*����5|W)�7�m����G��;町��J5Y��1��-A�}C�:��A	�L��?f� �h m���E]�W�������5�7�lSv���i.Gh~5x�G[Z���?5?8#֡�؝���M�,Ʉ�r�cp3���]2<<��a18MA��ɧN�[�p��vW�7�1m��=����Ʊjq"�����[s1�v��{[�����<dl�_�MLwj��$r<o��rN��:2�S8H@?oS[�zD��G��op_Y7���T8�x���)d:����,��#	�!Fea���_jo+\����Y]��ܢk� ��>#=9(G��a��g7+*�h�A�o�b�M���)f�O�Q��|*k�cr����܊�'�{��~�Ù�R9Ueb?�mhhs��Y@V)c���#wOj����9T��5��@�xL�7rH7]����o ���̈PE��tw��1NX+w��h_ ���ۜ��Q�t��d�����μ�EY`��r$�@ZK^�6G
u����?���`'5�������2E�=�T��:u��I�-�J]�vQq\�AK�O�c	4�(蝐" o�o���A��y��|�} �q_Np������I��Ŧ#�$)8���mP�*/~��W;:/:W����Se=7�~�f:�6vߜ�k��;���O¬a]�s�"�\���MOP�)lCY	�9^���H���g��`�����u2��a<L_F�,�t#dک�??o4�����@ۦB�9�R�3�՜V%���Ğx�2���GE���F:Ϫj��HV0Y�䥐Su�9����STO����ע��}e��I��g��	|����
�����N��]E�rH`��K����-o�%�<,��I����K}��&^2��8�����o$/�����+�s#��VGrF���'���A���ë'i�"7#��	
"�A����[z�g{����^wR���m�~[�5�z.�p��ZmI9>:@>8E)@S�gcϟ��3�����.�A���ӽ���O�y�-�e�c���������A��c�ˋ���Bi���+,�u/�9F\�k���8�L��N�ձ�fH�����{���^��+Ac��l�>J����s�:�[=�P
�����w��K�Ķ�C$V���� ��,�r�I�����,��d�i������5I��y)� �N]�!Cx�?��F l�6񩠄u�����qv���a��Q1�DF�Q��ś��$��O������|n*a���s�I���q+�e��0C?�!}��88`\a��>���VFu�'A\���;�2	�z]�B�TX!���~Q�M9q���J�7�e��Q����r�3H��V���2�X�Y�v��.:C:�Nd;E���X 5��/Q���Y(lBqk�L2y8�I� �⁆�L�@7���� 3X롉�妰�A�}Q�۰>֘5"|DT��=x&�VQ��CvG?b��7�S}��O��k*�����8����9�����r�$�G��	�B�d�����%zy�g��YT\�s� ��d�NSH}{o�]{o\�6+�Q��_���`��c*�ߙɐ91WMt�Me��J:-a�KA�g�����sR��Kڪ����*����+�&T2��P;�oh���wʊ�n C�����w�b��F-H$l)��N�����SE���߃	����u&�'7(�*^�ҤkvZ��8���d�s��V�<���\K�����&:y؃���s�}3�����u�4�#����l�9N;6�3�Uls�|��4I�<<�s��滢�^�%�{���0 d�P��Re�� �er�U#Ǘ�<o���+u���h�J~F��Pv���N��3�������>j��w����>�lx>��C�gk��6o#�|JK�Ͽ"�������۽�]����t��5R�^;s3�ю��b8�Jߢ�of�I̛$������1zv��FoP3k9QC2m?d�5�<g(���|��cG'
��'���)��h����m��գ��1
�r������]�8��3lj�bߛ�
f]��f;��
ᐼBfB�Gm��w��JѨ��I湾�ٺ���F���ýup���p}���1�9ԝ5�+�ӝ^�?�^-�e���wu�yP��t鋆��{�q��#�-���8ˊ�a!�(�?���h`�!i0[R�ݍ�*�9E�iUO�i���1�qՇݒ{}ZWmh������*{g�q{~�ک&�*<#%>��۫��b���x��$��%��*2y���[�g�|����L0����:�s���ܖJ��V��U{'���_=�J5��ܵ��螎�<i�:����r���͠0�@r��x�a��=�Ո$A,��3Kvp��|!<�l�*������zo�/ٿB�$g"4�9G���o���H�[s*i^f⊲���|��2/~��<�s�ϐ�a���Ϋ >'5UCU����+�~��������-!��|g������9��c'�����6�bɭI��3�#t����\��{��^I�mJ��Y�ﺳo*g@1�+���d]� HF���U=|Z�\J�G'"�1�b�����#Fma"q5����	��
��n���f�z1P�%���1e��K���鹃xa�d	Q�/p�GI��5�қ߮τy��;�b��X��XL��d'ŷUV������#�oA>EG�z8���7e͛�#U�B��vTWv�қ;QAl��g�=T�.À�7^ɩ�S(}�0IE��?K�-���U���$����s��T׸�4{k���v7H����k5�%u۷�p�5�A=_k�9�6����$�SG�.�^'L����|-/ֹ�$l΂�|�;nĈ���[��U'%��`���`g�i����< !�'�y0�ϝ`�6|?��#�\u�]�sH�9�;�Xt�㜌۟�Z��U���Q���4'\���l>��	ɈS�3yI�V���۲b���^�ľ:�����g;%&�Љ�7�æ��]=�5��v���ǧU��ͺe�?Ң�s����Y޾9���a2׏�����u��(ѻ1�L�x�fx�����N*�9S_���y6�n�\>���H�$��fD_r�Q��E��M�پ�<+�-��tuo���~��Ħ4����/�[����{�����\l��qP���k���T��{r�kd}��y�$N��4n�ɞ�c`�`a�D�w��Κ� ��JHP����+,F�5�R�ޯ�g�hU�G��Hc��0z[�7�)|�葼�u��D9��8�M�ar`,�Y�u�l�=�q��)�W��3M�VN���3�8g�Ҋ뉒�~��𜺣�	��{kfX�OY
��Ӗ_B1�4�+=���~J��\5��Z�\<x�y6�R�?��@)!B�)"�?����aU4ݔ��
��y�`��B�.��x�6�l4:�+���ɀk�5�N�sn[��^�Fz~��Wˁt���'�i�)�RW�m<t�;6�}{�V��\,&�}� ���U��d���N�%���B�ɩ!��YL엘�$[|Q�A���݊�C��^������:|l{Z~Ҳ)�5�j�Z+���Y5�|R�S����~���ӏs��Dw�'���g\z�L��< �[S�n�V��% �ܬ�Iوil�S:g�Ԛ�$'-&+�V������]~�Tq'��/v]=���
�=l���>�x� 8�/�c%���(�U��3�`@�ך٢R�gvJ���Ɩ�����*�q@�f�JT6����\�ߤ�~�Kn�}�W�!K2�X,���[��ߗ�s+<�ѢK�Z�M(�n�cW��"ډ�Τⴱ��|���?���ˉ����蟹C&�%�چ�W���R��7�� k���~c�׈_��#�H��X}���lM���q9��H w���meI&
�@7!�q|�� ��[U���!���|yS9��rWw��Vh4����=�$9� xR2���0�idB4��-�^��#�%�S-���Ac��4���r/�S�]�l�^����P��=ƛ'�+�)p��'5 �8�k����r"�qj��hC�%��L�>&V�Ԑ,�{7��m���nH~�w	ֆ� "��q�C���h���j	��-`H���\�*�:��.0�L	���zǬ(��!Z!3��ū�`�c��uz���f��Ubj�T�U �+w��2ؘ<8���1��2-'�lj�6[E@�o�	-O��sL�Cs8Ep��FZ��c:9c�#�<*����� �]�U��U��؊ �:O�k;(HO��oM3��?��lH/O�{#^��W@���b�-�g4zRRh�IX�6n��K'�VS+�ɠ��I�G�|�����%LYANjgq:6D=|��!lȱH�����N���������U�������Fu���͕��p�%�Z:zb<��/��L�'����ͩYDanY5�Z�s�>��I�p��+\gՙR)Ე�%� y�^�lȓ��a*��U3,,�\����og�ġ�(�I����R74��PRj/��
hEc�c����k9h�x�\��9�mX~��~��n����I���=�T�vw����hqgF�:��:4c�3�e@��*aG�|���>�FjF��l��ɨ0BO��/�k����3D�y�c���^vV���W-�&�Z��x�����/Y��1���+l��-U�:�����h�(t��Ӭ,�Qs^(kМ�8�Y-vZ?	�d+2� ��\���f~ݜ��O�a��<�3�@v=ƏuХѹƵ⢨�yY��W9:
�<�&6��3o>��|~�������� j�P�ݒ%Сr�m�l�s猱������%�����In,.~.��O�;P�����ou��k߮�y��y3k��7���Z�k ��M�Is�h����C�Y2Ӭ����Æ����p��p^GL��o���
p���9R��G�+@�� �I ��&]֌�}��U�E�X�{k<�6�WX��o���/2P�˨>q�;�b' ��M��>��`�3%?�N��h���LP����������R���VVD�knzn!��G5Jy����D�C8p���}m�ɵZe��� ����������g�'��$��}K��h�+t4xd�_#�oLZ�뤄��W��ٯ��%�q�u��߀{*M��h�>e֧�^��N�����D4D� 	�b��s���d���?��_�p��09�{�`n�}d�Fʕ|<��!#<M9��o��r9hg�W��lA[RlAfM�Ԭ$�?�b5
�����bޘ�W�_�B��k�*��nO�	� ��⊾Q#b�)$�o��barWBp���e��T�T!��5c��z�e��{��ۈ���?�h���s���G�xtr�wzLJ�j��c�)pĶ;������<F��'���!�k�ϊ-�YV���������tϩ~֨�+�H��ƹ�	&�Q����a�]uk���a~?Py�}s�ߣi�S���)`��@p�"9��)��d)j��ڥ-���~���{�W:��H����$�&ݻf�r4�	���s�;�%Ǜ�td���R�ܤ�r��ݩs CStf��ie�����N��]]Ҋ���K��`�U>�d�z��:���։r� P �`�f61S��E�zx�`B#��SY��H�'(�UQ^|9��OM�s�T���d6o瑭����e��.FPܿ[��7k�+m�z9���>�9@�a{DJ8��*>��JC�>�7+/vbN@��/}�d��ώWt?�=�v,Xl' \�؋����fo���e?��ٕ\����.|�V)^�� ����x�\3�� P���հ_>�}�TJ���x8��VD�T	��@r�}�~rUW��\|L��O��H���*�$�t8"!C��zx�Ռ���_\�D���ک���Ծˤ����R�� �Ѿ��"e�(f������F����fT��V��KW��T���0)�W�U�������1���B��ݢ��1;֗-V��"�qs��&��T�RDSU#g��1�l���K�ѭF�S�i�N���V]��f��f#}	W��r4���5����]�"]%�}�DG���W.����(�z�;~d��6[����ln�����)M{�abe\ �J�����=�u�jr� vkI�
�(���SnO�g=��vN��Y(��Up�O�k�JW.��-�����Ĩ�=������������y� ��ſ]��������`"P���U2�[�`'u���TN��C���H��9�V�V��m!�|��D\E�ˢw-{�yͮ��ЩM���P�xo�=���X֔��� 5�.�z�������5����n��$O!	�?4/n���$x@@��юI����1�/Ӫ���P���];A���k�: �ͥ�ʍ#T�)�ؔ��z�
t�=r���a� �ںN�1�;+;J��Z�����nx�{�(�KV��ؠ�?*m*VGw�b
i��{�Ҟc4�c��	��<��H�#e �}�g\�La/��	�0-�����GK"��|`">�45��*֩%����Cs�
��jw�Ji�ཆ˽Q��Qb��V2�\|�f�"-F��Z�乽+�A)sK^Ӧm�ͱ���hD�P9X}[CF�;^},���~]��!?�]���B*@`0�[��`�JT ��Ö�s�N�ě�� (Pu�8��Á��Js� �pp.����J�"��	����|�)��$��iIj�f�og@���iL�������d-5d�_&DҢR}4��{48S1�F�ݕ`v=�����<�(X��&�?̢��'��\Jk�w���g6�0={���4H��g�c)v�g���1��acUz�n2)RUϽY�L�DϏ<]
7�a7X���8�Cn`.x��aBⷷ�n
���o��k�+l�y�A����\���+�S�6�"[j�y8�aDk|�/О�	��Eһ�:�SN��W�n���aqTBd��-k�V�����ky�&��1D+T?�H��#��q��.�%9xQ��bʫ�EȲ�y&z���b
��p'�`�-��b�0�D{i���.=���
�*��
�me�z�X�U#������+�8x�0�gq��R�֡?C$��ؤ�����K��Mj	�Mn�ϼ�]8�m��q������?q}��o�2U��˵����1O��[���铃�4�OR8M���}o�x�S�Mf2��B��N�-��@4�c����9`�T|���Be$�z�	�<�*G��k"��fAJВ�4����{eS|׽����Ih%)O���jȕ&��~
2���s��=�̜�2�y�a�-��,���iPI�]m���N�4����Kwpb|�{�ZSbl����꬞��>�����\���;�8�Ӓ	�|�$���գ�D�My=��`�ڭ%�c	��\���@RA�W��H���]]��|0A�g1�zB}T��3/��H�]x�X��C��,ڪD���ϐy+�^�ϋ,�"K��uƬ>�?m�K�M!ϭ%����l��B��tq,m!r��$����L㣕J�v`�ui��c�LE���!�|
,��#���;�W�&��R��d��)�{~3-��^��Io]�:ӻ��ȉ�H�a���e>w�(�I��zC܂���}E������K���%6̤uZ�,B�n��/佻��1�t�}IF��;����T��x}d-��Hu�(���:�j�a��{Uz��C~Y�_�Մ�$�v@h��)��M ��,�a���#��ar�����M��U�ѓ����^5ޓ̂ ��^՘X=&߁h���|�~�/4���T�Dǻ���$_�'�0��ؑ��ލ�p��PM����0�r�T$7Jr+��Nh��`,F"�3\ܺ������ ��"�}��Ew�T�qm�؂sI��~���v����W�deD� ����5���{�%�����F��`��,;j�ɗ'�W�(r�Q ��<�]�`"Lcc�����G.12���9Nۺ������RĜ.-Ga�g�98(U8�Jsi�E�"�uObo�>&(��T�z�� �B,p�r�Eݷ[
�%�"y#1E/���:3MU��2��F(�f�}���!3�-�2�Ь�4�^�W���7��A:��׽��@��k`*FJh��`6�ߠ���S&
w<���h����;.�M5h�	�V�P�Myp`KYP�:�L�x��>��-P����@(�q�ה����r���3q��P�g�����5���C�%A�t�
�sc@���5e��o��i@��`S4���a���`+��H���٧����gt�t�y����ܦ���O����|k���D*v�#+kT]��	�!=L�0�����CIz-���uB�i;?�-jA����!l��������0�/z�b�ܕr�i��20��wnϋy��"�a�[��1�H��Hfɀb����8hn�� mp���'�W�d ɈJz��%'Ҕ#c\}A]0逽D��N�T5�pQȡ�ɤ]o7�-][�[W͈6���z3�C���ü^U2��*���c��pՌ�
�d�a9ΐ�ڮ��4��.d�9��c7%��;��V䫝�.qW�?bu�6@��/��*X�0:���t(��r�[�����4t@_F	˞^E�z1�ɉ]��pԝ��N�01����̂5�BTsH�`������!(wlo���h�7Q]��������"�O`�n�+&��NNt���Ld��5Z VO�^�KR������ہ�Y�����|;R,����\����8���[M��L��O�;�'~���5DלR9;g%��~c�X���X���7�]98�A�{�~���y�
�v�<1���~�o�PH|�_��qЉ�	k�P�|�5���lO�ϴ�Z��`�;���Ss��w�o�Q�栈�Xs�%j�gfh�89�V���?܀7�[���q�'�25�MXkN�"���K#d��Ba�������X	NS�{��9Sn:V�k�c2�.L��<�9ط�oe/�ڱz�����"���m�K��~�\��B>���^�z�2�NV �p+� �������', Eo2���U~>,�ѽ���O��:u ��<;8�����Lg��#h��>��5Q�ѱWS���&.1oi�	��d����̌�u&Z��+#&Ȕ��e�:������z$�j���I�#�%@ �j�nȶܹ�i�h�^�fRR�V�P��A��� ��>�Oud$��:��b��V����5�GI��癨D�z'w$SM��r<�ؘV�QVDmy�غ�����Ld`�=`�>��%��sH�b��j�����X,�^��G~ .V���KE��#Z�ۧ_�J�;����4�� ��F9�*����̏�J~��!q5�^*_�4g�̂�Ń��SҊ~'�ʎ� �4œ��"5�h�h�R/��W�k��av�t@&�H|Qy䟙�d�ps�k	�%~��9��6u��w�ѻ��*I<�w]�5�Dg6[���a�V����瘎���P��hDj_��W
����݈�
�d��`��O5�iH@�#Y�c��NG�v=���f?�����c]��d�f��Ռ���܁σ��ot�o�g޶ώF�t�Q~���r]�e�!���'Q��"���෭�>%�ޥ��ܤ�l�i{QW[1\kH�E�\zȤ��W��,�4 ھ��5sX�o�O�q��BF�	r �$E�b�A&�܀/�濏E/��A��;�
�z\�� k<��T!^I�F��r��^3i�D��*��2W��$+�� ���-�~��]�z+ᕁb��m���pNa���N��sava���Q>+y�ι�v��svL������w��г�U���?�{]��oZ���!�~|Ƨ_#]P��S4RA�yET���������8���yZ+9a�G  ����r�nƙ!���h+��Vn�%뜆7z�Z�6׃�4y��P�#P3[Ϩݼ�I_Ӄ�rh�9X����'�P�HM4[�� I�*V	�aq�_�m��g���z"�A�/���}���2���lK�8xI��&~	m
�h�h!a2���;�M�pD}�I�H�N�����c��Vj�$�,��N����sb�-��CK6� Z8Y� @����`��1]��{Z���fþA�Y�3'������:ѩ�Y	�b~[E;�\M�βSS��h��o�1w�����T�7�J�2T~)���HY�C�UcƊ�_K��]����; �sZ��6"H�K�V�����lW5T��%m�G�d���Z�'�3�}:�P��˥ E����H=�X�����-�C�������]�:c�������Z����Mr��`� i�z��d����M���=�"�8�0��f-8�sG1���R�I�R/��<dKOc�SR�m���g�BUi�R����m8�qm��6;9S9)�!���
*A��g�A�VL��h�>SG\��j�.$�P����8��/��*(+���Aw��J�)�Q��DXZx�	�E�-�j%!�8FbOfN�La��@�s���U8� K���3Q��m��%��ڨ��Mr~�KE	�q���%[�V�f��d��m�6�V*�a��E�z�k�e�����F.';�4w�����i �}^4�Z�#���b���-����M�K?k��u.���/4n<�:liV���UmyG��;�,{r��T�/ooq�E+Z�
�%]�|Z�w����;$?��e�h?���@���֧�:Nb|�0BVE)4����o����9t��Ŏ����߹l1�E�ȉ2�Bǫ��X��1!�C,����u�F�OWqbT����T���\�יì�l��8o���'w[Γ���[�'�	Q-��[>�<(F�K�ỵ��۸�$���5V�O-gp���*԰�8�X~��I�����r9�xQ�b���n��]�vp��z-{�Å��LV�?R�M��w<K�v *�[�-Y�ĿHr�}JwXyT�X�u�h$Q��J�!O[��2�4�3�m-0��N0'�9�N�W�4�2���	.�l�}�ea�Fj[�O��Up����zs�,5��՝#�08pų`��J+@U}�7)�D������B}Ժ��j�ESo��{43��
`$�Ɏ?�o�����ɴ+�����OK5����1r�z�ꇓ>�voI�j:�����V/����M�o?������r�_ڨ(ؑ�Gj�^�N�!���,'ii�Zuʎ�?�k~<�&�� @G���󨶐��ꖼC۞H��ak�H^����]M}W�U�&��Bt�C�u����i�醶��`0h>Fq9�q��[<�� 嵇Oů��m{�O��a0�'{bZ����ޞ�G(�Xc�@���91С���g�m"�3����m��q��'F��"��"�=͈<�`-f�f\XB�P�PȂ5G��p-��B�5&L}ɏU�T_��kR�A�ف~bv>�:�F�3��yr�hbC*ɕ�CR�P��>��w��)C� �UԒ�M��V�C؆ϑ�ҵ��La<��\�E=i $7?y��PqX�V���KP�X���ي�Xa:oq&����B�i�Ë�I�����=`��K���fcU�6�\Q,ƙJB�o8Lʎrq��}D�5:4ʐWb��N�͗h�1Jq���.ϛ��F`<Њ  q~�Cv�%��g��䲣�+�է�Ky)ƅ*�T�RVP��T�<��[�\�E��R�Y[5�'(8�������Iq�-��D�-���v:
��.�Xo[}�)�qA�~�!���d��
 -�ɓ�+#M���kr16��N��!U���Ja��
��,�m�N���k+HFd�v�:���եE�k�ǃq�bߪ��cX?c�o��N���9fc�eʗ��b���8���u�O�K�ƫ��*�8O�;4		�@(��ǳ���\՝��o6Oj�Sw��.cR{l��Gs��$q���r��q�(�q�<G������f��.�7oB;76��I����Xl�9�(a��)������f�l���x�hdV�d[6�!��Ƣ�o����TD6����b����	ބ�ǒ�4&�K��e �ޛ��%�H��d$9�'U8n�"��9�-������K�B���c�[ ���Ii>q�֘Ac���0��d���[|��M�<%�2Ϟ99��4��)f���$����d���m5)�m4���=��Y;h�R=��W���Eƪ7���Qc��5/@��?�8� �٥��ZfǼ]�i"J`�g.���Jf��b3���as_,��,��r�E�\������y�v�7A����;�3�ٍKa>�j�~�)�1֬t� ĭ���{�F�b���Og�����e���n��m�e���QMP� �O�B�a2���sUR=��d�K�N�	��4�	 �#Zp/�!쮏[c$<�ɔev⼴�{�2�h_�]���x^_�Qb�N�vO� �k6���s�WGr���!��l{�	��Hu�������"��'3��$=�M�;����0�M���#i
)�D�ӊ���5�Uy�
4?��x	ЈP5F7����&�u(�ѳ`���c9��.P��9�Ux��D8K��]���>|��e�
�q+S�Y�sd969%!Ώ$��록3Ք�c�oc����g�p��������a<�%�(�gBt����+���to�I$���$�L��޲=V�(~˩��CI0z�����*�7>�ު{1o j-�x3(?��uI��TχۂKL����)н_��~�ɤ�f�����.��>�#��'QƬQ��Vm��ؗ��u���t.�
�N���Uz�����,-����r�p޼?�9�?�6�ܢ��X���G��3Σ}�bE�a�r����W��8^��K���	�B�����e���S�!�P�<�Bo�<�RA��__�3�����f*7@�n@�@\/����˿�F�EY}o�hwp� �w Y��[?�i��*�W���N��wm�Bi�M�����Ӳ�h�{�2c��q۳�&j��L_Y�Cד�U鸐��/Uiƣ˯w��6.ܟ���s^���E���n�zk�6{����=�xl�K����l����Sp|r�ܼ�9$��fݠB��(�g����q�뇦ђ��X�\ �oc�a��qN���^��ʂ�G��M��֍��{�3��%E#:10bՆic&m� X�l��)�D��52R�����[�7�yWœd�A�O�u66�����̙Fvo�E���84��jɢ��'����o�ܢ93��w���.˫ck�� �)�Z������CY�|��V����_��Xz���e��jB�ȸ���/�jW);�ʏ�V`�����A�?�T��T�D�CJ,* qeEioT���VU�����������3����s�8� �'�+D������gC���]莚��s׳^b�W1-ia7KW7�ʬ����q]�P�a�- W$ ��.�� `��G��O�yF� sao	vX8��!?��ϨA7/�6����л���2,�Bx*�y����6�*����_�~k�0ss�(ס�uB���Qn	�`d��랂����g�<� ʮ<����hQ��͏,w��o>E.Z{%��Q�Z;���N8��Fm1Z��> d���݇����|˔\U�t����Z�[�B�z�����M�e�w����Zo�f�p��$s�.z�DK���˪q����eN�pL|�I�Nakv�^H���u<fB�0N������X'�]Ԙ�p��̧������8}M��Rs�_}��fb��x'���{p΄�i%|���nA��ɻ��8����O�)r����%ǖEte��W+mv	����"�8�p��\���dZMt���?�e3n��q
V�1�|���(�nۏm�k�wF��/A��l7��Z62O�g��0:�-��[F�������SR}U6�4V�[c����{{C�|{#��ӣϠ�fNHo�k#�R�*pI�X�e��~Y��=����\�*9����FS�2O��������\�P�����^�I�xaK7]|H4��D��<���������ν�z �ʙ̲Y=�nΠe�z������.`�dp�����kѹ�(�Yt"����r�� q�3U�����`T]n��6�����g�S+����`�h��Wb�,L�D�[��q�֑D��@W]7�����q	HU ZyJf�).֗�H�
�R�kb2�ݏ���d9��e+ehە�۱�$kWEP����	^�YM}�:�ڙn=�ƌF�<rSj�RK�N�5�2��o�����1k@óf��G�Y��cO�`{  k^毪����imԦV�b�+�O��ݠ�ϲ��I�K�F /O�h{�����(�t�!�VCX�w�aq�Y剫{��'i���t8�z���[#i�����Ɣ;[�tZ�I`;�҂�H5�-�JY��X�s�\����%���z բusw�ͣ����i����#�A�i���5��Ē�t~6� *���<���9C3�iP:�p4=��"5v���|:����# px���S�K�2�qB��"B�w����a���o{گ�Jb��?��Y[@�/��k���R-����9Q�u��U���=ig�<8ե��5�-O�HP�%�n��U�5f��#�P���<�ﳁi��ؤ��ߪ_:�a��Dّ�����mb���ˊ��"A��1
+1L�3�!:)iM�8Խa%�B��P,�p9�D��Ϸ�\J7��� � Fr����B��Fa\h4G?��Gnն����X�� g�m6>n��h��_z������.�)'p��&��F�t���L3g��5�p=X/� ����_5;�j�}�l�<���`v�u-O��I�/�M2��]�(ZK��\�����L/�mi�2N�T��aM'k��5��k&ז�@�:`�Z�ƙ��=R��W��w��Ӥ%�Qq�I!H`�wn�գi�q��_�*>C�ҥꘇ�2N<�E��PE9�S��OO��bv
A���u��z����ȓ�-`"zWG'c�ކ�8՜x9�Gx���Q����M�N���a d\�v��^�4�z�X�Ϻ�amhS���7��L���ӧgh�\���"7���p6�G#�I���vs���"� �%"!6������JX����f�oN�Ul��slg�+@��{��?ۚ��+�#l����>� =��aG���1/�t߳�iar!!U!MO31�� eC���2���W>?Ɉ�6��In����ZH���O��������)f�K4݇�������LӅ�6���Y5�ѮD�l����hN.��]Qԇ:��5@�@��@4�lH@�{�8�w��)ʀ������-���U�I�����Z��0��Fc�y����H��b�����Y��k�7�5����@�Iڷ-�@3`WQ���b'3��C/U\#��!8��t��Lb/!Ժ�78�T������4��	T��N�|V���3�a}JÓ�"g���������z��$\�	33oJ���)1~�p���٩�0Wg�6��j�`5=&	��K="�_�c��ޛ�7� �6�\��6������Q^l�����Y��#�l�8�;f�Y2��Ň6��u ��/^��ΦKG�>0��)�9��+eOi/i�B�-b�Aug�NFޑ�{�}F�.�	���F���b���&��H�
�V!��>u\�N��X��*���|$֓�����`���&�9������i�b�7�YZ��nr�����U��]qtW:L&�Y>�e��GB9v{}���^o�����VL���=�5��u�Vyr2��#����2��ME�d�I?�]�N�����E C�O�^��� +~0�Y�@UHsd=�0��r�@��!�9aR�I�<'��#OK,���;��%X�0�TD���+�R�5�֭p�Ã�R���:`���|�Q��uE4���Bۡ٬Mt�+E�K�$ć���C�h��v1��T��7�B7�Z�cա�?ԲB�kD�o����<���(!���YS��5-r!<�wD���8���� ��?4�;d&���:�5��X@��K�w��X���$�y�C���*�$b�˄�I@��M����zm�N4
ꃅ	���;�d�o0Z��@�&7�'�-|9hq�5`)(�Ho/=y�{�����b$��\��bq�l8�_��Z(\Q��Da�P۴7d1.蚋!a�h��v��'�p�#� ��5l����J�	�d� �����F$e&��Ac�U�+�&t�����>���E��.�j��b��d����i�|i��
+u�z8H6o5^ hs#7��+��~o$��Ϸ��'�b̳�V�Y�5�V�E��8�٢
��N�QϘ�̪4�����]�-��W�H����'{ë�a���	���Xִ
�w�C����mp���,I)�*��jD>�ܾBC��Nu�@��;(H?d��J{��+֦��,��n���Q�⦪��a��HQ��J%�:,�_��z
]l$�n�k�φq���c���!�E�:�D�8���г&�ه�������k8�8���n8�~R�V����*V��_��HH�����������R�B�?\�=�4��?�y�=��Z����:�"��L䘍8�7 	e��q^���#�N�3��`ɛV���
_��Pb8~���+.�����������ftn���@�?��8��!�P�X]lxy����i?��ZT%m	~. *����;��c>��S����n��~#��gl�t{M�
���{2L�$b�47M�{������:�)��J>�@.�1�ԯ��ig�,0l�ܕ(���w).s�!Pe����V^)��0������E��u��cSz�]��sS�V�H��A���=��sѶ=������Gc�����*�sfn���v�Y/f־?-�� E7�ݝ���嗛"��e���^O��	a��[�$��2�%�e�ː��e�]CUT$,};<�w��k06H�>��;�ݏ��ȈVD����x�B6%L%L�h��j<c��3DKd����괘v |�?�
ӡp�#܎���l7.w N��Q膖�	�wמ��c���!ZL��Ă32�;	�TfAP��3�=�P �O%
��8���fK���v���\�4�Z�r�Gf��Ұ�����l��e"��ݻ�x�/�0u�S�l����$YP����8��5q5�
;e���u8����.tD�J[k�lj��S�}�b�1t�ːY��k���t �H�$����:Y�d���Re�Io�qlx4��c�V
y�9vֽ�Y߄����R9o�� �A���"�{kZ��;���q"�B��.�[(�҈�%�� |��= ���m�l�E����͟�	v��:&��M4� ��G `��~���3B���]�ub��������Z�� +j�̄WI��� T����Չ>���o���l���-�S���q�%u���T���F�2�q�䅋8��b.5�;ў(�2A>��9���#s�A~�Zj��¾ME��Q[���͉�W�����ƶjE_���L,6�KR\m�Hf�-�g*�x��~�_N����.޴I���>lq�R��!I"Pr��u��T�>�`%6�˕�A�D�.i����@��x�_�W*��}����� ]�ʞ �n�T23 ~_8�������p�%��}�+�����*<�U��wq�K�V�����z��7�_������9�ub��iV4C��-����OC� ���6�}���LB�N2��b�5�bч]C��8.4�@��, ���ZOEз�U(Um��\5��W���>�~����x;�u���Q��gl��1U �.^Wd�2���P��L%L��� k��-
e��s�:���U=A���C7���U~�����c�-PɆ6Uq�!�A��br�`g�
+�|�$�$7�'�6�����s�u6�Y���]ܤ`�3���t{B.�291��C��OS�Q>�D"�Dw���;8ג�լh'�[[�a䦱���N)%��S�ܲ�,�N�z'\�l�a��^�j�ݠ�٨�I�SZ��ΐ��!��ʛ�B��q�ͥ<-��=E�6(i�-���)1�̅��2����#4���m�(�s�1^�닢����ِ��G��/{���?�(B��,�{��i�$I�g���Fܸ�"`��6YY�8�F�s����w���~����i����u@件�ʠA}����������Q`z��]�-	q�
qͥ��b{=�v��`鷒0�d�?R��X��F'�r�l�Z!!^jk�b�4ʬJ���Vf�X䛃w�٩��7��*`�Ϗ��i����9Rj�a�H�zY��l�Yq�
43M�}7����R��{#)�@;��ܹW&1�NB����}�Gh�W�lO�����$�%�]*�,h��0j��T��Yc�
T������c}�gS !d��PT�2(
��娦T��5v1�n&��^!����Y��|�UO���2��Ȁ�o��ZI�x��u#�u{S�J���{f�Lبs-�I\���]*�ix�@&Y�*�#NYڧ�o�V\f-k�K�ﯢb9@su� �4{U(�E�m����G�!{�����O߁��M�
;��$qS�6����W��a�n@RR�zǵO�3�>'>HX0p̶�P�����	$��}����Y��7���}�G\ڄ�S��5�y+����;�ƽ	�~������i.n`���իoމdaƶ3�9/��Yf�
��|�-�W��|0sĔ;f{��J��L���o�8��&����&�NC�$&4']4�N���������5u!}2d�:�(��*:� �I���&#��R���E�xVkB!a�AS�䊢0�Y���B?��� �U���-���1�{:
V�-�pY�����1�-�haF|�v�\�%B��@j9,DF�hZ�2ǽ`�u�M7YCE���qtJk���Ǘ�(�?�l��h=��<��\�≅����nT���T!��NA�j!�b$iP�vÇX�n�mypS�������aW�B�`�7�����~��m������{[�����N̦>�9m��uw��;|��2k�D+�'�^b��6}9A�L��r`	��l|l�eB�-�@��:�d����0�ؗee��~L0�ڞ���OTl�cz��?��%�F�=EB����N8�/F�ݞ������Eș�g����m�f&0�ar��)u���Q�&��*d��dsa�b��GX�O�� �,PS�v\6P�,8���l�9c7��:�wҺ�`�F�Fq0M
���c��V`�ϓ'��Z�F���

Z�p�枳�X�
�m�CxX�v����C�J|:�b�U	�	�~,��O�ަy~���3+䜸�]L'v�������H����}�ȣ��=�a�n��d�a:����c��{s�R��</���O�$�t�Ϋ`q��(j	�R]H����8nx���/}�����a�����X�$B������屟	�T1m���/�O�M��Os�IK^�l�M���D"�R���6~����(QJm%1љbR�-C���hQN�<d+$[�J��u��O�ʻ�><�Y����hV����6JԿ2�T>?Z�2\8Q$-���ۨТN}�� ��Q��w��}j�ҿ��38�\�V4kk��.�b��mo���9���%�&���%������W��Z�,*L��p����$B��E�r�$}�
O�fPuV	.]�K��r����n�zx���\%�����"��E	�BR��N�\�Τ���bC�po?�;}Y���,��Ҥ[��#zB=GW�_�N�F�н�CuQ�ћ����[�g<�r��a_n�h��ڸ�l]�s0���LŐu�N4n�������hjS`�6����ӆ�B�)|�g���Z�
x��2v���T��*%��9V
�qD��_8��V>MJ⁄
�h����v���SWRc��f��3(h�(�h܆�=#gj՝"�G�}�w��2/����t����Y�R��׆w�OGĚ��s]k���ht���W�����4��b��؅R �|Y
`�,�E�ʎ��t���~L����}Yp<
IXO��I?��֎�u-w0Z��{�C��N�6�8&�?+�������ݖ�LW����0P��Q/��p��Hs�}�{�C���W�ǃ�9-�
W�4-b�-`�`�'�n��mA� �~�o9�o5��,E�r[�j7�b` �[.�2`��8�|*����#�ܶ2L|5��˞����7=�⢲J�V;s%�5����Z��!���#]�@�#r�!m\|��̪��de�Q��K�ߴH�%6t�޵cدq�I��č�����R���o��^:�2�2ְ�`�g���R��VW?��ƀY���@�1��T"H_�4(r �� �p���I#�q-���A���Z�f�)x�T_�u���+��n�R�J�L��գ���yn�ƃ�����f;|�8&(T��[��ܴ/����ĮA�C?Ձ5Y"�G_���G(�M�Iؽ�n}P��!������Yb, Ꮢ&0��Hǂ�򇕭������+T^��ap�_�8cu5Q#.��~�b���'	)�3+̠�E(�'�_2q��)oz&r�=F�d�*��8wmٽ���a�2�Ŏ��}���[�!{�C��b�ao�7����B�v�r�#�Ț��j!��L�A�Ύl�D��/P�m���ccm�I��k'<'V0�wB�z&%��q��D�<��lt�|OA�H'�r�����[W�xW��3��GV���%: ��i�Ї'�C�^��Z�αpn=>�0���|�
�s��]����タl4�Q�*{��-c�$=��1d3.��+����ќPZsb�Aߛ��7�5�b0�g���#��o�༱���U��|�Z��O>��&I�K�]&pc9���Yk���P|��myǟ[8o5��Y�e��/�������.��
�?��d�`f�_R��	��y�zE��5g�%���'���r�$�����r��?H>"�7�C�H�E��V�Z�@�ܾ(��c���e��m�����"Ĭ����R�p�4Y��r)�ve|�"`q~�Lw��=����(4�5)mLu����dd9���H�,�lT��9+.V�#`*V�D.y|�x�H���B��C��F� (�����+����nC���ّ��V�Z��a��[�͎�6���|��>����)n�S��|:�v:3.�|�vd�:��E��rȭ[��9��$��Xx������W�$m]���}|;^-�2�^z��a���L6�E�0 ��<I����Hĕ��*XO��n~���vӢV���cS�@���ʹ��T��E��u&b����iU�2�Q}T�R��=geq�����1p`I�{� **�_8�p�9'6+��2L<�Qw��;>o��O�i�w��s26���*���e���M������$��q�1��?�Iۿ��^���-����ǒ��?iVx�� r �2Ğ�<s9tf[2D�wZ9`V�ͼ+�󸵄Ǜ�R��{u��5���v�;K�K]&Gх]
�p�s���Ѹ�����͢p/�t-F2�B�ޫ�w:�䩬Yg�q��{��D2� �-�󤟻n�_X�a&vh�W�����4�����i(����?��B\�k�)b-��1�#���KO��a-�"������@���։N�a��,�������~��Bb��(̦<ƕdb9�|�p�%N
8�#�L2�gMrE0:îEn�ߨT�*02�[�Y��tl@���z*B����q��z`��<�y��o�XW�Â�a D�:�u�|�;A��rLVF�K(�[!	�E�C����w���$9h�^���@��"��[�1OL`�c9��*Fkzr��#��:U�@���;e�uc������B_m/6�~��Jh�
�-NK���T��n\OU��{g1��#��Ɠ:�������4,�ep}_�=$�Rսq+sz�7�ְ�3	q�v�[��zWHi	�4m��jZ���i�8�|����X����/��N���jk:_u힔(�p-������Z"!�a��bl����`� ��h$[�nՁڞ�2�6!�
�K�c � f�M�_�^\&�^V^�I�\�.vpI�p����$����(�VC/>.� O�%b��mUY�s7Pq��G�Q�j�s�h_5+�Y�+/�]��A*�!ö́�����t����(vD��)��I��j0G�zo�K��1��N[�}c�s	y����.��H�� �O��98T����N�f��{�Wk^v��������Ruj崌�R�#038/��5�80S��Zӓ��FϠ�> ��@�E�M���A�HhO}�i��M2��wr�`�K�ˌ͙07��M`�7%ǳ�C�%�Dc�D!Wo>��}z>�#�Q�VI7�\���F�gu²W��y�D�M)�x��B�wǯ��,��t�y	�	���!X�c
V���䨌���ퟙ#J��ߟ'�ڀ�7�5�L8����ܩ����u"N��n����.�;�A�����a40?��-��%�n�ڋ׻��(_<��S�Z�{�1q���4����F��3-��]X�69�q�n�WG=B��1Vf<1��t�M9~ڼ=Q�@n���s�z:�}`Y�S9�-��7#���Q������׍$���n�V(��h�3�u���jd��FjG"Q���~#����K8�S_�s�w6D�t����]��*6w����
^�x�G��%%d&Ƙ�����+|lf_
l��|�j'c��ח��L� i�C��ƑR������z�Nl��|�]��'>��:���ċ�M�ን������wV�yc��<��� �UGk�=�~~R��eXI�����Ȝ���_eIu�l��)�C#.Y��.����2�q Zg�u^w����Ș��>���=gEc+nd��ҺR�m��w!C2���+2�~�,�r�U�cG�i<Slv������~�6*Z�y&�
 ~�$<��
n�)�!m	lQ^�O�n
3���k�~7��g+���~��q���g2�N
<U�
�1!q�;��߼���j}%��f����ލq�Aw�#���K�[	�q�����<n���w�`��X��0Wj�5���p���>�#fc�m�r�F� לq�l�@��KO"s��#`؝�'?��Y���e_�@�	�.��b������>A�s |1�I^�K�M����}%�tz�v��iǐ�wЬ�������)�8���	yI�Q�ԤpNE�nd�1C�fP�y�l��c�9#�m��Zw�%��hH����bE?Э"yF��%���5X
0�l&�d�Vv��k���Y��j���3xaG�ca��7m!1�� �,8����8�%:������E0��b�bFD0<�z5ٛ��D���+�7�˗DP�Э8�)�|ӱH�ǿ�X ���C�'���K��0���4�c���&�ĘhJP��'�QgW����[㖾_E02L�<]�׶���RK�׽!g>��_O�[���׋����nF��I�/��r����RB�1s�Q��*G�w{-��k���g���ڴI��7[YZ��Di)���~�RS�����¯�t(^*�Lӳ&֩=�oj�I�4v��.9�a�n֍�ʹT<%��P) �ڌ�k���������˴��w ���D�k�ZkU��ƀy5�C	%�0+����5a^�@\X0����~]����t�:�pC�P�aq�9O�B�4�j�)m��7���������&�5��2�>�t�-�Y��!,�S1t��ڇ��K��J5O. .Dv�����z������"�a���m_Y�zo�]��eGK(�f��h��{�K?[$��I����y�;ЅQ��ޣ��T�� S�t>۰p���,
�)�,:$��l�n��ͷ�d-!�p��#�/$)�Ӕ�D+H�q�9v����,���f��
=&�; W�z��T��~�j"IUm��@�]�t���a�y��ʲa7��q�5��8l�T5HM��G��p�dᢞ@̎S��-������������X��V�쐒\�%=�xvD D�Wí�B�sZ��҂��G,�$ٸ�$!��ޖ#ߡ�	��cN�P�/��/�}�B
t�����q���i&���@jXX� �;����B��1d�e�)&_>gE�9<M�Ҫ���mS�E��?����$W:Z�;<S���z���~��F�k)>M�yoPl��)&Hʪd����kdH�%s{W5x���a�,�2r[�f"�W��ߗ��;�������P�H<5�LMa{�yy�#�b�%F�L��r1�b�<�Њ섧�Y#D��^�*����a��3�f�,�[ѪǤW��?��W�*K|w+�����=��j�9�x�L�]fg+�P�R~e��}���sW�.��{�pX�R��O��dU����;��A�� :� y׿��:��<���C�r���k���F�$I:�{]�u#�Mm~�"1�J*0^ϿդZ;������J�����ڢ=��Z3���!D�l��8�#�(
<B�	|c�2���Xr�r�=��t�X�i���^����
6��Ġ�r�'vW��N�f�РG����;�e7s��>'1�eP�V�|2[P��IM�_��5t�K��t'>:�T*M>�P|���kaˁ��ī,��lߤP�k�:�v���:����F[��D�z+��ΓO�.���������,��.����8wa.�Q�U��P��td�bt]*n��i�B��0��1�{t|\����g�ą��N/|a-o��}j�*�f������tڀ�������S�Y��C�A5�}�6ك����K19 Z\Ba5��/�BQ|EY�*���g��=!���~�T��{�}`r� S�)��y���LbB7F�ݩ�W�t���|��\��v=��Zcb������1��yb�=����br��
7��UX���_vR��k�o�>�bG:��r�Fp*������� K]���+�G[�ԡ�~��$o����oU�H�@ǹ2*�g ����(4�Io&�;�~���2%�]�D ?p�E�=|�ǧ��d�����H��:��}�e��3�r�};i4x'�SvAED����&��X�W��f�= �Þ w7��P�ז�Z���i8���"P����U����\��fbM��Zg���Q�@�0.MJ���Ʒ�f� �!��E��W���Kͮ��U� w&ذl1x�e|n��(�[p\s�i��?H�|��p1S����v/���h��q�y��r�4C���;��3��*��ZC����WG{�zCdLV(	Pc����ᅼhw#m)~��6�T���,e�>a�O����P����t#<&"x�f����B ���nhN�8�V����]���)!�ci�ci��XhӐ8�k���0��`�E��he��b��118!'� �c���À5p$�1}���M�5&גLxܞ��~JL�K�U}n�|��D�ҙ�<��vB��O]*�u��u�qM6~�mB���x}�j\T/����"�xN_�K9�����}ƈ:���T�����BB>���o�& �d_ɅEۮX������v�"�AJ)�xA�;���2%��%���H8�U)�� q��pS��q�9o�v��t�A(��~��{��Z+�(�