��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1���e}ʲ��cg�t�ϙ�a�:�KR�%���ݧw���ȼ"~m���7��e-_dA�� ����Ԃ_��ia����Q��p7sB�Q;�P"��a|��|y�[�0�9i
+�FےE�~�[*
��0/S븈'�)���}SuLq�T���R@�`;��ZEei4+��C�����HU���
*���n������4��Y�h��}ٰJ�XJ������b
BI"�M72�*5e	p.̂�h�1S�%���!24�{a��9�0ہpF�8$�X����˪��V.3���#k�6��2�������D��	�p�v����-�(6% �?}Ü��=���p�S-f	eccm�,�d��Y����9��}ucا��	Ttu4���0;a8{��F�w�*���z����t�+��V�X�Ů͗��j���t���ɵ�.��U±H:F�<!Ꭽo�V�:p?G�(�a��R�g��4T��Ww�;wUk0�f�{2�|)m*�a��T�2n#T�OFۈw"j\��$!���&V)6�2Q�����l��0K�7!��ei�&�c�i�z���]uD��]R�OqR ~Z)k`Qo���(�k��ͱvΒ.�Q| 쾃;*���{�\n|���1�&˞12ϸz�/Jґ����A�,@;��b"48��Vދ�k�{}>�Æb�A}��I�de;��t������� �9�sj��h���3c|Q���}��`��g󼗈����$�g���x�6����+>�ǝ^��aY�� 4��
���R�� ���	���Z\�MM��4�Sk^���A�`2��5�@�����^��:��������t>��}���]�:�i'�ˍK�%�(�@A$+?��ȔyO�+T�J�-�5N�:��h�?o.��_���3����6��U�ѓ̯?�T� ��,7N��4|���;�)�C�u�j�N:��39�Ψ!K!�}�Z��UV�3@�0�˽��0֨x��U`o�ny�t�;��iן��|L[���Jh���GI�+�,[>��չl�Jִ��(�Cy�]r`O��a�bE@�M���R�i������!�p=N)s�*��T������	6��S�E
;PS>�ɘ	歇�������-@tX	椺����zG5��L��h3"���6R�HM�D�K�v�ş}�]�[��?}�ɡʄ)ۧ8�3���E��p��Y�)��# h@���s��Z��,�2n�&��7,��8j5�]@��J ��U#���AC�_Y��Z�*u������]�v��jgeO�P���N(6�:���eǏ����HP�6llN�O:��eQ� ���Q|�ڛA�ͅ�R�{/��2Oڦ��AQ�Y�����G���\�f��T�눌��� �%m'I�-.����B���rU9OJ%,��� �������x��b�C�߼�wk?�����J���>>g����BAJ��ei����ߍb�(r^A���B����E}�V�S�x��D3��u�.'��k��R�vX����$]퓷�dÑU�J2x�$�r���s�;�Kp�f1�d��(� ��]�=�2;X�T�Y�1F}�A-i�`\��6�$�Mw�])��p�q�{�:E��K�Nt|{N��5_���l�I��\;ϼ�\̦@;q.��r	6�G���T~s"����Tk1pwK/x���q?�^�~�sw�G�D����j}��/�=d\��dϢ�͑�U��E�綼�1���]�{�� �;������A�o-7��P�ʦ�C�{��ն�!ߘ��9�t���Ћ�J�|�jPv�Ŗbk�*�
���@
Gޏ
S��Ec�D��y�p���#���#U^��YW�X%���eu3�P�`Y��bHQ��P޴���S�*.��|^h9e�0{��7�*�R)#��h�B��)ĕ��0�}�*LD�W5]�$�v�p���Z�yeR��ѓ{b21��\i�۵��U�^p����,��H��B��#m�9.or��Nt�)��<S�c #�'�Y�x4�A+g�>VA��:*h�)c\;?���&���,��?�B��A2����B�'M���1[9ֶ�ɭ^f��K�ZLZ��v��g��>�����ʛ�>��I��x�̃=��@��p�Yub�����C���}�s��vws,JoI�-/�wD��U8�U��Hq�'�$��c��{0�F
YOR�ޟ�H̀	�F����U$	X�iT���B�ג����?r+V��@Q��;@���=�T���������7k���D-TLR�����r���Yqr��r��LD�3A/��-� �:t4]����'�}� #�V3;&O�]ND�K;i ZN�$����O����i1�<��� U3��@��Y9�cm��C���`U6g?��S���H`�&�~j�y�� A���wk8)�ոw56���G�|�L�["�>qc=�g�n�h��IIkfn8�����\�D"w1�����f���@,>a9e�aKXI1S��{�
����(0�{��m1f���DƮ�PC�q���ս,7@�ÿ�=jW;{��mc��{��lˡy���+�v �5�Rpm��3��
_6��b�t��I��٥Z+��^i�
[��%��8�F
z�NM�A�/�_S��ݍa�(��E�n���*�����:�$
tS*D?NLa&�hkUo2��m��
H�l��tvT�%2�RbOu�,o����5���/Ӝ��t�83|Q�Q)V� 
�^(�^Hl�RQ=5A�JX'� ������bP���^�����7��!;��2�/�>��B�o�q2c��y�EqMBR�]3Hಒ����O��O`uNTij�NL�y���
q}ˀϏ��r^�g |�TfJ��Y~����.K���Y֎�$s��"c��h~�R���VL��R����.g�s��S2�ơ��"m�7֤�l&�iqȴ@呫�x��[�jGh���˱i��ku*�|��LTWb�P@���О������Q��*_����!����v�����Ѡ����l�D�l�_�鑗TA��������/�Iu�¢�b��h�&��F�����Ëb�h�o��
<R�)z:^���Tk,!%JI�i��B����XԿg�>�5��:�G��З�k��hb��Q&�M^���n�Y��nrl��Bʨn
1��k"�]�oK��Pl��^A�n�؉ۗM��BMÃ�GOp��d��H��Kl)��VX~P� #���)
m�gvH�z�"�^c��P]UZ�;Wő��x�6E?_���~�3��`mN�	���$��MR7N����ò3tc5�)��h��"���s���Efyu!�?h�&�"�1�?hbA�g�[�ȓ�P�`��i�tlO`f��u��Ŷ�]�
+?��s���A�@Z����M{#T�:^�������q��^#鵫����ʈ�遄�^ħ�5�]Z(��PSiU����BG��~�v#O���Ӭ�Y�(~E[�����ۻO�>XS�q?$�T��J�*��bWw��:"��~�V��=�i��{��Y!X��	��ޒ�*�[����|�1�e��wՠ���fr���%�gw;�Y���i}����]��l����x#���ø?=�8'�С)�Z ����@÷��-CT�dt&�7�i��c�
�T�ſ�e8EuU��DmHEeP�P��b�����L�M������
�/�
6�x
���qH���F� �O���,�G��Ɍs�p��О*/�g��,o�f��m���ǱV���(�b��x�/�����a:b^3n4V_9����� 0r\˶g�3�CE��=��EQ�1����	.((2n&O`�D��g pJ_ũ��S�dw�U�u�5�����2�6��~Y�t���h���cڣ�`���JLB{�p��:����{�,�ۢHl���9��!�C>�)
;1��u���^ϝ1���#o�ˉ(��jl��z}�I�ۉ�\�&>犱A,!W4T��$.o��j`���T(Јlɳ0�t��A�M��	3r�#��c��;T-���~�('8�@*7����o:;�'�|V�l&�����N�Ӓ55�p�I�gJ�11�V���y!���z$�&�*��r<]����`	ɣ��-*[;��J_��(�&qxE�F�t����G�x���v�YB���k-�@~f�>mT��0͉��k�ف�|�ŋ�B�S�A�5Ց�7D}𤝹�DA����i�̽六�yi^��,ܹ��~ֹ���)x�ia(�s��l~=�8U�����)f�h�_��r�U��t����k����_�P[��ۿ�@vwC�c�㾖G}��	*W��լy�j����/v�bk;���?T������i�s�<?�V�"X���3β�- �V�Sn�;����Dʶ*�K���<�}8`K���8��ԣ�(�_F��߃�*���/RؙO߶���̔�~	�>)i��o�=�>��>�R9AO��h��\�L�;�}�ڱ��tEE��PE���]s.�՞ǆ�PBV�8D<��<bj�/���)�w��Oz��	��"OϷM4$ �Z����\��� lxy�D֫�ھ�Bw��YZc�;ϸ��R�V�<�ߝ��)��	�ϵ��#>�����P�64���Խ��C:��$+��h'(����ՠh�v=���͝��+D8-	�W�O*��|�7���v��G����l+|�¨Y�YF�:��Ի��/.]w�2�S�{��؋�.��m�y9�t���K^���F(R�PK��Z_�/���C��Ap�N��dػ��Bf�T��y�B84�|�P��&�c��\�d���X#G@���\gf��̓�殀�HsM���!�6N�� ,�{fɝ�EL��H4�M�"�?'�/F�V�&ФP��\h��������zH�a�+
Ak��ɷI��hޞ6OT�B�l�&E��'�R ���?�� b�*�������D���x��Q��ݟ��޷��yG&}K���оM~|�ccIV���F��k#�� �H���O	=M�h�����i;�40z�6!r�5���y�R 3�r�à�m��1Hd ���Nn]�����`�ʈƏB��xX���H�I�5>�S��Z���$���*�6����
���+E}�2Sm�o�&��
VD�n�<�a�M;�(�/�;6%3�+�	-f���i���ڵ�)�����vI$n��gc�'/�z�"b+���t�^����a1F�S�q�����3�h��2&̆n7�9�yM�����,�,)F7C��p���I��A�:&��d��H��K���7���>�:� h�GJ�){�p�#��3�]V9X�=���n��oXn1�1j�L��GK���L�ߵ8���q�=�/�9C՘zF2���m`1��)`���f���گt���i5Iq��{�;��^��6e��W���6�C4�Σ?77O).��[/L��]Z���ke��k�T��CT��n���y�i0L#N!��9�Ȩ5�iWMH9ӻ	]�-��߆{�����!X�����\�@�4`/O'*��[f���J��b���?��x�ћ�tx�$��~�a�B����s�ѿ�.����������k��JK;c� ��B�!6�z +,�����~F��!\"vp�=�����i���z�Y��j��~��8�#�����q��>!�gKX�6������L��X��H=�
Rrf����"O���:
�pG
�D7��ЗW��*�j��z�wQ��sw�X���C�x�S�	2��2�,�[�� j36|#�$�GD��y��h�iz㴣qvl=4���ۅVV��|v�>��Mu45$���ǿ"���a�]�ti7vR��l�,NVT�3]宱W���CJ���^&�i"G]FL�V��t��r%D9,~Ny�c���u����.X��8�P��	$��mo wOc��-"�]����b�kH��p
�K  ���s��l�ty�ύ�K҆��r���\1 �*F�7�����A������֏N&�ye�y2��.�RǞu��~pd��`�K[T���3�����(CyDR|�k��r!Q~,7<Ŋ��`��O�7t��t	�:��������Jڜ��W)��ܾ���Ԇ�$M�ڮAy��A�w2�����܉�
W��!;n$4���2�S�lu�DD�����H:�f P�U �UE~���$� �n�k���T��GG�9C�]k���q��y�lץOώ&<��f�o�1N �%aܭ�O�Ф�����>l��Ϛ��	������G32����V�[3��ÿ�� �I��G�ŋ������ f�7E'�r���`�Tc�Ą��U�S6w<|�?K���!4�ӯ�	9�_�V�-z�N�1��@,EY��%�I{Բ�)����̜��^�V�Z?U�}~C3����q>�i=-+������wF*���;�-5�5v����:���%qsp.ؗEf��!�S1�P��_H�X@�t������5�����@Z15Ā��+��1�?r��ϰء_ZI�z����nq����g�ݖ��Ժ�<D���Q��c\�De8�]�� B�F�?�(�;g�W�Cv�p7y�hNĞ�-o�JE�ae"w̿,Ɯ�g9����h�/)�̀>�m�3���$��_|O�}��)���va��HȼIc{��-��������1�yJ,)��Np�_5��y�Vޛ�y�=RLI~õ3�A/uT�j���cd`I[�8���;[SFq@7�J܎T�$Bq-�(F�y$ez�i�8ϸ��u�j%�/;Q5ڴ3����i-	����`K&3���Vv#Md����9�*%RS��h��B���`�v�`�H�3�D��hش1���M^��K^rf�>��u0��{)nK�P�Є��I�K�=�� ��1	zY�mBdM5`��%� �����͍���	���a϶]�4��2J���A����k.��"��R�q\��7���ߔ(�b1�=�?$��`?�0�!a��ڼ�`n�ߌ#"�?�!ӫ<���B(�M#� �ƽ��0�q�?BJgk�5ݎc���>l�F�r���g�� 5.�	�����a ��-�wQ�?Kt��@�n�c6���-��#x/=�
��������AؙR.Hg�f�h
K�4˱{��[�C+�W< A�3�<���t]���PW�������ʪURY�TX��LB�3�O�|�����;���aL!T�7\B{5��,q-N�p"�����_��3�4�mt�T�jQS��n���!�U��
-ˬ�1���x���6�6� �TM�4cC����S�[E$���K�Y��6�|[�ڹ2-Ӡ��>�k�u��V;��������[L�K����:�̬&w]i���]��� �n�o)���:�
��6���L��(h���ط%�n��V��$�T�ڦ7[ϛ6OG�R�"��4a��cBB�a��b��܁Q n��|·۟��濫�J�v�ߕ�nZ��w/�Sy���:%�5�l$�r��:��~�n�[�\Oך&T%֛`<�&6�3���֛������R�:ɉ`5;��J}8$��a��h��Z@v�%����!'ڀ�f)ޛ�:�=W�����Cq>ڴ�d|ܡ���.�zh�L�����g6:��f�?�O�O�wz\�V����P�MY�A,�+��+;
�I�Q3�6�T�:�R]s��-��z��g}\��>�]����yu�����V���	1�:��v@����A�C�޶p�ˉ�ɝR�L*�:���Ic����NNi>nAg�-���Ѧ�p֘��s�����䉒)��K��
�{��~�:�t�5��C�bOus���v�Ռ�O�mAV�ԁ�L4	_��VeӼ@�o�<'����]�lt�H���h=z���W����Zp<��Ϝ��ݧ:�`�q�(��
�o��|���w)�u��	���ҘC�ڢ�����&��weQ4���v�M��`�;���
x'��mJ���i�W�lU/%Ɂ�o�=�G��-�P�����E
��tZؙ��-?��0��$C6�hл�@�Og��@��:T��} |�l�2{��Oe`;J"w>�R
PD���V���F�̮��\��7Ҏۮ��*���g�ѻU�2����Pgf14�!A-!ձ<��y=NJ�_��ʺ����`��9�7�2�Q��nGP`k&�d30���Hh�w@#��~�Snދ�S��\��X)��sπ��JO�$0�vj�J���0I&�殘�\6GvC�����,%��n]%�|I�8�V'�z�M�h��|�U�6`���RDJ���)���71EX�k�����>��W�)Y�T�$�C�q��i8��W�ꇏ�ME�>�.<����\��LT��s���X����$���О�la߿Ӣ�قP��L���io�Q`���w�xb�3���*�F�x��}E��91�'��P�����:e��V����աu#��ZݭW��_�<�1䬼V���3�g��*�4h��