��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�k�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������H�W޵α���N-�`��6����ݾ�FF��eF4��_}<�ےA�[,�|{�?r+-��ע9�!�"��F�Wnb� �i��a��c��v�Ϗo@��Z2�[�Sh�+����,��ơ� ���P��Κ�q&�&=�Β��<Y!�������\����$|^FBX9Lc�A-Y�N�U?u�W�MZn��Ĥ�1ϫ��6Tw�P*������O���W�v��*�8��^�a�9M��
�ey��7�^D���>;Z�{Gү��[ۅ=�J�z����)�;�Ů.֮�B�5�z�$]t[����w)��~m3<'bU���I��j`��!M��6�żU���#\0�?YMX���/[�|��ϑz�F�[�^�F�T�5W]�W��2��њ�D6���R_~gɒi�d��*!�B�ߎPh#x�~x��^�{9�<L�c$L����J�ޗ��1���UO�xUy�
>09�>u�
T���NѻΩ��R��'&d��+�|��j]����S�ma�=��\S|��j ��0����t��o0we&�%'��~.Z���]�	}}�k��#���f�qm�����t'�X�+���t���l��4�]�l��E9+���R�^��v1�0�Rɍ�4�κTUp &�,M��)�z#����;x�nĬ����|M�b��I���N#E�0:�nߦEj���7������Cԗ'���_K���mL+��UGm|N�" �ͭ/$����ʸ�Μ���{���7�S 8}-T��
b�e%��E�5����!�#���hO�Շ���Q�TнK`�$��u�
�+ē�_�Е�-{Ɖ�.�߆l[�#@�
pQ��*<Ʊ�s��a�h��c�0�!s��HZc(�x���f�kSkS�~ن^wzk;m�E�)� 0jPr7�� 6åR�x�b�9u�uC�q27_��CH�J��.ӿ�Cy�
�)���q�FÍ�a;#o5J#��BDf��E�

=#���?��-jPKW����W ~*���}65��x��p�?���J�R�Ju���G�>t�;��FQ��]
��E!^/�Hq�"��:�����nȯ\�Q-=\���ރ<s``�(7�ho�,���
�RNQ���ᢎZH!����K�Jr#��4]���g���s��O�ۃ4�`���{�.�,�����^����p�j|	�W���,���"cX��tA�L�2^����v8�}V���%0eN4+�� �z�O�+�G�b�vP�"�&������7j׼bG����7P�w��A]����Yk�� rf6�4@��(�Ab�I�O_ߐP-��d��j�;*��D�[%�̑����h�~���(�#��X"x^���I]X��h>E��r�9�[Rs��ÇZ��5���No�q�;�zxfwD3����r�mt�h�Dױay�S�(TU>7��Bpÿ6��WA���5%p��u��d��w`�������JU�����8 h�jX��\Z��WE�<v�Ժ�"|��l�Ψ����>�S��h�.lc	��,�JR�'�7�u�&�Ǌ�f+��O��@�R^�,0����7��q�  j���`���N�/>n��������H �J���8AQ�adt����y>:]Nʨ}���&��qr7h&���(�N_,�����I����pר>�
u��7�ξ	L�E��9",�2�a�P�A �2xA��4�K�@[_S@�K���.�ywQ��h|����~���je��5^�eXŢ����?~8	�]�]G��FxkeKw�rw~�ę4�^������sj=w��tX�:8sl�t��o���Iry*D�����(c>�0��ޅ)�ٯtQj�Z�|��H���|`�ڱ���q���|Ǡ��$���.���ls�Eh� ����VV�?K�H�!���iD�!��BV�Q�t���VWǳY:���+�шJ�'㎍?�6������q��2;ge)b���⌛(ؿ��]3�����j�K�j`# >�!l,!6�o)z+N�{%��rd�ogB8��L���G�3I�q'�l���D+�ǵ���X`�^mE�є6͸�͛��V�h�_�˂�[�J9G��h�_�-��Pahʟ@�O(�?���w�E��} h
o�a�T�Ц"Dm8$7݂�����m�RZ�	a�kUP;��u��DG�=��sO����~�s��9O�_�X���,�K�m/�x���+��D�N-j?�ix�������<v�dM�d��������2��<�Ѳ?��15��1��fd�(�B�:y��;����3���j�������(Q8v$�T��z��3B�w��$�-��9�uKa[��)z(_��Fu �X͠�ֆ��W����r�Z���#���n%�h�)u|���t*�J�C����		m�-[���������ۤ܅��
f��`�}�/�7�hC��+��^M���a'�������]�a)󚦱���:����D�(�%�)�X���j����tB�Ǘ����Y�|a?�ӣ�llz�UQ��Na'�'��}��F�fk�=�
#h��Ӎcʄ�w��#����5�q|h��/9��r�Jd߲h�9 ��7�Q�^����g�F�"��u(�*��&I+��M���f�*-�>o��G_�}�u������1�ߎ�'�!0� �ӷ�}����G�u��;\�3�����=��x�BXNǥ�Yn�\���U�-�c�5V4�h�������aL��D����uL"D<E�y�c�΄��\\�ߛո��f�5zZL�G�Do�x��M���^0�-��C.�������8�&����y�6*�S��b?�o<�^d~8?!��_�WQ������:Bm�&�)m >d���7�V��.��ie=i9�i,�ݜx�.
�.�t�qJ�����'����]~^��c�7\����l���-Ѽ_�C��U펎��o�bE�gv�9�|���'oz&��r0��!���2�Ц�D=>����(�ܪST��)��:�7�+
��1�8W(xb�����iLH# {�8Xi��L�y���Lȏ8e:R=�6e���Aa�4�?�IfbUq�܍�
G�2�n2�{��m�c~��le�L�}��B!�K&�{�n��S���5�H��S�3#��i��G�V��:yAu�ٲ���Zίͩ��x�L������ 
"'X�q���M��o����vLAc�5ﳪi�6�&���9�0�%�����'��D�Gj�#���f�9�xu5�9g�헉!�O���w��>0M��1]۝$A9�'I��3�1��"^���0�]��$i�>\���E�0>pA?��V}��0#�o3�LBC�AJV�'�[S\���q�{.�w`�%�������#v�w^O���!�Ë:�:�N2���b���Zɘ���Zèj��1��䗬|Eg�?gS$�$�پ��Ǖ@�S2��n���t��y�m��:�l�6ɝ0���b<�Ԑˏ:�2&x���dtn�0[��K�e�����I����V���Oh��is�Ԛ�@e_o!��m�Z��^��7�]˙"S�=820I��w\�7��8+b]����R��W7��!,p�\+��p��uġL��f,'���8���[L�_����2��@r�kV��%�����2-��ڴg*p����Y�ﳔ��.�M����-�wɅ�����u�{�dG"�J��X� ����V���U��u4s$�.���k _ ��ʖ����iE겙A���xO�=�o�	�&Q�X��t�o�~�;6I����#}���=�M��<x)�ꠥ7�S;]�����-�[]_�7�ᄫ�3I�x�Z"�ȿ8H}��k���ӷ� f�,�帨�^�v����D �h��I%�1����+�(�����w_�U��%h�r��x�C��� ��\E��� .��V��7uBv��7ࢰ��_��ӱp�!Ǒ�������Hs%<��Xe��b�U+���}(k�f	m3r� vt�I��ݣ+�/��`�>��?�d!�hۓv1XoݦF{_�J�+�,�$���,�[9~