��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\����q�?��e�I8�b�Ǽ$��"����ׯ1�V0���)Ny[�g��V�uiG�nK9���ē]I?>�D���%�E0`�A��J��>>�C-��qk��G%��F��n�7�wVf�p�o����ȓ��nB�~I�-�1�N�����)��ړ���H��ǣ�M��`Lsj�do�����O�����-?�P?#���馑mN�=2���;���kV��pp�#'[:����{��G�4�)zz[�.'�.\��( d�,�b����Pڊ���$��(X�-א�6j��#0�R���k~8��v��D��ZJ����l��0"��������lw��6T��~{��-[��)6�/|������u�h�� �T"%�֒H�E��*�_|B�w�=�+L��[bH���M�����H5L��Yd~d�o�-�$��h�zs$��6�Q���1כ�@nu��FF�tk'�4A5Z�n9���dɹ:���Y�����`���5�C��}H�E��XC�]��a�߇(v(�^�����9Lm>�8i����������H�U;W-d悆2����
�rè�5��jV��A��з$���"�l��9]�yg�����g�B���$�k��b�s�z�C{<�܍\�#?�I��m�)OU{�/�ڲ�I�FPV$����,���s$Ul�|�f}����m�TN��IR� ���N�;��y���<�1��<LQc�#R<.C�]��
�̬��׎4O��U��R��LʫO�j��L�����H�� a̗�$��I�����R$d�H� �n	;%�ig�H*N�l&�v0C�t�Q�k-e�hHjf�kD{���ۅVΣNB�J�b�Z��J���I8�e܏�}����S�g%A�R�IzC���d�}Vh�
�$���� 7���s�X����	" �U�,-t��Izz[n�9���ڱ�����m;�v@�c��c��dJ�Yˊ:���AK[z�����.[��,< ��S�M����;!�C�m��P��5hR�GgDG�U�j`�����EK��[ j��/����@�� �K���Y��_�Y��a �r�s9�A��m^���[C!=c��1��q���{���k��9^�8��5�;	M8���|I�01+�����yƹ�&�lTױ�V���aķmr A��\Q�M^�A����D���{��p��u��u�=Do��H�����0-��_(�;V'?R��YM�A�������ŁΟ�a��i�zC���*<"��]�ĖQC(�J|�Ku_Y��! PĖ���2ݨ1,t��7���Qp�~�Q(a�$F�������a�@w��H��Z{@9���A���uWt��^A��aFџ��0�"��i-иԉ<���dr[�#�"��1�N4y����BD9r�'��ܽ��tw��E%q�e�YO]��X��o���- ~�������J�����ևB����-��|�I+t��	�(-���S�'�&V�w��R˼O��RsJ)���pLp�]��* ���2�x� �3�2�6�ٕ��EZ`
 ������Tf�c�Qgs����_����\|u������{�rV�H�\y�+��:�w��A��3�sA*���-;ڈ���Nz�E��j���>����(�u����ab��t�W'��Y?/M=� p�)��A�`�@�μ_�A����hu�rrȬ�}BՁ�|����%�Dz��.Ѿ�พ��h��Cs�hȳ��%Ç�Zۀ{_��`�%����֛aH6�d�+���d��6bf�~~����+�k��\��-�ЬVa��"�4^��#Jabq����1�.������6x�k �O�$�X����2�J��$�	�%N��\C_�r�k�����j�vW��YT\��ր	'���{�z��PH�����<��t�48�^jkH�|dD�-��[Q�&n�Bzx���J�V�����?��@ŏ�L���q��`ŏ����o�Ih�
�v�ׇw��V��1�����.�77�����X�|��>z�@���ZCyR�~m\g��m���}X����@&3����)m8����{�z9�(gv�j�z����A�Bɇ�,0�t���S�G���L8�G��e�4�u����wU���������nk
!��$��KU���&��&"eW%؏����B��h���H�M81��\Y|_��k[���<"~��z�i�ec���Aq����-�<s�n�n��:�����c<=��[���gaV�U�(��QLIs��f%ht��B4�m�Cq7r3'�
�[�1�8Խo�acMQF�Lf�ۍ0,s(ߖ|ѽ�v����B$LA��R/��AXaC��{�3u@��� cD��Pff�}�J�u�=ab���ῌ��p�+E0q�kN�1���u�[�]u�?3Z���1��g���=%�Km�Vs�n3/h����5�)���ILM좂��m]Oo���;��YLc j�)
{2؞Z0;
��/)%�f����������Jn��\��F$*_$F�P6<bk,3��=Ҽ����- �C./p.*HG�u��<�E�d��۷1���A4�=���UL�uJ:����	nQ�=��I���A��N-���?�H���R�L��o�9I��I<NK&?���vx�+� bH-�M�I���r�n)��_h~6���Ъ��h�A�����PЪJ�S�B��K ����W�j�>�W'B�W�i���A��|Y�[�}l��I苭O��z��yû	|�Z�\SM���{x�v?��Q?7���m~��w+��<}b_oz�>N�����8�ľW�[�i/ݢ���.�d�r ���MU0�hb��=[|�R䨌�JM�X���tL�Q�'r��Rb��Ė�M��oG�ߒz&�T<��*/��pn�o �"D�\�"�k5dT��yo	�sE���ѽK�Ye�+��o$���R�D4��^����=���������Y_0�3��Gu�?{K��tb�o�)�l%V�꽿��>"<աa۪C�1|�ȴQ4"�'�X�~#4�]�bfBW���}�b�B��-�cΩM�&�8���E�j!�2	6Q����r���}��T	?+q~���c����ݬ^S�!���>�[P��E�O�'��	��)�W��D�ݢy{T����%ځފ�z���[������wk~5��-���;��gԼ��M�����w~!'^3]\;[��b}���v�����)I���aG0�����o��P�
e��
�(�i�5=㉁���nh��i�����e�z.�γ�y��OG�( ��Y�>����m��$�����c/�2���	�s����u�B5֪}!�@�4�S~N�9�C)�H�y��燦EEj�W��ɮ�L�b�pF���}�c�ûD�J���yW��}Hv�u�������B��C`2��f�]���{�S(��/��&�38��D�$$}�/,���
v<��qn����*ө�D��3�D�G�G� �$��:���ޓ�e�2�Տ��(�3�?�-:Ztv����T=���z�1��P޹�Wv��y��a�����!��B�N�o�d���)`^�!���{�|��ģ��ӫ,��ẦF���C���L}N�Ϥ7�� �-���%��y7�u�>��gs�Z�Ed�ʍ�	Z�������5��? �!��@7[�� ���vKk3�����I����Cd��#\I�VB��nMF��"\#H���rG�n#B��4�#���mn?�<Ea�ϊ�s3x�A9�:�:9�<�E����2�ҙ�A�(���r��a+`�y�'���� ��O����n�O�^��.{?M8ͅ�4��i��H�x�p���_iwn�^��*�Q��(i��̱ʹ��y���B 2�^r�i�<��2�i1y�0�W6�t5�Kud��c ��^�lݲ��VT*���2o,�Z@���ݯ?ug�AC
 A
�6���ߗ���� W��<���W=��",�ú�V8�A+%���vq�Fp��% Z�[m�<��P��.�u�L5eW�#^w�׌+��0�Q��WҪ٤�,��#P��E2����Z�x����֟2 [/:�n%4r�X��A7A�!#��#��}�|uRe�<L�]i��8"�X�k�y �1�*8h�K��!*g�QR1�kD������n;0���A����傚�/��b�s!��H��H�7�{���ls� �=�"��	�W�͇�KoL-f�����YR�>ME H|��x�b��j�Aw�ϟ�q����7	7��]'��{����c����Gng��8Y���ҍR��`�h���]>�tX8��Tc[��6��K3�-��
RW�F�Ϭ����;�VE�.d�1ER��cbY��6�CS���ܧ�{z��S(#X���cq'�_�و�hԐH�ηe�����rs��|�Nz��u��Z�4�>� ���ڥ6���".+�\�^��,tm;�m�6�_>;Ṑb�J�6�zeuMm���,՞C6�K�An2�kz%�3%%-w�uw�T+��=�M����;���C�t��s:5=����L������1>�JK���Y��v���Aj��%7��	s��dv�nSd҅�����T%������w�1R�T����"#K�)bǒ
I���X��U报�p(�Tl�덬��Gq+l�?
qs�0Ủ��΃]�������y�3��X�����~���o�d��V�S�V1i���J]��lB��{�-���f�c�.>�!�9ag�]�l�Q5����1�\��=��堯�2�|^�}L��4��q$���?�QV���u2G/���L�0��ŢP8�A����m;��-�x��N}���gѢU\����:5��1+Y��%��rѽ�ݥ��@�rڻ�1�b8�� t8���[���$E�P�`���Uޑ�悙A �SiMē�R?���F{KT7c3�����|ޚ�Ӭ���AU��${���G���X����K����s$�����U�J}��ٱ���� �Q!G�5��
u:zW��V�Xl1RE�V����rˏ�ʬb���(��-*J]�cp��e�}:d���[�)�M��.�`��)X����o��_� �_�����oL���z̪�홡�3PwNk@�e�c�e��V+�j�a�u��(��g���B��z��3S�릚Y���9���S���`�E*�lbn��3�}d~�A�p��I��gnKtf�c�/�����_?x�|�D5�����p7|�_S�	=_!>W���_�[,&�o������~��Ӱ�\L�a��jxT]I����Q�m�!�N����w�Ǡ�)+���O�1�t�V��ք�1�:VR���κ�sJk�(�]<���)?��'�$4	��kK�O8��3��+bH?�r�>GKӐ/�W�Ơ���6��=�&v?Mm����;�+���A ��63G��F
�¡�P�l�>?�K؃��G6r���8B�ؾx{���?��g��R~��C���"ώ-ES�c�Ԣ�OXq��[�u�������,ؗ��8$W!��{�CWфi9���DO����X�ɞ~�e9��>)%y�/+���w�)pY�ɭ#�l�T�������!�܅�+fw���9�%���
[��7��E�X�P�wO9�o�3��32:`�����24��.b.*?�8Ȕ/���@��e��Y�_m2ߌ\�x���&@�=��\/9��>«6�o�2�R�ބ0��9�|��u/M4?�͹����7_�U��y��xV��:���[A��4�!~'�[
0)�/"n�7���[T��_�ԣ�b���iKf�N��!��%�i�hc�u^J&�Rm���$N�ވ�sɝ���/�k!.H,t�l>G^�=���l��+J��4���9�O���6�2/ưJ�G�"y���>ziuj���-���jl�\��pB��I��,3q����	a�b��,m���D�?��4�r�\Uj���Owk�G���Ǘ���~Sž�8�?��۔;�rGUEi���'@��}��|�\0$��6+�R/�gk���)�(���b���� ��W�M�U���Pw<RI)-�3�F���
j�=��k�SÙ�{6��W� �8$��O�`�3k��+U���D|�x��iʖ�̻B\m�2."����S�y�ш�l�S.5�p}\TE��g�^)�W'�jJk�������#��O~�G��.2�h9Ԉ\�"�4�4��ɞ �h&�'bT�I:!*�}S6�\u�HE�^J�IiLP%B�P����h�	"��K4�>"E�ΠDߠ#{n��l��x��7��� ������RȰ),��D�a��.j�6�o�ڗ&�`�$&�#bG��f�7az�$������.������Y߷��;&c��Е�ڒN~y��e��	����b���L���(��64���t���e�6���h��������
��!>T)v��,�����1�u��'�ARw8����z��jk��/2X<7A��v�%܁���n@�����mr��YL �o|
i(����R͠�畧��C�c�%L5ų�!�}]�h}F���}>+�^�<:�Y�BW��/A�8B�(	�� ��#���dK��+6]::##U��\����S���h��������r�����+�-?�A4���o��Zbo%�JYk��s��fD
,��m�<������`_Y*���ad ����	i���3N��H�#�::��>�N]1���$ݮ�����:�ݓ�d7z_�����j�Wn��F0�|I9P�o���~�G��)F��Hi(v��)m,�9*���5{n����������1���%��xQ-���X£��R�����j��B�~��9)��:޳x�d��3�92�߾���-=c5��[�\4 ����-�<�I� �ޏ8�c*�#��0�f�.�k�]��!%�kn[�F��E��׈VC��? �����6��2�@��K�l61�֟��`)^����-7�\S�JP��I�c|��r���#�\�՚�S+e�/��1l����8�' ��|E"�ҋ�R0}j�s�<m��TT�93`k{�����at��s�N���?�{\+*�A���E]����g��o�V迖H�R�(dZ��߬�{GC8�]�r0~����D�.�*��YZ��!�P "M'��&vd���91X�H��XN!e����_`�{N�F5�G�_X��Q��x5,���x�y_ȓzasI��v/в(���)0�K���S�h_,�G���PLځ�����/pe;�;��e��/�7��Dޮ�|*�+E��U���&��ps�I����q�����M8�f`N�E�Gd�]�t�Oy��Ʊn���j�UM��f0`�J0f�����<``������*&x/#��,:���% ����>
+����-#<�*�Oc�R,�ވ���C��� N�����e �\�=��q����xeI]p0am� �ڐ����w`�x��¥�V�Y��ձ��q��2h����0��ˣ����,4���8�x�
����#Ł&���w���{<�+{>H�����bf�^ʋpA,��e*����UQ�(�n�K����5�y@�w=u��\��z<E��/���(H�K�n>귞��e�]&�a`ћ��ߢV��9�� #~1� �(�]��mKߋT՚@1^���

�I��n`��Ҹۙj�[�`���9��*MBЮ�g������TY�=W(��ӗ�֕t��R��k.6c/�р݋�u"0�Di���9�h��"vĥB�q�$�*i �X�r�J��ÿ�O��l�3 d;Q�`O�G�q'��q��0<�3�bW�M�U��^̔k+r�;ɤ����X�*@%',�j9��7�	V|���dA2 �����C�U
\�{�7$;^D�wn�=P8����Q@ ,���PܪŘ��,�ࠃ�� z�i���J�١|[
��^=t�+J�`{�y�3(�J�c�,���~�&�ߖKk�r��둳ڷ�a�>�H��v�KOY�l,ji��u���C�Uw�]`���l
�����؀?h�>�y[��mS=3��A��Oƴ�@_9� �� y���� 3ź��Ƭ�-CX�A�J��g��u���kЇ�]�W9����vPK,�h���N&n��Xi��ܢ��#Q�M�4~2
]5G�4�5����B�1Pz��kՀ��Q;k@����O�;bWN1/�إ��O�[	&�����z.'�"�r�Q Hn��)��+��X�c��W�h��Y����P�_"�Ԇ��9���d�6 �ZEAԵ�4�H���{��t�x���6�b�Y8�__3tC�Ѩ��:�����\��ñ	��>�v�P��r��ƪtO��h�G���¦�"=�2D'��Q�g� C�le��m)����R��mH�D]���2�8���/t��ojxY���ca��OX���X�5BϬҝ&.�+���acj��IS�q�Td K��W
�#�	ܤ�g�H��tny�ゆ�^f�e�ӼO?JP5���ō���~O��lםEQ5-�����2���M��6��#����%L�a2_`�b?�:)��]����;l�����B�E��"
�!�·�xN�7� �g� �a�~��������˺���~x�,�~��v�����+VHF)��gu3���"�;�y�`�ȡ⩞kh���z�D�۠�/P�>F���~?���t<���ޔLmƪ\7�m��$K���_�ᷱi���Hl�y-�G"2�����08�oZ�N��6L���ŋ�m�!��Ʉ�K��RS�IY�=��ê���~W�,d�t��^��dЁ��3������R�MV�=�CBj?����ÝHv��/� �����2j�~�9�g�&��7�y߿���\�B���]�oS��	A��x�F�4GE����GG���E�J�*]I 4A�8�����0l�+�����{GNk�4��8x����v�k}���� C���m��W�� #ˁJ�`�pu
P�?De�# =�s��X_���Q.%����o6�"��/R(���f��n���+ʓ��؀�8_��Mz�&���9�k����jG�ߏ���x�����È�=u/~�z��k/rh�LK�	ho5�#�[�~���s�yh�s_��' ��k��)6�Q`�9��$Mз�����?Q�.���kmô���ċ[�+?^����8��n�Xw�0I�쪷^?����W�˪^���ce�]�P �9V�������+|>�����L��� 5p�	N�+�B���6�f��������"):��!$�k�k�}����(��T]j��5�w{?�|��^�k+{�tA�nB 5�l8�º����x'�æ}���f)b��0K�T�����k���GXh��a5�5� �mϻz���g��o�uu�G݌����K&��!�xb�s|���� -�Kl��ml���H�u�k`����z��Nv�F9RY=�@�a��Σ�\(p6}?౪W��	�6���|�>nvؖ0f����{i�SW��VȚ,<C��R�ɵHl�D�x��@���}�����	L���2O�M�\
��J��_�m��@H���p����@C5\*?d�0�$�@�M��m�y��1"9�_ᦾx[�Q�0���{M	q�HD�j��7�[�Zg�Զ�W�?S����${�3����k!���,�m����BQ�,�ci�'��"��6��~}7qy�>�O��Q�EXҴ��{�k����k+�~Z=Uq �~?$LG��~�<o����m�ϐޗ�>�wQ*��X՞VĢ{���%X�L��[��:i�w��qDd�^M��/w��g���E��VQ��F��قu�[���[�?y~��68�q��+U��&{< ��Mi��U�>h*��K4����u���4�£�ig�e���b-���PWH�qd��B|����>MM.��0 ܇CCR�c����ߩ�|������Kͥ&<ޣ�b���O�'u�r�����),���V�����eu��	�W�E���Ø�D��s���?�C�&������~M��n&������7���)T��F7��| �]T,Cݨ(�{[0� �#�u]��cV�y�|�6�
���vlL8����B
]���'�}����9��s�i�}�M/���m��}U�pJ����\�MiÀ��nZY�����yN��<�"��L�}ٻ
�L�=�O�L4��RULHv�����-��R?��	������7x��@D���%G���8�Mx+���u�o` �p*��7+f���<��
}��]^��mHOc����O�2`rH�O�7".�y�Nm��zܙ��Gopb��O�W���ͷ�^3o!uDA���a]�-�z���89����
`C�i�y�{Q.Y'{����gP7q�܄�(?<��֫:����|�yzw�2�nށ�|�.���|1@���׼Tg[��SH�d���mprZ�Z=-�_����b/*?
!�:,FVjy�B�<�eW8��{-SKR��a~h��|d�rs�`׎&�=�^+f{N��M�^{�'�w���b&i<�i����>�ɱ���*b��'��WF�F�?�v��k�YU���Ԕ??�ܧ<�r�E��Pt��Q�K_Y�j�24pz����#�!(�M�R&w-R�>A]�=�)m\��-!��?6jl|j{����Q�r����d�p�Ti�+��.���b��_�c���1�s%Š�1K�"��M��X����zY]7�Ȏ�F�7C�wV��{T2�O?I4����P���Lߖ��b����o'?I��l��3a" u�c�����9C}��k��u���X�<��9�9A��ԕƇB�&��IV]𚭉����Ӱ�]����"�E�+8�i��p������+��dзG ��=H�����6�e�i��<�� �9�]Άe�����?c���fPk�\���gs}AV����ʖ�(�d��Q�s�$:��鿰��aNL	tn��t���g�~By� S��DT��ɼ�_�<�)o��-�m�\�4֚;��p���#
_Df�#��oC��%i��@s@����A�{���`]�)a o�,Ɩ�?��~��y��_&��TGq򤃡�闃H��a"+MA%*;�B����UJ�̹�0�*p��HrM�F��Ű� ��	E���PJab��(%1~TѾTJ� I�����V�˓h6�&���v��Б��lM�t����82��.,���=S��l�ߔ�ԟ7Ϝt$o�����k�{��ѫ�P�>-��!uh�{���k��$1&��Z����$$���$�48!iG���>�&���k٪�b�ύX�R􍝴�/>�fo��}w��kOP���Y�S��6#.r��h�TZ��E�uA��Ghy��"n�-�̹Ƨ�C����=,A�f