��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|ۧ[���~�(�#��p�f69�ٙ�G$������
�:/è��S���)���~!���5���QZe�Fe�Q�u����ꦠ�!^;C��uZ�Z^�m����K�����O�����"��IUE|�7��1D��Z�� ���x�)��|U�׵`�F,�?|��  ~�B�����Ŵ�K�.j��8��7��n�7���:�SU�?���<�ͦ�t��&�OJmdr˯��+�f�~�G3� Q�ގ;���׍:É�τ`AZ�p=z���R������vڨ����z<�~`73�vs�s���Q�	��O�Z�����`wݭ�F�,a��'c�Ĵ�8;���PO�nO�C��y�F��N&�)�[K�U���|9nZԺf�k�e�f�ME��ڊ�x>�*���ތ�9����{�#��d���缅+*���íY�[h�*��gx~�7?���b/�(�,�5��E�xe�5z o�p"N���;Hذ�BJ9��]��^,Bܠŀ%
�kn�e+�e�.L��Uhu�K�Āp�Z����<����I}��h��7k�V��>ݞKiXʙ�F��$s_.�V^1M�[B���Xճ=f�M�s�P��ly�͔�S8����fh�8��D��P��[u�N%���Ө_�A4dU��Ҫ��	�}Z���{�H�M�P��兡d�cS�u��6���2�WQof{�j��E�")A3�Ai��7"�Q.���?�^�	.gBj�8�z�ud��\�A��FGQ��&�a��]��>��Y��Eƶ'��t��Z~��iki�x�jv�8����H�щ,'�
��(Pz%0K��eڻ#aV�(���)lφ� KT��Pp'�wШ���Ҷ>�X�S���t��C�NF���_~�G��
؇�b�Mx���=��D��:��KF4�S���s>��JF&�v��>��>�<`��$��)h�Ֆl�Ĩ3_zB(�L;�&�n�YxiZA�IK�*A��Q܃+)5�'r�����M�K;��<���?��,��6�a����]9\&I���6��]�l��[�P�k�8����3QLh
;Y��h�|4~��4���:����)�C6���뒭�����]��J'�l�ۉ�h���<x��������Q���a�ՑZj��J��B�z[+�3h��=��c����B�U��"�T�Rτ�<K��z8&��7�둖��f�d���`Em���Q5�A��ʭ��$y�^L�J]����PR#L'�����[�­BO�}��b͵��[b�@�k�5>z�=l�~�Ԍ���G��Uɝ1��R!h�q�پ!3S&�,���b�z����dp[�Ԓꐶ0�P�PT��q语�f��ܧ~un�u�2�;���g4�"���XXǊ��-}���Vd{�]�_&��l�	�� �	��b���~�3��_��ǿ�3M�⶿{#h���ר�RA*��@�F��1;��.��" uĘ�h;�H�]8�8P"M�	P&���>b�4�mZ�K�Y��e1�A��Ԧ���m��@ T)�L����*`؏z�l�&��/�_�4����|Y�F�W�<�,!�	�ʝ�fe�⹨߼�+��/ɖ�%�lh�ma�ΰqH�a.$�[p+5w�%q�Qt�N�)ȔA>c9����>P�pT��������Bd/B6@I�M�SmZ��6�2�$Y#%/���D�}�ş!t�95g*�Lh��=���c�����+Z{'�k��rj	aI��4{CL�Ʈ�n+p�N��҈U���h��`��œu��-f���&�$�Y���:V
���]���~?��Yڽ.�W���JTl����8Z�; $k�� �2ɵ���!�2F�z���/M	ڌ���/�؀}�?�n�֞~'��YĥpVi<t�L)J�v/_D7D�߁���fx���x,qf���s���*;ɽ@��gp��0����4�+�/`�R�FA�b�t	��%Po���"k��O[*��D��H�qю&�c'�����;wc黑��Z���ꗁ�h���>l"�M����E#�r�J~"�b�(�F����z�[�c'�Ԫ����wQ'pVw1xH+W��jHչW�JI=2[7�l��a���]�w]=�Kv!��D�n'�	�qF	P���3~���g�i�/��a��/�nǰ��'&����VN�-�Y��"��W�����z��Q�(r�v:��q�����ji���HI|94�`+3�<!ބ��Gl=G���Zk�Ò�eH��+�{R7Ç������w�:	
N���~��콃N���Z���W�Oj��<�`�.���o<�z��e}��V+�Q��_Ǽ�Fógs�o8#8%�C a�ID�=)�;�@��dW��&sC��'}��9��?�0'�	{�Lu[K2�������ʿ}LJ>C�6t�������-�+[���l&��ܟ� L-�r˦�6/����y\���pB�`m��CQ^���kࢠАk+��C/Mꗼ��q{�l�&�V�Z-1�f,{J�vHa��2�t#��e��3ב�8BHc��B�eѻ`Ϣ�lŧn� gA�"&C8/�E�; �N�JƣN;�R.Ȕ_����pg:��%��f�"�|q��1 �`~oq�Ҧ��������S��l�\R��Px�.|�\�[�O���M�:3�X	X���[	x�>5�x��ǒ���TQ�4�W˯!$�.����Lx�F���F��&!S��:���w�����Q�D��V�޵mƽħ$>���w>�{�����o�{�<�v�(pk�-b�����g&+�F�=�W���
�)��Ec����T}�	��僜6���:�WnXEfJf��i�!7QW�e�l�y��k����{�N��9�
�4�Ν�M��ִ�-����Do�zJa��]��	�Oz��E-% I}X�>Z�0�{6*�t����IPb�~�ţ7m!A}{L96�=7b^�Ҟ��?L̹���b�(��tڽkC�x{�d=�V�f�DJ➥v.�M�iMu���CЂ�V����2wK�7M7@5*��zj?*F���FTu���yhe<�b��3�}kipYs�鍎��ڔ�qv�H3�������\y�ئ4ۛ��eЊ}��u� S� ]W0M0�i��AH���9�E�ܱ~ŔEg�zL��f����RAZ��a��ϣ����oM�C�[�6/s�E������l��ѧ'��5 moL�T������E������
�g��#սس��qa˷���l�s�y�	�-s��ދM�!�j/Z��%�%_gr(J<5��$��<8��̑�L��/CH�����k��iv4ɯ�a��9�Diۯ�t����'���^����\Q践-Ǚ����̽��e�@�������/�C�>�h(��:��+����%�˲��ފ8Yz�'�(�.Y�`��J� ��P���j��OM@��O�N���Ye���
�y�P5�\\D��JE��`�#����^�D���)����iP�2E�j�I��֎^ }�f&�CLa�<��H|f�c`��.7��F9�Fwnq�#ݸ!���'m,�Y�	Ų�����E����˱Q;��[�m������RZV�7���U��_�O3_�
k�	��,��� Hy�0蛷�Z��|�ߧ��Z]��_%��v��1l��&7s�a$RDi�%n/��e$���Q1����po>�N�l�_�fC|��	�˹S��j����1��~i,�'6��(,��k�v�>ƛ�k�d=Y�_���|��gh�*���#җ$#-�~�v!Q��&"�N'rJ�m2�r=��J�R&��ٚ�w\�;A�Wzٷ�'������l��S�s�|w[��O��Bo��oN�N T��u������n)��b�e�-�����?MPJ��S�ҶS�EV��-L}��y3��yj@��G����Di8��S_y'�^�
ϳ�Q9����������A��-�Pv�z�ə�О1�r�!
 ��@s�|fH��%.��:�q9|�w���r�-���i_�j��{�FH{ńa1��`|��|&T=�����48��	�wg5c�ǧ.�P	����`^�wݼ��c�wꏤj���Ty(Z0]�P73����}�����\��d�'m-��L��Q]ӯn�#�=�nd8����Յ0qX\p�cp@�H��a����ɱ�n��+�h�6�R�8n��,������M�����4�T6Q̎ӭJu��Y/����6dul����{�q!��3�T��IF8�(.�O�q��N�b���O��9�
�Jy����"ཧ�T8�_ ҫU���z���.� �"��xAO�.�QbT�wu�r�nЏ)���C8�FA`x -n~�0h��(�[�Xϲ���m�#��ք+��+u^�ׯ'��8��!��I֭�����A� '����e}�!y`�Ƣ�;@�FNߟ�;<�k���{$�f`?�f��7���@,����k���k�G�&O"�����+_�-��u�ME���t��k6��!���5�&哧\�ZS{Q ��GAT47#-��"k��:�.ZUͽ���Y���, ΌZT�7f%��)2��(lӥ��CP
��N��_-��#�,
���{sv�������,j (t �\���H���c�> Xt4*X0�@��D�5
6������>�=.�r
Y�mbl3i�=�-�sO�b�Kj��W�7t0eUSNB�zf��0g����L`��N
��۶-J�����l"lnqꤙ��~��)�#i�#���~g&��5+_7�](�)�O�k����#��.��@y�IK��7����X�12�AІ�w�F�*�i<V 
N^gi�󳊩��28�!��h@�������Ee���}� ��&�QЂ
��$Z֌��п�_��_BE�}?��������ba#i��(O"��n�%�C�DZl��a3�BNWK��6�`�[̖ew��'oT~]y&��6���e����X/&�Ü�P�:Q�Q&\d`�+�v8ZE�� ˷\}��g���x�d�� 3����*�%S,Z+#?���m9@���_�r,I��1��a�p+��9E�+��E��Guv���Y��,�D%ku޽Hc�Zu���������B�����[�9|��@n���i<$"8L%�nOr���b=�k��B�kNM�QK�n{`ޥ�����Z�5���N�6�E9��z�!�ڄ��*��n핌WՆ��ٷn��t��i���2�[���V�D��
 _$�"�+�;9�8�-k�/��������i���)'�By�;#`6�����9���)��0�y~:v�Zn���5 �����F��F���b��Ze!
�SL)_^��>߭���&7����|�~�[,���G�����V^1��J�&ގ�(# �>dn�o�>��^�ݚ�c6@�	�$�9�_9�:=���P1������1����֕AY��?�q�~a�Ti�4�ӿ9�]6ݒ#|鷙
WuRm�Dy�cjs�|����;Od��!����WXT��O��l|�����;�cPu�u�G�����)�?i��F�/��'�9�|��,~��1��%OpE���,ۭ��F�����z�|�����ڢ?s�2?!�)�cN?�.��x���9I�NܔF��X���)�����a��(4��/�4�D�˕�;�ũ�b��p�Yl�%�< )�u�o��@K�Z<���b�8`�����hu�Жز��	v��Տ��\��^�궊��������ikNyb+�ķ���{�?np!,�egО����J|mp~��b�]y?��	�ԩ�<-����	�3�.��т(DxM /�-_�,����˻<�;M�Fu0;)'m���7���2��7r�t�~M��5[�ɔA����E΀�/|T���?N9�~��[qR��fgK=@P)y���fȼ�3cX�n'ޜ��@\�[oa���f�rl�rO+ҳ���;����0t��q�(�;�Ӈ�<��<�p�����1Kp-�)��1�b ����vx�Xs�`v���Ց�j1�}i9Ŵ�_C^%�
����wNh��
J�*(�.�h"�W�F�~TM�D�5��eћ��W�C�p�s7����Q����T3� �STP��xK��]�	�{E/�@�-Ӵ �Ҟ�7�o�s��LU��̿;�b���d�bKլ3�6O��Ժ�q�K+pLɎ
������{D���z�X0
������uօ=�h�Ip�f�W�fƛ N�#�Yn�لڼ������`�ў>���0�H�0]F �]��KE����J̵2讜<��� %ѵ*�:�¶Q���d	��ّ��X;f��ڳ*L$-wu��2��%X�fz�	�=y$�~�8z>ߖw�>��H�Rb�"|3�L�<.�pQɬx�q��sA)6�X�%�m�D�D����W=z�q���M	�B o� ��J����?��[���n�f&�*☒Ĕr��y�����g� $P�NmP1y���T,˽�L��5ʄ;ߠW�`�������E��E�����ب&-��S
���Ʀ=�6��k������u'�ouc�F�Je�������D}�Z^cn[OҰ�]� b����'+�1�ٜ��ʹ�~fE[N�DPy��R�<g�ǭ����m�g>�23�Ó�uϖi@
������-�O�����l��? �֘;���i��=�m
&8�0s]�󠾣��A���|�(��
���OBSd�S��~�S��':*�ꖝ�����0O�oY:�E}��>5_�H}��O���ki0�>O����9V�� fW^�)a
L�����c@\���gۈW� ��rb�\|�{��HO���/uͤ=� AGk���^���e �ի����aU�$��\C.M��Z����U�r�V&p����2��*,�%�b 圥������e��}��[���[,�%T_ލa��	n�w�-�l+/d�Y��tn*�c��ׯ?a2���G:�j���V�Ze����Dӄ���c�*��[��q��[���$1$�2'#=���5v�֍Z�=X{��v��hg	8���K!o��u��z�m�lR�D^[C��thݨs�3
Xa	�0^��&E�sEr���M���L������swNT�;@�)x!�p��i_gW��]px:1qQecDUo�O\�Nuo���P��$����V�
ZhA-
��g"�qO ��>�������Y��]��71����>G���D�r3'P�`b�Qy0���0]E���n'Y�E�䏑���Z�jSDݦ�O���c�<��g/L����s��D�H��EO��sX�Rw���+5����c���:��D�!�J4ħ�R�&}�@�WDE%�"T�~�8�8�+:#@jt��nS1S ��/���/%�ŉX�C~?�) �h��������Ib��D��>�f hT��Q���Ͽc��<G���J	��#�}�2�S�L��Z���i��mݕ܅"���v�E����,����W4��E�h����6]�*M�e�D�?�����|l�*YS�$&����L��]$z��7P�G��g6�+��I~��1�d;����	��r����hY�q�׫MgW-��:*�j)��aP�k|�`���1x������yě:s���'C�.�!ܻyy�l|�H���`.��@�k�FrI鄿�������뫲�m����fP386�5��X-u��Uwߗ�&u0�������K�d��6��&%�@ܙq�s�T�����h]�����sǽ4������E�~X/>�i@��8�kMg�T4�%zU֌,���疤:
(�r�� ���6��AH�hr�rh�S<��f����C/� �K/�?�4�]S~�v�bhYӶ'���k8A�m!��-�F�����W�^<�K����f�?2�#a�fc�o�h��h��O�Z_ĥ��@oʧ6ô��U���'��Z�)^�*���0>��L�k>.bu���T���0������N�����	;�^Zb���f5�>-D/C��&{��^D=�|�%&>Uu�Vrx��a� �>aR�/2)�MK{H�D��n�N#�ܦx����A�a�: r%�,�����G�M�W�t&}�H;W|vcH�_��{o���Y��W���b�� �y�U��Q**����� V��*��N������뽧Yf��ۖU���pw��9�V�Q�R���!�����h2+��� �������z]�\�!��,M�mg%�n5�r�GUWOY����v$�Z�d����e�E><���g �N�Sb���/�u�@ͯ"��|�	׬�8OG��ue���#p�Ft��65-��kTn�D~���l���!!<:��B���2���V$�x�Wj�sv�k�C�3������"Pa�L(�Ttu:ƭX����$k�[;$�~(��HZ�'��S4��(����p�TM/���$�l|��O�u�짩�Oԅى��$!$F�(������~��Y3������z�f(�������H������/��h@�*��h������H6\�\�d<��,e★k �6�w�~E_�Z���]�A7_k)b��f-�s�<��'9�L�d{,�m�9��QReLx����A06��8��(�s��_
Uk��X�X>f���ō�S$"�4J��ɍ�Rlx�nt�~�d��ǈ/쒞�Lʹ�~H)i����,.y����a��ǅ���O\B���3a��-�������r�F�3�F�.�8��3�&P��]�Ƶ7wY{�q4��{2��kҬ�3Ւ� �����m�n�@0E#��ģғ�H�V�9jvQI��+P���6��l��nm�������V���`��1��|��o�I
>�s�Z�}�,���IY�|%��l+�-A_�W.��xͲv��W��\k��-�x�Aur����;Ko��Rz�<~Ph#�D1��~�r�֙(��gA�1`�����#c��/�'Bw7q��� w�;j����T������*r��Ŀ���W����3�)N:I����Q�!��Z�3bs�P�|{l�,5�u�jH�K䷒���́�Y�ϡ#���֒�l�0���Z�9r��z���j��1e��n�mDA�L1�8�Z���J��O7��
?�5!k��ٖ2T�/�3V.,�F�S�{ӄ�6ن�+� �E��'��|��݊�E^QЏ��?Lʥ�Jo���C�J�e�g����g�a��7�*=T\�p�������WM�a��#��胚]X���m�r%^�7���+eܶW�$}W������~���4���?�e��)f�,Ǩ�{7�z:W�l>�q���y'�K��9�K��M�_S�0�^`:49?:�m��8,���I�҉@
^���ۚ��6d�%f��Yq�x�*�oJ_�}&i�_,��/mu�u�'�&��ĵ�e���Q����I�C@[�	��'�6U_����5�k�
̊!���{n���<.
�ӄ�s#p�����҃{Ӷ�8�U%b�O���?��4��.�L��
�5���E|G��Da� ��r`��=�ՂO��PD<�q��� �e�� 6�Qkc,i7�c�k��]��"�(��~/�������eB��V�L�����0a~Q��ܦ�\����C���u�<����,�FV�v,�R�zi�.2�Y�4��bB��ϣT>�hW[lS�Ъ��d�t��8�Tn=�d�AfLQ�Aӵ������g��y��b�$(��2�H
���;#�0֚?���s2����:�]��R3�<��d��D�:�SF>�V�>��%yx������ƅ�dxh�Z��h�"a�J��:6=�3���ɼ���B&�j`%�է��H ��$C����~#s�Yc.���9�f�gSln͞|�Gr�*�'M�x�TV`�������n)���׺~��g�!�[lDR�����wG�]���dl$1'�����3γ � }��^v�89p!G��������ܵ�S�ov��ju��/?��h�&?_���D�����ٯM��q>�v\��s�ڀ%�<�lQ	qݯp(���x�hp�qt��l��r`�Ap�j��$TYn㧼�ݜ��(�q�gM;�}����U�l�RQ,�~�D)�o�,Ku��}e��(w�&ՈF���8=T�;��d�����_`W9�Dk{c���?�K ���D�\t�V9�OoYf��d�?� �}/����D[Z��T�|���'K���O�v6�X�\�^�4��7Y�rӾ�H��f�Ws4ȴ.�� u�jE.���xni�8�z�u"��N͘�7�
��o:�@=�ѝ謄#F�������9���j9��%an�eT}g�Bf�zr���,�����K@1G��h�}��h,����Ư[PE��d�
0�3ڈ.�@�\/s	)\i��O��K�YYT�yb��q��k������缄޸�㦹��X�I�ӎ����t��M�ǌu�-Θv�|��=2��M����cHX�Z"y3O`h��[�6�ɿ~�]�mQ�����n�q�&������M��ٮ,��Y˔�mB���`|@:�&�B������e��r[�×7�j�Id��̡�B}C��D/͆`��������h5��L !/�0�@�@�W<ҽudϘ��22l�,d):pD��;�(�r���^}�lU�f}џ����箔+���Sh��XU� P��\��|�P!�*jMj�S7/ �*�k��+�
��W�"P!�l.�Ns���,7�t������d�n�W��y
�dի�����R�O\%q����e	T�����*z�&,�z�����O��� ]K'�\��NW0���R��Rv�D!���nī���fR$��0(WzQ@��X��:���-�ڝ��Q�lX����b� ���٢ϼ�:ȧ,h�Y�j
��_��j;>�f����O�����ep���&�� �Ma:Ǣ@��?�ջ?�M*U����_��O���C�I
<�dn�zo�Ɗ<��a��)�O��j��EN�H��Lq4�N�ƙ������)��DAit�#޹�raN�`A@�N-W��%)�fM>�_��D��f��{�A��Y��SR;=1�v���R�C-�q���`<(4CVD%x>��S�߿4�xN�,� �H݃B�H�;�jW>fp;.�o�
S�͆ZY�"JC���h:�{sVՑ�Dݯ��X��pҦQ��ا�3�>��h�܀;Α�b���a{e���X��|D���Q�|�iٴ�a�d�?����E-�$y�ϼ�
��{m�p6��urƫ�:�6)%�e��� Vl{�S	�C9��|��𦙇�����e��]�ԝ���X9����-y���;V��ډ���I���T�o��mfF�*��T�j�y?< X�Cx��n���x��p�4����cZ3��,��?�ry�5���o��� X������V��������=�{��F�2�+껖C��l�����#���P��o~�Z@B���ڦ��o0zP�4`����e�ȩxXV�dHGO5;=�է�~�Q�cBە��M��I��(�\Y�8W�ebI])=�D���`m�Fg<��x��:譁�8f�AC!J�u�r��KR�F�	��3����KIY���w�wW�3�5���`c�����ƴ�塄� J*�k�����YZF�0�c�<��`;��W�wo=��hv}<Bˎf�����ȑ!y ��z�5���\����eǗR�R<�����gPtBT�]��|�P=��I��í ��L��v�?w��뫏���q��'O���O�qGjmk��z.�-������XkY��iQ�sܝ �k��+���z���A��R-z1�7����衅���w2L$�73J�6�i��������Ջ�6��.8����ߣ`�||r�#,�����[�c➎���w��',�\HW���[rD�粰��M���`g��5�Gө��t����Q�ڽl�j�����~���E�S�}�c�QDvJ`.�-�R���D���L��@@���4ahʓ$`NKWo�Z�1�[��D �^O�!.�^��A*�,:�������M��������Ϣ��DÍ@i�+�ǿ�|F�|�W��\)鋥��B��E"��8ʶ5�K�+���EugFJ�v����cP��s	;�ý٩�d����F�� D���X**����E�x����!Wൟ��+�4�b��H�e�DevΟTN�^lY�L�u��[�@��Kt��Y�[�7�gP����~�����<R��NW��B�C��b������ƔC�]~ F���J�i��'w��DwV���_g���D���g�/Kj�f�N���s���	b�����������m���F�{\��;m��n��M#��,мAt�5N�q��^ӏ�T�G|k���c8V��b����i���a�J�e��B�aȕ{��\e��J8��T^9y�@�9���3�7ʮ.��_(X$�f��(9BșK��rh�%��k�hZ��������.@�z[�����L|bF"�az������QLj������0P�i��r^EX�qi�Ӝ��-=��U���q
��TM�D�Hd��n�8�^"�v�s��H����v��жW?���z"�5J^Z�*c̠����w�l��7CE�<!�����9��0ǁ��tO��+U�K�^���?�ok-*-?�+UY�FqRuȈ�Y�8��
,���cZ����ä�ɏ!���z�P�&W����b��[�~Y����W�}���Y��3�S��<�W� �K 9�P���N9<;#��	ȍ�b�:r���L���Z�UG�,'x�Fp<�v��ڲ��+��ϩ����Z����أD�-�R��cǚ���s�4�j���g]��E���J����}�
�$�>	G�'R�t�|@$;��~�eE.��Xb�-6("�����ˈC�1���R��`r��4oW�\��Wfd�2�|�bN� �ɷ/z��N]@UCE܍�V��p�he��V�!�s.�Aầ
���^P��%����n�o�CI<�'t�}��
�z+|�ks7�Jڅ6lh��K�5?V����|[��2W9˿8zj+�!x���d��_���&-��Z��9"�ޕu��L ��a^(6�}q�����uU��( �a�e���C��ABn��hI��
}�>'�Ftw�i@�o�އ����z�w��>�+N�>�+��1N��7nR�k�OR0����-ʄ��m��t�5���$?�V��Ǯ�����cP�q�ė'L�U�8�؍1|J�7�������ps�D�>O.���IgA �z��-���d�?�5$�l3i��%T���*O��fcH�����U8���]{��4ڐ�'Zڣ=�����pm�[���2�^vF��߮:�?hP�[[y�ˍ'�b��m"ɫ	Qfüӄڠ��60���q��Q�K�G��KӶ˻���uD���U}�C�wux��W&��jm����o���Ǝd{Ed�=�`�̹����b�� ����9]�H?lԉ�&5��!+�^t���*:��3��l��^}��V!�A�t��z�Ģ�ͳHRr�ߏ�O6�ؤ;���ſZ����ӋA���K�;Y|2I�.}�������n/�IM�V����� BV����^�0ܜY$O�N��ͅxc	��W���h�ԡf��>��_�־�2,���q�S�0���d���#3�>A	M�y>�oa��s��U��r�_�"��i��(++�+J)��m\��d�r~1��@��`��g�W��ǧ���`-�zUmv��I埰��;�Y|Q��0�:}�x�?;�]�)uBa}Y3�����P��d��&�w�+rBF}��I��Yк*?4����fC�ZT�+0 ��@�i:��2�5mr?��9\@b��#�dG�!M�	^�f�8�Ɍ�_���Y�\�%�׊�/�?%�C6�T�aN�2t�i��Α̶�}*Se-�>���j`­�l*�9����<[� 5K��Nƺ�8�>������P����h��E`�)Kh|u1D��U酊ֶ�]~����uX��dާgC`���1���V�p M�����^������4vҮ��+Ӆ��z�Z�i���݅��#���q����.���"��u�V ����p18E���x!��5�$�������B�EF��4�������J��)���(����щ��ý{Kxm���I�A��ԉ+SlfO����9�Ӄ���������~�*��=8�c��D�|�4lX�g0F����RT�2�g^5�o�|�jLB3�9T��F�����c��9<����8�R�ƅn)�a��7u� �v;x�$�W��*)���|����]\�����������"���Abl�C��D сW�͞���+���+
Q[�3�EI�ؙ>�>��[��B���&Ml��Tqֹ�i�'���������2n$_GԦt���*N��Ϟ�oZ�QRqA��͗#Ws�x��/_#Ԑ����
-~�|��� Fq'1O�d�)���{.��cr��Z�X���+�=��9鳧�h.�g`��@�PM�cbU��NHMw+��=��O`7��|g������wg�OE��*�sa��/ԟ����T,FR&�آ��d�P�{�&��3I��2�Pm�����<e50�1Z����O�9mQ�m�����d�VX!�oMR�}|S�|u�U�ϰ�Ɂx�+�k�<	�J�(�W5��T����oXqɁ�Ӑ3]� l��?�-	j�ՉmU����0r\3{V�x|���PΝ�m���W�È�m�@��R��j��𶉕Yo�r_D�:3��zo�� ����bL��}�� z@9ؓ�X�
�*F��YJ�1��u֔�v�*ɢD1�a����h]��~���	V�8��{�R��8�/!��t��[5(N����v�'�ko���?�G��S(�t�@G*@e��Y��񠳘#$�|������
�K���H�<���j<4� ��:��b��YhK�o<3n�3�H,�A�,OQ�E|9��x/M�R1�j_Y���.Km۽h0�d_�&�.�n���2��@����I�}\Y�8��(dH�����x����q��&o�^DEA\TA��jx��l/�L:*��;���w���/k��	�)( H�
�<Ka���_�*WRi�#�į)��B���� ��'r~�7��)�!ݝ̯u�*�ǈ-��/�>���P�~���t��5W��4H�`�M��.��L�@�Đ�����d��e��g=V���ܚJ���Wo�+�[��z��R�91����Bf�yh���;�_���t�LU<G��v��`ж ��N����zzX?��u�p���1�v�����<dC�XiY�[���"ɝ�N7x�~l��P���a�9�8����҅����e荞6���:l<-�[���M�_"�.,d$�d�i5�]�[��d
�[���0ҋ���<�����=�`��PMK'[�Q�5���jQ�P,�L��J|���=e�^���B�Yc~H���4ϛ'�;(N|�_8��t��#�ln��z�P�%5�{����*�Y��� �x�(X5g��l�FB0�`�G�Eo͈�x�6��ŅBA�KR��Xf~`'u�����>���JR1�̣��9��cQq��z��vBh%^�/�e��(�`�{���w"C�/�1.U�ŎR� 'T� ��{�)��<��4�	I�,��#�R�Y�8f�>�#��P~�4���s�Z
��L6�J�+>®i �;���F���KZ+n�[6f=5!&I����ܽ�a����I��f���d
*չ�3�oF�����{�N��Ot��*����h��'G��m�v:|e��Y];�׈"����2�z��VJ՟����b=1��3����q�~�&�Dˬx�_�	1��y��l�j��;�`b�m����"|	�l�5GWͩ�uT���$�H�J����W,]����x�l�&��_K���!�����TQ���M� � ���T��q�&�gE��ԩ8*����β��ռ���3����K�?�?���b�G4B��+�	�_<�]���S�
ѷ��O��x1}I��{ah޿�mʕ��@�v<2�|�d���>�Jǟ�/ϡ@fîM���6*	�#��Vt�;�殴9�bޙ2��Ze�d��-����ir<f��z/k��9�P�_��?*<���T��\�m�����[n�>� ��H<8�W7.�����N�*��� �2\= �����ٷݏ�Ǽ���j��O�e��%���NT��Nc�����GԚٵaR��4��������$~&�����`�hŲ�G��Ag揥�7����0K��/�s��Kb����1�S�^�73����0��[���R��T;�^�1Tp�@����$�=�%�~�8�HD�~�ܜ��<���f��}4�/\K�6)�����!=��Ql;���-�<�b�o�^��I��aف�`)��4{�)��	z_#K�2��C02��������?N �Cg��9;�Ys5m�\�"�E^���+�
�h�Ff[f\O�軌�Bk�H?�jD� >'Jq����^?��"�&Jݣ)jJ��q-�-��˩�ưv1�jXWE$�.�k�?�q,t�Ws��9xm�8/�{�y��0��7;�J� �h�B+�W������^��>��m��0�'e�}�h%��V#B\�q�9B9��2Rt��o�L�%^�c3P^#����<�9�%䙹�?Y���;�(�o*����`�m��)i�O����{>�S �<Y�J;p�wBkޫ�U:{�%;ٮW�܉�l���BpBG2����� 6���+�����h��ڝ��ƺ���-@��n�7m&sTN^�=��8�9�W?n{��`�U����&*�7a)��,�;tW������sp?��aX���ذ̣� ��Sd����'�a̋Y>Ü=D�6��d��\���\i��nA4l�'S���܉d�ͭ��e>E�<������iƍ�.�R�c�s�Z����d$y!��>:�Vj�٤���S�����NE��uXA�e��	gY������A����B rm�٘Y m_��~���������;��:���dDj8���)��.����o7mU!�s�������-����S�V� P̋��F�REWph9����Ɏ���* ܰ�e�Lէ��i-�-kߚ�_�X�e�R��bJ����g����aN��m�`�����͇b`��T4ggx�<g)��%c�_���Y�fT8��F�~��9[3	^��>�:<��f`�����
M0��ٞ��ߥV�O�����\-Ĉ'd��V�E�����)?WlLV�R����-@F=�ڪ<�_װ���A*�uMoX���}@@2�C��y��������
U��8��tP`V�E&T�m�䡿wF�S�(m��M���;ɼFl�9�G�$A�^������|�U	k{j~Nj�٬sq�6x�����I��)�._���y�.ի�IٰGX�|�D����ɲ��죥/���Vv'Ǖ�F����7I/�e��J=�݅���7[?Gc��{g����ku�ۨ���)8]�;c��"H�Ky���K!��CL�9K��J�U(�S��TV�0�̳`��4�ey01\Q�x�W01�1� �ӫ�)~ ��yJ���
��w-ɓ
�q��.�[�@:*}c���eh�D�m�p����T���S�no��.��"�,�ܮ��گ��)c\����映��~����P5x:
+ơ�Ht>M�SX�ud,..�W<�e� 1������;<����%���5�|b�~�?�8����/��
���9����|d��
U6o����D80��7+��ߖ'��te�ё%V^]y
�dWӽ���U���id�@(����`D��0N�l&S��E��`��~H�/�-�ѝ����6��D(���]lw8g��`_*�%1�\���VnKE�/_�ZI���P=b�i�L�}~g1�]��\
��Q�.�`�1�{L��΃;I�8� ��Vk4��p�|=s]M�3�P�⊹�<����b�|�v3��M;�e��>��s��y8���s�QGsU�k(~�1�&����/�z>��U��4�,X{��mH�ɺ6��_W.�M"QN�SL1�|n���~hq��������e���2�����R��jӾ��z��Ԫ�d3����n<�7��k���a��(���T��G5�	r��4x�\�Q�I4d�C�C�6if�%,�M�Qg���l�L?nڢ�O�B����)xn�`@�hF��yK��(t�5}��n���6��g�i��Zg��a��w��� q��2�t�.2[�;�������9
��Y��69{IOT�Mٖnv[�ͣ^�mē�bCK]�mz�T�
o�~]k���7o�.ҞM@�_i�Kw!�tG�����+p8�T��>�b:	j�g���#���YP/��'p���u�����$ƏBG	%W�5�%㋳߽j�z��c�����B6o6'��	Jn�^ E��2I8��uE�C�'�{}��'gQ$��
����C5\;�`�α7���/?#MI/~��HV©g�lW���L�B�����n�T�kz��;���ܶ��iA�<(��+�%�y�<'�����s�9@�_
,��MF�k�\�5�qCJ��R۸�y�cd��?��PPz3�m`�C	J�f �'H����Qza}��9A9�O��v�!4��+�J�<dwj�E�_�H���A-]v��Oa����6o2	_3�����8<��C�
1�/d�������C"�/�t��v�����ԃ�^�$�O�5��wpW&M�����A�T=*�<Z���@I:��"gZ��#���|�n9�M��L��H��T3�Ⱦ0�>���S���o��Bk�d�?`ц�e��ߒ�k{�Iy�b�D"8���f���!�T�2s�)�X��=<�$���d�e8�r�y���]�Y��;Ǹ�ډj��Z�)�������݊l��C�B�������	�����!�cDi� s����=fbe��W� �����m�d��%����f�����0Q&r�������4Č��/��n1��k��Wfo]�����JB�@���?����=���L�^�΅�p�ɻ����n�( �R��U�`0�Ⱥ�ȑ��qQ���g���Hp���\2C��v�&&��8�&�7��!w��í��L=;yb���Ԃ�/�B��<�L�à�e���U�e��v �A�L�Dg��Q�[G���Ag掂�"�0����y���3��q��������x�歴z�U/�
�G���	��km é}0���o�l��`���8<��ǚ��v����M$��{w�	�
���շJ�,�Ю�ЍE�y��*�uĬ�?B_&�4Ao�w�J�\�zݠ`�z�X�Cw�
�Yp�]��,�/wW$o�>���o�k;���J%W��Z4M&�O#��q-�J���;1��o��/<�d��oD(�Jo�om��MAH~{jC�54�o�ZNM���	%���!�C��s�뿧ec���`����#ka��q���f�1�������wc|�t�LU@�%s�3/P�R��1(���]��&��%-�6��O��*tE��"Q�F�:W�6�oT�`3Y7x�'��\qc@ *��B�(r�.��_��Z���}�R�[ɹ��&�~'y6)%Hh�^�	(�h�>z�1f}�]T���P��0�W�߫�����k
Z�y����4.�^�� :�M���*q-Uܹ���������ǣ��wЯ��Hy:��y~�{nFY�ˍ�F�D�} �?��i�Pv©�R����Lv/5Rg�{%q8�'��[���'l8�r�FzT�����{߰Y:�,���%͢$����)Lb�J% P�sf�7^tu���02 .�R��z�����+��M]�[��������v��o��(�8����e��X�@CIKB��W8{E�1tc� ��N����dڎz��Ӑk�6��&���u�aʵ��*��9fu��9�)�	L}3�R\"�$;)M����T��|	P��T�����%m�_�-e���C�9�=�b ��M(ʇ�_����`��w�Wr���n��T�$�3����<_�r݈��5�,�ݖ�Ǐ�?����yn� A`�\�~lC� �m��"�-�,Y�:����4��ٙO��`)�waM"��M��pl������*��Hcw�׶�J�k�&�|^_��?�i����k2���ib	#g�gs��H*�/�@����USƠ�^�dhF�>cK2`��P�����N��������,h�A}��]rN�DP7�Q
�֗9a��-����iÛ��f�@�@��>�&�W�Ȭ5
<C��4s 2�e˴���B��M�/;i�R�;P����1uQ;w��ݜ�JB�t<��"��SM#��V�a�]�_`�w�ߥA��xڽ�[繽�5P�9-`��I��_a'�xÜ���#��w_�@r=��\Ĺ��ɚ3�K���ޑ?y�N8�fW��!�Ys��>�&�)ж_����?��(lB�^/H��[,Ả����[��1Х?8)�1���':}2?�Ww�2r���L	c�Q���P��*V~ ��?.S5oΫ��O��'��]#`}ٛ^��gy{�@L��K�%4��fB�U��2������Hz�;�2=�����<zQ&���]��e_׎��L���צ�Qg��W�0Q����x��Wք����s(������S6���=���	��̎��wR��q�1��X�#f�\���O�~�/N�_H�ٓ����]ǰ�o=i�����0����Ǧ ��y�J0�U��z�ue-��F^�k�Nv<�6#U�G�A��Fz.s�\M�-s29` ��>����(�P���*�_���	/М»U,q���^�+��<���� �Zx��iCtT\�`h�>�w�f�G�0o�0?�c����=l��H8��l
QY}oS��v�KMCJ�b������˾�F�X`^�9P���X����^��U�=�����?!����-t��yG�%B��k�"ZBM�آ�V[MA`��V�����2l��{�x*��ho}��0��r����J޹L#ge_M蟶Q�A�x�o�G�:�{���|.�Uҭ�`��R���;�x�By0�lC��/v%|{��Z�im����P���Յ2�^�47/؎�|��MȪ�6�`��ޔf��y��$�	�hQd�� P,��p�eD=� s��o�O~�yتg������?ZJG��TY���B����
��ɺ�����d�o`u��?_'E���נ��}
+�2 ���������{�V��+���9nR���*,��}�³�t����Bujh�<!$|�Y̹nԂ����j$�_�!��0�sX5���s������� c�7���zsJ�K谚6Ԕ�n'/9�BI�K�Z���UΓ}k5f~"/� D,"��sc( ]����`�[�"a@ ���0T*<5!{�.3�e!��6�	mxAܿ�|[����(���2���g�r ���ȣ�����_=�kp��uR���y豝����{��m�ū̢�ȣ~��Z��'F�P�D�d �Q�p	�թ���{yE�Y!I�0Aɳ�![?1���XN{���
�2"��L]wt)`kB�Y�{��7>鏤��-�VG��Ά�'�%�[�n�<�C_B�CC;�O��U�f6e[���D|�Ru���mo�����Wƶ�.�v���5~�P�nz9�5��rR��tT�'=��@���<�guզ���[ѵ�%=My��Re����h�z _��<��,�'����Zڐ��i�u�ǿ����L3(:᝾ތPѼ�C@˳�[�1�]y?�t����F�����}����U�/("�vj ���7���Вj\���sWO��Dk`�~Q�q"К۪��P~�X��XZq�/�訮\� �l*@m�3.�d��&:k4�����@�m�B�;�D<�~�ソ��>���`x�J�w.���c;�_�)�b8;-�h��)&�\�WE��N�^�;T���3�0x��l����V���V�=+:������}�"~L���G}k���9�|��^s'��o�s��-�id�c��~l��Ir�f��$�m�����}�-E�����|0x#�������ߝl��Խ�+k}e�3%���e�] ^YM
G	Ok5��0ç�A[�c<t�Q�mBv�U�#���6�S�0��
�e�\KЎf`��ʬ����A���`E���5#�qս��2���pG�H��/Tw��p�*����wO]�ᰞ�	��N���J!r����|絃`1P�z(Z����!��	� S`{��m� ���u�D�|��s#f�}�����ƚM(��R�*��x�Մ��"v,�ƻ�����ª��c�M�������_�L"�m�߄��Qny�S�@Df�� 8F݀�����ݱ��c]�cP�3yޅ
ި�&��~3惙@��	�N���sϷ9'R��!�T�$�ҁDw�����T�M��d�5J��?)n���~A �� օ��j��W�b�;{��N�S)��}M�57�9p�G�*m�ڢ��N�d��({����7���������^��vT���qF��Ƽ/��;��?-y�#�xw�!ٷP]h{���9����^EiA~���4���u�f�K[��4�����uZ�io�/#�+�<��P[
f��HE���겱ʹ�8S����~�� kx�� ��ɾq0P+;�zq^����r��*ĩ�Ȗ�۔�/"�����~��P�s�Ģz�]�S66#q��N�e�%�D�V���gG��?�k�O�q�����O��R����M%�^��I�q���
�e���De�vv|�n�����;�$�=�L�W(�E$��i��w��G)Z�����G���񒇌�vo�>គ��,��8�'�u�n٦M�i����gZ$F5d״��jc���D�R�s����=t��jP�L&�o���V��������3�+5\��NR��ڹG�*�ґp�;����J�#��P��ʹ:�L˻�}��x@�^\��:���p�y�R�:� 8F���;TᢧA4c��TG[�m�h&��jF�"�Ą���>>[}!�nߪT��\�2�+�`d����'�W[�az*�b��6?����l�� ��.��m o<���}7	_wZ��Jb��X:����R �v��>�6w4�J'Mz}��Y�Y�c]J�`t�s ��c�G�η|�h{�¼�4"��Q@��o�ƵFJ���v,%\�t����[5��Üğ�B���Ԡ�|)��řh�LQ�.6���{��nC�̡��Ť�}���^�3F�F��D3��;g���6���gHԨ���1GH�d)`{W� ��^�ٞ�7jԄ�%�!� �$C���b�\�+�V^B����=�9vU
�� �V�����++��,�w󮏈�l�Ch��ޱ펜@6a��<|�#�'��3���z2��|%8��� MJ����cr��Ze�A�r1�ˆB��J��R�Ó�L�y�§�/)���]���wTvC<���+��FN^��όY@�{�����?�m�~��,�-��+�4L��O=S�����k)ݟ��ɵ �hɘ�C��P;��mn��6&D������^�~u�9��2�$�Z���ܝ��J(�;(�b�Gk��Yo�t��@���DЭł�%�z�ʮH}î��O�i���~ާă� 5g������e�*��:Ш�_9�����PV@{<q\%h�((+��ղ�rD'7�L4�"~=У�;,����/|f~Ů$(�ޓ��*Z�z>*{��;��s�)��c�x��� �CR�z�r�� ��͗��|Y*J�x���Դ m�(�4?����������J�C@�.i�\�A���s9f�k����/}�1������Tuj�K��N։)�~���9#8�(-�gյ�a8�:����ۂ��Y�H�A>��	������P�"��<w�i�1��e��R=ҩ'�FS�o��O4�qZ���y�����WL^�Mg��3&��j�ʜ)7����Iީe�L?g���^�Ґ��r��giR羵"����i����M��������ⳙ����5�H.�}w���-q��m��H$4e���.�/���;��C�>a�m�T��u3[�5���+��20�Ml�z�������z��z�������.\\�^��^���T�tv����$��u���_U�а�3���<���5����".��[�u��?�4H1,W�v�6�K^;_�g=�Υ#��)+wܟf�11~�K�	|�Ǭm�*��8f�zn��Ŭ�?vy�4����� ����O6?ro)��$�u��@ ��H�^�s,T��k��~|N���5I�ENfN/���z>5(��OwB�TU���D"��Z&Y�ڡ���xV-��jq��_*����0�,E)"�g���Y�q7��o��rTGM�E�V|\Ȉ�Pr �x�D�_��c�t�(�z�KMrZ����Du�+�����F�|Á5���s�5��)�g�)e�<t��NKY_�9:8t����΍̷�IQsebs�?җ�C����N%F�{��0'u�SY�	f�L[W�>tp�}"	J���w~{�HMgB����1�Vu4�%�N��	t{ �O�x��.?��:KP/6�\~�L�5]�5����-AZ�7�g3��g�N���1�/��[�[q��!��='�*g<y%#���{�;�_�z�s�:jx슇��J}ݧ�'
0�=ߒm�)$Np����l�0M��O�)��(�����6���t�ab���4�kG/������p����+oGe��iKI�$Q���s<ϽQ,�n��䤪6ƅ��������7y ��/��fԜ���.:�? ��G�x�N	�u����xb�CD���U��n��g�	i�~Φ����g����m��B�Y@���C��3�ï|���!t$C�ȸ_�#,/����6{	�c�w�P�1��=��S3^[�)�
�v'�q_|��S����}L˄7�S�'BS	��C<5�d7�g������+��ߴ��
�"���,�I�l��ƛ^Õ2T+|�1������덵l��jWK+����I�SP�zկoh��������$��Gr*7J F$!p!׭?|��l�L��Ⱥ�,,��.���|+"2x��,�v?���?k;A"�`����>u��HU7�}�9C��oɳ ƌ��j�u�������3Q��|+�)ӂ�v~����PK��x��Zo(�L*��Yu)��A���[^,Z��_*��G�AH����|�5^�Uq��k_�!�7�n58�����F5�K�����F"�ھ�S'�q� w�bri*u5ƌ}ӑ��5�B��/k��p��V���5�*�t��8�>%���`���Z��z����U��~5�	24uz��J�"W{*���v�ɯ���<ׁ$�D1�\��╼qG�=�<_o �>�2E����3|��|�H8�dn�s��sJ��Zj|�:��D�g��PcT�:O�h�'f6 @�z��8��s�9Ǩ]�w3  7�#��s&�C�e�fIs�J�0�&���K�	O��-�X�L��S�A���^-1.&�9�r�m�j��p���T�U�o��	�BoJ�q��
}��J��Ȑ*(v��~�7>���.�T;d��:�0�?J�̋I�;\����g�d@�NZ�=%|��0;���ћJD'�c����A������$.I��[���@&G8QTE���"ݰg�d������ 7(�JJ��Y:���+��}��pB�� �����fN�n>�O�`���g�H�U(-���U�&K8b���u��F8����4��&3vd�& ^E�DIRg���}���J�������I��C��PD�앗4�Ss���"4߯�O#ٹ$K��Re����y���ϛ����]dqJC�qQR���ծ�l�����Z35���w�����e�Op�CR5L.Ni"�0���g�"��tW[�A���8w`�#�k���q��}�?J���'K�ӣD��x�A�%RA�h�m���_��n-��F:�ѩ ̺�ve�o28�j�ՠ�LIrS+�C�wؼ3�A�"2��Em̸E����f5C�v`T���������tߟ~6x��BS�s���Kd �!��;P~�#��kv�ƻ,�=ㇳf`�`�ˌ�ͱ��Mf}�)1'>d�Lir�^��i��m\�	��=n5�K�2`ɛ{-�1�xI2a��|�
y(���hi�,ՌGM|RH�,Q���6I�h#�2G�<b�)s�'��bgGW�W� �5�V!�VS�f_�r0w1p��C��ϡJ�3m�8vH�g�,�X�i��]-��W=�k�g���ɤ��
/~9�s�R�hvW[����]{�<	!�I�����p��m/�S�,%ܪ����A�����DF�m:|��Q��%o����#�6��P7�	�k%q�#�6���^s_O��=�o�s�j��;H�}֤׿��U���j���H<�\b����?"��QlQ[���37����t�����o���I}�77��W7-�����wu�@!�J�{
�5{�v��PsS��Pp���|n�ք<��γq	��FW&$>�maը�}�6����MF�#�������vA���S�ʨ���`%V �cP�(�X��O+ K_��p�|¶�a�)I��Zp��h�.������F��rf��J��������^�6�e��F�k��q�@r � ��xz��N������0�$��Ց7��t�ip|��P>@�x�;&��S���Z�;Z��;����.y!��r��1/�v��{��v��h/'�̅���;����
z��Ҟ镪`�a-�&��9^P��������z���sI��)��h��\ϊ�2�4�G]�B(5g�ru���}Y��dי��r��$��z���,¨��%Y�~�K�ҭ�B���fH��!d�d�Q�k��ِm��$O��芢�|��^��o�s����Xa_'Mٝx��C^�^���{���\�.)��p���G潮Ei��֧��!ʒOC�����d���ڋ�J�ǒ�<���
1�G,���ZbDo�BR�JQ�3̑+vڶ 	���R��)�-�K8�MX��W��@�;	>��)cxdU�H񌛈�}ϥF�����e��m�(9����	��q͘v�A �F�$,"o&���$�a���ժ{�D{P,��+�c�9Po�ĕ�v��ʤ��	�e�CK\1�։�s�t�������D��>8}y\�>T^�o8%���X�@ڰ�E��yȿ�~?�6)��jLf�r���(��e^�/ay拢����ّ��O+�z=�!_ǣ��MGN�oS���Բ'V��e
��C��s��V�B=�~��o���GQ`_]oq�Oh�l���C�B�& ���M��f,�,��0-gt�.1`,�Y:�i�P,t��nRuv��Y���4u��Uܡ���М@��=��1�(�X�8�����u�Uk	���%�m֚�z��L��(�Z��R^	r�x���H������3?w^�3�>��}y�P�#����\w�(�/���Rz2�-QX���$�]�z<��10�70�&��ޮ�!j��2����D�eݳ�9~ JT�Ƅ��X�]4����T[��*�Tu���Rz��,��Xk��F�|���C��ǖ���:�N4�K���;�m��t	�4��#:�?�4w���\Ԧ�?Z���:J�2V1�Tݿ�p����Ѣ����
q~
��F����#5��eB�6����P}3�b۴=V�u>�VӬJf�f^�ٕ�15��)#�&|�o���{�q9�q����5�zc':�n���xh��(���eIQ�u���C�sŇ��S��}j�d�������W���񏠃C�GìU��ӌ��5�WG��o�a��MЏ�˞���J�^h�V��w�R��U��QuՌ�' �RM�J��ė<�~sݨE�0��
5Y�{^Su��UI#qA���`Z�\����\M��{��H�bo�3E�{����ɧ���uP*�y����C���B��K3�^_������1�zRrͦ��`K*[��25P�,�qu�/ ��ᴆh/��O&�%�����!�o�c�"����$����	&A"R���Xұ��䙱�%5Ob�$��մ����(�z�4a�-%|Ek׌���z=��++M��,��,u�b���yb��֞X��/�~L�<ƞ�F��7�y���U���I!"-�gG��\�tCX�F�w| ��ϘO ����卜�'���U5;��3��D%���)��b��vOQ���x��%�����`a�t�������M�X]��z�a�}���U��-����o���������7?}��M�����2da��~�4���H�@i�Vy�]0��`���}4F�[:c�|*�$�0Y�r��c�U�G�7�������ϯϻ����y3X��"��B�j�i�y#<����~*��_�e�l��!�J�'O?D!�7*��		�	8��b(I(����8ߓ����;�h����a��d���ҷ�H�JЇ�un��� �L���B���.ͱ��9�8O�9�I�%X^D�j�������7��	�J�̢�:���ֈ�/跊6y����S$IC}�L�t"嫺�6��A`�9
-��WE���I��ٺ*Oa$ʡ�5�U�/2�������>�ځy�&3SgY~T
�����k1�+���K�]r��-��3��1>��z�k�V�H��m*�e�x���h������b�f�W.����1#:��ݺ$7K��_��?K�EXǈm�\��/�T�(�M#����Ch�IA�fo�(��V�H�P0�-]x2Y=�	˶��}�}L�Gp����-�l���������y=�|L�9��c�ĺ�$d��dv���t3�f]Zfq�N)E��8~���9�Nd�à�9��F,A��2JS˛��W�v54��cזd��7xn�� ����>���?P�1����&	�o�[��߫T�_�FPLץDǲ�)i���K�	�EJ�։��;!��Ĥ��I��8L)e[��۷����V�����.=⛯�ht+��V\���P
�<�/��7D�1��-k ��M���F���6� �5E��]��M.�e� �V�E�={'+��A���!G���SJ�)���F̓.!^�Z� a���h
�Ӊ&�:d�4��Ew�Lt_<��{F�SH�+#e���t+ҠL4\q;� ��m[@r�*��A�'3����x�=��~��`W�����pm��Pۣ�̑����>*m�6=�'-���7s3v9�_�<�Pe8�?�m.��Sq�V�v�J���Bj�W�l\/`<��vQ�����fRA����h���݊�78��{�̛"��\�S&����� ?��ӆ�X ������ρ�K��ϓ:�o"��X��c�*� �M�..l�X�7�/�A_J�9D���A��n�6xh&��)���(���F X��� �U�/�������檁�x	�swb
��ۓ�z,T���b�I����a������}��"��n����S4���t���u��P���2_8E�[���h�����Ɵx4��a��%��hL����%���h�>�w[�M��U۷P	�y�����NIE9< O`�����c0�cm��ܶE(�މ��ԩ�#Ҕ�r$z�V=/a���2[@����w�ds�ͻ�"W?5�ib��L�5?��y�6�SO�(=�Z���=��r�,*�6Is-�|��_��?�TuA�?��L�7�|���9Ei�X�Q_�ѷ>�"+YVJm��VkV\��G)[�)��Yӥ��6m�Q���hz��Bv������\=��x[�F.Utp��'�dl��Vx�З�<39�th�����O>�+y7�����	��$�JH0��-�{��܆�8�>ih��W~�s�~ YC�e*	�ׇ�e�]w���t'�wޘ�AI��2U�N��?~�R���J�Ȣ���@G�@�짐Y�R��-T�� ����ϙ�\�\}�����ؾ" �Z�����b�gZ�I���0j�����9K��ץ��r9� l���b���6�Ɍ���'/�<�h� �Z:�������!13扁G��2����~9W7Ƽ�C'�,�8F"��٣+8M�7���6 �&�����$�ew�9��~�Ϧ�R5eK�Ԓ���I��&�ow|N�[5�G�s0ʈ|am�u!�2�H��x  ���?
X�R�S���*Y�u�4�Wދ�ݍ�:q���a��W|H���dq��"��9�,ך@?��&I]j�Y�\�^z��DZ���h	���0��an%@�ʧ[��{sv��5�c�9_���q��~'ӊ\>J���8��~ :iX=kA�Z/��giH��EW�{�u�B;�UE]?��"�����S@6&��>�1؀����f�.����r�{)�SK܃�D^���c�G � {[e��g�(ѽE�S�1�������x�OmH��
a/H)J�'�(I�������}��	V�{�AZ�{
����}�q�d�k��I�"ߎ����u�_�����e �k������:�a�m���rH$ճL�[a$�-�S�29|�@i�r�A �R@x�1D�R�w�͟�%�S���n�<1�@�V��8�ߕ��L��NY&�!��%-�]�;H������gB�K|7�uV�����F_|�,��E/v��]�Z�:NE7I����P .O����4Y���B��&�
䘫Д9��E��S����%~��5����8uSN�_�O��Kwn��I��S�.>͏p�b�h7;ʂ�rӚ��|�Џ�S°���7Ӭ����{żU�4��+ʾ��g����_]ix�]�t"z��å��h4�{�Ӟ�S��FR���L��\pˣ�􅮌?"ן�^��uw����i�px���A�*� �r�*Ui�!
:�$�9�l����m\�p�S�FHJD̎z��>���|\d���C԰��ȅ.���j&0��EO�&�������L��v'G#(�;LndRC������˃��]hN�pV�-�|{!���BE��2I�* ��q(�F��W�����sZ͸�"Ԉ�^z�bI�;��_bO���k-ޏ��1޶@�����P�U��tp&%����T�l
^��u�����Ɗ�b�3	9�+e%$���I�2N��rU�>O��"e�[��1aV��K\ZFp�H�������E�MF��/�C�²;�g��N������!�Nb��Y|���}G��7�����B(�:P�����<D��~cVU�m5LS�"�Q��=�����U>������,A�Qcm�q�l���_���Q�zPid<�:��}5�z"B�	[�G)h�Z8�٤��z��8�C����]�͔�;�F�ϗ'	w�1��i*Kx?sa�@ʺ��Vi�1��b�A\J���˨ג����S[���Jc�r9�Z�:M��Pmd����1�A� :���l�^�t�����h���E�jA�F�%-'�7���'^�{�'W�`�C[�}�5�9�E��gW\��*ڳ�%�ԛ�.*#�M���#.�rtnؘ`r�yOP��`�[����d[ 6�uC�K1PW���q�����,�rs�����s��`��*SiJ��@��y� F�:T�hi����*<�p���E��NP.:��6�f��3o����	t�A��� R������qE{����;_C@|�X5?TWej���賤='��CY�i�֫Z.�^��~g�k�7l���#�����Z�ѳ��'	����Ӽ�q����@�|g^�⺲�7�m����H�F�ϝ�E:� ���a�x,&�&��e�r��y�p����:c�� ��K�?-��'��O����+�a��qp�\�t�� ��0pzJR�%nj�-�}E�_�"V8�$2����
δĽ����D�8�v͐�\ �a�]$w׮��/K������4�E=�X�d]k��p�*BP,i�ߟ�?B�4h�
��ޱZ�)��Y ��ڌǀ��%%�B��+k� ����!��4D�%�ĺ�׀�/�vD�eg
�\�P8����EҕQ�� e�a�O/GRH!]��%��|����:|���};<DH<A�zh�/E�oޅ�}N$O਱�t��O����x��o��y!Qiv�
��'/&��e�SYh��b7b=��t�������b���Iu"L�q��<�VP%ea5�J��dv��yOo��A;C��Ѩ�%������h�'>���ǧ��[t�كmk�ύ�����;���Cz��"j,'�]"J��e���t�梞��&�+�ɟ��i�F���(�"@l�%�>��.�u�lh��K���R�Q�����G6N�<O��ٰ���#��c��"��J��{v��o��k�ͬ��m���g!�^�C�T��32z8=_�w���S��X�rw,�S:���\�ڛ`�^@�i͇*�E���-��n�� N�*�ӮGM�� x�;\h�I]��)/�Ķ��l����ruD�MHf1̑��׏��N�`"3XbJ��ݨO1ʞ�b�y�<p��NB��[�S���Mi��~��Z���1�\�m�����e�zܰ .>�
�́�4���Pb����7��hݚ�>hX�9���S���������;@�\T/8Ͳoj�<Pl�2�kq��Ň*JlįLڍ�rM8E�;�ZQҁoO��FS'�;m��p��������e�j�+��Q��U�D��n�m>3�y{���.&�	:U�[Z��G1�����='�_y���1U�����R�G�2�g%�|���o5� ��)
#�U���E���,��xy���)���{LgP�~�Z������Kڴw�ֻ�<u�����tD%��(w�I��Y���I�'��!lWe�5(Y�X�e�7�h��Y��`Z�+�c*�xQ���;q������ҫ��ܸ9hT+\��w��>�S�M�q:e���^Hrakv��`am-��6�=���rY��g3���&I��^׹�����::�E�c*wXX�y!�e#q׊
Fym��,`�d��0TMt.��Y>?�x,�@ZS�o�� ��m�!�!Syʸ,!~b������T�n�1�sg����� ��	j���B�c� ;!�r�Xj�)[`7T�)*����J�)_@ׄ���7����EN�;JǕmf��]�e^V��o�o�oJ��f���1D�{T����!9rc�?G��n������^��H:p=��Y�$<�7��~P���z����-� �]�嗒�S=׮!8'�VO�1�ֹ�%��c���Zi����pp�_�D���'U Xk��}�ɂy��N R�	�ؗ���`L�-hr:���P�����c~�gN�#P��.\��m.A�9�J��9��P��nBB���Y��Ǳ8���u ��Z�r����?���u*5[K�F�
[���#]������0���XeƧ�	�v�#�{�a��Y�^�V��<��\��M�}��+e�I�%��g����~�d��s�M�jo�q�v�~�*���8l��
�[��z{C�@R��VM4�"��7$�ࠠ=ӈ��E�7Gs��) �Ζb�o����$�]����1��\q�UM+x��q��j}8��*�^��s�t�ok���mO(h��σ�f��z��h�����1v�ژ@��E��mE�Cni> ���U,��7�Z:+3\��,M�ɤ�}Cs�:tĹ�Sp}�n��}��HJ*�QC���j#a¨yOFo=���(�y�SkV�,��|�|� P)O�o�t#��HM=�K�~����������'��K�zz�2	Ҳ����H�̴(��cSHTҨB��8��or� �ƀFʤ�'�9�S��y!��Ds>sZ��U�B=	�g����� 18���hM$\�I���;B�B?a-������67,�,��Y2��b�ྋ4?��!)^�r\S�>F��ѐM�nk���H{���w��L��e�gA�!�)�ۇN�"�|�����A�L1�����Z��~�׌���큣����%Z�5�?���e�K!Okh)��M�����!�>�]g�n�g�~�
��iǐ���U�
�����ت׎Ϫӥ2.תnB�J+�FrOUR���M]�쩷��%���}-S�IP�P�<�Y�8�1��d>�o�{|n%d�z��i�c���s�#��)x��2P��<��7*k�a<�-���F��ȔӖ����'�f|�\M!�pv��{#K���yk�V.���+(�|l��Ӣ�S�l���A��#��`Н�5�>⁠M���ua�ݮG�p�S����(u�t�9HE���ALN��~�'c0>3D���EOy?g�9#fg�D�L!�\��?��1���Fc1���/3����.#>�m��Q;�f%�!��y����(����-=�.
TѲ�M�I�֍/�EDb���R~�4�8���&M0��4�&�V�i�8^���C�y||,%��y��"�1��p�Q��������qYӶ�� �=�An�
��Aw����jj����,p����]<1v��r�n}dF���Bh��F�����0Br����^��!Q��j��2!�(g�j18�և̧h[�����3�P_w6��}��uW��d�>1X��|Q.�+�|~��1F�'���x�+$2V��3�u�O�y�s;��p9��Fg���)÷{��DOek���ϊ�t	9��in!�Eq��>E��2�pEE�����~��v
�0!�*Хp�����v�h��K�$1v$��_���j�Bz�?@Љ�_�?��{+e��P>a�����5`��{�K�NE0�ڍ�~X	�����?tʯ���p�|��{�*�>LX�x��Y�2�R4^�V�!Ё�'F��)W�9x�f���.5�I�#{U3t�b$6�62۷�a�~��#m��(y!N|c�-mO �f92�}�~�K]Ш�&D���-ѹ*"����VfH'����R����y���^�⊓�е	��oR+�T��n%֫�@��L=�Վ���^kkS�I�q�:9�F���η	�'Y�8�(��*8f.��t���s*1��k&�\ �N�R���4p�v�����"������j���@���X�u��<�!��ߒ (49G�/Y�[Y9.�u?3��m6<H_<� �U�Y�9t�d~ ÷�wwa�z,L�[^{���;�f��n=�Š���x4�:{r<��
����B,�X�t�"P\�o�xVkL4���i�z��tZ�=��'6ҭ����Qw_�!4�FDX�|��D�V򏎛�"�:[\������<�?�F���U6���(|�y�{���h��m�{�ie��_X��K>s��Y��&�������k�EM�;Q	�v���k ��2-g��1؍`���QX�Z"p�9�S7]�YS-�����@Z(ʝw��Y ��@���Lsl����E�wlYh���zS���N��)B%p$h<Sc��þ�3��2�j�ěe�<dR���J{f��]��ɕ�b-b�'h������n�+����USE��Ě�A/{?�ǃ�PA�,�JtjW�V!?΅�>��*�ԑ|��/f�_U,�����zgVi������\J�YX�u�֓�Yq.m�{=��6�y�����RG���eca�9yI�̑Dl��̝(��u���{�Ѵs$6��v*�ʁ�N?��]w�r��,t��uvo����)lsz*����?���d�b��Ms���S�$�쉣u�A<��y+� *�P-�`]�5�T淸QuÉ>GVBSoG�I9�׊�7�C�����;s%Ri��@&K���.���\��<�6�H�9����%�>�:._�;S
c�٬�򉵄_��O�֭� ��㻅�V`���7!��&B��Ra�Y�5:�;��S՘�C���/��zc�5d�1�����5U?�&���cƟj+�t��az�^5�-rn�%���'��-�]��]7����=ݭρ9��͒��g�6y�M����0���bȖ���A%��jnr]��.`��G�wd�b�Y��5��v���f6�Z��s�cl��g�i&.���HV��K�V[0�r�5���&�s(�o�0�nQ�i�%�@g��_���V:�����|�vp� L�[;|ئ��� m"�LՈ�ʅ�Y�� �;��b!Tf���KX�H?v�w ��ϼ��O��Ѡ��\H�̔�����6,���:z��g��:Trc�����@�g�S���j�[���?�8A�k��-�HnG�/��^b�n��fG�������I97�mT3����$;���w^��/Z��&���Ξ?-��C��e�[�a*�+��mQbUͮq��\���Z����d0�$�� �X����ڂj�ySs��&�U�#������̇�p�u~�d��IO�3<��)�{Oxq.��yH��"D����[Bf.��A
�޹���X��##P- bsnw�{w���T�k�w��.�̻�?z;��Je��}���Υ${���,�	v�[_E���ֶ��[n��`�c�jv7��!w`���8c=9���v7��Na��)(�({`8��n�RJSs<�yX7}B&*a��j��!�RC �+����F�,�.�+�=�{��=1)A�2I�i`���������\�j��P�&-e�w��Д��Ƿ��x"5�>$:y�#F�~7���B�x{]�z��%y��;G�(6?c��"@x�w�=��9#��RSc4\D��r����������&��T'��[�GA@#��x$_
���w�L���T��n>�`ɋ⭯v�"�y�k���
��k�g%�����Ӓ3"=P��]��Y�����!Ʈ�8rV�e�ņ�[{<1�{_��$��NA,_�����gG�L��%��K�H��BZZ��ҕm��x*���ap���[�f��\�+y�u�H,XL� o�_�;���'�(ʫ�H�'�6
�&~wtR�ֈ���=^fV��ּ7��Rw�ǝ8�*'׋�"�b�ΟT�eP�)�{��P7�g����G���4C�VZ3��!��'G�%]τt?fQ��ņ}<����ow!�`�[��q�0�,���妎^�~��d��GE�	�j�cI��Nܩ>��s<���a�be��dj�F�g!6i�a�t~�#�&H�ʖe�̸���D!������.�a�"�؜h��#M���U
��W8���b�ͻ1R��F����g(E8]�1�bs+~��hF�8�W��@x��u]2��� ҩ���4RcO����]����ˮ7f��MG�ym����'���l�P��3\ٙm���'߂���ɦ���4E���(���6�~�O�(M�A��K�Xj��Es��M����k���������
�W�Q�"2�x�RSk����c��a���?0怫#��t@0��+u?e�)!odm��85![�F�+�#Ѩ:V4� �ͤ�w��NT@Q��b!��M:��7������'|u>� >P��o�g4x&��	���u���4�: (/��k���4�6����Tz�6��c���
,���=�ǵ��n�P6��E��vq^����(u�[�{l��?���G`��m��XXmC* ��*m�iE�����|E�'ܡ\	G�rr�t�.Y1B?&`����,й�ʴ�%�6�y�'�Ta��UW�����?�V���a��͛���B a6f�{cXS�-6�]����ʜ��"NR�,�K��o<���S�Š�DjWXӤ-�o��z�W���C���ӪX��0��Y���ݙ���ҥ�ݐOʰW\�I�%*^��
]lw���G�U+,���o!����8�A�;���U�+�bm�0��a��>ڢ߸�#��s���g	��������y�7+E�����^��3�/l�;ڪd_$�(՟��쁤��a&w�2���{*Ű�&�i�YL�U���>,޺V����<p�
#a|`�vXu�\����~�Շ����f:����_�y#&i)��4�B�^�ݵcĈ�yhK����񨪘%UC��t�P��*?#KJ\�6�ް����B�w%�D�gB����\)������v���Ϗ��"�F!�xB��g<I�-�1@�QL={�<�b���n���p�';	9�itZ�w�?��&�[��`����9@(�8�i�X�I����(�P�����$:I�c&^9=�A79�J|��f�O�J0$�o
���/u7��,��l5�����ŬoGGq��dG�Ӊ}�	��oPI��§MtK�MX3����K��ʨu�3JJ�	~2~y1��h
؛ڏ�^�C�J�Ub�}��Zg���_B��no��ص�4�:�.#�.��U�-�l[y fH6����k�@6�Z���OZ=�,���wu*˲�S�IH?�K�*�4�QB�j5pl1⑿cW{�r��K�s� ��ͽ���Zj��#P>\N�9ǶM�o�Ӆ��/��BWIbU'�j�9���G�5��Y�z�N�ۄ�ߎNrn@��Դ4���a`��F�ۍ���l�Iݭ5ߛ�+��4�V1�Jܭ��U����߱SWe��~�Ь�"� �o_��:�i5�N�
wH�����Q��}b�A8�ȇ�B8;�LR;��� �,�E����­����� ��yc�VY�st �|�K����_�.H��էb�R���'����?&��=�� {�;%Z�#��PB��x�Ͼx����+mp�iKK�n��l��B#�����������X�\+W��gH&c�Q]R+.G!�r����\�mTL�N�랟��Fr�:.#�fҾ�	��aS�h��n@�͹D����b:�O�M�N�`��������[�vY�i���&h8 �"�1bp�#�o��|n3�g��Ŋp���( �D7䟷4�4G�qY���@;`j���ǳ֓	xG�X��e�ԧ��h�ʍ����"�u��Y���U�Q��&�[�iñ��1�k�!�I%���e�/)�6U�s��:�o�����:��v�j�k3��B�����x�CBB�m�ls��fM�t����T�4���4�(�
���������ƚ��q=��;�s>Q�#S���ʈ�kg�ؘC7P"�#U����y
c|U8*�Qn�g��/;����[~Q��6G �����M(�4�{*X����yW@|������h����5
��R&�s�[q�ʒ�3�ͷq�@�*!�&��Y>�b��)ď��ڪZ�Jd��u?�$���?Fv�-զMll��)�R�M���H}0�T՚�EnG�4f��]�����Mr�
C�ڴ]g*�ꨋ�mѢ,�@a��u�0�'L 2�&Y<G�h���̠�/)��ܔ�V�O&�����#���4󸍩�N�x��^76v.'ڽ�̤a������}Ρ� ������}h:86��g��{�mA�4�6�����{���Ԕ~1����_�k*P�ƷB60���r	�"f�jY�3݆E��t��3~��KjR�x���i60hu������s�I=���&�3�{����2�b�9ڞ�&0�� ��ȀW�߼��J"�U�K���7T��A�`��:��z�J_�W��$M�,5�U��%'P�`;����h�K%��mlt1���芝�ﬃFll�q����K��� <ئ��"X�*0\��U�#�-94Bߋ��GNbǘyH�H%�JZ����~Y��� 7XKm�&J_/�<�X1+'<�ǽ�"�`�E2`V9�A�e3D��w��1pI��R��p)��Ag�qx	Ҭ���g�1|rE��#Ț�RoFX��o,�%(Kܯ���}���u��^�H�^��L&�4I��UK�"����	��΍��5�Cx����*�!�N�_�
��:D,Q����;�Lx��V�92w�¦�W�$���q˖r��[2E��:ڞ�D��!�;�͝�bݾІM�.�sC>�� ���7��
w��he|�.��퓀7�M���|�*��S]�và�|X�L�N1:$_C��:qނ_�Ӛ��-�pQ�10irB����ԥ]��K�(�񲛈}���َa��J��xO��z���|r4�?��Cƭ�)���D^���_���-c�e�𥝶F�͓��YX�l2�����'21��f�-��q+&�N��#@a���)���$�_�B �#�y�ܯ�:���Nm{�KH�z�.����+EǠ�k1P�t�aP�~�e��
��ڳ���^{÷��&zJu��,�݃���������`*�y>�f�̮����b&'�����.ݼ�n"(�(���|���͹�!,���0���|�[
"4��X�aA���V�kَTӸ���K�Ҩ�����o����^������7��k�*���[��լ�׺�\���c�A��g�+}E�4-��$Ay%[Qg�Tw�%��]�
N"�p�q�[�^Ċ�6Ȟ�Lv���ҏͅ{��Xov,�e��yzcYZ%���n����љ� |߾�Qc�ǝ����X�p���e��#�|��i�$J�+II����3�h~���d�d1ߺ󋹄C�b��X�L�c�S9�[�k�@BK��^��u��,C�3x�E���̘���r��' q��r�-�C�z�y��ͥ��"��X�U��U$��Ȍ�fxf�T�BlI��ho�P�E��"`Rr��:@ �kk��b��l,~<��%I���0I!ہ}g	p�׸�pL�e蜼Q�Y��)�BQ�ɣ�-n�wuBl�8��؀m9+��i�zʞ��bP#�N!�)�J���׈�[0���_=�r!۽���(�VD�� $��n��wBio3�T���`�!d�Ϯ�P���P����J�(Y����N�����CrB,U
Ͻ�LVL����V��h%�:j�ۿ�Ot�f�(d�eP�.X]��3ɋ�U�gv͡��WZ^�SD�A� A���H�gEf)�X��7Uu8EP󕔍{�O�lF�<gW�����C��>^���l��HFqǜ�%�ɵ�i��	&�.�=�k��dK�$��tiή�Ƽ�Φx�~8Y��*}�
${����l�����	D�����H�d��5��9(*d��B�2#q^U�|���� ��;;;5��n�V�"�-��7�R�����)��՛����������p�}��&�yL���������Z�t|�>���㿤6��O9���
��旐Cz|��v�,�~U3�� �a���L~ �/�V���e���Z�w�k)k��ĈϢf��F3�.����zfgHº}	��Ճ�鞃�S�fa��p�4�/\>��1.pN��H�]��]yL��l�l:��S��$�֗��a6	}��lɳ@r�	.�����&�8#�͟4�������9��C	H|���j���
��vg)��R���#?��SD����'�Ѣ�5z��s��� 9EYC�2��w��[P����P��J�0�\�������9 ��9��"Xq�$�/m��T�
=yZ����Qs;�׮���qkʧ0q�-͎@sp�Z-�����A��%����Qӄ� [�h��s���pay-$fJ��7��_\c�B��G�t�r?���A���+��C1�n1І�Qi�J��ɹ{0�=3��F��IqMcs��u�E����yp�{�V�������q-�X��1m�َx��z��r���ؐ(���X7�w���Ё����:�Ȇ�+I4]�M��~�r��2v�`�ɊBBr���~d��3�z�l�(��o��0���7N��9�����^��r�F���ߪ�%��~��p;=�J<���B�V�E��$E��f�f45�@(�k� ���-��m���gN�~��F�4�u��x��2�A�nn:�]V(g���|�|�qY*����Pv+d�v�'�3���0��m�����Ҥ��ĵ���`�F�e��!gظ���_��"tzV���׆+G�fo ���C���a2�+���]��f��@ ��F@k`q�`�L��d�����z�2�e�1��^�+TT��J�좹��hx����.��N,�-��Ǣ�
���wB6ٴ�� ��v�)�䂑��2h�d���-����E��%�Y��=�:�6K�4{���a�:�E���}T[9�NoQ��/y�M��Ҁ��u��{G����VL�9��n��f��*������a
����Sڐ�-����8�5���
�|��>�'ɼkun�#.Ҕ�@O���]��;LF��)�%h`;V�4�yBH�Q�p�S�cʀE��*;V�ۙq��Rr�,c!�<'�a��pX�����O|�!��jd���"�J�cI�Aŷ#�s4�N�b���D���fe�"���M���G}Z`��^�P-r������ �S���P��.�5'��20fT�k���ؖCf �>�܄��}����`���uqլE֗P�B"8��y5y����jNoǊ}� 8�|�;<w�~U�F	�࢙��!� ���`�;x�i���1T9&�vD�����aWJOM�8sl�
������:���k|�ޠe +��](0���Nd;y+�Pr�&��X��2���&#R���]#4Ih$����.�-��J�ּ�)o:A�'7+��:�.�o7�x��>�J��/�j��_滣
�\�l P=�z?=G@���ۋ���ͅ��W`������
�8G�ŗ��.ne;�%	��k�>������:ݪ*3�ۛ>;�S��Yw�}�y�b�+�?D�%H�]�׮�&[-~�5�KK�C��Y=�;�׮�t��4?
	ا
�����<9����6��طE��3b\�.Z?ț��Z�US� 6�8�$'�j\�O���pj�IHfq1U�m�Z��o0.�k�)c,���&G	���k.$*�Nӵ��-=����	Շ�)�����UT4\⬭�/�+���M˱6c\|u�~t�����/ʝ���aZ訊���+�����U<<L��Q��B�TX�#]����+��L�W�]�Rs��3�p�֗BxyC��z���8<�3@HO�Q@l=�N�ͮ��>]4��:\�8�j�ϋ��Y�3Cc����KP�����1��VV�����#���<ݔ��u��:v�a��4��o�T�V8���s��q�N�fpVx���#!�=�B�r��i�H����y���P�ؼgr��1��3R�os]�ZP&�7�=jT�d�2��ysKU���'�xY;g������yS��+7n6)QM1�Ǯ6���7<���kB������e�²����,}E��̻��q��y��ǆ)��rlw�@q�@���8J�tYݚ;d�f���t��o���
�D_�~��/\�?�]�}���

���%�T"lB��2��r"���a��r��E2�*��>)������`\q�YXp*b��~��ί��lPV�����oAHz�h�}�����J� iQ�۔�	?�K�v�RY� ]�5�ٰE	�F;��V�z������C��C���?5i�XR�bw]�ev�K����~��Ϫl^Z�7J�X�ZX�-jQ���&�s�A�UqC���0)i������_��_�65�_�p,�*���g��*y�t����j+����
|�{��|�������=C��M;��܁ �OĔ�D0�?Z�H����k���	�#P1{�
�x8�/W_��/�<g����B�k�~T�ɭ���ͱe�F	�l3*����8��K�`���i�
���}}����B���]^tj2�(g�v�ہ}��$��b�%���S��h��H�aRz����X���G�R���a��V)��9h��݂f�B�#R$�F�.�=�Q�5���+KaΉ	hڧŴ��@%"�	��zm��ND��(n*g����/��M�ڴ=-�7��	������E5Tk�I(ɦ�v�D2�2��4���Q���c�w�BM�>R.$r]WR���$ ,��U��e~�_q����=����}hyWָ��P��u��E�Y4wV�f�gO˥�v��t(a���d<��rSv���t8n��y�0����ֳޜ.�U��wɘ�
���{)���E�=��-<{���tb�ԩ��2��@�oF5�|AN�'�[��5��s����^���F��EF�Q�#��d7��P����j{:B����x�v� =�"�]5h�����)_gߺǞgn�#�/LU$>������A�%,��]�t��j��_�q$7xz� ԅ���z��1���sl�@�2�ѻeOx�˸\\đ��Kv��P�%�-�ZJ�{�/�I(��:��B�z�t\QVG`�w>�Q�����3|OJ�E�?����i�6D�W�9]&X��M ��L��/�ݎ�Ԅ,������3e9��o��D�\Z�
g,������L��P�4�a�rR�)Ѻ(@D�Uϟ�r�h�pp=��:� ����Om�j�&N�e421�]�{�N���뿤�P*Е9��K0|���Qm[�q�
s���r��;>�����\�w��-J3�؄GQ �ϴg�\�,�����Q#��E�[�I=��rD���$��^>u��r�×����(��������^�&,��Q5����T�B�0����p�0��l�k����
T���6}g��j�]&�����ZE��g"�[<�;�r�H&_����7�e(��T���nl�pZ����R�굻��J8d�����_�<�t��P ,���F�{�=�`��i��ۣ}
��� ���.������'�zH���X���&f�͑�&v�t~ěϦ�Πy$��3o��-�h����$�i���N=F����D?`7r�ʸ�I��-�$opdG�{�Rd�����=�	"Δ�n��N,�̤}PɐͨO�!3G���k}lc!f�ɇ�`��k�ŀ#U�CJ!��z֦, ����|�S�w����D�K)�L�6�U��~�.9u�-�r1�92��,'[dD}J^�~�b>��6�X�1�}�-�r�T߼b\v;K��m�ڰ�qn����̞IYEϵAm��1K�9]�G���sFd=��&fu�6��`�Է@��x*ׂ����"4*a���B4����=fI�*Kn�n���/cԟ(bץ�ϐ��8Tb��\;%��b�/��4̄��3�̅E���@�HZ��<�,@��_�o��D� ߧ7�_��_�^����&m��K��ӢF��i>���=)��v�|�| 0���/��G}ǫ�a�5������6�<��$_ߞN��w��]��([s�A* �8#�@��aؕ�א��G������ )��tD�P��,��N�c��L��/?=*�E����R��	j��У���&H�h#�K�Z^F}��14�EfK2U�-���)�"�2�r�S����J<��Bj'@���o�}B��`$N��7��`�~����ԋW�T����D�������)����[��o�
����e���,%�����y���u�*����!�ҬA6*��7ٰ.����|�ݵ�#n6 �{��xdؼ�Zo$Y}���$�N<�Z�I���)o�[�^�[�'�X�&|E���������ie�
���{ ?�Q���O�LI��*v#~Ɠ���xUN�:=�Qj�U�t���>�َ�W�	g�ӵ��ay����g��h�w�>�q�� 7�<L�6N5�|~lWXz���.�VK/�Ų|�K�CZK�p�6������ߞD�G7��e` �N���*r���,��C��SIT\=@[�G��&	�YqXjE�6H�������0ˍ�(R �jm-v4�2
`��tcPJ��A*͊�_�阄��Ԓ�G�� ���ģ�H��w���A~�$�RB����5�?�={� N�AM �o�@���"��j�Ss�n�ް�KxO���Qc|��EM�=!�&�/�C7�ؔ�q���D <���j�˶}���_���訩�H��B�fw���6!S��KS�4ú]o��٫0�[u�/C���M.�=^%�Dd����}��m�y]�C"4i�����K9�.��@z+����(���v�-������D-�
f`W��X]�㏻S'R��$�{w-��?�-[�y"��7�X����.I v�E��
�vr(���
u���3�� n�2{��}�6��<������A��^�'_����^��ɴ������; 6��9&�0�բFu���g/��o�o9o��
�$��S�eew5>1H�%�]P.
E�B���}l}��b��
l�)e�tM^���)� �u��ED��_ףH������+����94H:d]�:�!~�tjm�=EE,8Z������p�	\��p�d֟&�6�AY�/Y����旾�ߞ�q�t`�����l׆�t��yP��Q����6\�J�z}�����dJH[T��Ժo,�A'���c$�g�O��% \~\���W����"�>�����!p��W��D��
١ީ��ٺq�! ��d\	�Lr��o����b��(gh������ODwc���O��Ȟy=L�
c1��ޠCɥ�y9�s�Kόk?��;W�JJ���|����7�|�m��I��]%�ɬػGI{�����f��F\JZ����L:6�xkR��0��h�ϼ�LXo�:Nh�a�����@�!{U���@�;��
&�G�`�܈�|6�����/���*����]E!�"$�LB��F�|;�qh"DkA�����p���c1��Q����X}��*zS�y�Z� ����47G�uԅ-���h��mOw�jE%�j��{�^Z?��ԓ8e*߹�<�"g�X��oT�a�ŉ����rM��4s̒��7F��V>���	�077�pq����}3�!�_�[�G��,�C���b�t�H�=��7J��۾��X��EMÄ��d����t#�*�k�e�"'�a<��(DyŃ�7qz�~��;�i��4��^n!9�Q2��+t����1����+��oؼ�)\�� *TDHT���2J0���@��i�f�x?�bt��\ŵk�i��g���CS��Q�0���i�Y�~�;UbLȜhrt�Bx�^VJb��TςN;Xģ*&|�]f�='��ii8���%�9ԗ�hH۸�b�?W������oD:s=>gۺ���j���Oa q��	*=��Y�nH =�ZQ�I�,���aT	��>|	C?�BƓ��o�;������|h����)<��2@�_��o������0�`P��y����6&݂͐D~�*~s�E�W<M0rF�55Q����������h��Nt��-��n����k%)���^���,��@����k�L���}2��8Oټ|4/[�}�i��*3����Y����u��G1�D�!s�h�Fk~|Bd�?����R�-��\�����Kq�3�O�c+���:C�����>Mﭹ�ӧ�x'\�Y+;0�՛�|��B$Ya�"�T�u�I�4��|������u�R��7+B�(:2d�a<Fsa%w����>�w�94��_\ P���s�9�U����̃�� ����m��v��${1�`ꆶ|KS*N�����L_ݚB3
����V��T�% s`��/�^���:.�
8��Ju��qF�a�X�4� \�8/d؊F�h2�F��� PdF9<���,ρ�<S	D�2V��,Wm�#H�{��f� A��u����	����ܲ�E	%�^C�M9�h��m��O�⭳�H+2%MѢ�Dª�E"E�V�_mF��dy<X����@	��c]��&��H�~����n�1-�~Ԑ`	@ׄ�֫�NB11I��7�2�g-������ ��χwV�}X�Qh�[Z���d���^a��]w�;xzn쑀�i�p��:k��M���d,�k�-��e�9.�|�yXZ���:hlE��)��K�J���;1���y�ќْV����g��� +�&��"m��X����j߳B�_΅ګ\�o��J�Do�ac$�	> �y�����G^$�#����y����d�IȌ�)Č�����������U:Vz1��K]F"4s�:��e+ju9\�\�;�
L�ð*"]��Ѕ��Kx������X\��sQ���r11tʕ��!��9����G8�})����3�c�O�tMI�UAd�~gl�':���G�D\�� �>�'�ph�߭pn��lJ?G��t~�|FXv���h�vP� e�h�̽˓�[� ������ӟ��)B���]���W�
C��&�~��v~V��a�:���M)T�p�A��*��񻸐ֳ�->3��>}�6# Y��h��(�v�v� �TތR��y������Y,m&n��d��l�RJ�� �@؎%�77f��[�����m�q�����,fwm��c��������?~b��#�sJ�c	PqP��rH'��$j���4�n�yE��pF��)����XW�]Ka7Μ?���kj}��K$׀�V	G1졇�(��`�Yșq?�+������f��S��@�ޚ0����%� �OT���{czHW���*������o���u�]6��i���ػONՑ(��.J��8[��E���k�l���//�g^\[�b�����,Ӈߚۦh���mʉ1m|�.gS�,�� rap����̈́�ج��n:����"ݼ6�T�j'B�{Z�o�lu�� �kޟB���3,�����r��<���ã��������7G��fOj��y��ӻ����\9�����o-8�>�>�7U�u��ۆu�㨧�����Ē^nx&�0�k{�+��m���|
+�$���?M��-�Rx"�N;�@V L��\��컒���!���M_q�]�;3��Z�|_��}zH5«pƘ����-�9���U����9����	A:�۩��~���*��j� -�-��fx���蔥�����HTf���:H���ъ^�_q LG��)��	�Mj�`5�.�5@�f^|)�	���j���.?V�pȚ2�XT/Q� p@Kg�*.P�fP�%�j['���.���8V$	��pS�b������&��V\eq5.~�$L��-7bI�{��ao��F���Cj���[�ش���-�hM�_Ǵ��?ƺP��R�1�d��ӥrt�ހ�������$���v�͌��*��i?������^h�#���6Ѯ���N����|;��M�"1T��������+�J_5��Ɯ�p+/~��AmhjcfQ@���.�?3|rI���s��Ç��������g|���rL�����g:�>VR}���?E��K�r����,<�d��RG�9�����$��~l���Vc$��z^&�5����?��{��(�U�!��f'T-�y{,�g/S�
��bϲ;_�g8�_�M@V�Ha5�nF�P�lٞa�s<��N|�OH�J��E%i��&,������e�n	��#��L
���UB�2��a|��ף��':a#EH�5
���<x;2��,�!�᱀8����6���q3�i��/y#��QV�z���-\���S>w.X x�7zH�����5D8��ʹ���% j�/�;$|��a���׶�u���O-�	Ē��B%.m�����q�f�fs����T�AEK�L�sul�~��/�	ܮ���Y"�jp�D&Y>B{�Vs�Y��A���UJh��M�6�j�ȶt/�8����tA�U��?i����͙�1b��#�H��b�Z ���3'�`g�D�?�!`8����.nA&J۠���������^߿y}`
hy���r��h��u��loo��2c8R����C9�~u��α�/�����A_��k�u����]F땚�����28�Aծ�=����R�6_�=�y�"%4�̼Ũ1>� /P���Ô���7��
�s o���^r�@�y3�jx.S�;\;���f��P�~���t�������=7@����˅A쥧��N�{��Π����������
��fW��9�C}�S�f��kwޢ�$9G	��o\*�O��E)�B��l��|�O��6
��Е�q ;]Ϩ��u�Q=tb�;s.h��i_�v��,�i��
�K���c��<�uf����4�-�G9�*��$v
�RË[�ח���h����b�H���"�F��	��l�(���;Ǒ#��z ����I
����>_mHג����h[���;d���@���_�	��`�ߺV<�E9I 8}�L���"���9I�s�/B}�Kne0�Q}� ��T�e�zR�� O�����j�@��������0�{#]hP-�Cɜs.���M��y|�Z$�������;l&�E݊�}�V5v������ծ{���9��v�	JM9X�<M7�lꑍ��!R��M���.���N�Mn����_�iK�w�rL�J�'�����r��4��#miN|p8\�����,��֓cG�%��md���&۶��l������}S���nDW#��̌����`������8U����7H L�̡�gܖ��4?����x�K[۷91��a�4y��|	���u���ge���~ҩ+~=;�J�}��:�4�n:g�L�ێ��O�!Ƴ�[�1�<4�� ��Y�l�9`�s�K'�|Y��J> PR�H!�;e�,#]��5��H_�%H<��$���S�G�1�uݚ����X/�A$�]j$�+W�kGx�2�b"�A��BOxr�^h�����<Q�i&�xԶ|7��>�)ۡ�bwt�b��5�G��p��崇�-�@��9fW�s�sۡ�
�[i�ej�k�kd���C�U�/-I�W�D"��j?4�t�L[�C2�n�+&ؗ�ů�M��p|��]/a��"�-�`��.��x�T&���֕F������;	��\j�T�s���m��\"V��%V�2Z �#�u��)jk�WL,�zk�rpK�=�QCV���\�[L([Hf��x�����w�c�$��SԮ�����"��9�R%_��e�U�=��n�}�\�d�&�"��:��ɻ���؇��Q�n��Y=>kU!�4���A�`�P�,Q!��6G���eP��`maf�Q�HdMȲZ��>ʐn�>�GV�:p�o���.P��%ZZ��O���Ө7�q�jm�o�&;q��񒕑��WU���^Lߒ�L2y��[��`�2txIrj��oy�{1y�G�g��o�h�R���EcW���=�S�s����
5��Uh�0�_X��A���>�'�7�l ���%�a2ҁ�΀�k�s����yJM�Fh��-��<��-�h���wSK����0�������h9��]��N�����hͯ!n b{b���u]�ҝ�ܰ	Q�W�oK�|�����g�t��m��cz���D�6�}Y�r�o���#�����aW���.���QwUa��"�e���*�t����M�vc@~+����B��;x�c�,����^B���̍2Fu12��s�� �������Tc�|�"���q?����sc��!Uz�TK���<�O��k�����A�܂6�����%�+zZ"�_(��$9o'{�3ֿV�����{���-c[5$��e�m$D)b�9�I�V�1k�a���M{}\��ZS|�j(��;Yu�3a�H	�b�Z���x����T�m@�ȷ�m�͛�W�*�NJ�Q�tOwA�iZk �����v "9D@T])�Lu���1���7�=��̤��b,�p���9�G��Cc�E���4l�H��ȾE�x5�g�~N�gO���@�.�2�D��x`�u�]��α�Ȳς�Ѻ̀�lO���<aq.�����51Y	�OX�\%�͍¢�	�Nӷ��*%��']�@�oz�=��Ta�Z���M��'��!z����29��ND,�o��WP�=�	
��h8N̈�P7&/��(q-�	�l�F>*��l�*�~P����n�������s߼s����F������MN�����>Ԋ1��/r���V�#��È{0c�'!�6r�khOō�*�[�ש�gɟf ެdQ 7��V�Q-��z��a|f >�-�l�"���v��[醫Y+g5)�E��'�����}��?�����1���<*	+�i���ax�N�G�ܷ��n`~x/�j�V�mC�p/:p�$�ﲫ�]�Ѡ1I�$�&�h���y�}�P&����f����{l�O�=����c�)�ڈ8d�	:�<v%mv5i+5����f��ҔT�׹�h�#�p=5��@$#_O�PK��(\�y�8W�c��KN�>@E� �B����}�l�w@��cd�f�q�+�����oI	����ò��W�^m�������r�h\u�R{k��hbD��C�Ǒ���\�>�V�rV$���F�8�_��3BB��}(�!p�{p�z��6����VThL�1�\��R�3X�y�ΜJ��lV΅����ÿ֘1�S43nPA7m�����{:[ӱ���[�u4�}J-�ۯ�ӑC���ɱʶ`P~KZ�)��Ty����=)��	��-��2Q��ݙ��F0 K��Dy�odtzw�&�q@����º�O
��1U_ ����vJ ��)L[���A�?čO��0�]��N-��@k���'�ɩ���k?�K��0�F�}��38�m��`�������`�8��h,NȗK��.���SK&�9��hs~�o)R����7�-٩n�9�Z�y�x�_~/7Oid�~���=2uU�nn�P~�[%sA��]g���Zf+�t!���yPN�i�uTٶ�5�:U�˾������δ�ey��D_�peN86���,�o_�x��̌�����xD5�nCg�������/]@�⯺�*�3H�̎�$a����y_�1�)��ݞ��Q6U��H��x�_��������Di,�r���©GZ}��ڀӠ[Z�PUT�vZw�L�tIr�\q���f�W��Kc�e��^l8�3�������Q������\����dم>�W;;>|���,z <��΀�ͻ����p�K�Y�Aw���@��<:�b_��ȇQ�
NT����[�A�iMK�uV�5�r�&��/�X⅟v� @���=�TM��y%�xh;�>�����B�]���m5��6���8jn���r��[�`����=�b@ �>y�Xօs"fy7ߨP\5YG2��W@f&�[�t���(��gB�kk�Ԑ����w�1-�i�h�b}�A[v]��[,ʼ�<v��_ǆEk��cꋨRs/��:M�EEL�N
��z۹�ݹ�+�d/�K4ϼt+:�m�NN�k�uG�g�f@��Ǘ��ۛ�� ��2�Ah���3	��@�ޑ��9{�.�2dj� �^M�ϝ+�΂�v����3���L?�.�>��-s$�$���q�@�(y�\X�q�G/��W���\q��>�#�ߌ���Լۢ��o1���1�E�r�Hj?$e��o��4��i2��0#��^G�e����P+}�I���YL��\`8�����y-C�m!J��C[���V^;3+�����0J��dq�9a�UU6C�����Y@��CHzf��@-�²�����k��it��0���I�P,r�?�l�+̸��xQ�k>��kP��'-�=ybq����C�7v`�fӎ܂�[�r� hA�i�o* W��0R�7qؿa��~�JNMe�w:�+uMHm�\���r$5�S�C�ٞ��J�m�C���t|�-�������<�v������/�n��QhC罨\�6'�?�:�X��8�����q��Z��K����Ṙ�x
�:�?��F��H$rW��Mm���Ad ZY�|L��C>s:?v�a�6F���ˎȽߴ�_ ����Iz�	t���iȢuE�C9l��v�6��	�c�Ft�cn�����I9f��&(���U@�[�(J����ی���o�|��qۀYtK�@��&O�M� WA:�XX�ww�QY�+�Z�xD�t�Ó08�l�1�
<���V�_�1�)SUi�^�ȉ%�9���n����`�>k����+t�MN���%E�0w|��p:)�N���d̝�(��������d�﷫�S/0kc^La�A���¢��V�3�h�n��/�er�_�'̨���7x�[�\���䌧rTsL�@uw�$��0D��Ӄ�)���I_̓��&�:!�6�s��p�p�q��%�3|�i]	�M��|93��k���S�>4C�%����Xa����s�KD��Y�/� +��{=��6�E=�.U����ϫx+0u�v°xw��A�z@�ʱ�㔃�Q%����7$qݍ�wq��*�	t�I�a!�=�!�ľ~�k�gJ��n������K��,Az���!]3G	Y,M\�
R|&�`x��3�l�� ���R -���ו��e�����x�X:�!�M�+5D.����b�� ?f]�M��#7�(Y�ʼ��ֿ)b%�4�)�IN�GStW�)� �AֳĲ�Vl2m����,!>�d%OpC���)R�\��9��e�<}��K�/�#�X��}2���{&ێ��5**���7Ǎ������m9��彛'>ٻǦ
���\P1a��g�_������`��p��/��w��cK+$ox��ٝsJ�$IE7�3��zH�{Ѥԣ]ğ[d,p�)B,�Kk�C��I�L�i?�&�.�#<�7r9q�Ģ�V�:
`Uς�R/��k��P�RBYX}�EP�B��3N�a��J���d����0�떺�L�I)�B��!�vjb��P:��Y�t��d��d�������O���N��dB� EQP��Z��$'�i���-Ӑg�x�����p=z
�C!��6~�v]=_%��"�P��v<�g��m�*���D���zz}�:~���@������Ѩο��@0ه�+�}�|V��!�<�J���}�sTw|�Rd�w��'��������ŝ��vfU&��7�Nɬ���,�k}Ҭ;]n����>�ޚ�slA�l��u!{�	�N���)��2��v5ǂ�XX�c��"��"u}��8JSi[�߲����䔷��$I�T��|zM�R�B�=����v��)pZu�٘���_��$&".nB�z<�#� <��
X�en��t�}�����颬F�3��/���l����[Vx��B6z!�V�#�	0n�����������k̽��#���5��/���؈	�W���DM��aJRjn%����ݣ��Y$e^��N��A����/WbN��Ϯ�4��`�z��x��?�} UT:V�٢-�E��$��1��*K+LD>!�i4����b{�����į��\k��� K��}QKh��F:��i����J�:5}]Y���#����*m�~s� C�{-8	{�Oj���E����/<O�q�F�K��"s?�_�ډ�b��\IYS��'%'ɧ0�s{�B]���O�s�=�ӭ�7S?u��LT�=�_O���Ow�gk�vJ&kFeH�K�~u����h�;j�P��W�v�"���$���j�w�z�Dp��N�jF�	�$����s w�"ȧ��n���K��:�;/ y ײ��&�G�A�v�\j��,���_	�����p\�?
��2َ(��:�}�K
�u�zω���V$aT�R\)9�6����`�q{(f�P͠��Uz�LR.$@�5���,'��*�"&��V�F��r�h���'�o�!b½�\��T$�(%Ǫ���M�4{�D��'���%�y��(���1�v�����ȭ���qi$�u9�4�����`�J��@O�ϽƝd����'��&
vit|�1ؕ7W��O��1c1��׃��ߡ_A�s�V�c�p$��8ME�9j&r�e��:�\�}��1N�Ѕ�l"���#��:t�Q�"���l:�x<��[��.x	E��E/uP�����j���E�7�Y�y�;�q��Q"����m�;p�*ȧrG���|&��fldP�0*�wz�5I�o���Պ{/11H'Te�>Ԙ'z��� LHwL_t��n�m�ղ"�����t�I�--y�R)��硝�.��̳.v�+�E���)��z��˯�[��$��
p������P�m��\�/t�|�0�4�t�Gʶ!�(d!�]�?��!G�W�����ߙ�Bʋ���W*�4U�!m�OS�O�a&&�A��K(j���3.ZOW�N��J?w��=���T�:�U�Ƴ>�����b�ߐLP��h�?����B��<�┯��d���T�3,'Yy�t��'�G��/�n����"6ўl(ܣ���$�H��Yb�,��h5�5�vC�� |wP�8�]��_����V3=�.�|��(y ���:��fg�c�t����֟1/#�kD��xG(J�H���R�~�^�/Q��-�W�,bس���W7y(�Ü���2����9 ��&���z#뭞��5����^C�cM��M08�+Lz��V5���y��\<	�#�$��)7�_�Ҟ1��CM�ʂ��X�u�����'K�6��-���=�������*_n<m�~yn.t0��:I�Be�q+�)N���e"�ߴC�tV�9�[�&�^#����;��[��O�L#�~6&C�{��N�3���iN�J *Ь�n�$���:��c�_�tm��iz��!�&]�q�l`Y���Õ�)�b��� ���mF�uy��+N< ���T���Ui#o���O
 ;.>C���Ԅ��_2���>w%��L���d`~o� �ʙ�Z��dt�l�(v1��lL��i�2��6���n��)���(
\��#޸��v�����.��}���.e�0�8�3��UbϚ*щ�=�8ZaT�r0��ܒD^ɒ`o��itip��5?�P8�,�į�;&�٣��f�ԋ&63�k� �B׫���=��"����m߬��pD�ŭ��z�������p��x��?�U�_�v�?���	�M�3������+�.z^���8I҇X�wf�k�.��t�-��<p��w%��y�������X8�1��A��hB��V{�d؋�0h�(��� �8X�D��H���O�DM���q=��sظ�4Y��Ǳ狮�� �c&����pi�)cGG+ͺAB)1���6���
`���#�H�ckWNG.�$N����:��K�b)6���"s1�F]�A��xuR�b�mF�6��H ��*n�1��^L}�;,�����J'O�W�}��h���U�5($�OnH>���G<>�����k����4�O�e>��+��Q#�E�8�?��V��3�s�4�k�n饤�e.�����uC����2²B�a0@���_3zl�����6.��B�C�mt�9�H���d�H��Ų�.c��7p20(�c||!�1 �1�%!�_|�?.�O0����7n���?y�R5)����x�9�y9v x����i[N�p(/�H�6`o�;޼d���N�����0kƤHp�?gň�9�7k�eܟpN���6IS���Y���)G�C׭^�d�[C�n<j4F'q.D�0hT�'�/"@�F���sO1T^��}�3[���o{������S�:kc��/7:������7ʺ���	�$)��ʩR�HT�F�	�TÊ��>6P����Ώ�t�ں�L6L�L@�\�>C�y�y*�b	�3���6��0���i�ޘx��U��u����o?B�#_Y��=����o�W��ԟ2v��m��v�Xv��U�,M]�*�HhL6î|�_!+]��;b_V����cAw�����o�HU��tW�f�V�l#U��[(Du�gϙ)��6A_����O�ґ�4�]�{�G�]��L�RkD h��0�O ��"5���[�qsr�=}/�$�K�����!��o 'P
�[G���*Xi���J��Pِl�F��iո�r[�@qb-��� ����#��0f�~[mEr؋Ol���L��Y&|�y�M��"L�[�2�-K^�L�� �����3���ծl�f��]�����aL�kTs���5��vN)�Ҫ}��F���6��8��Kd�� Daq7������O�#h�vK��B-����M�֙�dX��ƃCl�`���B�M�I�����������\9T���x�:����5[����:�*g_4��o��)�����}�]�pRI�?�y%[���[�z���ʅ�f��\8�R�;r�q���(�Q0L�C<�*U�=�-��_����Z� ��O�
ֺ׺c'E�[@�z�����h�w�|�b�v~-�Ƴ��u"tmkн�w�:9;펔��?h��g����Y��ϙ��'�	o�Ϛ!9m�Y�#�[��b5��TG���
 ���0?�'�����w�������-5gl����	��8��	G *f0�a4�*�9������jZ ?Ku�!���ZY���|��Y�9b�]�m��c���ǡ���A�s����\�ĕ5,�ʁK^�#+��xw����SΡtq&�`��,��*�3GÃ���>���4���80��.<��)�<�~r��}t5��9ۓ8k+�^#�֟��i�r�b5�X0�r�Z�oGuV�N�dB��VR�f?�3'���B?תϓ�k֭��}R��3�D�����:��r�L|��	���?��i�I�����U�a�;�?6��y�����Cg���P.k$Nr��h7	����iB�NE�����ś�v[Z�W<�+��P�:�=>^ɶ����	�����HQ�'QaI�_�� |�^��"F���3b�����p��D帰O;���T��7���S����I��qI��O�������(^l0>�hC�5�6ڶ���������x���8R� ���9����[Ă���[�� ���d'U�~d]����#}��3�8Q)SxE	����k]���_i<]_o�w6���
G �����؞;v�b$��p''\�P�� .�w����R�5]��c]����Զ�w����!M"��7�ো�9^ggb94)��ȿ�Qή�җ޹{&9�`�7����A��?Z�Xu^�Luk��!/������W;2��(%�ԩ������q8��:���5R�Zqe �<oMł �>�1`��
-ږ�:x�Xs��K&��r[�� ���M;��W��~���(�?�S�̸E^�c`D樗��.V;�^��w�M�
C�t	6�.�������s�y��\-�/~�{D*��2Jwf,ٮR�"��������[	��r���o5�����|�G�ϼ���_C�z~��Ȋ�d-�úa��B�j��>%������~�(ұ�Fv��hX=��"���	44[�SЀB[�{�P�'�-`�B��

�5aaڶ��I#���$��^�]��g���ʋ5~Cͅ��I�R���&^/�`�ss1{���{��L���X\\^�>��-������RW�r]n 3����5k��7�r�TWMh���|�`8�%;����\w�:81��e�ݬq���(�,E���w�i��8��S	�ځ岗O�m�����8��2�a��?dY����6�� 䨁��-�C��o�JA[���������t�Z#Ï�j��wC�$l�vȶ>���''�	�M#�+g7�`4"��I�}�	}3f�R�0Hjw%�7����Պ�[��8I�����đ2(��b�),9G]kՎY�'m�Ħz�����X
�Ւ�ۇ�&��u�#`q��{ғ����xj�؆s�#%� E��
}�ۑT8wo�;lg�U�ͨ���&��B����V�U3�o!#�%��ޛm��ؘ����Ykw���T®�s<�F��%�Ù����o��*��%��N�I�*�����l���$�;Z�j��91����6W�$��{9�i��k����L&8M���	������4Ja����;e$(/bߚ�ԛ�0��T��-��~�,�"�Xژ�����ս�?8�����S��~���˨�Y%�ĪŅ�2�T.��'j@�4IVR,:L�>�	�Y��;! %Mj+����0��EV)`���kr��T���!cNp� ����XP�oK��o�'H�z�{�8���~�z
>���qq�`+��7x�L���!�����_�̑�6t�G�I	"L#���y��"�7��2e��1D}���i�7���?C0���3�M�7�ˡ#�|-}p�9�����	b� �'͔~pd�;��$���B����n��%�Ȩ�؟ڗ��O'��o�Z��ι�W�>���"� �J�sߥ&��R�����:Un~�隉���,�b������M\n�	o��T�yh���-0���˯ac�z������mhD=GF���ɘ����h��qD����Ϡ���1�w������(@
4�L:�l$�Ƴb��^�*
��At9Yd��{����=����/�����M[_���O�`a�@a 0 ?�������{���Zcƒ[�����hȼ9T����KF�x�L�uׅ�����1����5�[Tc@ȕ���L�"�w�A}-�qx�5�0��Y�f�Ɨ�Nas��m�����E%>�<ve0݌2��k�&�H*t�[�M.P�Vy���?�]���.���ԾiD�!�i�^��+$L�ֆ$��r���uZ�/_{���uq�l���`�I`�C�Bd�Ѽi#�^τ�I2���;�?��e�ƤF���v��κ��ƲMd{�&c��Vi6-W��-�*B���U����3+گ� �pz��ު�y�]��C��q�ྦྷ#���ň%�G=��5��T?��/У����Y��a���#����E���)��"��}�6_����K m-� �E*q�K�� [� ���$�I�bn@� %#w�;�#����l��� P�9�2Ь�J����ߔ�������� ^��'	�_������V`�S.�R���t�2u���%)�Z��zP����R����E���l��r�<�~/�[�5��Raq����=��kj�ԩh�\1ԫ�B�a`/*�s鳚M�;�㙚�����ICMm�O�w���[D�x<�ֳ-����П�vF��O�
{�)b."�wӧ�Zͱଲ�y}�q2�G��h)z ,[Oנm-�T�ƙo �A�ܘ�.����x��cM��<��y�BK,أ�DU�a+ $y>I�3�@.��S�U&<�Q�����k>!>��[g]�-�!H��*��`2�4�H���)M���&�9i>?U�%Qp�3,!v 3j���t�N���<�]� )ae���C�����P�����-e�3���g6#yx�/�W�a�:��''+��Ζ'��m'������0,⏝v4���Gm~�Z�]�wֵ����}J��r]��L��T��!�t7�4GER1�ƹ�ʮi<�7�@è�a�=O$���Z�郆�M�Bש�S`�pAn+��9�$����\�dv@���ϧO�X�Z`�.S �_9�cvL�⇈|VD�2=�"]�*Ew"��n�en}KX��$�;�L(��@�N���X0BM�w"�]9���P�;��)j�榁@�&�Q�����l�Qd�Pdl���լ��	���WzW������L3��F�U�`L~oP�:C�,�v͞����z�"�T� ��$~��߸<<ziL40F>�_֋��(�y�	��@H�f���4��;F^�A�2���n�f�3D��]/�2C���ڋ������u��OZy��3d��q1�Lۃ��B�t����&�v��f�(y�� �(
wѩ�e$��Ȟ$MK��OL-���[�C�LPC(mM	��\��PZ�W�E�1�;\�x���ӭ`�7���[�?��^aaͦ9E"j� :�A�f�O�������K=��IV��i�-���]�P�:&uR�1`#�z/[Ǎ� ����)?��rp�o!�
U`z
x?̈́qg��d}Nޤ���~T�~3me��ݯ�����㗋K��+V(l3�b��.|�h���FP�4���w�z!�xZX��({�$<#k��n�6�H�-_��>�����x3q��l�L����yJ|.�W�E�Nj��ĩ�t�v$qX#�1* ү�2�j⡴��l�RȖ�ޖ��ʟ��2��c23$F��Qz$tH�|��7�6��<�C
��;��h��a��J�;1�7���4�6��"#�2y� �2��2㟾D�'��7u�X=O�Z?r�jB^&�:|��.�h"IG�H�Ny������N�c���@M��=>&����w�