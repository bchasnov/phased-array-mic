��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1���e}ʲ��cg�t�ϙ�a�:�KR�%���ݧw���ȼA�����6���Jt�߁&g�h�R�F�h�rӀa_����Œb1�}�,t�-]dY�1�~��9�aW�W�b��8ln���r���#n9o2p�&:8�h`��g!�}M�{8y����޲t�p��BzyP�؎L���a�*��eDЫ#;�8s�c�}�I�<6 ��.��.Xo�9��%�Xs��b�Xi@�}��ݓ[��Z�fʵ�琫C�l#Y/weqq�C,E"ȗ 7��K�?+W��]1G�ǒ�H��:iE�k����$�Y�������}��M�X�&�FtVz��D�7q�(\| t�� �cFH9�i�DyY�|5���*�	����f��������2�ĺ�"ѿ���S�� �W��d��I͝l*�b�-�0"�ht�i��SIA:T!L=��Q�1U6)��������r/�2�**�!��UˣpG���L��g�v��ߕ�vY�_l� ���������I�A�rr�O���&1LƼ�$&�iV�7(��٭`O���A9�p�;)ð�. 퀬�
P��L�ʯ�N�:�d��w1v�1�Z�o�+�R縳�0���г���7��0xś�4)w��.*�l�l3`��5ȔwV��1���n��x�z�A�sd��S8Z���Q���dD��B�a���^�\�r&SA;������8[�p(7�2�H�OO�<auQ�N�}\v%�|���;���D�I�(���Mve�F���V�c4 ɉ�*�����k }���.eT!b�<��7��9�BЋ��b79��j�˞�Se �Y��O�߀W:7Y�� ���{�|���=��س7Ʈ��?������b��::�(�����q���3ޔ��,>XA	�m��:2$
��
�x��(R�E�a*0�cP�~L����9�Ywq��n6Ҁ�8����*�T��D�|�0q�c������{����3p�Zk*h�0��?�dw���)�
1Af���ƍ(�0 P�պ*�H����ܖG_����f}}ӣë��Zc%��P�#���V��#Ab���pm>l3��n
�푂5H��������l˧��XO����OJ�w���ϧ/��:��˺����,l!��b(�E"�d�?]ko
���ܪ?x��O-����d�����{�����1`��#	!T^�=yь���K`��o~ZS,ѵ�NާXX������t���-d����%l����|/�h�u�*9~��W^�3Y ��朰�"�\�[lNZ4miUͧ���Å����<��G���������B>`�A�(Q���>�M�	��2?$0~ݟ�c�	�漝���pC�0m҃喇n%&R�ی��D��8��5=5\-jDc�J�!=:���Y:L�8�1@%����֕�ş?Af���r��zZ���a�jɜ'@�6�RJ����Lp)�]1�����,��g�&�w<�w���eUP|��t�|�&8Ϳ��RMu�z�������!r2t���I��H��)�D�y��F1����"Z&_A=>B	�VhB]d9�����L������<׭��,4 �)�f�VY��=:]�Q;��.
���O�N�]f��
��^�y��73a�ϩ��颡���Q�	�t�%1�,*QbQ]C
C�(���ߠ�I��>7#�K����%�脋H%��g�Eާ0�UIs-�-,a=�U�GΒ*J�m�/ Ĕl;�kG��э(�(4-�y���f�-#b%)�z^	�&HI��<@�X�1�#=� ��ϐj���t�)U��̸��<|�\/��0��Z��*��5@�<��D������_���4w:2�ӹE,��1+��N0��q�R �a�2B[�VU.�c�ɻد��w�J,�������Ra�1�F��ă��7��,a�h�(k�܌.�?��C�(�y�8x�����Z�O��H���d�l
�?]�Ra���B����ܞd#>�m~ETg]e������^s�Y����iԛ^�'p��D���0�u#|��u?j9/�u�2�p���fA0�J�2�de���ęH�� ��^b�mH5CRdoFPHώ1�L8�2¸3�k7A�?O�
�R�~ޓ�+����lv���yf���.2�Y�tV���wL�	�	��K%,��2�fpMg��NRQ�x1z� C�^�(H�&_(Nv@�HJCl�%��x��RC�(����,�+�9������t�k��)0�A�c�
��p���@�FS,�A�(V�����z�1�p�Uax��n��~!b�L
���jm��[W�
�D2f@ ��T5멣�|�?���x;*�)%�<��r+��}�X�����@Q��m����b~�ҷ> VPe��
�
\��I������2kL�?>i���܁��\IRd��N��u�����U������E���U��u8����4~���!�N7o������*q[�N�m��P�����fW+
�ﰮ+;��`O �bL�2]�IO�����ٷX���T�H���L�l�-|t��|�\"3ܛ�",�( ,��Y��J�jGk2 ��(+���^ÉzKK� �n��n�'��GCC�S�^��$
��O�*�|��G�U���*�Zح�2\	N4B��B�Ѕ�Zi��h��p?e}$�5�74�	�B:d�Z`�=�P����#s-9b�n�b97`�l>��Β�	���
�uFb�8���õ���O
�S��
�N�)J*1�)����t�e^���&�4�e������.�,�<��6��O�PA�끪KgbXa2CHF ʎ_}��Ԗ�u$$�4�r��/F�1��X_A�Zy�����D��B%y�)o0����)B�	k���mڳ��S�T^}�]9ԝ3]$Fi"W�������V}� �t�e��, �W�E��]��r�O��Syĉ��'��)M����a���~�/�&�4D3q/��^����=�+�/��8^�i���s�"�!tUNΰ��qBց����E�8�{D�+���mD���l&Z��@�p��:Ÿ�