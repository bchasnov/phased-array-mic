��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\����q�?��e�I8�b�Ǽ$��"����ׯ1�V0��������2|��&���)y���]a�r����z��p���\w\w��PZ��RqS�*�
a��R�,�({�]�-���"x�����/�ָY��aA���
�`�ˈ"c��C"�¿>П�6_nq��+IuR��	���~~�!�{G�[��G���K�t[�
���s!Ͻ��¯���ÈN�A��F�Z�,@�p�RI���p2X03]>������"��hه��)�W�l0��UYRz]�l�,_����A�z"�)e��ZsŶ��#��<�0�ľ�t���f�ƍ�/u���^���A���9'US�ںK]_?r��'��3H6�[3�l��l��W��w��nv����,>�ea��~P���N��!2IrJL�Ԛ�^������^��&�H;�VY��{TT�H����x=n�;@� >�ui����8[�J]e�K�ͣ�ZY�+^��;�^�}WeV(Wh�6��lJM�K)&�?��p@�r�뫣��"�йv͟v'�J���7��*'�;)e�K�C�[��r8����At���:Ps|��BP��*6oԒhv��m�o:��A�:� /z�}*��� |5�ru�5$�,7B�b`S�iLu�3���j�qJ�_�B3s�M��2k*L	��ڛ����3'T���F�iķt^~^��WD�E�W�[r�͍�g�A�z�
/��ʡ�,�� ?Ţ�������j�O��I(��EP*�fI�q�����x[t;�f����L�R�-��6^�ˌ��rhp���r�����A u�'	X��[k��'f�#��n����y�k?������1��؋d"t�&i!��,�Sݏ���.$�"���0Ύ�%������@U��W��0����$m�Mn��}h�&�7�ݱ��yQv�~�9��2y٥@j�&>x�S�s��b���5��eр���Q�K;�1���\P��:��g�@ݠ�řu���d�{�<k�#�Dn�h<`t7�Z
V���p���X�*��@�}�"!K��U~sJ����L&���z��E��)(G�5k�i�z��/���A}'�"u_T�1�֟�W�D�un�=�9ʗ���h���qb�W�e���.%���*'$ 
Bx�~������w�zpl���<�ҹ� ]q�"Ў4Q?&V8�
�T����ākh�t؝cNA�c���S=����ޚ	}�&`o�3�+���^F�%K�E�A�������8n�i���i�;km���ϭ;�/5���Wp�>��vC��s�FFRa��m� OG��6�K;�Xs�yhT�'q��T!xZw�*�8�	���z���g��#��'�÷�Jb�m]�	���H�/$d��Ɛ�=# n�:#����]D\��!�.���g~��篠Kv�گ;�@��;�u��l���ql���M���Z�
>`D3T��3��-\���ݣ�;>1��_M^���<�p��W����g�a�kfd2N%�l�˦78���1��p��ڸPz�"
��5�9�B�M�V���#O�;��"����j�� ���p���71X�+��/�}�P,�"�ax�8�:פeir�#>[B!^|v�b�^�&߿�����C��Tu���Z�M/�*��6��zwx�m��X���,G8�g\��~�]�}RI�җ ����3��
��q��7�1īV%S��EG���n�P��<�Y%W0z�b�ᶽ��˔Hi@g�&T����������M���l�I1.c�N 9�!q��K�n�hM��:�# ,���k�=�G�B���h,��N����4��_��[��sw8UY�^=m[�*����;`�*]3�8*WP�w�d�<hòڤ|�R/��ǳ��e���	H�z�es���