��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf��4Oᐢ��\���D艛_o6h��!���g��t�S"Ň�d[��A��;�i_����������ʠ�h!|��O�ʩap&�j`Ky�����M���1D%�w�_���0�t�v���,��(��W�
��Z���ꪅm��o����	=�h9�?1p�o�El��`Y-(�,0#ǥ���'ʤ��>�*Rτ���!DwOt�U>���=�y�i�b�i�h��@���4�N=GM���P�{��-�M�f6��;��Z��5��u�l�Sڒg���k�n�S8I-W���E���w������ l��0"��?��]h�f�ZL��^�*hӷf��˖a�4, �a7ƤR�F��+y�[.��PŚ��E�]���&h��k�	1�
�9e�+<�`��4��E='�/��1IB\�]�
�46+ͽ���}3��SB�%��	V�i��a��LV*W���y6��~�O}-�T�~���L�b�X��!S5�s��6& �l�ɗGea�s ����0D��<��=1J�?S��m��-���Md;I��w��Y�{>!63$�s��������{�������R��N��}Uח����"c�^#^#�W���5��-�������5: �;6Vo���@>��}c���dt�ڍ����x�E��%�M�
=�q^h�!�}E�:��`��]�t�����J��y�ΌY���)td͐�:~�/��*YKr��O�$���ٯQK_>Ĵ�&Ic8D��<�b�⹦�bhj?��10&k[�����#�v��k�Qo!Z 0�HA��s��.W(�$�#PW*������0@�L����3�H�f���-!	$����(ܺ���Y��^��V� ,�@yqR�Sn!wl����DJ������u9M�^��`!&:뿐S�o��Z,���g�-�c,;��8��H���	�x?�o�����b� �!�&,�o#5�WY���󦑪�ژ�W�Naܓ�8�ys)��f<�Z�����C5"Eֳg�=˟�:�Z��hR\�f6A��Ak�v�I�d&$Uܫ���nL��*Mn���Ӥ�H<y��^A��p�VB�i����x8�ICT���^X7_ܾ�F�X�e	&���ĚRO Vܮ�F>"S�Θb�&���䵟Y�x�7�@���*�5���o5�Ci���jwku��:*N���PG����YZz���q�(Q����O�����%���P�ag��/C�uP����ė8�� ����3E�5�7%�����j��!��Bb�-e?v��]aF��ra�:@zɕ�=�_Lݐ	��EB�����������2�M;�3�]R@�ݙ�� �^��w�)�������:r2t �5�@/���'��۬wF���,����R�/^z�G�E3��z�G��P�Ԋ��HU%$�I]��O�&�^�P)����(ͫ�®�âs�t\�rV��"s
2������2�U�$�X>���gE���!֔E�Bn���ŷ��8_�3��U����++��� ��<S>��a���%�0H(��_Ik��������,
a��X9iŰ���7�N��kJ�6IQ��ج�1�2��$چ��^�G��M���Q[E)!�V���h%�� !��}m���gBm�(Qr�
v�#���=j��`�:,c�~����)L_��`Q\�� u�!��2�"=��]RG��9���l%�Vj��Iu��O��azKz��ө��:*�+��CV60�	� L�h�AS\�u�b/a�ߑZ� ���(�cZj���Ɔ����ǉ}��֗)/b�Yyl��+lix��ý��xQ'j��<[ ���.;/mt2G[�h��J�|���K���bB逈Cb��*$>�M&+u����C����e<�f ��D9> -�������S��q�c���u0���Pu���2��b�w.WT2��@c�@��������љ�ؤ�g�%��+x����C���p�]O�2��ߋ�X�=�)
�~����HgNt���J��S�	�;? 6(t�� �'�Xx{��Ou�����O2b���n��ZAw�!��5����b���}7���4۾y�*�}�/��#���"�I5VF0]�O�V�V�C��?V�*�W=IcSв0����g��$o�����5J����B��@	�xeI������kBA���,wE��D� ������-pws0���6�(�꒾:MwC�Ru�5aL��لȜ�2�W�Wb A�N��YȊc�cQ��x_C�+m��"��w�}��u��#�1��C�3�"'��Ì�S	0\��|Ҳ�.�c&V��.l��@�Kv�Z�W(�.������u�<#�RR�˱��*�C�J�@��#�<�9+e���Q��m��m�^H���B
qj����a[�j�9#�4.~|:`��?�F�����/�K�zI� �S�3W%;���a}�AS�c������9q��s�7e Qg�=�;�-�Mo9��R�绮J%�L	a�jP�U���{�XDPJ|	&"��w!���mΕ�l]=�;��Aw�CS,?�����q� �ݣ~���d�X�N�{��E� }J��.ռW+&�q�o���#�����uo6}:gc��+l��o}���?�eh�L���u�4�T[���E��R|��E������[c��3qG;8��!�КJ�7�NZ��6�j#�-��rH���m�ȝA!^V)t7�S��SJ�[±�+�xx�����pg��H����˵f�,+1��#�|�9�T�����R\���L̡�����:}YL��!/s��J=V��ؘ:!b}��ǚ�qH��>/%�]�n=��uo��*�@��c��G�z�[��7���BJ7�Dq����t��!��4Y�[Sc=��Y�a�p�AJsE�槆��И�y���"n�8�Ʊ��	�#���m�3=Q�7Ͽ���PZ��!��Α)|q��@��΢/@�"�Oy���AE�W�������P�-S|����r�+�Hl�d��s)���?�U��3�?z�����T��|8buz}B}�|�&���>4I�c3V�Y��iOoyd�Xg�z��ńD�WI�gB�6}��C�2e�Y�q��b�27��ưӫ�%yt�㫀�����f��ɅŁd�=����%��)���$��y���!3��_
s�L�KS�(r3���Ts>�- E�\c ��9y�'�HK";* �s-�^���Cm��<AKw���7a*j�=�$��TP�?�s����rRu��i}�r����4"��������қ�D���/�r1�M���2�r��$b�|���t�l]�~B�=֚��&{��=�'M|'�o��O�E�� b��V�/�z��L���'%~�˰�E�m"}G1�LeP%~�����{]�8��~���f����q����+�\5l��D�<��dN/��ԸF?2�ݨ.ma#+Y�G}}���埰���t�npb�����/đ��+
�6�xOȀ��{�c���n�<��J�W��#2] Ƴ�C��G�a�&b���J�5<s��^�gO��ɕ#��6W�eP��d�L����YTy���u	�M�|�!��!��I1'+�̈w��T9���g�Q���	����c�y#�����b��\���@�_���+������5H_���1��8h[ϋt�0\Sx0w����ܘw�{�.�k�4����j2/Jz��d�x\������*۪���S�Mj��M��1�۲��)[Q�N��@CZqR&]EX��4�\��
OY���8Bl)��6�x�@�;	��
l�_�ս���ېpɼq$��fI���Eul�<j��8�����'��b�`�����v�qO�J-�ȼo��,��p�	���ufƚo_��5D���a	��T���AӐ��a:�Df�:p��y�xK}�]��2�<�: WC#�`�[R�~����*S�iaG4��"?��i�#f�_Y�n�q_�X�}��������ߍ�KX2�3P^��}�Xl����'N��i�S��>ے��Wk��Ԧ�{ݨ/Yj"Tei�xc�nm�o�|4��$m`������y4Gi�b}��v[�E��EjT��O'��v)�����������9�5���Iӳ���U�<��k`�8������@�]of�|�7C�P�}W�����ק��V������vӐA�
�4I�Ә1�d�ݠ�rᆭ���c����ˠ�w-׋h��[)�+��,��c�]�ܿGc&�|bwY/�����WT,ۤ���uw���$��r��}Yg����� 1���o�~٨���ĵڶ?���<�:r�����ZT�O5�s���v}���8V���?���9��hi�Ã�Ƕ˨���?vWx��C�S��=C����0G���B�S�	鮂{��k�ț�j�����}{`�Ycq��?�.&�"�a�'K�U��َ��~����)^����iJ'�x��Mh7�=J��~� ���If�@ǟOo9'�͏�့Mxv�(�ѡ��e��$��Cu���?�4��ͮ�n���;�����C:�a�Ց�DrN����lH��Y!)�]HlN��r5�o����Y `�0eǳ�4�Ѿ�|6G�E�y���؋����3� ''����)8	I����$άeNF$\nMU�0���I�Q���W�o�_Q�?�Re>�Y����A%m\�u�9��[!���τ�r㥘-Rl��U��zŰ#�p꼻~z��������gyOs��U$��/�v[���L�gR'E�_�fv�F�T+D��u��ݮd��NwZ$�
��2�]���o����]~����c��C��wH4��b�0�&/�!+�~��ˊ��1�����^���STՁ�ݴwa�@��M-<��W�6���z|�\�bt�h��A�J�ZPv\�,�F[�m��%L�s9/�� �9f(`�,B�`���F��x|��%��������9���]�D�u���dS�8�QAχ*�ją ��lmQ��HA�=��N����%)O2��w�3�Q�c������e���lq&K�ش�c�d_r�b�"�əX"���~��t��vC��`��!��׻�D3�~T�N��}��Z2n�(4�_�D�.�y7Ӕ�8���������iD�M�
��C�� 8��"j�I�p�s��aBD�B�`L�
;+6Yr[p[,�9U�[��֎E�`3�b��6�k}󠜘�h[l�xY���ߺ�[ós�'T�{�zW��ޭD��Lw{H�̩^���y}�f��[�b��E>J����q�F-Ry�3>O�	��v���[�G�Q�Ugѭ�2�2�mgN*\ A��Gbb[��]��H�������!Ac��T����&	�h��K��`J�c8�ĳ,��`���Y�f��D���!������߃$���O��6���+�gK�̫c�>O�"VR���fS��KUG���m�����#1>����9F���F)q�qG���X�@�;�,>���O��v)�·)j�	�8��g�.$�l~/,�הF�@J��'i�=395׭�dx ��u^SQ}���#�efs�aA��E`/k���x�l�(D���_�����#���wy�8�9v����G���x�	����=�+��ف5/R��	J;�o�U���_<XO�zʓc�r�����9�w�������k����<�C[by����f�}�؄�Gr�݉hC�XK�5�S��~h�t;F2K0A��نn''F˖���C�P�XO Z���w'MC#8��v���F��r�5$,�θf,�%�5OB�<!�.yղ
��%�Ź7w�[M ��yPtz���&�	W���e(ͼ+Z��ʊ)R�璣�<4�7c(��(Ѩ��?���k�UJ,[�D:{�����w�Y��y������eq��I�Qv�o���Û�˯!k"$�0�13��i�N�A�Omk8�	~|�������_- "���B��Jٷܠ���?v����	}8�L��7dj%*c̔����	����geVv���g3������"���� 0x���gg���1U� =�5!&�bQ��G�^����M���l|����쭨I���y,WZ�W7M�V(}���fq��X���΋�1
�A���`>:Ǜ?_&/�RH��y_kܗ�m�M���Wg�i��.YH�h��E���5�jx�,������>�ƿ�;�Gw�h�
�Ǆ��H(�ǖM�h��������ԅ�Ch��TΕ-�G&·���Js����?�K��甔�sm��r��=0�c?�1���J�-c�2m�5Mm�{٤^~��4�1�4 [b���pZ��Sƅx@��:1!��!�q��x�גԝ��>�|x�q�A��nѢz({?�xN��b=Y�E}Ş�C_3r��̰�b��HY�%�1REBZ��������
�D�g���?juZc9��#�۸�%x�^⊋*������R�=�ʁ���Ú
��N[�k���x��c�?U���y�D%G���!?�̖I��dO��k�M� ��n��y'�H��k7|u(D@�8����P�rߌ��t9h۴d�Y�t�w�4�^Ɯ9��+f�$��K��:�v��T6�������I��1�0�/��/hԸ�_5=l�=����뛆��b>�2ׅHС� ��[�À�L�fJ���|�:T�E� Ņp�B��	7倢���'�`d6����=lJ�ŵ���Y��Rp��S;�vq��qUa6uf�'������&v{�-t�/������E�����N�� Gĥ#���[�@��Pw�!��f�n�7|��XNa�F3) FD���&�Ҟ�&Ŝ�mk�y�z?��#�|��ߴ����4h��|�	��1=p��z8��(.�0��l�*�d������[:�Ӟk��V���ڌ�
^��V����ɀ�-E�]c����߅��%��d�	���u�>�Y���Q؝l]����B��"!��IYn�{���؎f�}�0����T!��0���H�\�*�G�<�t���i�����ն�yK�c�Etz]�^���wf���z�������� ��g Ȩi���e��L����̔F}Z��l������ �	&����X~�}Ad!�{��q�p���j΍E�����j��%�ͅB� ���]:�S�Z �)77s�TT@����e�մ����l�.��W>��2����X%fd�g���:B5f��\^�)Z��4o'��n�o�Ƀ"L�J��%��5!(��<��Qa�s����X�կ��xk�f���l&�&�V�����Ĵ��=]T�%4��/�j��A������s�V>
Y��^e��h�\�x�l0*D[�(�d������F��$�0I���� \���	DZ���ϥ��1�����!cO�'�A�����kk�p'�*��-��/P�@|�w]�e�a�CJ�v˦�6d�)/�Њ��g�{\6�滫�� ����:9fS\��M��;��Y�4bIPe؋{҉�[g!G�d)��Dg3&�j�-NaO�׹�trghx�#�R'�oZ�
�	��.��D��a\����O-�	L^����A���^'�؉��so�(����[�<(�n?1��_�:�}�7O5}!� '*v�d5~�Woyshu烬��-�A?T�
��:�� XqԩDJ�uAaD8�m�`o���+ڔ�x�l����Q��$�m���u��t��.��\��ܩj��I�A�h � �d[�2U]�Wcp\�ٓ�ս����^�0zB�H�MehC�����K��#�����#�WP�m�	5ϴ�	f=�2�H��p����RW;fTlZ#��3Xn{�ы9�����т�����\����A��f�\���K�?��w���ϦT��G��߳�1������O�����6h^�@li�6�L8�ч���jP��,�����y��<n���'<�E�d�nk���u��Ne<c��W:tVa���Ճ���tp�!���_B�z�\�W�2؉��5�N��s���K 4oQ`+Y�/���bڑN	�h?�))[�jqNzE�<�d�������M���/����^^nU!�@Yb^�����:^�	�{��L\��H��W޼���!��br��h����זU;+�V���¿��,�6�U�c{�z�R�ӥ�rn��prM6G�і��:O���ܫN�[�er +t"2}���Lx��:��S~-a�(ش��:v-|���Ē�R�5��X�D���s��IQ#�ٌ��\����B�I��tF;ޅ�:O�Ǝ�LBڀ�CYYo�~�m��P�5�|�?�?˼x�}�r2���A���,�^I�2�'���{��|i�]o�iA�S�_�h�4���Oƹ�.iZ��_P�������\Mdx��wE�k�Xl�{�Z�-8��
�}
���Nm�'S|7\\�ǒ  �ob�x�L��S{�D{ĕt���.~R�}�4�I~���f��������d岷-��z=V�� J���'h~��V>�1[��?���)�1�@����9������y��a���pD��%��2��;f���Pۿ��JEH�u��gw�,*���+������l}ܭ���GKV������yK�Bg,N��HK�z���Qn��|��m�N����Op���G �
�F��9^�r��Ո���%��̕Y�� ���F�{�Sr5��]x[G����LD+�GE�TӃ�Zyx�Pi��)�/���z�G���Ο�#��:+iO�s�p<�#��)�X4�!��f�ǹ��L�k�$v��K#W%=]a��+��,�����+5�&e/6��đ��z����O��/-�l�wHp�ꥹ��ے����S��� �e�_d�5��Zw[�d�x��1�[���E�����h�.]�7�g	��&��%��-{%�(���Y���ҥ�iLK�S��~.�;�쨽�:�m�(��m�j�Q���^�6�+��1�Ⱥ��{aR���K�f�e�9o�Wx�2��1b1�:�]WJ�o�;������z���`��\���Bw�����a�M )�#�H�E����R��f4r��Ǳ�t�[&��!Kv0'�n����'�ȩ�ˆi�e�m����c�8�W�@}`բ�M/��s�5�mf���qaxN_W�{�U_�sP6�;���W���MZ��nj���Z��f�fW�`��GKn��}�l!��a��WDd^�ڸ�mC~k�h?0x��,L��v��G9���}���;���;�y9�3=���W.��X>���I�!�'�|W@�D��gkGE2��<��&x�,��p��ʰ.(��;�z��y�bs4��Sf#j�fV�H��:M��[-ap�}�.E��f�t�˱��x1��q&�{ �M��c~�o�v�1pY=�b�q�
S2�!�)AXTsJ�.gIe@��a�-G�#l�|U��ў�W8	OH-����z�!���QX��W����}�x`���?���A�A��� &�W�Vŷ�Ģ�c>��������M&|�[��`����7Ú������0)vekۼm[0�c�yt*�uG���B��O�A�B1� ���n@�["��j�u5��2�8��)R����0J���=�$��xC	"���KD9�/\� O��ԁ���8d��T���|�1����-K���Y:�#ijꁁ��J�_�Ģ���F�`�?��78=�	@]��dt3.f+����	`T]��U�������6$h^U3B���v3+��χI�"�c����	0bl�uά����h��޽s�;
�#�$:�"��~�!��՞�����C�8@Y�q��3�e1�U�٥��e�U*�QA�P9\��|DJi����dw�s,=k��^2�#��C�����O�^jܔ�6�ǧ�i�^��Sq���!��#QM��M��^DuT����Q"��=?���2ԼRML����Æ�ŧˡ���=d��KWX�d�,����T����ua@!�͚���wv�F@L�����,�']ʭ�jx��%g�~��R`���Y���_�g@;��c$!,��5����T	XՊ�ޅ�=�~���cl��Z1_�6��T߷Pv���U�i��Nm�o�k���_,> T+�|˖!�N7'����N��6&j��B���+
S�����g�2����z_�My<�8JJxǡK��i��X���Ն��5��@�
����f� :����ݮ���G͕R��t���h�Ñ�
H��Q�ܧ����"'��޳WI�F�r�Z������X�* �G���7�r �-�T��-�70�I����M��U�z�;7NCnD�xT����}��uH�1VF�j̝�4Z\dK��@�)�pb/;�\��;@��Z��N��� ��E���3/�_�� ���\BKka+�̬'����Ĕ�LU�SꙜ״P��qIݩF�_��� |��\�@��SF2I����d���(�`��f�$8Z��[��X�~�k� f�A�[)�ǻy������m���B�5ʔ̴ީ>y����Q�?p®���������b��$�RI��#M9�[%��FK�9�Sw
�(\..])��e�zUֻv����Id��o�T	�t���T�M�-�,?*S,�O=]�g)�Ӂ��(�hn�� ������t87��̠"0^Rl3�(��}k����?���j�*���0�i�ԇW��vt�la�2=�Q��PcH�*�HQ�KO3Lt]����;�غ����,f<�5��i\�PY��7���;�~-�9�Y~�V�u�:'��跳���EH�*%K'�}At��A��"�T�Z|��z�M���?r�$m����+�1Y��>#�$�,^ܗ�6Ԕ0���}�v^bx)|����I�PU`�Kb9�L��) �2
8%z��Mp&yv����N2����9�#Zj��- �:�H:�����u�_owiӓ��������L���NKi�$���,���2ޜ��wp'1D��v��uy�l)\{i��H�� ��D�C�#�+�LebJ�&��1�c�Z��\^f(���|���s(�Ca���º;2~�&	������"V7�Y�#ۀ���ӆ���Vb�w��ZC	�Ċ�}+��0z�_��V�9ڬ3=�l�g`똖Q ɿb8־� �o���LM��8��H(���sP�Q2�`���8Ԥ/'lUW��$w�����&O�����l�NL\��SZ6E_�fckhw�-c|�u�|��TKdO۔ ��V�d�ž8c�F�bM�����ϰ�f�{��$s�C@�o�Q�v��ac��:E(I��Z����vba*$��E�{�5*̗�b[��Xӛ��p	S ���(: &��>��+� �a%�D	0���m��?��N4� ��>�ByE���=�{5�G?�-��>���7#��+hc����Կt�BʳՋ�����i�p��j�0��v������4�7�r��@K/#q���z�:������̀� ��>j�d�Bc�2�`]��:F|��u4�W�m�T���=����0�{;I��D�:�Ĝ��OC�����X��]�ar�݌�tS�I��OhNE�n�L�z��Ao:׮��"���If����i�y�?�����b_��\FGJ��}��O��t��v�ln�w?���.g#���M�|׍X�������|ĚT�_��4�4�^z� ���8��b�q����rޓ���Zm��iŜ1B�;�����2&_���Q��������	?)�?/u��&%&LV���N���q$[�'NO��U�J���)�|�XOX-}���%_�^�����V�ʣ&Z���)��A�R��s�6�E�8��X�9X.$��ߠ͂�uiyN��RY�d�d�;��������5񶪏�y���.�[�X�yyL�Ag���,�����qQn��j�8]����-��8�4շE��)<\��s�mCi�с���������j�;�U;��E`�y��L8:��;���5��˲W�,q���3�c���w��uYL�O�gA��� t1�n�+�j7���&�b���ůb%���3U"��N�ʓUo���;�T�`�5��qt���� �f>�f�p�,8�u���m��qD'W)�η�p�)��--�6��ɣ 	A=����oyՙ:����9;.�Zܿ�<�wg�c҆DA�J�������-9g[v4�Ph1Xl���-�!�AEh&\O<�!A�i�>u��}���!��b��{��Y�z�?���&�-�h�����M,�_���=��A*�,2�}Ƞ�,NN^mp�x{���ُ�����A�zk�ʫ!]� Ϊ��x�/��ZvY1Q�i�Z���K?o�g2q���s`�^P���v�D��ς�g)GӷM�󺖝K+�.Q �!\t�B�./Ff�����&�ܒI�LgܙA�����բ̚�����
Qz�J��yR*�4/��ei�����U�/f�Ń��`��;J�<�ߕ7���?p�+�{��8 *= Uf��6N��ا�Sz��4��)���l`�uB����X~������6%�O.���q\�C
Gdތ{f\�k.����Ǔ������e%3����>f%LL���@ƅ�	����9��D��Gc��)f�)�yRe�p[� ��b�WP�k+�R��^�WusS� ��d3��p	rL? �؟���>ha~1o�Wizl�����S����̽#��&����*m=�#.����]_ڣ�P^T��{�n����T�0n�Ո�Ԝ"EB���ݍ(x��'��p�h��o+�~ �^.=�øR�Ȱ�p��x�v�u[��?�u-j-%	$���4m�������_u�օ�Β���fOop��h�� ���Y���'�>�h�ڄC9k��Q/"���9!Hd9x���lo��M]Z򽖏i֫N������B��_T_�q��`߅7Ũ5Y�o��\���Lz��"�2�೶���Ɵv쮎�}bV�H���
K�{&.5*�|m'���"�.~�z��P��8��ĵ�cx�ދs.A x�l)��u�E)f�3����o��"9� �y	sR��0��9����/��a�4	mN>�Ii��UZ*WƼf�r+����?�-��Xh��]�kA�iɩ�o�܎f|��8̓#0��Nٿ Lړr����K���.5"��ɥ����K<߁y�E ����ly�߬����f�)͌~�oUn.ߒ�J���H��ޓm$Fxee!ú�$��|��B�(�?��9O��ׄ�
� �v��#�R�Zσ�b�  }* �Z��jz�:Ck1���Mr���r��:C��#��z�4]�-���(�鶣k%��?��-sB�Z��m@��ٓ`�*�8�\��ǧV�>E[��s�Gt�I��n���*��n���P΃'r�S/]��;�Dw<��@₹SK�3iQiV\>�a���eeQ"d\���=t�p|��s2pz����o׭����>&�bq�SH_YW���e%�
4RU�P��9�F"��->�:[�@%�=�0�i�m��j<�����U��E�}������x.�!�����M\#xB��*���)U8!?!ǀ����>�'��+�tȂL�*䘳w�%/��y:1��;�`�����P�r�2�����>0��P�Wޙ��j9�L���l��ʟ���,��Ha�o��,��n���N�(4��ލ�'��^z�ɵ�*����[s䪅r�DdW�|�b6�����xH߀Ygiu���lF���TG�m�6���-!�E�i�瘥�E!H��Cc�jRD�3AH#�^�f��%w|�[<���fj�D w��o�����c��g����\��	:#��c��F�]�++)v�sg޿�Y���7\�f�;3o"�`��E��2jI[w����҆��9�{ݎ���ߵ��ְd��/.��qU@�ne�8P�e�zA��.�����C\�%|����w$�����TGB�Z6�U^��Y�6�� ��o5!
����FP����Wm<ף� �Q��'� H&��&�vC�]���"d-`7i�k�꘬L�R\�4���
�򵡨3M�A�ND�_Zc�ߨ3ݫn�01�I�Ԋ���O�'I�5פ*Vy���s�z\��F�ѳn-:N6o R*Ĉ_dm������p�6�L'�h���u3�l�^��������_�;MM��ERS��U8 *�ޮW���DKU���3���'�c3|6�V"�����D�k�f�n@Q	�k�N_����põ�u�ւ�S��`�K�"�����(Bu@�u�Ǔ�#�#�)�*�G��c*(�<����mĒ���3�9��3��S�_P7XX�AJyB0�3�)��(��d�LN3\$�L�w�:-�_u�`)ې�(Y����F�.���Ny觽�ڈ��n�VƝ}�Ч�ZNz;U�"g�H� (���4��c�%'NH��~`�j{�%]"ai�����ـ��[��Q�����Ԓ�g$'�u�ďje���+zk�8������X�����V�T�h#@ߨ o:��͸�}�&�K�m?����mc������,�l]#�G��L�ۅ��{/�'�ܕ�����Mu�N��@m]>x�싃6��LAb�t��TE<�U��kHQi��P��eV�i�]AjE{�V�ƨ�!��Ċ��C~��A�*<T|n��"v���"�jh]gY�e�$����/�Qy~g�yF.W�R�[ĵ�ɭ�`i'7�4dS�ѓ�}�~h'�mN��;�����X�c4
�O��s�J6��aI��O5J���6~V%���W[���H�/�x�0_2�c�NM�,b�q�i�8#o�g&�d���0�P���ѧ�V_��O�a觑QѦ������6,�����Z�p�M�C���?p�R�w��_~%V>T�׵b�b0�/v�SL�IAOʈ�0�����i���gǻ���R#=�
�.�J�p�pPܲ<;�v����Kh^�~��R]����VVaP�\Pp�y��i�~S��:�|����DӶJ^�R6&ai���f��wM� H�<B/�{,��cݽ���S�t����P%��B"D�.p�4�P���SߵG
M|T�6��w�Й�`��2������3����� ���X��W�=7�y]j��f���;���g��w&-LK��~��%G�T�W�A�����13��@T��u�h ?�$����^ ^���Fiy��@qo�~�<�G�5����M�O#�2!�X�&�s������ϯg[�cw����i�t��u�(	����8�U����_k��S�տ��q���ǚ �@�ח�Q�S� ���uO�[1�2�^?�$8I���o��9ƀ��s��Δz aw���*)~́�n2+|�Ҍ�Q�n�!�yC�$}`6�1@u&Ύ?�!�ӉX��:c���}��z����������Fy�ݹ�_��5_�E�L� ?}�8��7�jS�$��{���!vV�E��#�|*�ke���d����_���+0�,����ˮ���n�k�$��J���85����;��e�w*H/:Kd�1Nj�|�iw���Q�@����p�H��t��-a~ҽ���QGñ�e�(O_U��rn@Sߦ5����3�c���'0h��ɨ?��J́H�Bh%�8$�2B��[�eQ�&��ݑ���@Z6���Y��.�OI���p7[�C���r����4��'�a�<�i�q��4 ���� �ɏ���ގ�[�ǍSV7�ab�Ğ_�4�X�oYP���\f?�'�hHa�Ͻ�+<|��>j����e����
��.J��
AO<0���֑��	�i��*��77XEs�R%�;zz�k[�%�<��e�M��f�q�P y��`0z�+�@��X�p3�C"�xk��M��7�� �oێ�I��!+nEdi:�$>�'�%F���^*��䣻k��3R��7cOw$���e��K�]��-t������"�a��9�N�\ΔW�̈́D�ؒ��
�T�٠*���88���]4�j{���X��ѥ�J��;����i'���$}�pE�V�W��,x!���_������b�u@&Ғ��C&�n����1}BJ�v�0��1Q�'�i�t�ǷQZ
2
6B��lsR�TI +Ӥq�Mt�3��\**���8�\>��V�cĐ��EқQ��8�R��b�yK�H�EI[v��U������W��b�򈑧6�&?��њoL"讶��dN�Gp�З��q �>���I]��~�0D�x0c����e��I\��LV��+|����ww�C�8��©��N��yGe���2��k���8��[�"Rj�Τ>����庮4�� :	4���/\oę�x&Nɉ)�ҕ�.������Oд<O�R��J�~�&�8O����@�&�&�
a���&	�1��=�enat�dWA5_�Շ�!��d?{~��'��t�? �C�cĒ�i���:/5��Z�Q&�~���Z�I��]M�T�p몖��g��E��rʲV� �j=�/���ȫ�]�S.���aר��NV˵AU�,�)춱�'����CV�߃� �	�/Bv�kJҚ�ݛ7������H��B��v-LF�R���1s~��y.l�k֏m��=ٲ@��*�x�>#!�t]w�����h`�T����V�@��]�+.TS�g�+����!�EX`+�xqs�Jj?w��[��T�&��fh̋���oҔ� ��={�B֫<N�zֺ���e�s@�����K+���z�Ut�̥KI=�⊣�k2F��������P,�<�L?��P���|�����Z��X��~��� �������c�������ڼ���F_�q4��UX}Ф<���^9�����B��4�q����V|�����b�04GJ��t���ɾz�D��]��S%�vfv��?%`e^��+N�H!���ݶ�