��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\����q�?��e�I8�b�Ǽ$��"����ׯ1�V0���@�Zr9�����|l$A�c�mw�0�{籪������̼&��Ys�_y�2o���Ĭ�o�b��e�hf���_���i�ԙ�_$-�������M��>�zYD�i�⎺��(AQǉD�j���$p�c��m?�BYfz�r͋p��Qe	b��^C�D�mpdi�����_8<b,9�	�N)�F��d{n����o�{
��|�;2Ni�����_�@�"h�
ܜm�;�I-"��g��)+}L����#̶��)G6t���P��b�!�wU�R����	�V���pC/4F�J�|`@Ÿ_�������m/<�~�b�) �F����+U{:{��vt1}�7�*�0%ZL��°��&͏C�Gu~Az�U�aV�5�(���G7��4ڼ2QNF�;�W�Z�$� ��l�E���?������V�	�;e�3� iQ.h�б~�-��$���3���V.O5HjF$.Y�w��Nqz������ͯ�EM���d�z1ϼ�^�~���a�t�z�k8������-Z㲀����X��M��%}���I�D6��y�8�����E� C(W�c��f��@�kxh�r4e3�~ ,[�rje�P�&�J�:�eb�;��Kd�Ǳ���-mSG�b�vgUudY���
��y�-#c�P��O|��ME���f�(*���u����Q��,�-K���aG[{|1� ��X�q��Ez�y� &�$�N~���� �O���?�����Et�.���%:�/�z�G���=�P��L��`V恫��e.x~���$��)+���=�q�,t��v��V�^c�X/+4�+��[Q�w�� 8�!�Z�/�[Ô��!��HNJ��]��zW8D�h.$���ְ1W�_X(w���b�2*Xb�\�΅a�]�6�z�1pѺ<5m��@ l���S@�8)~�X
|�������R�t}惃��+٫� Ί�w�����X~���3,�j��'T�L�ݾ|Gi��3���U� P"�\V� �gZ��F7��E����������}�O�#��xw���c$��"�p:#�T�O�� Z���Tp�> �#Jv �.O�=�v(d��N��B��Ӟ}�M^��sm���W�����G_���Olm����p(58��U�gU�H����̼�CQ。f����#�57XLVo�M�!�t��e�ŝ�w�����;�Z_�'X�簭�LlhZ����3���-M�Ȣa~��A�y�ZKH��5�Q���\u�������l�9��j [56�h�Fw�;���4�C}0���t:_��T:��%�'��(h<����2�rm���e������z�I
��g��m�$�^�R�kޘ���������e���~�cr!��7���������85:��\E�GB��f-SP���٠U�8e-��$ޤB)>�[9�ou��%Uu�֒9ձ`�����N���W�)��7�{{o�:���u���{c8@�� ��+�����HӜ-�8EV��V�z����ÐP�>�̌G���ϘO5��wm�	�c�K��2֋OMǲ)B�	)�H�i>���V���F��}�0Tw _dc���3��!{�tMW���p���o;bQ`.k�0�] =`	�i����ȿ���ܖ{�x����J����K��6�a떐#b���b���0�P��Hm^iϔ�|񣅬δF1 И/��(�;�� �U9�o�R�/M5t��`*��J"U����������.&�M+�A���Z�~$o�dR�8����҆w�Kl�9��X��%9uy.
㰰�.}{GR��P�]o�[>�(��8�4#k/;�`.�ǵ�#vN�ى�^M'Z�Nm�Jv�{q,�J+��S�$��VU,���������Nܘ���Ȅ[�t��۹����ׂ�?g7�֛�Y�U��=��*4[���Q�^��l4{�<�]j����X#�E�L	|����i��&�PM�#�?�q35�٬�&�y��(˴�	V��$����i,�0rޫ���׋[G�\��a���uK��16,r
�An��@vH�9�r5E����ۏ�m?bg��ăk
u���{�]��	Ļ��Ln�^QD�|
l1�W��<�^����4���;��Oy$i~��Y�%4 ��9#F�t��rq����O UQWm
�c��y�f��	�(���L R@����0j��<"������{r��a�0��l&5��Nw��)�:��i�EE!v�+ɿR�y�	V�5�S;�� ����Te�4ʗ�^�qnL6�	���#����;M��j��Q�y��:p���q�2u�4(-������;�o��uپC��{���j��;�+?��|1��Èn�Sh��@<])Jm��2���8^�W�z������M=�s;�H`�+>�ㄔ��_2���8���%E$'��:��m���sa]mN�a���㉃�����d��qTɉ��/�1�f�Ã�}���t-��v?��#�O�Opc��q���/��&{��FGs���r�i�Q87H�ɬ&��۷	y�Z�G��4>'FY�ٵ5�A ���4р��C�=Al&|_���:���>���Tق�N(������c�R2��-�����C����a>��v��4�q0W�)��-�鞉�k\���_�My��(�����Q����y����	��]����{f��!a�Bt,��y���{����[��,��4�bz1-J|>o��KV<N��	���:Ug����iW-<B2�ֹ��%xޝ��7����'y�M��n\z0��8&H7��#�t���gO�z)%��Y!���$�s�k[��Ȑ�����?�E�Mq���UÝ��	Li���wy��>Ѝ9�����Q�6��= �@H��%��N�' p?|�����@�sֵ�N,q;�"J��OB⻮*�z���}�x��3b�K%	��z��P�y�ǧ�Gغ5��@��ͧ&)h�=V��6cm��O����#p$�� I�|#k��т⫍N�,�~�[����e=��ۯ�;���#�mǢx�)k��8M5�n�(�L0DK�D`P(ӌx	|��ȣg��0��q�O���kL����e��[.��_���,u�+�P�b1�ޫ��G�j�o�Ռ���6�n���� ���4ڰ��]��+�o��`��6ֺ�%Յ�&��Z(���m�X~�*�4L��Vc�J}:�v ���
t��6xd˦ϋ�G�o��Jv�ݕ>g!�A:<Z�m�d�  �%~���S!6����c�
���&�c%�`�\2ҫ�^�e��rAi��i�P>	�"�XM��]ҹ=������4�JRC�8��v������뵔�p^u e�����{�rt��r�7����,aY�>�?��.k7��a<���wj�nS�Ɂ�\D3{���$�s�G�-�q�Iu���t��0���bN���S����l.�%[�����_�.tp�L�e��v�������} <]���<ܔF.�\=�9����nz��!�Ә�Ԑ)P>B#�r�i<U�l<T�K%ᔡ�^,)���Fe�K<�����H�>t���� �t����?����f�b�æ��3�����1��_s�_o�X�Q���L�[���C�n{^�̺��3�v��`ã@
*�&_ρ���`>���:!#�=�Aw����؅�0�0�pGhhrMk��b7ZQΰ�W5����:x��T�s��A-4Q��yy�]� SVO�;��@} ��O����k�K��H>�R wBXS��MQ;_4�۬�តj�Ċ?��;Іtt@˲������D� ����|���f��RΚ��Vd�(�-ݳ�Qh#��xm1�gjZ�Ŭ�S�� ��W "|�4�=�`���x�xcX���|����7�����F����9dc��K�}nG�Gz̧��U�ra1�`�� G��_��}��	8g���<����G}c�P����P����굩1�y1!'�c�w�t�S5~ny�����<6���6�!L�Y�����1[-wW[_���8u��:,�¦&i�Za鵔�ݨC�@~݁��a�MYπ>�������s��HK��u\� �*�|(��pP��:����xK��bs�n�)V���"b��5yvYv��� ���(�����%��w��Z*�򇹎��_ٯXIR���~^Os�p.��g���X����,o����|�y���4��8�ƀT��x�U��~J\@�wp�q�nb)r�}5 �t#�7��!�<�й��uL��8�֮v��|�<�/��I��% hy�5c�4Ƅ�.S{,��@����u�)2Qf�%RS����(�2���P�埕��W��}�}%��z��b����pP��a �?Q��f��ߊOn�0/NZ���e[�����o6�X|���?p�&��q�o�ܣ*�L��MzF�Q�=�Z�>��bqc-T&#U)�Nc�99_����ZQ�+�")�(�&���!@�	�C��=d�b��=����@a�Ĕ��
6p>^jxV�C��0{O=�����t�7do���A��L��<dRBC�_;_��j����VaA��n�`�b�+{�6�,��.>׼��M�Ӫ"*]���֊S��ΐi�
ZyS��t0��/z	����*!|��e�����V&�R�]�q���D�����1���|��b�82�OO�m�V��xu�w��n��S*O�����_x�ǩ3G3��E�����	���a�9�hբ+�p>�k8pY���d�'7���m��{��fIy��A�����OT"~uV�F�6�ɾ�A�f�oxK+��f&���:9�A�߄{�ʌ��t�W�r �YvV���=u��m��#A�|Imgfo<@=D��_g��R��B�TT@���3�&`iX�v�`F��#�S57[	�5�͙1/�����&�_H�g��@���P��T�>ԥ�3��>�C}�i����<x�b�|�{G���}j^կސk�����2����^�`��~���d!���)�#�A?pߌA�Q�f��1�|/+���=�vR�.~&#�5���]�I�X�;H�G��qF�X�|Bd����KGy�ͤ�(]�ƘZ*H�**RT�jN�7��"m�%	٧cV�(1��A'&���s�M�2�NE>�^�d��5�t�e��F7W\ڇ�`W�o3y$�/���a�<���J��-�:�����3n�#:0/��n݊��ب��/!
�s���-�
�rIny���++c����[�L���_��9hRځ�q$�6���@�3�Bj���Uf���j����{SxW���+�������\;���P(�8���=���f
�}�~6a
��4:�`P�|D�-dqh�f=*��l���$�v��	vSf��,}��'p����G�?��<�V�<���O�Jj����-���'ͬmN.����C�](��
�u��4�t2p3�7t��U`�����q� �S���#�X�/�K(`���t�D��@9��C�~kь!r�F��q��Xǯ�zEȧ���x䝲��w<���r�@���.�a��涰��z:Z���Ƶ��l5��i~/'z;v`��`{��}�~{Y�3���ju|��������bճ��PF���]U�EX;9����D��-A:�I[�W���,ފL��_Vn����=U����+խ�h�>oJ����CG$����h��P��Tq�\���1��/�i���T�E�QH��5��_E`fȐf"��v��J֞3��_���5N
�V9^"0�� k�~���G�"vJ�֊������o\r�	4��#q)�$��9�rT��6�m&iy�L#�TS�.���X�;��N(IQh��1݉M���d'�P{��Un0je�����kl8�5�^H|���h��*�Ӡ<��Q�Ҭ4���flD�����T�C����* �$�����p��\JV`��������K�ƶvVz��+)i�o���Dasv�����0wX�"�s���`h@�(���r��#�� Y|2Zx�7�yTMrw���p/X�B��n��mv�y�݉�J?������K�8�*�����M��0�¨�:h�&.��Zе��^%��=)�9>l�/�T(��^��1HhsEn&"�D*�6/�g��ṾGRi��'�k����ޱ���/�W)iOl-H�n��z�M�𯲕�/���^�
c��$����TK#�o�QQΌH��
����x�[o>_���@���
��1��i�'�D��Q��O0Y��d1�>V���5�ݶFu�����+#T,* "�ڂ�w��8|�_CD�� �zݫ�_j8�r>ڲ	H�ܹ��,��4���Ln���}�Մ f!���BFhj�}����],=o�p��X%+�/��F��VE�,�=��5��q���#��?X�*�̵�3�� �4��ї�̍��su��j�:�1n8k+Q8��rXaw�@�aO(Н�/�<�u���V� ��E�tH��׼=� *r�� ���LV�2����8��riV>5���)1N��B���/	28}5��#�gzQ,#n޷��C��=Ǣa�3a�=8�t���4��Q��u�>�_������_��/�L�>��U�����m�T���q�"Pt��h�}��� CPfah!SI~��V�ar�&{���z/����̗s]-<�vC`�	.8H\ !UY3Bl���z�y0�;阇��a��UZ��7�0!|v��H,�{��w��޳���>+�R̥�d+s�:~���b_���d�ks��r�p��x��U$����c��\����a톐7����d��;6Dn������ׂ]8gLݒ7߃&	x ��=�E��~���b�ś��t�}ӰS�3���7n�pó<�-Y�� ��gS4�Ij`���w
%�d��}���A���u�+A�G��u*N��Xߎ
���Ua��C�y�Xx�hv��L�2���B�[VM��9��=8��VL≃h��e�^"W���r�k,����.�X [�:qV��i�@���kg��q���l��=iSHJy�	E����`�ٷC�
�^\9n1e9__}�\�M3vڷ��?�S�0�׳pi�8K�.W��t����4� ���M�e�z+ףa�!��ߢ�մ���e�T�@M>�&jZ��0|�c�p��R��h�D�]M]��B���0�n@����?�͞���'0LKC�ʳZ5}�7�Йgn h>ޛy ��Ȑ-U���O*��{�P�nf�������ySJ�[t��h1�Gcҡe����1��;B��(g�q*3vH �l!9rw�����2j!m�Bv�3�E�I%U�)p�,�%����7⦳!����"�tZY�8�r�ڕm�K�3e굞Á_m��;�<�BM�_^(%���z��zs��[EO���\����H�M�:�� �_�-��Uv�a�3�
M��9�¨'z1�����"\�r���C�m*�A�RT_=�w��G�+=$uW������.c.k��[(n�qf��noqGF������C�ċ���9e{N����<9�1���@8��9�H@G�n�zF����d+��{�Z����τ@��4I�h[��Hct]���%�\�km8�5�w=!!�5Ӊ�4�7�>����Ab��d�_pb�������Q�w�M�T�*�����?��fo�1Dr|	n'-�l�C�)nj� �ˏ8�~��Q�X<��k	��^ �(�<�~�r�'��$�D�}�,b����م�̛	0_� ����	z��x.֬�gn��m�c ���!Y�L�D'}>l���:08�8��v�����+���ɛ�	�C��\��R!�j�I|��SN�&F	���9ϸ^��s|SS>�~-x��r�Es��P�b�W�?	��( -I� l���� �e	�F�7����"�Λ���s�?_uj��V�y���8��s���U��-��Q���3�X��$����d�~⫆�s?gX��BZr�ױP^T��m���S��p5�[l����o����13�=M}�M�%O�D��n�4��ﭠ]o�y����J(K��VG�Պ��O�^b�7�S�0�ѓT�΄����b,�M�NK��z��K��O/L�RL�C��؜�Pˑ������+�),�-��?��N\��⃸"�W��ԙ��Xx�|Kb`*�9vo�NU����6���W����bC��h�1������4+͗��gM�)e���o4l�"���>,��d��豭�#�?3w�a��?���B��+K�2�(2d� ��V0cK1��Mg�?�E%���8��P���[�!�H����t �wto���������&�+<���p���H���56`X��f_^�o\I[����a|�ç�ö�&�f=�%�����=�`���F/hi&��~��X��)��+�S�'�~������=7
 n�