��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ��5���5o�h?\bv������Zr]�M�wM��a!��6���R�}���h���ƺ{K5I�*�q�p~"^g�3��j���;�ul��:m>s_`�i��wi��2������hL��ۭu�+U�u�.R��_�o���%�t�|�H-�*��I��x���yiI��`�iJk��B���e����O6��k��;�q_�׆�Y+�M���´}��E7!��J�Ż���p��_U띕Pݻ@�݅'"`&�1�`t�z��yE�W�z�Ͱ�NBi�YJ���VM���T�y�f�rf̟	�-M{�>!:D�N�9��!ċ��A(�j8����n[	��W�u#kNn�.0��$�Gݿ?&i�h����0�g�kq1�;���;���D�,]*Z���3�>YɬK��w�c�hx�]�B�d��ۈ�b���Y�C�.�e[�芬%!-�~�Xa7��ؤ=��7X���q���z�(��Q�P
�!_m
��"y�%��z���^�PS��N�T;������o�C$��No�qP75a�yHp.=su]�B^��9�u�oP���Y�VƎg�嬧���^ʑW+�C�BW�52K�?$#j�PXƝ�LGG�c�B�V�s��l�$J����*���1����h� J'HUg�|��P�������M�{@.YT�Jb�#�Bѓ�refU!�7��A!P-�O�Yx,5�u���N�Cي$#���v�հ��.A|:��Ec�-an����!������^�,3�"��ӳMp�T�֜K�� �#��/~�� �gvWRl�L�c��l�\Y�Z�'��R�"�>�<^���?�/3���c�_�]�EP#YDc����5@'�/��r-L�������^e��pH��G ���3vO�)��Mx�ܞT�z̀�#`�Ye}�8���c%�{����0]�����2%�h�[g�=o�-��nx�H��7V�V�J���ɐ����'�th>X�*?�-��6�؅Pe��\�$m��r��4�,���ҏ�4+ y����8��F9�oSm�~CԲ��LЖA_c+7����KCE�;�̆;[Jb�l!�~'%1�
�z�x����yd�żZ��mg��g����c��.��=r��X��m�1q8˔3���7�� �PE���u�?��mS��(�|1�D7 \��E�s���)��E���D�Fѫ�R���u����D]��;�]��R	R���
��kb�2$v;B���]����\_7�-�u����	tbN�
h!v����C���.��`|7��������^����()X�2�u�߉���kȜ**Q�����\8���F#b�,-d��͢�fH�ܭ��o��iLK�۩33"r�e�|Kwh\�A7)�^��ꩂ�UQ�QSXp������ v��о3�A�"��	��_�k\��]3Vdg����1��Ӊ�[�}#� s���2m��\���K� ����<�;�K����P߰=�b��P�fj��m��Ù'�˨�~�����ׂ���#����c�'��@bGJ�s�|>i_��y��[�����[]H���2g�ΑdO~^��E���k ��I��A�Y�B��Pg�^��g��#!3�{-e�
��P�H:���O���I4��}���!��e1z�Hg��[���33��?�w+8��ZH�X�֠2N�FЛ
i�J�����/�i�ٕM�#O*�^/)�C �������`���b�8u������g.��r�uU�c����;͘�y�WC�@�[;=��
�x~�"%N�)X�(��$!���d�k���F|�~4:D�����+c`�@�m!�OSh���zy	�'.;��	��R9ڈH�ݑ[<S����=��+- k@�?x���d�ͬ���k`�%b��
��ڤ]��-TD��J@������b
1Sf��䒰��<*�t��[w�`~2��n���^�[I�!�y����/�8�t�R�d|�>]�z�*��-�,p	/h�jfK.;�,�E���-c�?*�*�G"�m������!���f���yZ�idӆW��x>V\+4���@A ׃0׌��O�G{Yp��$M+�3��ݎ����ޙ%���sl��L_�����̲P�z@�=nj��jP74u�6xk�%4Ѥ!�'�#��z�W��v����=�����E��!�j7U���y@���v�j^������0������LL�M�o{��i���k���m*�{s�2ٱ���JI� 셒���wU��nx��TS�#I<],�P"�?�ϧ�(S�x�kA��-�Sv�o������V�pZ�[�{���m�`#-g�QB�v�I�
�����eqƚ���5eO�
k	�F�an�Ya)�&{�lFߦט��t�&(�S�1�b`x͋~�<�o�u�^�m�Ԭ����U�5������a�hu��x,���rM7��H�/c��8DvI�c�՝��
y�����*�:�2wwpm*�X~�`˵��'��,����[���k7Qyu1�SȻ�]�_��'uK��/�r�ǫc/�}�F$��?�C;e�E��wR�#Su��[�U��ǆ��YBC[Fks��:�������j�R*����R�&{� -� ��wT� M��d�uG���q��=�qI+逷b u#���-4���	�b�~O1J���)��W]�{�D�-J~_��Q��qi^��Mr}H�ޒ'���lE�.��EC���^�F߫HMjZ�"��}*[�� �yH��/�+��)���L*����;⒅�b��B�`H��u�0�$@�#�V6rӡף�E�ܕ�y��� �_�>����"Moa���M$�fc?��).}����
�������?6y0x��z?�p$��-yȄ-��3��P�kxN*,aP/AҬy�?ް-��t)�\���P��.��E0f� E�(Yv�[3���dy�ȧ�؁�V����3q ��)0~���"����$x��TSM=be	���qr��9�S�+2�|�ے�����1Gh�m���>�S!��WCn
����Ø�n�k?���i�k\�n�RI �����Q$K��׹���-u"������>Pl�[e���1�n7:i��T_�v;�6�u�	�<(�N9�DC�_�_��X��7\��p@��|b���kL�:������w���4?	$}��?>�@#�,�/�(�f�Hs>�q�/Gj�����5�Uz�؍:�ł�r۔ga8XMlh�N���b�j
�&��
�	�kIY�][��\���Έ����ǯ�G�ʊx�?.{��k�8�tT�R��Z�JYJ�W��a��&�Y}_<F��Utz;��a�˳SS�y��R56�;q>FB��Y2�*��9��{Nq�.���Z��f�?�{Q�)�Y=@_D��e�Ra�mUk3<�
E*<E��qɟ��Ң���(K4�����d��X>ƚB������dZSd��(�=�I�D�ET4��:�v��7%�f���l�y]W,{�����Q&h�j[T�a��/�֩��4�����()#��v�Q��
�-u�r��r���u5U�l�޴���6R�^-���Xj�5ڦ�+�1oY} �"�NTE2��g�(� ��%�H����t�iI��2���5��`���1G6�i�h9�i� K�
T��<���?Ft�������7�}b��c:��3�Gtؑpq����$K*.��e�hI�(9
�.2��������-�u�4����6d�F�� �p�T*3���:�k�&+��H �P���������E)J���U�,
��_���,gN��Ԣ�d��ΰ�c�f3����������h$}�܉�������7N�{��)��өr-9��mL"m��z������v}K���s���.S��j�T6��:�����O�aL�[��)޼@J�-H����}��)�K�����E�Ənt3���^*LW��w?v͇)bq.tł'Q��]_�������m� y2��y��f��JV��h$��d��)�|�����Q�;� è<�D�A2zH0_���}�
�PV�4DJ�q �t5������|�J�K�1�t�|���[avZ�/��\'�1&�����8m��u�G���ve=0v惰����X�-��~������\�����>��j)�c��e&�H{��h�eg�����l�_�F`�q{�S�8cl	JUO�5�f#�2y	
ϻ�tq���B2,1Uo�33B�4��|���UG]&E���_�G8f��,x�!Pt6��"�Z�
�EUQ�atd�eT����t3��(��<�c|6 W�Z\��<��;���C%�������C*����zy x�N�W]W�{[E��.�,��p��>�'�p>H�y���_j�-�gd�ړ�A,���AP٫?ϊ��I�*��n�jWK�NmW��qSΈ�\��q̮�p%u	���=��~fR��ӓ�p�-���#W�1*$�� ��W�����˃+��L�߫Ā{�k`>