��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_����m�e"kxu�Uٲ"#oB2�-g�j��h�p� M T�(�P�+M��&�[���+ۓmU��a�Z6Y�X�I*j�4E�#ل�!��0z=�^j���-�՗���:�$���_-CS��'�+;�iu�u�t���h�D���}�Ϣ��3ϧfQ��Yy��[f3�[aag�x/g_W�}�}Xw���8]ҝ�s�(�8���-��H�L�6>���)
o��ӽ����A���?:�J�dqO9��[���k�Z��QX�|��J��d����}�ǲ ��}~�LʄE
s�	�Z��I��u��N(�������)���X]Xi|DR�˿�S�>2�]��]P��(o���RE����^K����@�zM�v���CQ*5B�A��
�v�C�n(U��h^�҈�Lwo�V���ʏ��c]�4�����i[l��Ӭ��;�L��qɉi����/􁸔=�͇�,C���_d����d�zFO3��v��w�L,�qv����G��g�d� 77R*&7LT�h��q����3��p'|���(@�ڙw�=�\��^� ��b��+M�3H�^nn{�vY��-��cfV�h�_���6��n�v���n�|t�SX���p� �9?�>�P�q��<$	x<c˫b*�B�⑛��O���͘cOMD���ѿ-�Y$sVL�.t-pp�� .��,��N�J�(q%�ל�C~',fV�E�S]�E�\0������JJ���9>�Ypq�Me±"a������@'K��h�$�UҴ��m��OΓ+�S��p3��ހ�U;����[��ݽƮ��Ӑ�@��&��}��M2�lb�[iݳ���(N�����Θ3ۤ�k�7g����C�<`���rO������&����Q�*�P�8�DK�C?ඇ�%����,) D���'M_%�qy����ǁ;���V`��纅s�ރ����r8���t��p�� S�9w?Sl��������u��M����єW���`�����i��?�\R����=S��o#�,GK
��B�-��y }����.������Ʉ�p,x8�1�bژ;]e��=o�Z����>�-v0�
γ0f��b�#���{���L�4��ly �����,�N�k=o���։��p��M�>�'>�#J���&�|a� �~��E�����',�t��ef.�~�c�az�kw�o�3�$k����D��i�%t�x��1�����x[p�EE�êFL!l����'*g��r��#u��6��3�<@�Bi!�\�t���˓���AK)��qOΐh����o,d�A�&�ܭ��`#]ߊ�!����Փ"��1��rFG\Pƀ��05stW>�< ��1�U��'TFR�Ё:��t}��R��T��:�4����[[b0C���[=��o��T���ƕ1���5��'H��dN-�r�¸�ْ�G���n�Dݒ�)8��J�ʢ��1�K8@�� �yn:c�/�lc.���e���>����t�SL�МnN���6b�r��+JDgݣ{	�8�E�Ǝ�-�5�{�$�n�O?xt�p�����K�b��E6#��������{q�z(5��~Ƿh5"�5��t���Q�+` ��q���=�>��;�T@������)?�?Z��m��c40#��WE���:'�a.���Gg=�E�ĆP��?,��ǖ�
�`>O���۞<�1
����g"`���\ ;&w�Q`��dN�@q��[�LP��~��Z�<T��+|ek��3�:�_���,�n�ʏ-�9���OP7~���5`��PR�H ̀:h��6�_񰊤�& �f�M� �t��TV���CU"�@���Ax���i,�Z�j/���T7�i*Z��;�@v�%$c�x&��6���x�te���>pEk����ς��>|���_�yqu��Fԋ.t0�9(��.SԉT	����<����o+�"�=���,��N_��nV+�6xE6"�8!=��:N�,Ag��z���j� �n���z�QG�^�fTy�U����)�O��~�}��t<W .w���CIi��*���K�qN�/vl�ڵf��񡒫_�\i�"�tM��aT������հ��@��|D7Bˏ$���MC�^	��<�~��sז8a�����M�̀�;x��~q�ڄ]US,����7�Ց���P%�o����|D���#���&.	&& *%e��ف�&�&ҹ