��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf\�|Vv �|�
����:C�q{����B��\�e�w�s�v�����ē��ZzkTqk��A>��4n�pt�3�AƓ��F���$:g���2��.%�G�[�P��U��B�/Kݠ�os�ΐpBOd2߻���G�)I����~y]N�53���y�����pnGpj�Z�cF����/Ѿ���� ��\�E��7��Z�E�΃��~F٥��������Y������c� `T���$4��^�y���oF���{�vn�@��y������S,L����	�BÎ�H��[�I�O�,ͱ1�Q�b�:h�\��"����K,��rp�g
�����)��;�/�[9hqIya��XnFʯC�)cɛ�:o�J���H�m���tĖ�vp����	f�)��pc��F�}�瞐n�Ƕ�݈[f?����-�l^�@a7�q��. 1�=@Ț�ٗH1��b�rGl�bX�k�d��]��z,4�� �7P(����:��i����V��x����4�M�"��	�'�_�E#9��j��y��������+My][?��r�-~7\�gFbJ�G�I\��u�������@�`��vXBK
�$�M�!z��C���TF,/�͙�d���|â�Z���5�җ5�G8�n_�د����\yѳK�^��7U@�#1�U�`n���׍�RU��~d��bdv�y37y1h�g�N9�앩oݸ�Z�V�]r�}(��]́T<mÁxf�������c�|����H@�!��B[1�"�S�<��x��]�1_'P�8У��?1k�+T���|�z�}�W0F����d��#�o㸮����#a����y3�!a(�}�Y�p�=�B9��I�6�;g���x�_R�"C�ӊ�'��C�<b�$癄���6_�7~��k�྿ #F�
�Ĩ��	��^P��r�S��R&�_���3!��ȑR0�5Ll�v؅y�����ѽ�}�}7J΍YR/䳂 f��T���4�>���D�j!��$�Qc?�rn�sMw�R����z��/�<�Ԗ\�����3��JqC�O7&I�Ρ��lXEf^	��
hE�����]�����{�����y�c�oL�B���e�]�#���Ƚ�}�����<�ǌFv�?N�&[ȑM9�F�b���z;"���c�Y�&)���r��]��}���x��&9�J8@�UG9c!ϛP����ә͆��N�2�Y���S���3R�:���߬_z�wnɘ���F���-\�҉}~���>�&�Ȉ�ws몺{��n�&7�r'�%�4��r�tdMh;/�)�0Ĝvٺ�UZ4'�VK��u/
����epm�Ҏ�
��j��.Я����_�-�^�P^�����%y�ǆ��ud��`�m�q�]�7�{i�Lki��������C���j����a��_S�>;a%�{�k��Ő�U��Y@CV��TKK|z��2ѣ�Һ��xcշ�Mߝ��f����R�U[:`A�a+=���!��̺�O3{=�K�T<�k����fN��(Y����J�>��/I�ߤ��z
x�C]t@��h	�H�S$�8t�K�{�<k.B^�
���Z�|]���H$�q>�l]�"���!)�q�H�©�>e�5��Ĩ�Xu��/��
��� ~�4�@A��*D8䆭�V�k�L��B�Ŷ �msĦ�]�ܼ����u�d�x��4�V�	�6ne�`.�ݘ�6�;O���:؇фe��1�J���5iMq�`���z�)��Wb5�Z��_#wZ_8ҧ����,9@WI��:Ͽ�m�}�_Sp��I��S6,?�0|�ǫ�����I������6�Zcai��{I3<d,e�.k��·�A��-����.��:r����ϬA:t�rQ�ji�*�@
�9��$;,W]MN�G
d����@H*n=qp]��>�S[���<a���JIܻa�~��<V��Yo�aP}z���=�� �HߥBJ��OtbG>y�����٪���k��E7����* ^oCI�Y�p)�Z���U�y:����ξ��� "��uM��� ڵ/��e�.�!�)�&5鯚<�4*�y�����X7�ل\�pxΣR��rʟ�ςTS&m=z��F�x=����_0v�]F�o�%��'��JΡMP(��$LoD�C\�N����S���O"��L�F_�s|M�x�z
���0�`�t$M�W���@����7��I���B�6$I��y"��νGY�=�Wfu�i�f�������J�yEt��U�5G��A�g7�����˭N1aǢ�"��j�'�1��2��e�f��u� �v_q�Ijq�x�j�Pb�l����)WD��a#=_��ɏ��u�DE>�.���Zu��{6��X=����w���:���4MN�ʂ��b߰6����ѵ�AWL�4y�5-P�����jD�9.�5���B}���C�hֿoU簺��3�Y��&�_?C+�/ZἌ�Xtvn-�wH�>�SY��%_�vK*�]�G<����P���4����F'k*�����W��Rȃ����ɤ~�0��Eq*:��̼h�έ�rN�+��A.�4�E��A����x��ծ�p)��3�DB��������9ۤ�%���?Ԗ�h���f�A��1�W'������D���i�,޸����Y�:$7�֫:N�+�{�U�$�m�s��!���P�<b�$[_?��Z˜SI�h2�GX}4�dm��v.���ƥ4��?��>��Q�Xq�t{����'j+j\=T�-:l�9�*H=��q��˱��s� 4
������Rj��~�j�����R���ট��l�\ٞ�3�L4á{���L�$��M��R��+�u|���+�O�̣�P��r��� �z��v�@j7Y�D4�FW����HM�P��꽽�Nʐm��J��%�t��hq��}�9>O#^���p��=XQ!�gO�����^�qӑ
�����>��t���}���-J9�R[��ր.i��!�N���3��b-)Π��r��_gZ���>���>ь	�잜�Sf:1�֐ZƲ(�؊�ݠ�O����Z�`��'�s�J���b ��]��>�I�/�(�u�5\]�n W0s/[��������:��*�J�݅j@�/@Uz��o�	%��F�d�W��~� ��.�@�]����S��^��fW���o7�O ·+���`��	f۩B�C���t����C��qۍ(�o	0fGv�Y1���!|Q����插��0[:6�S���״k~'�
�3/DqsB00\�-BL����dN������Js��,�v�j�EB�6\ee����i;�n�j(�ߘ�8L���?� K����i�S��5���G����v�{��dv��~�%)5�;���jv	Q�4 ��8z7oT-꒼��5����&o$-}DJ8��zN+f����V;�)���fP��g�3����"{y���`��{�1I8�#�bn�c4���dv�h�=�j���\ŦC�
Ai��ފ��r��	xTr��b��<������T�:�>�$�(D�`��Fc�-9�:����W�tn������L��D��׫�]��S}w&[��β\.|��vh�>�n�x4B���^���<�Ο߉��&pކ���s��_<�R��rf,��-Z����>���ntӷ|�J$��	����9�d���B���M.��t�w|�~,C\gy���$G�����x�M�.E�j���,�c�ߙ�?�nH�R�؅��@��uVp��-�J���9�B>k�-6��`祖�Ԕ9ωDM;�HϲCh��Kڄ�H�zʤ����1�'�*��������x�
U��]�i�S%�hjR�}�)ג��[���ݣ�{���U��Q��t�Ԃ�����1d�I$�ΩĞg�	7w�1aE�A^7 �[�!j0��0�8�G�<ɏy� �`'�������R�Я34m�� �������d(�5c����s0�K
--pkY�O��_.�"��n���e9�~��!�N6u�Z<v�I;�Y�М!���H��O�̣�����P b����?hD"v��(�6��{k���4�v��:"^�D��u`��P�!F����
�2h[��Y"X���\W�$��,?n��-�~*�&O=��Ù���H�aIRǓ�Ђ���'�8ƽ���Wz�x�h��"J��i���	�k}Ġ�T�"e��-�ٷX� .��5�U羝��o*rs����L�'"��a���	�.ʼ2�X�Oߛ�E�Yc�߆�Uj�?��U�� �k��i�=:3�݆(a�����n?����¯S�&$R�9'���k��O.�9�����g!�\�#����V	2����9k�0i?������Q�r~��9\8��1�S7)=�lp3�}#C�MT���]�H_��CКml^���L�(��kz�w|�/'�6j��3nG7�q�5!*k��.�C�s$=f�YJ*���γ��Q/��'�z5��A�g�E�������f.����e�w���ʌ��^I#��8�V�ͺp�8��K&ב�������#s+��B%K��8���pW��R���Je��=:r�yba�o4w��^-�������v�5���;�$��0�>b.g6� F�2	H6����L;c�,��
�R��sgzH�P䒻�_X��x#���?���?s���[�m��ˎ~���<V��˿I��&zY�M�GS�.��fhPc,(��u���'� ��˱��͙���C6w�w:���E�&u�.�|H�w�p+�3�r~����l������_�F�ͧz�Z��7��[W�z���2j�w�������L����ʬ^�#�uU&Y}����Q#E	���OXN�U腉�B��Cik�����pa�?�Z���K���-�V�>����8��D�Q�(��G�%��\���}b��iP(gA�y)���D9�}H,��H�S8�?��YIΙ�Pl]W3��`��9����7�����S�# rL,4�d�%9��&�>�C�g�[��_)3l\��!�tf!-<{�"F{ڝ��y��h��uFZ�r$'�v�FMT� �VA#ݦ9�wIm��U����w@Rh�Q4ͮR��7o<y�V��X��O'J�׉(ݪ�.M �Q�F��ƻ�≽˩����A���o���=�Sgo�N�7������72�?�Y�\�Si��l����T�,��?*E����S��n.�(�!s�5��K��ޤ��$nw��#d��[���!Z���Ǘ����9
*F�J3��Zi-�J����M$���iv`�;C�?:���r�B�g��#���k�=D�a��삊\R���߸}�uu���$X�h$`����j�����09�+A����=k�:aF	=�$q��Vn���!��� �^;���h}�	bM �Ģ���Nk6a��27�u�R�<;�i���ÿ�n�8�TSv#��e���&���WGLt���bv��G��G̰�6�'S ߯�~|fZ�Gh����K]m������Tb:��BԈ+rK��?�ܥ)��~�f��}9����
����ƥ��%��X�t8X���L�G"D���F�� x!b����X6�t����<�w��p{��4]�]{Z66@}�@	ˀHɆ��hʙo��s/��0�i%�h����e�:v��7�����/�%��
L����S��6A�1���@��e�8��8����9�eo�CaAiT�@i�|�7r*F'4�ϷNv�_I:oc��A^\� D�OM!a\�%{�@�3���'��3�f�D�^U�����e�r����5���{�V�d�O�{4����g��P3��z�so��w'�~Y��v�Tн��3TN��+�o�ad�x�@���B��#�������։���|�aO��T�dA@g��1�'esɡ8���ֲb�?�Z�\��82,�2P��R9���a�j�����R'��AX�Y�귋3�s�a��E�>W�:���[v���xS(�,��SL�'���}5�$��n�W	Bƫ#�=s9�&�?щ)��s&操�6�v�ޢ���ݍ��D^ɓݠ�u�m�/@ܱ�?����#:`��ȹ���d[e����5�z!��Ƨ0R�����m[1.���cH
g�7`���9f�V�^����Cw��Z2|���tW�3y�W�G�-��D!ˁ��#�#~��v��ҭo�[��l��l�3�>�Yl��&��'��. �{�ڬ�%�+ER�E��reNi]�ma�[2g�u�D�HF��.y{�t[|q̢�,���s����xh�Sr������L����p����_�w���ZV���q�Y�x�n����Uhq�����e���q~ь�qŔ�t�p��`}a&R���j�<
g ۙ=�#v��B!e �a*��^cP"���81�~�C�:(���Z�G��>i`	/(�L=���_U	�)�YӢI�kYY�wh�T�7�x���eh';l�~&��j��|7�\vvS?�(�\U���x��@+�,�b7 t0;�^�,����#��3=4��F^��dE�[gz�l+���7�'�J��#ڵA�]��I�x&{Ԣ�	Wr���g.L)�Hf4y<u�6Î���4��b�v�S5S�Il�<ԓ�ĺ�|���>�b&�������>�ݸ���2���x,��t�%5o��}�1럷�ԩ,q;%,��)N�|��$\=&iv���[j�2�$1�e4�{R� �"�z,�r��w��?ӟ��\eQ*�f\��IF����w�� ���\�䡬�y��RN�Vf�T?^dFA����e��+��u�z�����������( h�7�o�,Ɂ�1?��$����^�D�>��{v�������7Q�K..�s�����1�B`�~)�v���ҍ3�&�׼��֜�$
�˝���Ws�{%�bX#����f���/^3(�����x{�
����.��LH�>n{b�(`~���R5T�]�IK���.hm+K�/"�>Eο�x�0�v���{{�3����VF�1��1���T�.rgq�f�R2�W�����/7l�����زγ�L�s�k.}G���1�V�BJ(C�	�J	��E��)��B4���ګ���l#�f�a��E�^D�dL����R�� �x�z�'~��I�MR.������/�4�k�{�r����l��ͅ:v��}�d��8P�F��ۘ�Cf�$��?��Ή����>VOϲ��H�c����X�/g�
�0���.t�e�a��O��Dy�o��.-6eҐ�;S��\/�GO���	���p7�v��v%����O� �ޖ�\l�qZ�*-]�� 6���K���%�Q;}��x��a��:��s�e�(���������||����q�b�ṱ!q*�[�z��{%y�#�^IΘRB"�����Ȇ�s>�,s���1�)�7~8v,t],�XvN�Q����S�����F℄Gg����ң�:�j��wȀuHR�G��kR����k� �B@�e������q��Y��3��᎕��XE_��,:@�6��f1�!����R.pO���?I>'�KH�/�p� ̾0%��`�G2=�A�3p�,F�0hB���]9�p�������N�G�w+��EN��]g6�����x0،���V�Klh�}3ʤYh�����x��E�1K@��BY_��Coz�ΞZ3���i��R�|ڇ��x�)�m�����z��x=\���!�n���L���� ���l�A�� V�2"�[�X����^��1��c����-\�p1t������	�$#��c/�:��A��0phgi�v	�ƀvQ��K��~p���ֆ��s������-�z+��N!V�7Z\.
*ʚ���2#a������w�T-x(�����]8�,'jZV�@��1��ݤ�6w�;����ED��VG�س����8���ap���(�Mq�Z>��p'�Q�ޘL ��wzf�EK`�>����2i_�z��2(��KNX6&^�}p5��,7��~u�@�hq��/��C���:�9�-��QD �B硲B�Z���u{�Zb�27ڲA�D܏?�Z�G�qt�C�J�	IX( ۚh�18�h��W`�����?����E������OG�y��V%m����8h�"P�N���!(tz�z�\?�B4�mpB�3bȯ�L�ʑ�iJ��j2Rr-�!�SF �<��5T�eC��	%:blU����]��`2 �?�ya�Ǫ����wW��Ĺ��Rԭ	\t�:��5! �(���_��Nh���o��pVF�4�Ubh�9���e�jZ͒G
�8��P7��f�����Xv�t$2?\���c�nQ���g��U�M�5AK��b��EQ�i�q��c���sX��3����} �����>��*���?D4r�G"o2�  #�O�X��5������o�,I�RؾBKB$�����GQx}��{bH�˧oc�XΟJ��W�,���`����$���>!��

��!l�-~',88�Q��8* �@��7��T�9�(��������en<����c�8�Q;g�:HQG�b�����KV�� �H�a��t��->��{-^!*^��"N��G��"���m�����.��/��A� [�(^t�0*�ӟk�_�柆��a?��d��1ˡ�Q�͆gJe�lI�pH|�0ߤL��K��%ge���������?�-f&�+�.��&�|8�[��:j�G�V]/L����G�,��e��k���x!yo+qW���|�c�y������iO-78n���2:)r�^��6�Rau�3�����.�w�<IXg���yb��%pK��kH��m\{J��`��B����=�����2"K�lt�l�n"�!���W�� \�A��k,(�C�R.���,���P;��/;��X�O�b�,��%�)-���_�GG�r��N+T[/���;��`��|N"��|�������k-�6�v�c��nᩝS�#C9��ѽXb�i��OTm�nރ[9e0����S�����t�$���%�9�qjZ�����A��P�*\���qtc|@�k$�6D���%�ڿ�{��T�D���0���跐ݷ���7�#jh�&ߜK�kX�RGR~�-&��U��V������<��
L*n]B�X�$֜�]�����~'�vێ�d�sϞҌ~�7�����3���p5Q��]S�@��4)#�5��aݴ��)lQ�];��.�N�<�<�S;L��we}�p[ɳB�]��&��V2��z��_�qWg����o�{Ŷ|���_<�P�gV��o?zΉ�B�~R�M<�~��(�ŏ�|�b�G�;^8��H
o��`�\X�ȱ(}3iY��%�)(8��F��R]N�*����s�����[�I��)���W��`�CT��YjřR�Łta�<c��D�晟W��p�t���!���G�ַ^h(��4vV���0�U���b�Ǚ��rڒ�(B���1��h���JO��J��ٸ��D�����_��{?�<���;�S��U�Ứww7maV#��4���З�W�b�M1�.����뭯��l0�p�&�ܖS�q3!EoSQP�k�V+eή֧�����K�֥7%8	1'�1RHz�2~r�,EY2\*���@�֬� lt'�슥��3����!��v̈M�V���P�5�Z"\��.���$�!�gX���ݷl�~ ��$���Ϙ0 砑��HQ��;9d0�gq��u�A�|񰃊�Բ�~�y�r��Q�_�fܘ����޲�ޔ7�I{|g-�J�FK�<CN㤍����W<��ʝ/;�>q�P^��Ά�����oG�տ�fC}�tL�Ly����ԣ$�O2��R�b,u3����,i����_�[7�O����P�Iw{��j�0�L�;e!)@��4J�92."*�o�w�:�A� �ܽE�!���@m�e�K@�����9� ���6E�c|��Ⱥw���B��1\���r�ht��@���Sլ.	ӡ�>!�������ZE+:����+�;>P����rXڛ^W!� Gv��K�CPi���H�I����X��m�6��;�K���6�:Z��[6
%*)�kY=q��ї������hݳ��tWP��2
����IN�+d�@Qd���B�$��g̎9<��;hb�2�h��:oxߡ	�R�y<���a'���̝{o�f�
��K/[3:6ހA�XN����"0F��B�i��
��F�Z�.]�����nG�+��	51|��+A��.��	SN<�$"��On9�K��)��Ư��-�/`b����~��M�'�0�����ٵ�!g�<pv�4]b��k���4˄��u�I�>vj���-�����Þ)*v�y.��x%80n��V�I"�q}�3S��Q� �(:޼_#��2p�E��֨��9�-}������"����:�<��