��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|��&���i} Ĳ?���F�v#�=��te�|��Rd�Ѓ��'n_�H2h04�lA�k�r���5u2����6*��>v���V����牂d��L�E�ͱ{"�s�}q�Q5�`�!���edʶ�_�4xɒ�,o��t*5��70�f�p2�pn�_�q0�Ǧ`i�[H�����x+��f�X�YW9�x�w�:Y��)�_E�k��G���f ����X���T-i�g����V�򹨰�$*0��k���:�$��q�W�+ӹ&�!_�G�&]o�׋q�v˵�/�ISm�<c4Zc�9�h��m�������-���V�n�O�'�Ҥ��Iէs�Y>��ʶL�˼�2������� ��tx_��&Ob�]W���,z���^?�a
�yI�\"�i���`{�h�ߵN>MtOݼ��{�p]a��݈u+�ͬ`s�ә���kh{
�>N��#��b��[��c,7���i�i�N��F���Eeo��$���r��dU!��g��6���ͦ�=�ki:5��,���{�*{k��4yDk��/�Ee�_-ݾ�q��z��K�����a��2֏�:��(�ݡ�<������C�(��T�@0B-W�o�f�6�w�V o�g1\p�P�%�jGt2�㵜=Roi\�ۅ�3~�����:�sҩ7�����D ��֑��o$,�{��bD��]�[g�s������J����/��I����8&s~�\�05���_�e)�2�vu����P�h����O[�DH�Qh���b6�gI����� cJy)?@ePw�U��`����Wp����	������ip�	�?8��hʦct�I��Ƞ D��w8���}��A%v�({�ޛ�4��W���qU"k�1I��FbG\��h�)t�k9�`ۊ�x�.�o�����ɷ��d��/��?����ͣ-��هe��G�϶���](�nmQ�sn��:i��Au�e(=�\a�)զ��ą�&��D�M�!�}�͗���퓥���s=��z~���X�<�����Q�"�D�Q��'pc0h�N�ő�H�3���{a�~-��mqM�!L�Udu�͵��;��du��L��}�X��gr�`�=�ӍƐX8X(�fZ |�5�yX�B���v���I����W�^��M�W���>F�G�zG	ܰ%�tn�5�O. y氃JgN
��q��	���&gTcb�����7�}=��I���	��3|\7zE���~B�X��2T��X߹�|1+~�JX,5l���|5~�/����Jn�zZE�ֹ;Dn����v3sU�q�w�5�ןv�7L���֌�=������|�_#]��9/��q��r;Y��b6��ec���pJ���A��J6'�ߊ@"<v�)O������j1E)�=�����M@�[�WOG�y[�]gŊ �ia4��g_�]��v���2�S?7��"�5����n�u%��e#���ض��ws�b&V �*]�6&�=݉����U�$w��mF�����N���kЖ���=�o�Q�Q
����-���l�+�|<9+M�7)�(
�H�`�R;q�%�pz��*� �k�[n:�ԎwU���(��"� �LJc�{�;`�Z
cM�HF��cb�� �_qv=�	����3z8�������1�a�{{_г䍆5o���^5�����{�C7�Фˈ���&b��T�V�:�U�r��񸭵�4Čt�V.cC�o�'t���k��Y�6�t�}�U$�b��*5���?�@�z=��R�'�r��B��G"���S2׭p���`���0��S�	Z>e?�q�j�z�%��r��1m��%B���,%�Z�o�*�ӅZp��8MeRa^��z�TK�[o�P�9� �m�w����S�����.�] �@"(U�XqIY��N��|T����"���"D���P�Ƶ����O���������UK�O��z�So[.��_����3 �O[��	����R�D���7�(z��y��u��O��������B���x�4e����{����B�4�����CG���" O�I�kJ���E��Lz����d����y��+�H���d{���4]N��\��[B��_��
Oi$Q���a��������V51�G���~D��L���x@��Ԁ�܆Ā~x���_n24	l ����!"b���T�,|fh$qع���M��4�/A�Gk���ݓԠ�R��Rf�H�w���=B��{�D-��f�h��*�oD��DKlG^�W8T��߇<���6��n}�j����l�S���7�\~e��U��^��G+f�����w�pH9��a9a�?�hh��D}I���K�Al������̱R��b=(";hx��Y����� ���v����+�L.5-�;���.��Z��_ Īb�)O�L>2`ɍ\�ӽ�����~���oN l&3��b�Rzb�-�w�8�WH��eBڀ|�S
����_�/�t��z�	�C!�x߀��L�_&>Isd����E�RCc����xW��*Z�
=*B�:��b}2��G)�F��|������q��P�]���rPR��r�6s�Lk�#�΋k�h�z,�hR1�Y�%{ž&I��j�B؞�xeb��b�����:�j�(����4"��k�9�.���Y����N�"�?\k��y�4�]���k4�4U�1K��L,��y�d,_�8_�桴췎f����GuQ�݆MTLG��E;�Ǐ_[/vKز�nj�4��u~;9��	oM�9��t���}q�7h3��+0�I!]�}�Q�M����mЈyz/+��l�����i��߈�>�1�k�4N�s�����0F����5tA��'l�pd�޴�j�ڥ\#���P���y�+aI�J\R�&5��+���8t)���<���$�k��sN1�Jt~���{û�C���U!Z�_uA"��7h�Y����8�D����Ғe�uW�P�3��J��i�@�i4$����H��2�Mdrr�ȁ��#Gor���DJ�t5��³ʬA �#�K�8��J�2Γ�@���䒄QV�^���d鞑�xg���������-�\?+�Nc���w\i1���v���W'[�4%~m���Wo��cn*1R�.�����^I-9Iu�װ�5.�5pp�Ʒ<g��		ܺ'I�Ox0cQI���a��t锬�ۑ��g����q�?�;"OA2�?��]�)��}�&���1J]�we�>�+�Ph�f�L��.C�cw����Zy��*R�#
�4[ӀPp��X��ck�N\��[r���R��K���kXnpԛ�y��Y����ZJ��7bN�q�)��� ~<�:08��w�(e[���_���6Q}�')�b�U>����Հ�Z���ɜ�NiX	��;&T	K���2�� j�=�F�%���gN�m~N��z��A4�x�V��t/�I��	�}FD8I��L�ł�\]0���x��zw܀L
�aoj��l��F�qZ�RL�_�ʉ�P��:��!�&u�Q��$�ʤ�����|�2�O+��^�!'>B�S֙ݒ	%	�c8�	ABSvQ�]��r��$I�@{�G_��
�i#��0S3<�A�� U��&��Y֑��u�Qx�B�$���F�"��Z���R�3��$j@�i�� ��h�M^r��I�6�V�TN���&g���)���#�޻�>8�5z�.ُG��&P��y��H��o�����Տ�&{y��_�����:W��/�gJο���ar���& �q�!�Cx�ÿ��o
�?�d�Sr>��I��䏔�W��+TTr����@��Asc��6\�hK~���>�LV�	"x�F��5�{�X�Ѣ��{s-�_6�����kI<���,�J�+���n=���M������t������Z��^
�sE�iו9�h@�ϲg��W8:>Ǽ:�dt�F�k�8??fX�AL�zŒ�����~�n���~�h��Fwsb��W3#-���07O�;��)�����Ɩ;ic��p`���ss*�
��o��h�e���M	g����gxa�I�P N�OW�B�c0��/$�㽠RH�-$��>��������`'SX�������=�Mt�_6eM1���4���R�ӄ-5A �	��M?��L-#���Y}l�_��׬����o��TZ�Xt��{'aMrp(�͢��d�bL,�,�-K��q��?�!��e�z͞������$����dw�F�(�U�p���h�5��4*	�iy;zm�o�e�w�~*S�����	~5��
W�����R� ^@{���f�<=_9�FڌE��c��Q���j�'G�d���y�E�!�Œnߜ�H��2�Y�)��c��H�T��-Y�5��)S�8`�<�����" �g0���~?�b�Y6�i۝$�����/��;���-b��!?XX����)$�Bܵ ���f>P�ԽTdd��r7�K*�?]1	PBr�!�yk<W�,Q� ȉ}&�v���F�29fh��'d�?����7��g��M5��o9���a_���������B��K��g�����&d��_�4�T7`u&p�EszR��Պ��,@&2u��'��V=��˴�`��^l߮{d��d��\#��9�s�rT��%z��eF�څ���N�Ō�(�Ro���Z��?�Q�S�<�OD'뢢�clѰ�(���j�ΠN��}H�;�)c;y3�E��oa�5z�����?��a�x�sV���������My��^{��'f��������gL�|^�ƮJ�ò��nOEN\��s���f	��.ś����㵓���,�9��Ne���^��U:Ʉ>�$����1��Q3�#�
�yD$�o�e*G(s���w����Z�̕���q��| ����ʪ��z�s��KH��T*��lw�H��jZP\`v!P;�i���T�P8�O����|�խ�H�m��S3{���u%R�*;`��J�����#��,`CCJ!�۽r�a�u{	�-~hA����ڵ�F覑�Ap��w��Wa�4�s����.��� �S�B�55�=?�����3����_�t�G�D�lb�>#.��B7����S9��5R3d��Ye�I���#��0�0;�&�]o:�:���c��>G�a�~CT/s;R��s��F�T6��,�M��U�Kk����눕�lg[��苻OfukYzy]��TcE�=&s�r��!�x���ۻ���������J)�n��Ku�tM�`��6�]��Lߟ��hZ��HT��w�P�$��9-~�t��v?�i�5_��w�]K����7)��N�d�\����ц�f�Cp�]�:���#���Wm1E)��kg��xEJ+�%sޱ1]yBh�l���Į̺�kg߭ٵ/���VhX����szSJ�x��1����4uF\�'
3V;~ �J��Ur�6Q�|m���Q]�s�M�tY�[�����2�W�A`�:2�
��/��{6:�W#r015�@Hr� ����{���S\%1��,��� �i��/\�s�7�u�����#�hCH҄���E",����ᇪf��FL��	���p��W���x/=Vh��M�{����!ؙ�D(�A��'��~Ċ�dA�u��xWTx���rL�ґͩHY$�V��x��)D�#���>t���-����x�5����s;��璝�Z���Yc�$�b��_ߖ8�(��V9�6�c,4pWkC��'�_��O$yc����7>W�Uw��(��B_	 wS�?:T���P],ĲЫ�م��k��a���1�yK��ڥs`)~oe��Cx�ʈ.��/���|m_�fÅ�C���&^XN��^¯4{���>N2��̵�q�b�6�����%���{-�t 	~/V9&�P1]2���9'�tI3K�&�� w�h�Y�8i�Sg�/ ǒ�O#����[K�@o��n?�>���;��]�߿>�M�������D���<ιH�#��v���ʜ���-�N�JHyl��vns֑��'�9��hi��@#O�����S��Na�4F���IC�izBn;��N��[���Y�;��F�6I�	
m]/<5̷I~����ν'CP���OR+��f�$7��v�5���?�|�8
�s���r1�ҨJ^�I1$�F
Ĩ}w���6ϑi*�ƚN�7�/�:�	�l9� �T�v��̜�N.�9��������8�jS�nu����zG�3f,�0��Z�2��=����"o�0�ޗ�V�ʸs��<�;�ߤ��a岑p�ê,S�'��)�#�#8��E~����6r?s�> ��r&�؋}>9Q�X�k�����&v����t�`/0{�~�t����ڦ���㎎0�7�θ��3z��Z �Xѵ�i�>��SU@q��($�����G�����8���Ǵ?论4d�5�F�j/ȯ��$_p;�����kR?��S�����A�K�A�E��o~Ōn�")n%ed�Csg8Tٓ|r��1O�1�#K�fլ�{�4��G�
ñ�T:�IYLSm�Fv���$�3���N�q<�h����C�0�`_�>qv����A�_��eN@xt��\q4��i�k��l�yanx((��n���A~y�d}����i1�����v��	��,'Z��'j��do' A�+	s�jA�Dq����m��0�KaCi]�/��o�:�A!�&��M�؄��`.F���rO�ô2�Xk���v��\�y�����l�f^ 3� ��r�g^ ʬ�ȘJ�YQ[�5]������� ɤ�2��B���82�%����.o5,�c�=P]���p�1 �������ƞ�>����;�=2�'���c��$��lO�o���Z�Q�������{��7?C_�;u����˓���%C�6����e���>�� a��Q�o�S��c^���I�Zy�ki�q`�{9��B�	�I��6��y�ڦ�����S!m�4����}���P�{=���:ӌ������!�k	N�ք@ �(q�8}��R	�$��|O�žSOV�ohI% �/+��q�lY}
�L3��^�QQ��FC�๩Aƿe�П���T����7lF �G���G|���v�7g��.��@�;�W_��I�ɽ�g��L@u�����ڳ��?����G�bI�������k: 5�,v�xki�%�6�'�zjG�@[�?�����N�(6V���'Д��aj�����Ҥ�ү�w-�[)h�x�^^���~�p��|}�5���[I4�e4'Bo���~�~ު&��r"{��2s�״c7xJt*��)�Ur����O�ۂ�e��4�3��v�9�9$�������{/�^�6s�z�Tx��R� �[�"�2A=���{�4�����$��ͳ/�����)N�1E+"�S��YTǾ;�T����:�g]#>�9�bEL��H�5_�R����L�&�D:A�� 7`��W5;1���S�rDet��D!5(��)#�y�����E��1Y�,�_��;��u1V
��j0��7�M�O��Cj�5�z������9��YJ��Te�塰�~]/�IQ��\U5h�O�t����E[&Y[yjݲ���Hw}��B20<S���f8p ��\��G��4�[�c��٥R~`.�����CM�E�](!���Z��|<.9H�?��w�a��#��;t k�!��LM��FL^�����7p"=VVp�۟~A���;�Ч����-��j�ɣ>�Kq����Ս�:�Y��P�������/[�GP`�N��[2��n�)Fl�$������	u#���u���� Cy��u�쬔���Sh�D;
�����N� 3G>�� 7NGC^=]鸚E�7�]��e����iש���}���0��kN��ym���Rg"���i�ƈHX5��=�'�i��4Z��}xQ;!=� ��@]��wW냋���级�-y��I>2Сc������$�����l�#5�IX������ߪ�8�vR��j�����s*O{��:��%��iJ_Q���OZZ|�H��JÆ���۳�&��6���̘8�cp��иx�ޟ���6$���v��|�]�{��4�Τ�R��p)i�/�6�p��vw�Up(����7�|k��b�#x}�%5��#��2���ͣ���ꈳAh���jGrR��[�#ņA����jc�d���jyu\��Ȋ��m��i5a^�{6�^��>r}�lu'�<�>9fx5'A�����lC�Mm�\)o%#+����g�����KH�q���#!J�3�c�'n�>��KU��{VL��9[d
=zi����5�y�/� +jWiꋻ� �&��u7G?�k�����,���'=oi��V��c�b�����&�q�ʥ�� .Z�[�pp���p���}) e�Ɛi��K�G�G|�Gkr[�`�2$C��Z��3YJ�_�׆���Ii�)X�5_�O����oh��6ϠO�؆��M{�[Ew��*fuUZ�+6��$�N|l���H�*'d��P�qse~��	3���U���f�d�7�/��{���WQ<��t�;uqG#} ;����z��c��皇f�p�LQ��������q);�D����\�ڑ�6�e6�YE�׷Nc�&�:�/��U;�۾!�� p��}d��A6�t'�͆w����t?��##�Q���&��3����%m؇�Y�禼���&��'�Ɵ��&4JL�>_���fd��퇣N��U����� ���j��F�]�H�V�5��m��xJ�����5\����:�����$���Pc�6�lP�l"���ez7S����̥|��/⬲�?���JN�ݞ���s�ݧ �K�S1�R�,��#���.�UV)��p5�#��`����v�YV�4^���a{%��)	u��� ���9&�֡z� L�'���yߏ;�����%ċ���N?2��[T*���� �@���e֠���o�P��rܜ��wP4��2�u{E�d@�+�&(�:�1�+p�#��]?��0�������OJ_M�Bɀb�āX2<�S$�`�+GShM$|�p���/� r'�;����%��� �	cvH�(iZ��C-�裛v�oW�|���,�}%�I��I�*��t��q���҄�h�u�4	T ��/�QI9�R�
�Jμ���(#��(gm}�\�YQ�&aH��I�5�`U�G�-_quc5w��*J���ET�K��
e�����B��s�y ٹvP���j�����)$���
o:}�#�vO�S�
�{`��|؈zp����� ^n&�R����mʻ4���r�nQ�.\H�>&�='�S�7Ң �����t�F�'�Ŏ#Ξ�=���S\ꟻk$���%Q3�+şԉ�m�������[����k�4�s�q�ƍ�0+�%��x�ayz|�n}�Y���KZ՟i�`%�U�E��~/q}���/����Ɔ����%�ͣC��_�~ �O�jP���y��Wg�� ����a��LsJl�IY(�i��	:{X�/�+�HA��(����l֐p�9Y��%�@Y�V �g橷��N�3�'!�*���x號��	z��hW���׫�|��O�"����"ۖ&��4���۶���!�R���~�q&�?6��J�&]g�:H��6�#\�ח�D��VR�<����8�h�Z��?qm��@C)V�xX@��
i	�W�%���%w+�j�QP�R�$GÄr� K����8P���H�g'h��,�� ~�Z�q���~7վ���Ԩ��-';g�t��z>!�0�6�yX�`�7�gT�5/a'h$$;��&~N5(�dC�x�`՛tH��ޕz5vT�czɣP��OGȵx�mE�\`d��q�H����p�o>6-wU����ka,'�g�a�'�������%LȊua���E#7PÛS���
�`������j(���28r���ƍ����mK5ǥB�G��!T3ı��b,V5?�D�l?�\b_��u�*

Bi$���h����,w�[�&�x�������߃��E��G���JL��r9=D��3�5L-���)�V�+x�EY�2�,L��y�F�C�e��!����$}������(��2��j�t*.%��W�lJ?�R_�/�K�+�>fC��Wi����ϵd	j�w��mӁ]�����}���"��ݭ�UP{�?��T�������$��fQfk�d��3��i�3�`8�\fAn�>M鍼���P��\��1o	�ڶ Q�f�úXc���yB63D�
�1XZ$���~?t��0Ff+v\<��\��ϋX��U��Ӻ�Vv�B���ʒ"$#/wZH�̌�����z���9��#y�PDr�����\�k��"-r���a��򧜎3�nh��7��B�B���H��H�u�){%R]�#���TjN☚U`9�댏�G
���Y!�r���?X5��`���%�t9bme�+�_-�ձ�o�4(ݟ���)�P�$)jͦs^�������^����]��h4&�3��I<�z���e6�e�I��flB���zM|SHa�3^2�Z��.-P��m��Y(���g� �����?����%����3o�}
W�5!ϖ�H1W�K98�������ɬ������� �3�x�b8�z������Вn�\H?��>��D�-�=+��d���@��ʁ4`NbM�`wR��y�x؀}i��@��E1M�j��y�$�
��Σc[��`ߨQ A8��X�3�S ڴ|9���1B��;3��wD�*^����w]��,ה<����2at��=��B�8t�:w�F��S�*�j�ݻhmk}��z�P
`��ָ���w�m��\���z$�𚢇Uc�t�E�'k?�_����)c��#�6�Ӌ
���q����*t�I���Mp��W=W�3�j�x^Ǝ��iA���*���\��*0�}�F՘͖�'7V�6�ɾ���7���B;$��g}s-��2&�	��f�^�)�em�q�����/���g�܀T�ec�e��w��314/PC�a��l�h�߫>J�n�ZgZ^[�;&U�{bN��w�LJ0�����Y7�2/N�Ֆ�	P}�I��̗�Yo�'j�qu��4vYw�R`$pdh�`��`+��<�q�X��&8ь��<3ꄤ�}F˽���/�B�h-�ޡ<�����Tk�{?��m_�!T��������k�0�h�=�I:۔g�t�&]�?��S�T��Qg�C`&�X"�����8} ���MZ!���5_pQ?��?Y{�[``{��̃���e�M1K,�v7������
{�<9]��jL��V��9�s���i��F��^�HYNP�wٔlfR3�^:u|O�|=���iB�r�=Jj=��O��i�t��9�-�_�3�w|���aP��JX;[���dAD�GZ��"Y��%P凇}�^�|ւc*��R�ۼ<+��*%�������F]���y��.6sZ�b=P�᪓$���@��	��b;'ʁ`����<̖G�T^���p��f�Dz� �J�(�6�@�=�0��+J.`����	�/�Nb&�ٸ<b��5�^p"?�#��0n����̩w3i�g���g��3EU��!�%c��j��UP+�x�+��c���q]�S8���8���w��+�㓭�s��d�7v�J�������h�L�,���i��Gv%����a��S��o�	�m�[%$c}:�z��+l�^�Щ2�^��8r�Ц��-h�BO��e6ǟ'd��cLz��4o��wH�[ؼ�!�Ty�k���IEQ��	<������(h'��X^Q���'M<ﰇ�r��""�(3�G5���[ϖ��H-q�
Z�(/�|�I�*0��۸`�8�g��C�5
��Q�[ׅ�-1�?�#p.�JmAܛ�}_��1���MP���E������i>��^9Z�i�7���]#&kz����B�����#�#�5[��_�x����;�_�򃒨즽�>%���&�ںP�����Z싈ȍ',Q(�	%+�5���Aw,B��ynp��!������ͪ��D4�!�`9O-)UyG��0k�k�W!�B
���Y��cur�=��L@_t.,��6k^d���h�_l�j��8��h��8RCdZ3�wa�rXvӠ��Q�x@�t�{�a�R���{�((������N_�����ᤴ ��k��l������7j��;��c'���h�z���˨�կ�&L������Fk7�"��6� �.S����h�N�vĳ�J;+�{	�K�I�p������P���P��hX�h&,�B\�k/e��T���F�����`����
2VT$�>(���(�_�F�~[\�m@3Y�1Y�u�]���v���B�G��\M	
J0���\r�̈́����r#9��z�Q]߲�宷?1V\��mg��I�`�/׳�!���LW�LQ8'��u�ϩ��:���*�8��(W��Lw���Ƃu(�h�*v�?�*5⚼������9����m��g_��p)*�����$6�p�&,kۗ��xl�I�#�w�Q�G�p�_��0U��wN�4�dwsz�G�*m�������ڗ"�V#�
%�oü��I����q��i��xQ���/²�|���>vF0�-�4��h?�za:� N؟�!��e)��ڝ[	��_Oس����A#�D!3%<:�o4^�����<n������h��E$��ĵ?�0����V _��k�
q��`.�R{�}�p�
4H�HEYE"7�ܖ���?!!i-m��zW�{V���Ϫ�ط�9o�"�i�ގ_������8]���J��<�C�Ke��i�4x�*&1k`�<!��oL��Sl�<�����͓p�񯍎z6k?2��gy	�{D��@=X��s�*��p�X��l��;���|�G��ytChQ�N 9���45? ��e%o��_��O�_mI9���\$3�)7,���n����ֺ���oG��g34\1�L����_��굥84X%��x�&�C�����B�#�-�f�8��1]��ͧX����펨�1�� e|
:IE�Qu�L��WX/�<=Ɉ�!�_���ױ���@�(�_%$���8�bni�M�>����6�b�k���!�	l�9���]#���.����#��_�<�U.��B~�3UP��pl=ӿ�%��e��ܤ���S���qՆQ����{�o�Й>�*Cem����/��<��H�o���F���#eC0���tv�u2���:�3�d(�l��������=3�T���}a�"�6����Y�6Ɋ���Y4����`�;�lP�:C�6
'◪T^��^�<��V�(���t�}.�k�lh�.y���n#lRh9�^���g��t����e��)L�9�@���<�e�e�Q���
>C����d����b���uJA� ƅϾh�`i昚m����z���!��c�I��78�`�n5����q9�X��Xꑖ�y ���c[��vVTB���ڮ2��)�`��j7MH��g����	7��2_*7���P�����*-���=��:=�tl�\mVU�������Iq,�:�}V�E����[J��j�Oj����%��%�g���w뒩���|D<��	�n�0
��d���Z�*iS ���`I%�-Gø��n�E-7����}�&h�`�]�kH����G�,c���ZT���b�>"�>4^ٮ���<�dk�T���\6��Ҙ)D��� +��K��A��3��}���b7]�>���w.}�6]g�\�b�@]'#�Y2 j��J��&?痕��1Ωp}���q]q���,֐��j���DFH�Dܒ�|@=������
���7o��pK�檎�*b���Q��f��I����of�6��m��x|!��ȩ�2-����1���ǽ���W���w�Q'�FU{�e]_!=jq���|�	 lެM�]�h��9�􄱕��8����:#+w��ݾ߾�!����ь���g�[9�vHTY�"!���S$+^\�@�8����5�}k[�rJ}�.J�t��������9��o�(���Lk��϶���Y"q��݈���>���<��Q�p�'���\|#�"f�����<=�Nܥ@��0:dkO߼Ӭ������+$��^
�.�lȤk!A�ːO�х��@�U�gq���>\������*s�W�#x���;���R�X6�xf��?����X&��V����e�H�P���ƅ�)N�uH�ާ���5��WF�#(No��R=Y����z�0N膲����_�_�zwG�mE,��"]��J�����H�����^���{� ��?+9�����Y���Y�Tٵ!�yC���+Nj~�,R�Wu��n\��L��;�)\���n~��04��"x1^�/ұ��i�Wy9�;�p����Zk:���"��V�zj$CT�"���/�3��qr��P�S,�P�~B%������JuP�r4r��A������d"�_������@I�z� MF��
���� �F(��:(Ǝ^����ɺ�f�37h{^�zK2|п�hS/�+Bl'^`�%#�B;�sMG�pZ/Ĥm�?���&S:x���]D�-����]����q���sd����34�k� �Bx�`^��m���Y�����YP��oӆ- h	F��\,vxAΨ���$�?����4�lջ/�\\:� �$嶑�}��\^�����O��!��~8E*vH��r�5��A���_!�>�փT8n8k����̷˳�1:(�/�(:��l��F�s�{��7�S�z4��5lr@S2�k[�t���%�e��a�&��v֨.� ���~�=�G5�Rh vD�Z���`JLVBBw�SWm>DVp&��"����ơ�=p!���T�Q��d�a��
c)��vR�����{6���F*G<����X��,��j��'&��k�`TӰ�Is�f�%����/܎7��&���3�D/��E�#�Jj�{��� �%���t�N�/:c֌�l�Krʇa��_�����	qS1_����0�'ڳ��L=��P�� �F3��(�c�N�����u~<�� ߿����}�L�D&q�">>El�v�H�0�^Q�gI����א��I �a�J��r����P����U���� ���۵j"�&��"��H݌La=mc�z���`�~k\R��6�4�W����`��#�:ب$uq�r��z�d�/��Kf�ۉڤh����֨�>�]��"��	=	VN7]�H���W��h"�)��C�lM�v��`�ؖ'���xA�9a��F���]�kVw}G�/��}�b�^i1���.x�T���4���l��Y���M*���
��*�����x��O!�bya6B��)��Q����x��PKzHw` �"�R�a?s�Tx��8��e���a�aս���֍* ���;�L� X��ػ��D�şi�W�υ8�m&�&6����r�}F��i��W֢S�^Ɓ/���~� �?~����X��>tnA�(����g!!��8�8��v���	q���o��&��j��X���2֦_�
�[�]@�q��@��ug�d	c���O�?@Z� hDJ��%����g�M��'�bF*��ʼi_���.{ ����9��tI7��.x�m��E_��ε��J h�h��>���/�pO�c�,�#u��,gZ�ri��M��Pr�m1&�����5���%8A�u$7�xp���Q�o��5Ha���}�������B	&g����e}z}��[m9A�纳S`%!Iw�'ס���n�VE͆�� �zVE��k� 1s����{��Lk��6������v���x �Xb�+�)����|H
��uVs�19ᶳ| �|�����MJXV��:��m	� ˍ��M V��4*@8��j]��Ғ�a���z���d����_�
�Ȉ�	?�P�`�Ո=�TVլ���/Ιp�E޿Ix�wj���7q`nf��&��ܴ1��-9�	~���>X�r���B
z�,�)�[u�X(�U���H��e�����Wc�tI�����-����;�Õ8N�R$�?65UB�K����yx�V���8�'��xy��кOJǆ9&Lg��r��yXd8U�S�Pl\�Ӧ���C
��_0�=x��IS���trlݱ����r�ꄫ}�x 'S�S6޸nh�P��P�}���/�&��_~�ӝf��;�>�PGx�K�:��$b��q�ETc���"�L@�ڇ޼�����	���JD��.����	�;���@�d�kt�ԧ��	��s"��7w��*�ڃ3iA(�n�7��C��B��K�ģC�:����"�|d��v60P�!�o�t�}�%�M	���?[����I���<��"�ףb���&���|$C�(R�rH���>r��މ�������(�ִ.���[���B˕������iX{nDU&�I��9�{���:�v��3���颈�t�Ж�'�;ew,���ڻ8���&�O.?\�
b�����n��ψ�_��o����h�.�������	}�<�ŃVj���H�E���=�)�a�e\}�"���<���*q]x���R-�@��$��e��2�˖�˻smٔ\GW�!O�����8A��7a��w�5��w&�j�Ʋ{4W�\��a�w��|�{o�j��K"9�ġKfm��!�3K72�q��wԉ��*q����L�� ��9M��+�$Դ�$:G����ø4P�wV�c���P"q��;��v�9�����`
Ѯ��OQ�ȿ�#���Ap��j��Q���I���T3;\_��Fȗ#��X�.�B]b��<�5Dje=!F��X4a
�7Dϴ�b��,�c�@�x���]�%<28��-�e�˛�g� v(�����sa���l�p-���� �SL ��F�U_⍎g�]�Y����dN�H���]
�ؽ�� �n��
���V;�$�LP�p�{��RW_x���I��iM$�5�ILz�by��O��bch��(�x���h�pCF=G�.0p��e_C�	j��@�"]i�W&_�Nj��n2a5#�6�)�w��Į��G�Q,*�
L{�Ё]T��jv�b�Y��^��+�hJ�1HL^���mBG�C�����E��V�`"B�[J����7����E��Exw{߶t��Cz��3�{�Β�RW�3� r���7���j�F*m���v
�7
b�A3?��#�h�W�K�4�����3h�@]}���E�<��M�iw*v� `^�J�ҋbZw[�b�n�p'y�(p�����lx���
j���ϊ?F�]F���46DX+o�A[)W�+�>O�Ba� ���{˝؊!���J�x��|լ��v�y�E��38<��n/�}���X�C	�]�p���*[�@a�xţ	�x�/�kK ��{����0]w�qd��Ȍ���=�q����y�)[��d(K).[��?"P;H�jq�5���N�����x"�tt�[ ��v�BA;����,��u�a�Ze�
�~���?�YI�j[r(s�ӪsF���L
T���iZ;�^��S�z�a�h�-W��-��6�N�l�HQ�RwH͐���ceN��!����"$����q�����gN�$�z��88Ģ�F��k�>NL��'���#S���
� 8&`t�E�� 5����.��; �;G��GZ)��W�]w�j(]w sw�	t0�)�K��4fr`�+ex�麈C�\�+��d$�<��"t���T���u������_�?B�P���>wq�,�M���/��V(O�YWƭ%�5E��=���)�2��<Q�P�"�	PGw�0-B�uBm�����V�T�<��9�ӕ4uFͥ#|�!0�.�x0]Ϧ���
,l����(Oi��Z� 㿧���a�]Wؠ�Q.6x��O���GG�+��l%]AMod�.1o;���F�Qv�/s"򄻓�wS/@����;��T����ݤO�u&��I��ǐ�'�o���3�S�\��'_��9v��RO�9�SjK�n1zϭ�%�@���B؊y���` ������6�0�}gz����T
�6Ս�G^�O��t�yk5���<y�MC�#F��L�c��.I�x}E��'����&s�C�Evޣ�Xwi���=� Mp�V�d�3'N()���s'�C���	����T{��Oq�*�ܨ�Y� ��� [��ـj,�]��/�H��]%^}�:�^�챉���-����_�"�O	������aQ��]1�s�&�U�u0�oy\�@�7Ǡ��P(o�^�Ⱥ��#AG�Zt]�PB��8��D1��W�-�.F���ԳSհK93\�-tk3���7/���Q�qQ�T��6��� �I��)��q��Y�����L"H��:���B��^q<�7a^�bK�X����r��61 v�����{{������Rܽ��E�b��\O*���0��ɏ��y*�`!Q��(^�݁�2
��ʗ���m��ı��K��RX�od-�	eu�z&�J'slV�Lܗ��X[�[���^�Fn�5cn��S:~�m{ʲ��b�η��ٵ��|�Ņ8U/�4ΐ�]����|�(�)�-ˑ��K7{x;�v���^T��Y/VX,���z����x&b|I5���Pϋ�v�7�����O���?�����J�x�
�y�����t�����t�fp���%>W>�e�x�J���k�`~��G�ӄ��̿�i��g ��#VMW���E�x]`��q��e�y��߽|X����Oê�{��aH�W�U%@':a�^}%�~�M��L���ތ�1&u����-��qѝ&�K�y��'���<�*��uxƂTI���gXο5��C��A���Sl�2�E���ǵK���ב�UnS2I�1�2�H7�TW�1؀�AF<9��Jhq�e�v�k7�>"�$+�	���
�kE ������suV���
�}16���gu��2~��k���9]�;� |� r��:�k��D�tO	�ğPC{�=�J���u+5�s!�B�k���3�
��6��r�Rȟ��K+��?L�2j:�o����k(����!
�&�
�4=�24�ى羱����|%�>�#����o���ǿX��a� p^��Yo̲�?t�9Q�_�`^����[~Y񎕼��A	gFq�����u���?�Z��r�����W�6[Fz�і��� ���k�E�Xtg��s��7���RJC����I�������,�-�Q�{�b���67\j��P)R�72�G�(��
9�JCM���(�yE�	���EC�-7ś�L��wGs����(k��V�>�#�О��9�	@�Ź�cP�Dn������o��N�A��(��[�0����M���tJ�D|,�w��߸A-�����v`\�6%���\�f�����Uiـ[�w��|v��P�fe�KM���^W�Wy�\KՇ�}�Ɠ��}'`T�$P�����OK�,N���"!g��.��� Q��Bo_�
���1�뮘y�&��w�t��N�l��k����}������@^q�f���T� 2lw�l��܅0M����r���~�/h���&�/�����yٰG�2�(3��3tU�Zɡ4�cփ
�xQ,����`S���az�ԥ��,N���\�Ք���/N��Y�� D
0hCm��6��p��֋�M���iVI����Ǎ��_e�֞�h�������d��B��bDVY�A����Q�H+Ց��˚ƅK+��r�s�]o>,�a�PG��<�q-���2Q��p�g�vl�SR��x����=��̮a�uy�C%~$�����H�	���2ulc�x��E�#L��0T�ɠ�W2���㲗/�ݓ�[3U�t�@-�t�� ˂>�S���1,#�տ�a��s���Ie�AoF�z_�t�1l���2)addbI
e�<����¬��(h���nZ�8	
ޅ~�v���~WG�b���^�f�w�pc���u֘Z<mD�I���bњ.���s�o��<$����m��() IW�05����al����x54�+WE�hp5>���Xp�y� 7�G@w8���e�WO�ׂ���v|Փe���1e���QT�`�4��.S`o}�Ըc�}I_�,N!���/W��|v ��Q�+�R�p���싲m>���$�c\ҙZm��e.X&��r���I�;/�
����D������q{�Xo�V�W1��-v)]B�����^Y}/z���.@VO���U`��m�F���"�bWt��.���Ogz�L�y��t����0��⪗��l\��:����0�PL ����~E��E�xޖꍷԸ��4]����Z���:cV�[������ѸY:3��*�i���3O9�I��+^���5���`����o.�w�A[g-�V���$@~�@�([\&��k��Hi��Z9`,Tp�g��a���uSZ�~SB/c,���1ݍ�M�}�Y�e���}�h���o�T�l�=l?���e�/^�%{H�y�r�� ��� �DM�h��D ��Aj��ʃ���%1�/�Ǻ�GȬ[h��:)��ֳ���Ic�*�d,��y���n�~�y�l�w�v�k�4��n�R�Hl�K��;���Y���`����'���9mj׋��jTQo��+�Yyeş/�ֿ^9]�X���cL��� �8�2{i<v�ñ��ymL����b�z�U���	�4�6Z��m�=R�,k~5�-��s ���[]��H� ɥ�����#΁���81	����a�khZ/%�7�M���:xb1�����	�.���!mh^ꯔaFY��96�Nd���n����09�)AX��T&q�e��O*��� Bv�f\�#WRۏss��V0ﾕ7���ժ�2-%��z�6\��O�)[�j,�4����|>�wL�A������_��F��26"
l��b�C��-(�?�3�Jj*����)�^����)DIZmY��"����!V�]���fsX�?���7����1㲴&��?��e��+ޘ�h,���:\����:: �6M��z۹S���K_�x���G��BL_S�������f���m��WKX�h 3��ʚG'O�0��u}xf�k����5��-���ڼ��Z��ؒ��!J�!��b�(G���o�������*2ݬ�qa�m�Q��]Ҏ�Z��=�ߗ����GL�����_���~	���ϓ�dI���W^�����\`V�4u`���C�]pʃPN��ǬE��3ĝ'�ւ�+E���Yׯ�?��t*��o�|f��Q���5G2h�D|@y��C}���M/�h���EE�<��°�х��q^��M�v� }�m�i\�^�?��Sr���Ab 1,F^4��g!�|�)����he�Uo�d)�C�4O���:�1X��U�r̡	�:�����N��L��}#���6X7�)��_0��|��}��5X����� @b6=t�=���nj����`���FW�b�J�L�[k��8'Kl[ok�������3�p9�M��������q-A�"��~�e��i�8���5�f�Jr	�srqk�o5x�h��'���J�e�D�]ϧY�fx�c�e�~��<����c�M�h2s�_g�K͈��A~aC�����<*�RQ�6���"�$Y�1C<t؛#y���f��wXL�(I��c�V�
�u�9mG�%�K
��#���h�u��E5���EN�{�qO�%��߆ijJ��ly=S6B��KAi�咕2&��#KA�az��� lV;>�u'��e; X3�4�e13��Hw�K%J��'/�m���#�T����-)_�$r�o�<Ϗ�v��hC^�ٍ��v�Έg $����F��Ia����2�8[��5{s^\��yq�Gt5v�Ƶ�@�"N�V�Us/�y��֨]I��NR��sFV3��/t�A�a�A3d/~��A��w�s��|�6�B񧋁{��Q�oHJUWj�%�/���"ZT���> �{ ���j궅&��s��*� �KK��5����Am�q�(�C�*9��U	�vD�o+�y>%ck#�69c� ��M�tฒ��tn�'�u6�͠�^��",?�r=Y�>i]��E�f �d��Rm�)](HZ���3 �Ld�o��w�yE��߽�PV{ozG>�>XZ�%�hP�z��8�s���G6�C8��d\�0�5��1
��V�Z���@x��{�]����b�2��i'/�������3���J�D'W	�R�[����XP�5	�Of�o�<3Q�a7�f��Ĩ)�@����	�i1��'�5��v�raZ3l��z>I�o��I��N�R�h������e!����{R��	��?��W�zv���g�DF;i��6�q�#�O@
@X�'5ݷ��aո� x�lƉ��>��=d����W|�9���S��6�3 �kgI1���������g�9����)v;z���K���΃t�Mٌ�PO��,���]] ��� T�������,��nc�ƇO��$�<Q�hx� S>gX��r��qZ�Ia�a�1�h!�����bu$7K
X��y����5����p]�ڎ�{f��Ѹs�k�@��Ƞ�@��0���G=�ߞ��[�k�	�ύ^i���W��x&[����|"���h��>2�ː{@�1��n)�8%�̃$?���c�*�6.���Ȳ1�E���q	)re��d�f��?��u�p��a�ou��ߚ��,9�R��8kM˵��"�4c[C�𜡧�#=�����Č)�Za�R�3��9�cE��r��G���!�#��<��i� ��dH�"��F+�<�uE�ρ��[�;�^X����U��(�A�@�6�%9a�ŋFu�j�0Em{�&���6�^h ��3;et��Q;�h� ��o���N(��MԴ]V�*���&������ҳ|'l��E`,Wx��wrg���Yy�kD�$�s�d@���]aRz����m�%����gU��<}K�����&��j��Q)-�l$��nA�"ZB�����m��U�=�"p��4�aT
*|k޽�VY�\.���� ���5�7�M����y��	C`�Ք�ғ�Ƀ����+�s3�X��r�3��4�o��b��ͻ@��/E餫�hx��np����A���������!��$��/���y$����y�ܦ<�#��k��g��c�Z�y<��wM��9b�6�c��ެtK5������z�4���?���K��=X��}���P)?��G����@�\���f�P8g!7s|�:�ͼ<S{��K_@X���Z��seC�A4	�9���J"�Q���HO�/j�Io��:Lr���H>
W��4�_V�!NS$��c97UK6��.�s�#e���#1�k�$dY�