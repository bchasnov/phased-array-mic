��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�k�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������H�W޵α���N-�`��6����ݾ�FF��eF4��_}<�ےA�[,�|{�?r+-��5K�z��!��[��S}Σ{$Gx^����c��Ʊ�U�I��}�*���="����s�(S�h��
a��o��~!)!W5u7��_V��KeU7+M�^O�m��tR?}���}��f��S�Zo8��	
���G.��1d�"�E�4`��=����K!��NkW��<<����#�e슘�T�"�#�ݍ��M�֏�!�=\9u��ڐ.=�#d�N:A���qSg�^��k�o��E�>"&�p�>��π6N�L���sUW�Gm�,B׻� ]�Ǵ�-�M�[т�G^ӏ��/�����>=�0�'҄,8��zN�Ji�y��,j��u���0,�Ȕ�	Z���aK�h�6f�9�IF�)��Z}ǡx�e� �&�}�w���QݡK�9<V���'�d�ց)�v��¥��x2g��9����6N�
1ܨt���[���UUR��p�s߮�5�d��&F����.�6��*���X~���;��TΔ^�D�V5�}d{�����H���H���G~n�ׅ��̐:��<@q��>:�+���ߥ���"r��V�����+�� �c^���I���y��ށ��#>��b�$�ZM��"B޷�BH������DL`=��AHf�|�� ��l��Ք3qxPA(ly aT���ə:�%+��� :����l�5�A�?�`�9���V"$��΃���5�sǿ�쇊r���^83�,�#�9�_:����������1S?pw��μ*@��r��M6(��6l�a����7�	�����@���I3"�% �Ѱ���(��
��w�oH�7P���|:��5��ݳ�UI���/�oƑ�x8�_���[�Bs4TR����4�-��>�,�L/�����9������*e����N�$@`t��`�؄¬ �E�&�|.��b��i�{�G��8��Bwj|�:6^<�S��p���ܻm8F�����Ƣ�C޻����C�1�=�vE_D7��؀S�b&�(!���~��I�:S\�31GЯQо�Q����=�� �Ⱥ�EN���hE���ܪCx���͔a��Q�=���ߒ��"����w����4���:�Uó�'��ِ
�� �����<L�X�Z�oƸRH����M���?�.W��I���m���Z�._F�����ɵ3��������ja���
�m����{O�����|p�D�Ә�I�+��-c��čA��`m�T��8��V�<`�� � ux��j�'w
�4�ˆ���'~���hE�ԍ�&�Ѷ��_�΢��Q��Gyy�����Nj����=q�FT�e�R���^�W���Y<;`_'�}���(��iY��B��Z'�:�'��L��i�\�жү2XT
u�Q�,9�p���q��ƭB+��U~�@�����0��	Y�Ez)=�=IrE�jc�<��~�