��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\����q�?��e�I8�b�Ǽ$��"����ׯ1�V0������ڹ4U�<�w:�V��5����B��}� ��(�GD⮢V�Uix�L�@��L&�X���V�k�Tz{s��O �Y^�\Q����G��UAk�t����Ҙ%Gv��|0�����6�@�gcI���an��J��$�gR��s��	,��Pz �τ2FFL����`j�*�9?V�]s������v�׌�8f��n����=���}w�'Ԋ��*	���#�56��2	d���c��W�[�b2-�V��/��
i=^г�Q~/6�׌*΂B�	q(]���A?�x�fn�_�t��~7	��A�����|��>�|��яe$�icy�˜�?�d��&w�!OW�v�@�t5���[JJh�\����I�k��٩x�	����mu L�M@�"9���i�WD��ɗ:�2ˤ�B�Fֈ#fm�|/�42�Z)���"��v��o�p/I���n��>�ΆbZԦU��R\c���+,I���ӓ��w�!���D��i/���UM`L��V��G�Znw85���G�� ��+�9�M��j⹿�$�����Z�:$d��c�ۙ۱!Mv���w1	�%82is<]~(�8�VDk���6O�Cv�!�
�Z��T߰�a�)ס���X�wf��1�Zbi˔FFN�K�Z��19P�mv<��S��a�M��Vp���b�V�=�Pz)�$D�4�i�����`�����ĿJ�ä�^hрF0h+Q���6�U����ܹЂ��#'�{��a�VB�IDw()���r�;
i�:?�����S�r�};�i�lqy�q�=��yW8��g(��=�ӂ���p�����'{���ğ��t��If��7w�kXn��Y2ow�S�yL!�6����'��	�g���K�4��uN�Z�۷��,�V#ep9�:�B؁��o����#F�7��X�C,��\�UD����q���^�Q�st� T��A������) ��!4��W��"�)��cג)�-3
��\�}��;�a�;�si�߹���P�W+��������BY|��~֒�GC:ɨn��]�\���_�'v:���
,^e��[V�*е���%]�ݐ�@eMpB*u��\a�{���Us���p�cw1�K��Mg��	<!i��i$����Y��5�:�<8�-dc�j^ٓ��-��4o蟢��ף�Y�	�eL���0�-Efsd�l3
���n�D�#�^�6��s���o
�l��T���ᖆ%���>V�h�X^��5~l�m�����
*�\��VM�r!��J<���K ��+t�*�ԖҎ��5ǌ�LgfLȼ����-`ii�$�k� T�kjg)zufDd�c�1�^�`	_�P]t �p|;v>IF��ɬ�fSh�$b�
W�4��>Z�����Gis ��n�
 � �C` LS:�����p"�>��Mt1(EѮ;]�B���gP��	C�0����E��S�o�?�m"���v��*{��lP�)�-�\��ښ���*T�lR:�A�j�q�E�]Άn���ȉ]��ĨqN�bI)�{��h�'1���?�B'��y?��� �%���Ybw��M�O�� �,RY�=Y��6��''��E�V(�c�u�I�K�-8���Oۆ���h���<PIéf������A�!"�-�U	�e��鸥
�y�s�S�^Iކ�QEf��>�Y`�~�:d�`�)=�BTi!�C�[�NfMT��8o�m�Ms_+�V��1���6�g����_C�J_���ʜpܛ�%s�ؗK^�)~���hǶ��m���Hz�3QMܐ6���` ��Y������m�`q)]<s��NE֛���"��PCz�ۀ�A�u�7ߗK��;T�K)�6:V��RIQ\�[Z]�ݯ��I���]ڃ��6�_�d��s3�A����^�>,��M94C/�s�G1����*k#cw�Q���h�&��)$P��m:���5�� '�e�kɨ.�4�s/��)���`Hi�8
1���bW�ٟ�+L�U�g��^�-���[)�qg�\�"�V��v�׀��~m�K��n����)5"xql.���iR�;��]!�-�LoT�\}�- ]J�)�MZ6[ j�+-H
��ZO
)hk�l��v��������v�j�(㥂U�X=�n��x�P��%@O���Xܷg�W��A�>�iHU�-`(b6ey�|��E��m	��r:��8�$�c)sc[�<�lQ�!�zлR���6���F1�q��Q�q'�!P/�J���d��ؾ��1�8FWX����W�0�!��&&rz�SJ�d��|��s�WE�Q����G;Izj3Of\d'B�տ���r�	��M�,������C[��i: 
z��!'���E;h}!���L�z�v8r�4Q�r��R�m{ �������(p=/�P��e���k��I�SU>���p&;iI�m�WAL��x#nc��'P��� ���� �'�1C�"��>�1�/_�I��s� @�&!��=!h2u�"��d�T��fp��|~��������}�Dz��r�dظ�<�,���v5��>r=k?�T�k��շ�*s{�%o�n��藇=��ʔHB:.0�����>�Ǭ���v��=�#(��C������R�Ⱦ| ��������b8%����D�0V�Z� �����y���^�_���B�\b�Il�KkN�>|���瑟�at���J~�
�X+�'�"\a�����"�BR���]�L˧U^����9�Î����V��>ۍ���pt�P��E�����z[?-E�-�}0��<�q;{�>�P���fA�j�m rX3�|߆���qV���N�_?+�E`op�B�Po��5�t&L�v�n�W8,�<w|9��_S�428k8�P�/�9:>ep�炤�DӤT+<�(Ō����&�<�"K�G��,yc�?�s�yԅ��1����m�Tq�@L��գ���g���^1�ZL���}23��D�1�/�.��Rь̒�]��Y�^�otw��QxF�{�n�:��+X@E�e?GZk�5�8(�H֛]�aL�
 8S�4U���&:�!��Tx:h�ٸ�yn;���s�˒g���T����h��~��S�.�]}=�1�5a�Q�C���g�̀�8S�����:�����K�-�|;�6�b��`�5���
���4������������0+����wN���}�E�bćs�_��^�t���?7��qwg<��^���`��/p�j���@�!�O%����l�6�@�bf2����AX������4i���\L*H��7Ӻ�K��-m˔��&V)xy�(��?�{N� �x������χ���ʢ�(�O����_]|*Q7e���
�{U�:퓓��QF7`��T�n��(�L�� ĸ�P��s�1�k�Ѡ�q�32ɤ�m�[���94�a�p�9���bK9B�������y6@C\EA�([��*ϣ��b�Z?I��G��'��q8XL�ح�B�-�A�3��W֢�;������S�ȣ���9A�[����g؊"�AS��)�314�څ� `e��lr��֓0x$!�H��.\�c	�h�/.�*}^�/�bl�Y�����J��gp��9���,-�٧0Lu�2�� �51QU��;�!:?R�8�ԣB�33}�U��K�B��V�D�ЀP_7�j�D����т��?��s�1�xKs�0�?�
Xc8SE��c1�uK��V	�βƆS~��ب׵�1\VF&]������G�W��4��X�d��P�U�H�>��鶋]����y���v]�i׏9.�M�G��Go��|��e��q��k��m/�E��Ɨ�8gǊ:k)���W�0���b\������f><�úQ��''��	@;Γq�n4y��ǬB���G	��ު����Oƃo�05�����/�K����{�@�x�ھ�J��7�	�i�m��(�
��K��e��9c5?�X�0o�h'�G,��$����	���]K ��cU��Ǵ]��B.�	tT�����I�Iw��?c�LQ�l���wΓ4�m?z�>����DqJ��i�!k���B�}$��j�� ��c����j��Sq!�S���)!��|ڕ��)7�s��.�v��R��bc�#[�ط���/r�$"NL�C��*tրH
u���O5n�p[Z��M{ʻ�����뛞V�-]���9W9p��:Q��w={�����e�ޗ����ŋj�v�ɭ��#@�C�_z1����e��Zۚ^�Z
�ࠋ�դdZ=�Xol�%S:�{fU^j�a{�g� ��1�(iz�"y��KY%���h���Q6{&ߠ`���N�(8$,�"�J�
�ҿ�d������(��	 snam�i_��A�g�M")��q����B�N����&� =EM+����_���� ���7N�ŵ�4��2풄B;�Lb�>��µ9)�(�=�����?ZX��]O`^:J�"����鶍�}H�>A�ڞ����DZS�p6g�r�l�{�6w�����Hjv�!����˲��mO�����\��/@�~9�s���p�l�v�ft�XdJ�n�� ��JI墻2���՗ì`5#=�9�E̔�N3����ز��b��Uźm	[�7�w��p@`С��j1�m�2{�F�^-�1�K����J��q=�<\��4�l}c�Ȃe$����A
l�AcR�w��_��U �"�_~�T�B�0E�H��!�i%������G/�1�P��Ռ��?5���d�.K�FC@��^}�/�o(&�A)��y��_����+�+E�<4�ܿ��[�?@qy��N��?>���H2��u�'��*��[xуT�r��h��!��U�(�mk�s�F{��d�ݶ*R@���d�� ݓ'5,�z�?hf{�������=���R!5� ^~sұ>2W��3���I�'�����k�IɃ¦�u�ʉ��Cg��c���K��Nť�����5�|-��o�ߡ��'�,5�����~-}M���b���;�KL�e�-��4������e�rM��#�|�
OC�ik��V��6�'�KEE�?�ʂ�$휎�Ȕ�!}?��t=��SKYP�i�;�����*�ьd~����pK��P螗�Oe�O��r�G�<�K`��zί2Q�|�R$�u�}�Xh DӁ�Cw��sJM��[��E�t&eV����>;p[�����go��E2p��B���R ��|ef~�:h�Ҋmh��+�%�,-�\���P�kpt��e���D~��2��ӝӐ쒢X������j�a�]*i�I��V͑�k�`%����p��A���e�2�-ċ�<���vt��\9�@)��i#5S�Z�5����`��4Q�	
O F�<��e9A��N���{ S��o�ӛ6��b�c#��A1�q�Kl��K�j�dxE5�&���SJ8i�(	cA�V�E6��Ve+[���Y�Wȇ���$X2�0��6�r�J��	]O���Cw4U��3Jk� ��#NAD�ԕ�_CU���j|��� HR��o���|�e��]�������� �o��O��3�� n1�=����w��Ld_	�S����	;����Z�e�te<�l�;�d^-`c���-�>���^�)ZV�os]��3�I���f"Bѯ��������f�/�$�r`��<���}����y���G�~��a�w(�B��Wó垭�7D��߮�J�&��(�&#��@�����D�⏉+�SQ-Q�x�,:�k�W��C�_��i!�C	Gf�uo�] h�RwU��x!8*,�E�$:�J�X�V;��}H~�Vg�9f��>�����hp�i��r'ov aE���{��X�iU:�uV���b6�^7���CV�q{CeRv~gj�͏�<���V�j7��P�!�+�0��BD�Q ��'<U0S���3Q���R�x�ؚ
�d�\,�\��Te�h@v�l�3V�DiG��E���BJ�}��9&O"F��^���K�0��0ສs�NH�x`�O�ٸ��Wc�\��!�{��s��+s����&ΓЊ���lN������G� l��n��O���I��a�{��gL�]���ꉥO1)0�b�Lɓ��I{�>=��D?���<��I���<h��\\+���=� UӴ.C�����X��]b[H(Z�u� .tU�dC���#�:�ZXz�*�3L�;�|<�	��e<E�UG K}T@_�#u�V�X���һ{������3�]�[
v9P>a��y۸��o��ZVM%e��S�f�D��<b��%.sR��c�O!Z^��O�V�� ������Թ��w��D��h�<5����W�Y��QX����C�`zI8vf�y�P�|O��;��n�00�r�w$���%i��+H_������Q% ��� ;(t�"�>$�g;��_Se�浤�%�,�ٗ.�^_��@mtŘ��@�Ċ}(O�g�D�|�dL0e�m��*�o(}:�Uoj��c���C�����`���BX�R�أ�>3,���O���+K��k�(,kOq��KW������Ԧϳ}���P��[���M�FV2y�*hZg�Wb0�E�z�x2�5��YW�"S�]�y��̒%��������ee`]yѩ���-~��+@��Ħk�)�b�%���f\K𑒔���<��Q��L�n~J�R ; :dۢEl����{���Ă�s���ѧq�5<ʍ�y�����8��qr�C���'�h�o�V�8���HZF�����/���H��-�H��z���=V�������fe�ME�}�52d
^|��I�¶�Օ��d��a�uDm��ig0;�B��|zSÔ��ܮ�����a��2�2<�:qbg��������H�$�]�n�ު��z�� ��$���W �6�lIRhc����x�Җ��WE^|o�$�)�=:6p��a��|`�4W�<ծ��>�
_v�}PυFEQc%��ͭ ��v����R;���6wrѠ¶�I����ͽzm8���@���g$��!X�A�4���)�Fp����/{IY8������ڏ"�ʶâ�(ʨK1YwJ��4����@�V]'�Dwɶ%tyɳr�1�����$�2���\Yd���)i!/��!�(I.S4�`�#��r�c�����ad����P�HN���~����N<�[���(�-�F�]�'<��[\�����%�����(��ϧ l����-�����E�N\ti���p����I�����.c#Ҡ�ه�ot�oj�ЅM��@(a�g�^E-6'�?���'��V�[j;^N��w�:��4F#���6{��bL#�~\���F5������l4'�)���ȉ��|j�\�rlJ�PF|pS�6�/C�/�=1��J́��C�6t�$�&�����7��ϕ�	��Ȭ�;o(p�~��|(k*Ч22pOn�`����U���;d󗯛�eZia��T����'�4��L�ZH:����L�����r��T�Uh�b8*�391���hzP��a�����c��T��Ew ���j/�8�O�f���w+�k�oT{ly_��Y��W�c��^����q��#�/�����2�{�D7�ڽ�1a��ͧ]�ſ��%����$V �_1mBS�X�oUɴ��541��n	of"�ۈ���7�f�����]T�:6ffe"P������U�p��1ͥL_��Cc��m��	ek�kW\�d�q3#�j̺�Ǐ
4�D�I�9yc���Z�f Qy/J�����zU�k8�0�B/m�à/b1U�6gX��6u������V��zͮ���?��̳�����d���}�$����Ȭ�DnI��l���Ec��I���v�j��lT�+�^�f�W�%�U����g�[���x����'�ϓ�,�R`�:+F�q&��� �z�e¾p���O	�����?��q,�t����E)%	·�6��1��[҄+�,�L�VY�P���u�B g�n�A��������	x9Q7Ϛ�9�7ӎ�M+_�Vȃʿ��F��4���,0y��
�Ǡ6���d������\�^�cr���Cd�M���PҲ���Oo�
�%:�����_�,>�h�0[hy�y����6�IYj)��_���xώѻ5y�'����4�y���
���G���%b�IE���P��S
!S�l��d"�v*>�0X.X���v�_�B��e�`��(G0��EB<�Aʠ���*mM��%��%���,U( �K;�&��3T��л���f~*|���5S_V�B\{Ѣ9	��h��^g��<�r	}��tQ��x�R�g �]�L�+l�����!��靵b��&�TD�W.Lf��3a�g��e�=�&�^�&��5��b5��v���_���?�,a�󞃎�������G���2�K�b��o�G�#Ќu��,ɱ�_ /��(�$����*Um	��GX`q���ِ�9���X��V4ǚbGy�u/v�9fZ�繎)�|�b�-�V2� /z���\�i@���[����1t����6��qf����M����u�*��V��Rv��IC���s��5��Dئ��{+F���F�E�z����X�)Iz��D��C}��E�Ӥ��ꙪqkmԻ�S�0���JcÆ(oԻQ��f�!��� O���Ha�Y�����8<.���9 ������eRV��"E3/�ZRD��m��1}N|���6����^%^���~��X��-��c,�Ȁ�5��Acߴ@o�����"I�y�hp�/LTq��Fz�� Aq�8��NUY�n�K�Og�5܋�P��v�g�s�B�L8ɱM差�{B��B�L�����S�P��z4H+�^�!�!��
�i �j�`%:��n���km|gŀ~ٷ.�0A��Y��X�R>��/��R��QѾl�]�o����B��猁-<���0\�d� ��;e^�����sA>������B�� �0��tX���nf�ֶ�e�k���ǜ� lV�$dw�ܷ���!���MkK��@B#��>��GQ���_�l���3�?0��~�9>,�6x'�[P�hI>ц�i���j1�)d$��,�b���xT�
��-��Y	6��-���}��\\�fL	#�xӑ�n��óu YJ�E�c�Ɓ6w��;ܞ�y��J�'��SɀN�F��H<U��;����O<��ԋY����xN��_�u�)֮h��P ����%n� �Q��'�/}� ��#k+U"��������%s
��������>o��4�<�_�Rf@��Ԁ��b�ߺ���	��8*�f����k[���_��j�a�\�q`Yn��=�r��)�S✁�Y_R~?�囹�q�(Bo����G��v�� �9��w,궮�k�B��<�|��\�l�(~�VU�e�A������	�Os��@�����6����{fc�Ӫ�$�X���:�}%Q\����š��2�p ڶN�A�-���ċ �Qu��xyL���~���zf^�,�7�����}8ӽ��5��
�Ұ���椿Z2,�����V�- �j�y�Gݗ�͑xk�5���~	�M��fiL\��wz�x����kT�&U�A�^S4q���'c��v�	n�e3�8i�\y�׎�L�����޶��"9>Ǽ��_\B��_����PʈsN���q]��&�A����ߤ�pF �f��>�l�#j�
2�1L=N.i�1b�O07ǖ�� ��k�B@ah��	�r`{N����Yr�&v#I�(��j�n�~D<��ܧf��;�.����r\��M���o�U&w�Cŏ��,�DZV�>[w���~�߆��z�jʌԸ/��\l�M�QF����q�ku��F�A�OY�񀌐9̫Ďu�q~�Ն�F�c���ѻ�=����"�ʡ���^�b�k��T)vu�v��
P�5�����V{��j�}�`��J[�q�~��X��;������,�UHn��s�{By?�ɿ2�ء�N���sԮ!Ь.�5�-(�F�"�p��V$)Su�ڔ�7�*6�[���rR�wF%E>\0�v�%S�#f���W)s���'hyXs���K'�L*:dNi��mo-� ���`iC�9a̮`��S�լE��/��!����h��y���=�:JF��:��7=5X�Y��m��;���	@:IOUf@���b߷=��4��H�Nl��%?a����M�S��+�yκ���7YVM�<�`z�]Zt�nU�))���|t�!{@�<��̀����%�f������r6J�^l�+*su�$s���g��F۔�Lh�+U�Vl�@�nI�-'��Y=r��U�+\�*jϙ4k�d,�]���։c}S2��WtV]2d���T*i��6���#6A�Ht�{{Bű�����h�:�[��Mb���I��������Q����o���_�����(F���l�U�
Њs�`~<|{lq"�ݎ�Z�3 A 2��E�"�鍌Y�g(nS����n�8��f���QJmzS9U8�W+��&<e<� ��vri8$�Φ�mԹl����a�p�B�7���t�����=>&�G���f
}q=	 �\�Z��z�B�9T���^��%�WC3����5��H*�9N鳾���J�q�8o���X��k�J��!�4+�g��:����0�++����x�~��Mc��
-p�	��b�\��U�Dh`��\�.cTH�x�S{�A��0>�g��18.�s}�.}�к���Z����-�2��U(�s�&�%�gT��-�f?ay��,r�͗�cF�cX��-M��ϗV�� M�)f�6�#@D�ɡ#A���!��,Kj_āyD^�0@������eA�*zcDX��!xܩΈ
��.�d�zqj��k]
3lj0]}���+�#\>
��V dr��:£Բ��AN�G�!Fq`�:;��*C���7�2+���1/!��5K��==���٦Ɏ�FFx xA!+�m?��e;1!��U�:}���l_,�M0O5�	|T��Z��[<�+�1[MI�@-N���q>k�U����	�T"1���gL�Y[m�`���݇0�B��s6�0"����Xa1����IOB6蹕���˫�qa� �A[��_0͖����x�W�&f�K�������y����i wٍ�.�g!�Ǣ�׽HX�٬Y�)�-�c	c�g6�3��@��V$&ٝ���3��⟾ف��G�G�����1wL 	U�6��],�Xu��.|���NN��Lu��\�^��������G�E�c@�/Il�{^��"�r�(h�P=\�}+�'nr�nN����S�]�L\6�{O� �n1��&��H.�+�	K�� �����"zMX�rEg���g�ĕ�gȤc��3�������7�#~�͟k�,��g��S�{O��fi�!�R�j]���4��&���2�!�J@5nl4�]&�2'�F��5=8ӫ0P�r�jRg�( �)�zC��hb��rۧ*'��s�!~�Ctl!w��8���P�!�@/џ�Wz8$Ԧ&2d�1 _e+��#8T�L���# o:�DR">!��.��Pf|��`�|���ޕ-7a|z��uU����A��1��=��f��/0l�o�D��eC������)"���))T=�G���U�Y�
?OJ�vDY�EȅW�"a�v��߀��S#��h6�8U3�������[=������"Q�tQ����|�Q��*S~�-��v�U��3�+�C�o����}P�f�K���
����p&y�L;����S����ŚEs��W��Í
�p��^�5�+�������-�+�T�b֢��;[ꄅ�>)"�h����� ���eܞ�W��V�||�'�0���7H`�j����^�t�;���\���-�[Ԣ7bfB�ʽ̬�CH���&��O�!�m�۶�	����[&&�Iٝ_c8 D2���(�4�M�\�D]hd(@��\D婶A�5����Ckņ�G8s])�/�L9pS����hA��7�z�Ԗ=��.;����AH���2B��I�O����rKaQ4}hehI��O����x���Uy�w����Yw�#&������R0�s�uT�K=�0a�el9D/�gq��Ahu���y���v�A~˧��1Q-�����!��J^���r�Rc�.Q�i�@����k?-�"��49�'�!8��|i�����G2f�ʋ�H��/2j#��)��L/^^�/���	 |���ZƖ������~���2��}��eV���1([?��\��"����%�&>�R�CEC8�A{����a�`�&�A%�F���F�U)�����;��&�<��ī�ox���2��V���k�U�����S�������y,I�W��+<��@�˱����3��]�K$��w�W��@�)f�eT���$�#�XJ�I���P�١ �����U��`r��@.;hq��4ߵQ��(p��/d�5�]/%˄�V�d \-�pٕT��P�奧d,��˘|����Rt{��~6f�<4x4f�Q��PL!Z����x�B�#t�����xmdV�Y��cG��ŸXR1�M?�AB��ZJ"��T+ׇe/��S`<��WIzpVT��9Z���LΊ6߫L���_t�3�����x~-�J��@*�cC/�b��2b���	3�M���2�6��aZZ������S�Oۘ,�e�<����Q�k���E�e��.=��=fz��ƅ$xw�9�7X��f�Ug��K���9�~)}��\�c��-J����$_����c�]�K���z���,o�}��;���h�f�k�}���H �.�j�J?��Su�1��ˇFM~�6����:Ydm�?K`e�=E'��y'�{<*����%@x�6#t��mg1�-�-�O�ulC��H�p�v�̩�!�9_���# le�Ry�MN�����^�FZi�A�W�Y���0�������X$�C��
�`R��J@�5�?B�"�;hbz��V�؆�[�n�НD�AH��4;x��T&i�X�6c%p�ZX�����څsI�v/��AK�����)& ���}��P�)�8W�u6�e�ww�@���ٳ?0��Ob��-����h�=�8},l1Ȳɿ�I� �c�w�Tx%��Y{�K������y'<?����=0�$\����ģ$ҭ�,�.aMS���!������Hj7?#�;�Z�el[�� o�{�_H���f���͟��5�SL�F�q�g���n����))��
�JK�+t�ɾ�)�8Li�Tp2�$M@]�LV�>�f��H�y��n�jY�?`���S��
ӭc��t���tjMc�`�3�`�nQ�z�x�\�o�>�WD�o�2���7z�^��O��:R�&���!5��׎��J7$��U�����E�_�������ľJ���p��k�6���5�͜x͐ A\���J��)+��h,��x0�h2�2�Ù��⭜_�F���	�7W��3?�־mk�E��F��M�v��.iX�:%��N�M�.�h����ׇ�(ڝ��$��F���K�iJx�-��{/v?؆� 'ҵ대w��n�������i�b�9��
I������&���|Ga�a�:�`Ң�}}흳%���
�%,d($ ��H�vM��%Q��n�4�?�.��oG'P�e�ؽ���'`z�@�m)��mW%��M��J]��I0�$$B���Sp��oS���K�9%�k,e
�@�[���c{ ��0v5L�ܞW���h�6��lh�Y�4��w:n�� G�(��]?�svm���=Ҟ�r�´;�J�+T�X��i��7# �[�X���-�,��O'�x>}E�����s���<��
�=�6�[�@��y�v`�����p:'❲���#(G_��W�Ьad|&���3=|���=�A��+E}���x��Ǣ�;�jy����]-n����7�#�l��_�*/�Lj�T��̏��=�l��0�P�-�1b�z�C��`4E3Ί�2��$��ǆI���X�(����Q���O��|.����G���|)���d�����ܗ�aVƕ�E+�$�J�T\���
��	�˸�
����WD�k�Ys�Jp�B��x���t�D`\;ґ�Ulc~��E�p�Q�)D��n��ōy���-�E�!�Gx8���FW�^�e"(�&�z��yv���M[���[�+��ƞ����4<�O��FVr��U���˹/;��bs���5��5�t<��J��p��Q2�XT���@ߌ7�'����ߑ���s���y��+�V�{�<E��QZ)ضw�"8�.#0V!T�w�lx�m�&E�E��!J3K��&��a.*�ۓҴB~���k{�
����/�E��+ ʖ�;�#N`�>~.��^ �
�Q70r��K^�;O� �B��b� %֥�%jv���*��QQ��R%�Ҷ�+�c�,7?4��У�9�.����8�w�k(�|;�N��k1Z���
D
Ď�=4-r¹��<Q�M���Vmc� r��ҥA'�Yo�4�<P�
�_d�D#�/P	��k�}d��jଚ�z	'�����Y�+ߚd9�׳THJ�*��4�����D�M��UA��\X_�Jv{������b����(f���n1��-�L��T3���+h$3�}W{]u��KA�Ѩ����*b�oD�YJ$I�[Ԙ�P��e�ۢ	c,�i��v8hW)��RɁ76�����6v�n��^�σ��<�@�5Oj�������0$Y��]�ʇ�H`Fn6t��A�F,dtix��*�������D=B��6y/�B�7޵���%e���~�{*.��dk�nt��#�:�]�p�oTym4���([!^r�������x��p7����O��t �s�F�
�C}_�䜔�	�3�xz��-c���l�krHp�/u �0���F	�,N�Ǧ2M�|�I��c���{<t��G�(3�n���\�3"	�[F�C���Iv�4�౒fR-4J)kL���/��YBwu�?�����MKC�����.�A+�2���rqK)��V]BE`4W}��#U��#��$6�% 
�ՐE&-֤PpE�pKJ6H�f<��Ўݲ��/#��-5m�|�3�i�&�(��#����A/j�h*�Y�8��|W������2�d%�ϝ�U0]�Mȱ40��¯$�,Ό8cb�;��ZS^�2������L�@������7j �T^?���\�Yz�	j���2��5+zPj�����	��<�E,]U ��v2�	��6~a\I���d��O �j��Wz&�~3�t/a�tǋ	���vt;�[��N��0�G�jp(���<�-��HB������T�����O�+7���R�XVY!�9��	�*g��&Хg�+�:aD�	?%�c�N*iM!w�*�vP�>���e
X:s3�'N�wN$U�1FߴF4�5�WY8x����$�)��׏��M�sZ�F��9Sc��l��OY:2)1�P]Z�`���Y7Lo^=/�)�FP�<��K!'Hج�s�*�bKE���G�)��<�.�W���jYK?8AF	V?��hZ	��|0�/x|D�B+h	T,���猹��}�K��aHV�=w��#f��k30-�ex?7�H_�0�-���2�O�!�;�Zo��7����Xh����Em��l�A����pVK�U���F�|\L>7�uP���x�*��"Ŏ9����W�_T����K֓���j��8�S��[�1ݟI�m4�7B�T���e����y���a�s%�r��v.�:S��|�-o�����Ew�$Aj֧r�CI�W�%����rѫ2�k¹<��J��w1�=��a�1�2p��<Ɲ�����<۝]���j�׮�6x�%�-��h��-�"7u�,��n��\�b��мYW��� �3��	�
��J�(X��?��'��CX��:Q�AEn�z�bD[	�9M�f5'�ߋ�1>��^-}�u+��JY����3?�T�����j���U�-7��P9`��.�u�ɾP�!�v_}R:7vv q���-��\������� u��|.�k��l����@�x�ɽ�QiC��0$����-��DѬ���*о�`p�!T��{���0�=�L�W��u�۔���z��>�La- v$��=�������^ɳ����T / o
��8��2�"��ʪ{�J��oA��y:�*�������6W�V�Q��dib�g���g�8)М;3�m6�7'Z	����🛘�pԴ����qho��<��S�&-?!4��=�V9� �PSⓥe�u{֙O�4����{P`"�]l��N�Y�^�7l�݊L%]�(��S�7��T�ṟ�5R�^S:���ȕ�T��P��FDa��鼃�+��|$~Rȱ?�$Y��+��U��g!�3���L�^�S��o��g�S`��[���n[�$c��� ��G����B<�{�#'>''V���T*��5��T~�|P���0��>ѓ��5b6B��Vj�����u:�*V�#���d�^��Q�`Z�>J���?!(�ފ�7gV��+�=;�9�)5�naL��č��{�������_~Z:��r&��i�h[H@�r��QI<�?��Fg��rb�|-&t��%���W_�.�谦����a�E�Dw����	�SV�p�X��,�������� ��^D3�4�2V�@�H$q�d,�1�i@`5���4
���&y���� X%-��z'`�-<<{ڀ{ 7l��^���Ϛh�H����D�Бv����Ed�/�$��� =�Jj��̰o^,�BC@hŶY7-	`�]V�A�����2�?�'.@�8ܒT��q����f�D��U��rߒ�5hhv���*�3�.(�uyK/�3x�H����AO ��d�+3L <!{K:{��{�������(c5�P�C:.�R�Z����F�Y����=l������ٗ�M4!S�1���iZP�N��>�F|����"�3������y�7"���,��^r��	ぇ�3�h����\X	z���&.@�k�
��"�m�� ��Y��c���>d\_??vwA�_[-ƦE�P���~���dc��m3�cO<��:S+���4^l5w��Ϟ�)ѷ-6U�T$J�|�B�:����Ŝ�.����������)p_'b�MR�\e�z���:dG����>Z����E)V|�Ϋ�%��Qb�J-8##hغ���R��X�m���`��h�;@p߈����Y�!
�K0�;_���K�J�z��p���������^SY�����0��Cێ�i����e^W��=ѥ�YCӾ����l�*���p��&�m8�ð�������H�����A|�6Č���&�C�S�����eh�{�y�<	�1~\茥O@ٱ��'�{8����qܑl��"	3E�Z" �=U]��Q�7�L��p�f٥��Alf(/R��uڰ���F_��+����<�Y���=͵F��GNQn�B�~�Q�8�1M�nAa�Go�R��$�j\�`_1�~���8�FB��p,k%��ʍ���ֱʔc3@(�q�x�͐�.�[��$ܽ����=5�>���b��x)}ϥt�u��H(QԒo�蓮��t8�O x_�#=E~�,�8���?#$�I*R����J4e������$����G��:��
��"4-�c~�E��A�>1�HPtØ�\	+��I؄���4*JW��e��4k-սq�@'��E���4��쵵N#�gy��k��V����E�7R{�8�Łx�
�S���]~�G�N�j,�vO>�hq4��/�S�W���ޜ�����^���}8�[>���L���4�/���b��M��R���ѕȅˏd����"�ם$XD�a��*qy��l�D��C���6�u�
)��#�y��p�5^I%Z�f{�����/~������Zt��Z��_����ڴ]e�����I���q�*��2ޔ�(���k���/�	s2�9���F_�&��O!�3䋬��������G��Ԝq6�B+�l�ǰ����K��X����4w3N�����Xʳ�E���:�����^���·�2���R�X`�Ա�� ���>=�G�D�XdK���)f'L��}�`�3� \���.�,�:ܙ��n޲���l2���kplc5������a�[��G{Ӟ&x�4&�!
A�.`�Y��*<���=m<��ܝE�:���"�m}��d���Z���:���;�\	����i���[`��"_պ͠$c�Eez���My�|�'�g;���M�{�&$���h�� q��V�b�z��M8��N~	�ݵ���/M�Ah���x�W@2�d�5�D��T�xA�����L�"��BV�����*WNQ��t���T��ҿ�dk�e���k��5ѿ$��g:�zퟭ@������l4p������n3#nH��	5oa,�7n>τs
9z�� Hꇵ�QaM��6�T�`���%|)�vHE�0�U�i����Y���k'�'侇�E�ˠ���p���JNP �)�$�@T�:��~d��!�5��+�.��,����L��@ͲH��{�8Y���m~��\ź�X�:����;�)�#����ް�=���֬���Z3��^�s�:67,��tn�Hg�ْ������]�#�Z���-�S���ٜ
	 CX�ʸ꯴��]�'�L� . iv�z�=�\���ީ�S����0�M��a44E�e���������>�������~)�x:��-�E��G�����UQ�L3҈�!c���Bj���l�h|S������GhS�?��-fzt�s���<�b?f<l�0�H~��-��5�3���<���V�)�O5jK�x���";�������4ϥ$K�:k(�+~Imn)���D��׼��v �(���F��A`����\�G�(,�)��q�����a��]{p"�R�}iKp���$�K!d�����Q����$F�?v��K���s{�� V4���H'���qM�#a�]�˘�
\b��<^|�yPxZ�wɛ��R��o��:��8��_��� �T"!V����`O�i�Փ�f�1����#�	5�⏳ȝ1D���ނ[�,2����y�����j�`�"��2&W@��>TN+C؆9���W���X�t��U�>�#��Iޭ�^���m?��)���{���=Y8cz�N��9�}2�w'ˠ��-dn�a�}.��ҿ�����J����� ��_���\�ӛ0����=-*w~��S�74�͎���c�
��\��q���� ���R��Ѷ `VM��������6�D�����\^�4�γa��}f�����~ݚp��5���l�z��%����ir��y^�3%c�\ߑ�����С�����PF��/KyYMZ��h�̘˰@�y�V��:����Ҭ=(��1Z��˙q(	/Y-���c��RF5ʌ�u?�F�^�o��pqޏ�y�����
������B:?5�r�j0y�F}6	fBJ�pη)�dE �S��'�IM�=Fd�5;2�:������tUЫ~�I��E��d�\�H�㣀?ET�L'_N�SڇI\�"����[S����/Ƌ$�3�'=t�K�,$�f�[��ů�a��L+�U��j;�l��-xg�"@
��\d��hyiRF��SQ�}*�e���7�y�"f����a�$�t�Y��+~��_K��(Vw':$'�����}�M�D���k�N�8�=�]0+v��,�}���7�f���0A���k�A����_��ISC��wG�a��D��i��l	�Z���g�/���g���"�g��a4�����d���t�;yy��ƙ��֪��b����L���r����^kZRQo�o��9kԩ�5�vw`U�;��g�kQ�;��������cȐ\<uj�}[��O5-W��;n�@��`���3 m0pǯ���?rcp�I$��)�ϻ�s�y�%�#��F<���
I�e���5Ԑ�l7�C���1Be�Z�q��[Xr�2Ʋ[ !)Úy�!��g�Cw]0���L)އw�{_;8:�L��z��_q1>��߃��q�)�z���#�`ʞG���s���%?��$�w@h���pZ�� �y��f���|Z�t#�&X�U�$9��7�>&����PM��>h����V���{Ճ$�a���4����J�"���fE�^��Ŋ�1�~O�}��� ٰ"��%�����@4m��/r�Z�T hW���^���gj*��yTqڻeR�)��/v"ˁ-�=���!͊J�١��F��`�Gt�c:y���k��ED�Ѡ�$ ��=#�rH^j��{|X��.�Gi�衕k.a��� �wBY놙����/!�^ ���#���^�xxs�lα��reh�oH�7_z��2��>�޶�ш^��\�Z�W?U��Q�Z�}O�ؑJw�)�U���(ť�w��,}��	
@���G��UӪ��k�0+����_dy�� �7���si���i��c�~�,�O����k0	"���E�tr�p�;��/5C�)P`1��r������H�5���I�����:�S˄=ra d����s�B���[�m��� �&�4�	#�o֕)DD�~�&ǭ�Y�Ku���x�#pR�+��O�ئ�Գ���-���Hp��kpY����U��[t�P�agh����u�{^���/x!��A�.��P���� UUx�x��ĻpK 
�r!��8_񹛸�Ⱥ9����Rj�ܳ|����f�!�P��j��������qi�zJ��C�-���|��>s�U8_�aC&�Ũ�f��!Z��L�H�ݺf�a#r����Q]|�Pv��`l�O!����ax�������o����}���
;W��ى��gy[Q�+����`u}�gҹm
{0�����++r�P���blG7�=�Ts*����nm���4�+'�І��@�� �z�����<���Ƒ�WM����� �<�(/9���j���䉖A��/11�1O~����X
uAv,� ���W07�ӻ6��a)Mc�Gn��j�R���,H�+W_�g���~l��<�
&�N�+ �1�A�-��b%|�.jd�R�!�~G_�~�l���V���2�^w2!��ދ��n��jժ)9�/�3�3Bf�%����*����tB���W��q��6���� �����9�3��ր��j8�/�ol~��.v�%�F�����`�?������O��'A.j�x;��$�m��6�k��~R&c�E6I�d�Y��qï, A�ҵ�ⓠ������)�0(��D*М�T�ެ����x�/�Iim"�!�;A�)UDd�fɔ'��h�Bi��Ü}`��d��Z���+o�6�ZR��4I8���?�,��;��坐`Z��l}��`��$쬉vxE�`�����w&v45�)��9������X�b�����S���(@�Q�W�'Cc����7K#�AL������J�H�I<ܗN�+5�s%.��\Z�����1��$�K��:'������F�)�	�[F����2���Ɇ�f�����GVő��M3ڬ��瘆���P����"�l�ׇ�K"�'��p���בN�s1ٛF��t�X�U4���+�Aw����/��+#�(����9�ܦ���5��	KgE��������a����ߥK���7�Y�-~��$?�p�n��f��65X1��h�s��Q����**	heM���p�E<�J�d�qϾ[P�6�ੴ��th��b0B�������zӐ�4I^�X�j(��xq�юP���L������Ɛ47��Ϸh����^^������<
p��;۵�<�d3J�	g��A����q��0#��^�F�RQr�w
Ұ�ҫ��X~���^ߵ����	.z�m���xě�'��fSl������Z� 
��+k��ԑ�ԉo��ZN��G2o��x�|&�d�&��*Щ�H1����j���x`?$�vQH9MZ�r]��,ۗw����iy�.�t�ع��¾�:��Ӎ�֨I�:\.U/� o��=� �}@��p�f��a�DS�ˠ��'aAZ`g羣o70e��8.ݻ��?]�^�W�R��t9PYC�=�P�����J��-Zp�䅃����]�|��P�i���$z�t�y2W���ڻ��X)����5�c�9��r�=�0#4����� �a�l#l|��AO�_��3���v��D��6���b�	����s<pE�Wi4*7�p��QɲԠiw(\.�`.L3�<'�߬��7@�߈'#u��G��!�iE㨯��i*6
"V�g?}�0�^Ƞ�IQ��1Z��1�"Z4cE���|��#4md�M����tEb��B홿�{��/��kw�:M��I�e��W���h�*�8����mk����%����-����0�z��h��5���.�����Ö�Thn��M^�%x���.^�i9�1j�H2a��D��}� ��ΝW�n0�<|��L܏ëH9�:��B*{�T���%�&q��>v��t���'t�%�w�����ؕ�l����x�W��w\ͧwo:��2z��j���\K�)��p��gH�7�¡���|ԪdU�,�f�V�����\����u�ש~���[��T�~�	""R36v�g�,��EuRg!����m�̑�[���X�o�<~�Ao���U:��Y����ﾫ��w���#������*���.�ﮀ!�״�tB�Ō���_�!�=��B��2�!t�7�DЩ��@�`�9�k�����7�� |O��A�Nj�TD�&�u)���mɭ�M��b�=�_����m@�'*��"����	Q�}��O;�����i��s)��p�E	�{���a�L���CX����ǉ?�C��UM������w�J#>�(�]QBe	#_�t.����qS7�]4E{�4��	���^dM����)�R��LUb�K7Fzږ^0 SM74:[��'���\C�Br�VK�@j�qO��n�C��Ј:�����i`��2'u�HU����j��)|T��~���]��a�e�����Q��I1N`X�z�����x�� PV�Gfe͂&�MW���� ���E����`fԞ�7Z�*i�@m޺6Ӈ�[������0���I�VI���1{ڳ*/V���.����E_h��e$���L�`�%�����D�_�~��ө��6�y�HT�W�X���5�B��;�Q���ʣ;�H_O9�T�5��.��1)�h;ۇZKpG>���ؿ~hpV�0��D��� �86�&��=4�1�"׏\��f�唨ю�};�E�6�ڴ>T]�+De[W��X����k�Y+0?{\���~),���ݷ'��^��l*�<^��I�[z^d����H�0w�F`�F��������F�A�Y�'wa%R�8V�i}��&AYΤ����HU�Uq�f���;y���_c�)���1�$���������;�r�fe�⚀�O���[h��J�7��;*��,�3R��D�$��(��4�:�����G�,&��z��C����%8nG��@��	�if�s�>��� �t��eNj�X��l跢��8�>?$��`෎�[ъ�K+�p�{��{�	'��LO�@�J�LH�K�	z�ti�����Η֚�:�ꆦې|T�=&�ί�@2V�$�&��|bso��?�Il֑7ax��&��4G�~�#?��@F����k&O�?�0�c˻}��%���ûv��d�鎗«��/b;%奭� Y�#��4/_Լ57�.[�]D�ǽ�M`�ah RV撚�n�pٝq��ѥ�Α�l���q�e�Z&�m/_�hV«�u�)�)x���ZT�B���z���ڍ�9b�2d�g�2�= �1�}
�
���RT�H)5���|:�7p(m���RoN�r&73<%��b�@��&�`R�g��)^��(c&�� &�|'�]�b�&[��6�Y��4o<
.i�@哔M,!�\�����$�x~�+�%i��[J��4-���g
�H��,��f¬t�0U�@y��ㄵh��Z��Rd�����@4Z���F����o��?���/������t/z�����+�$z��`�C3��Ph�J���R׿>�>�3x���#Fr,���Y�hh�z�|h>��ho|����E��Mc��<H���<*�����-#ce]��Ӎr9v��j<C�;F�p'dy.\i�<A�i~�ܫeGq��{Ǫ�]x9�+��R�,�w�H�DF֑�޻�\Fq4���B�b�Pٙ
ūujS ��Fɕ`����Tx��
��/L��rʈ�_�d6�?=����Xd�L�������>���u��!M_����Me���X~:�E��ʇ��l���(�Ko���!'{#�Q�@�d:Ժb�z�pR���8Z	[�:���O�`�Vw��h������� �d�U'�^���kL��t:�B�PΣc�O�J(\�ij}�St��U�l@Û���� ��BBц���aЦ�*���xM.�Q����Qh�P��<�Q4V8���]KD�y���ӜG�7��	\��^a�dƱ���T|�^��	���YS����؟b����F�f� �-��:��Pi��@ @A FV>;��������J<��Y{Nu�C���"�'�4��5��{��k���Db�8��)�&	�-.��m�+���~fE��n�Vz/&!EhцY�田���(b"���aa�
Se��A7?���?&���[�|�4�;�-c��8JA�?MH��RǨ���hg�m0�#q�T���M����ѐ)Qܱ�_�UR�[+�	J�lt#4�9�ц*CQ�����_�
O+���~0��A�,��[?�N6?��|Z%�:��F"������������Wh��5�.��w�UNx�?d(�	��`S� ��!W���+�2T9�z�G)\:L2n�[�r�K���N�!O�n��YC�f�l*��h$�T�u��&5s�%��`.��cvA���l��-3�Q�=���e��4��"�:���RC�`kO�l@��������aaO_�4@gǽv5���j������τ�N��k��K	@�/'g�z͜�&j�p���mD�8��^g��"�[F�}3Y�ʲ�������ѭ�K&B� �ќ��+1}&3�R�G�����Ni�Ŀ&�8��;p�\�l���%�'|������k\TYڂ7E�UD6����\l$���^��v��o��Mi�4��/����Z��7�,�x� @���-���-��`��b�F]��5`��c:<�����@���ͻx"�@Klh�F	��^���0|�. qⴄ��I!��C�0��4�U�B��,F�XC�߮�w���wH?����L��c�x���٢z�&j&MgC{�p%^��M���ʪZsiYNv3 |�@��Js;����&k��a��Q��ZL\nGʾ���^�%$��v�*.��w��H_�BgIK�wI��B�u^�9 w'a�l0�8�&� ���`r�7�9
A>��d�w�5�(���j����\�:+F���H��`�kl����ŏH��L�e���{9:�������W����Hɕ&+6��������������0�S�@V������&?u��7�5�8�o�ꒊB��/�#T�p����:�m�P$!��������ҭ�A ������ɀV�!�Na�|�$c__�f���9� w�W++�qm�( ��
�'v���ڝ8���c��O[$���l+/�I��.ޒw�����[��Y�,F����r�S�#R�����Ԏ4j :>��um�:��f�>~��ʎW{��G��7n,P�}j����������Jq�*;dۇ���Xz����ەR2�n�3+Vx4՞&���ڋFX���f�� L�³�U�u�c�C��w����_1���u0�Nʒ�Ȋ!�Pe�h�L��S�N���E�#��U-�]%+���'��7mw�6e�j>�ҏ��d��w�)N,�����ۑE�����Y?�V=�\�y���J�+� \t��35�,y��0D���Kp���+F��; N���Bhig�M�T��c?H,�i�兌'-��O�tY��YW��:�-hF�'M�=�d9\�c�������рZH{t>�3��h���7ks���O�&�%]t3��̃���_��M���nG�G��sG�V��9G7�J����Σ� b,ulà^]HǷ(�J�;��t��|N}���e�&$%BF�(��C�?Z%�e����0�׸��L��������m?�I�Z��b��`5��sq����r�KZ߱�*!`�M��ҙOmJ�XD�79�3]���;y_��t�����!���X[cxx+��J�P}���g6�y��=F���|�����9��V ��8I�u����g�1� �U�����z�I0}U݇tnO�V��+��#��f&2�O�����1��i4P��}i�ϝ�hE4,�:H+F�vX0Y�1Y1��n�@�Cu���F�<w��>(�+��O�n"��0n��$��n�U)
��ˍ��z�|��t0���QO*�{�ѥ
���'�T��
g��W����^��{mi�Ĳ��f�%�(psv�F�fIK^xz���^�ݲm�g��&aiQ��nܺL�WZC\>�5��װh�qt���3��O<���u�>2�<���?L�j�1Z�P�_�fqL_C������LRl��.3����*������8=��
B���eب^U\\��ü���f�$�s.2�=�81��h�q=d��]�k3ݤ?�8d�H�?UZ�[X7N����|�h�(-NZ��M� "X��q�&�ׅ�ʊ4�HS"6�_�E{��%�m�6H*GW��v���#Ⱥ-?���p��Y?f�f�E����sI�c�oY�aҴ61��� ^5_w�F�Rx:_G�"�1�]5��A�8{o$1�mz�{�raB�t��m�%��I�&khW�U2P����fae�����$�䂿_hi}�/ 7�	[f�8#|$�3�ՇP��X�(��y��^��hնk��}HO�m�����O��`��LR��7ұ#�R�w��VMμY;~�N#� f��٫�R��8�<��%?�׈+�%��H��a�5����U]��V�� �uO$��$��o�Z���K?�[T��Yj��>��UF�Q�@��yr�B��;%�r������c�]W:�=&:�Nsĸqd��Q�:��H|�b�K3�Ԑ�^�M�vY���N�2�j�ri�4�yr�N.̹��(����XS"��0��mě��m�`������ D��0!�ux{F�d�t ����{�%���U�nS�_�����h��G3�si�I�D��2�)k�jP\��A�mѧ����L"���ϙ���,����*R�M��
QP$���>�����3�S�O"����Oz����T��M>Zpc�ۄO���G��cJpwA�_P?�K�pwX����G&ƽ�*ߛ=|"�9��,��b�̯�o}��l]i?,�=:u����W-	�8	V
f{a�6y�z��C�E��hdHԢ��ڑ��� �(��6��p�<l�i��Na�o��E���i��nƟ���T���6¬�[?�F_C����W^�s�R�E��o�
G"N�	�qo����𫀙�Ft�sLn^ڻiN(�)�������
����o��AZ0%uUo݃W�.Z���U���3�����i^��F�&G*�Fsϙ��Jsu���:�,!B2�'��+�w����}ݮ��8!��p�0���j���w�"�ԿS�ǘP�n�/a5!����%�)��Б{��=ַS��&���	}�X�=BG��M���]}%�X8�5�n����n������2x mj��O�����np�P�@!"s;/��eI��	0����ѫy�w��ŭC>�������7Q��e���9Q8��i<�Z���1�|�0�7��]�L��a�_�-T��^�@��5ⵐ�s�a��,�A��K
�8��р_�D����d ʁ�XJ�鮶%'z��;�/��^;���|9�0��d����vٸ��M��I*��`���,u��_�P<��C�5���$�l�P|�@�D+�6�Q*B��s���ŉ��E�8��=ڧ%w0�k��0J� T78�����2�q�X��������j��Z��&��y���*ȵ8�
��kÂc/<��cA�����~�b�%'��� �D��3��h?�󁚣�o��Ƭvgp��W�H���-[�P#E��C�f�a��)�D#����_��֌kJ����y��9N����R�4Y�a#Z����0"��G��_�v��қD����Hwuf��hInȬ ��c��~?�(�Q��[Gņ���i9�c�J�P���=n֣�SrGQ3Y]����;��>V��?V�p�>�dZP*T�~���_�D�c��}.Zֻ ��DE|��B֬�֎�cY�vy}���� =�L�fT��>u�i�a�r�X �M��V��2/����4�sm6=�Bmo��Rl�w
9�b�9l���'��Y�H���6� �u=%�O�V��2��VZla4�}T��_x�)�&��7Wd%�s���$3�å|���`�h��sX��ĉ�a��r4�U���g��sҩ$먊w֯X���_�Z����T
�ÂԹ�z��Ym�P���u��u�#���82�M�;U��H��֑;I"�V�����S��S��҈�\;��ˏr#�-L�/����Fm�d����-"Os��B��/�Y�ګܥ$A��֫��[�m��k���'�wu�k�AZp�a��?KK_U�iW�H�L;3.W��@5��\'~��#]�3C�F�0��"�
\>x��Fc��A�ܑ����L����.�tRF�ˮ������2����Λ?�&m���4dq-���ܓ���u�RЗ��ջ(��6��&����-����32������L�w�|���m|�dm��"�RE[���0o�{�hz~��_@m
c&�F�9��K�U���
W�/;S��� �48�}��I�%}l��_��}�Ȋ	����H~6��t<:A�����(��=��=�"�){�Է!�=[����c�'hf��8�)~�C/MT�Ȼ�+�>�=��l�@0���a@o
f+���n���Z�
#P4����o��K������A�1�O��dj5X�t`�8�~mȵ��)л�a�)�#!�vs���g<y��߾5M4^@�$ �)�q�}&�W�h���?�.c>�\o�D=�@w����4N�i�ծ�W���,e'��! F_1�A�����)�Q�5�����A�k����G�j�m�B8,I]�3�Ңt8��|1	�!�0����:|�Nݣ]���(����Sx��l��&m�H3or��[N���A��\�h>�(R�z���1d6���E)z�O�ߙ	M(�l�x�I����!i`���g�����L�6�P���x[�u�]��i#x@�'��#�ljq+��Q�@��C���񵬂Bt�MB)aԦ�U	2�\K�9v�Ŧ�oű��w5{�̑�u:�Z�O�����Ñ�<��dq�U��n���r/Qq�EH?�gI��;^���p{�m���� 20���R�Js|C�2Ekd:�!�iA���М���6o�@��U���G���{/��iQ���@�
���@�]�'����ԙ���W�����]��k<��2� �r�>�`g�J�8�<��j&Q�R�:��nһ��<�;��?��l�ԥ��Z3�~<圏<�>�L���w릦Y��1��Q����b]
S��,��'_�:�а�Ѹ�ξC��%�Smm�@T^g�Fm9�r}�p|fS��Ԫ]�>Z��A��B�JO
%�O8�C����i�EJ��v�ʵr�x �݂�R���p�u F���S��؀˶����F)�sU�LT�9�!M{)��˱��ns���&��وL�a����O��v���Bi\�s8�[��q���-= r[�n����w����NC�9�4���J[���U��
�n� ��ߔ��%zKU8���V���-wM��\�/�S�	`/��D�n�|w��� h�I�d?�L��wڲ\�3Jߧ�ߝ}�\0e�&���ž7itזF�F������>�����<�_'iI�	��;���-q2�5��$wl�E#�=�
��z���>2�<��蒙�p^�d��u��Z�J$Ȧ`����O��� j`�%��'�Z�1�g��Ѕ�&�%�m���s���telQU1�w_�%���dD��'lk���rE�c{Ѥ�8���r)�J��ݩ�k��)C��xE�%�V���@^-���D��B��}�b��9�-0Z�t���i�:+Z��ګY�ӞŇ�L��}4뙯��qH����Cx[��v��nྮsIbHCvսN�=�PM�.���.|�����̂n�z��n���A�����P���Qm��s'XX�;_$����{,D<���#Ś�c�d?�Er���r(�(Y��+�Hrof���<L,Ȏn�{C[Z��'�n��?ꊑi�;�����ae�~`9U�g�}�*n���RU�ihfļX�\���燍�L��\����F4�N+_�١�a����	»~�'�E#�j��ې[�3\4�9p�`����d��s����_ǸB̮�H«%~�I�.�~��b	Vйu������oF�V�X�(����kk9cA��P���ۼ��@�c(
+t\%���؆���i����+}?����ʼ����,�3��H���*��%��Ɂ�����=vYX[:���@Y�UPc��#v�I�N4?b>^7$2r��#fѮ��O�U��N��@�^�g��� �6Ջ
��>�=a`������#�
��G&�fi�OkP��^���3��(�:U���}����f�v��(���Io�6����i%B�̌ҨW��]m[1U�RftEA�Y��Z�`o�G˂Ag�@[�I�nN�_yK0�q��ˁ������`ʡ�1�/$�s$��f{j΍��yϯ�6A������^�k�����|���MD��P\BEz\���ݤ�`R�&��5-DR;��ح��{��r�$Y2���*�v��(���dwX�Z�MD�w���|N��  ����F3$�T�m���'���4�q!f�%�vs��
�Ұ�qJj�q��Ot.l�9 ��X!<ޗ%~+��`��o��Q�m0��;�v�*��B���(N�S��<�)�K�B'U��ҥq�Y0���9��ny��v�[Ӌ���ފ��ǡz������{y�!��	��`�~Y���X!3����]$R �a}J㚬ʮ�xi�n�@�
U��;|>��<$���TCk��s@-�5�e�ʋ�x��<�X���O�g<���p�}��H��.���X!{���F��Pb��~<�����T���H.���^
Ň�&[:u��M`���I� 8�a����DqA>j�坙����*ڶ������c���t����;�����)q����� 9�L>���/_W���!Y0�в�ã��ã߲�_��l�n����Tp0	Z<�K[L)���"=�[q�Gz�A�$����B3���9e���N�t�<��'��6����*���߹���i�	�%�dY������Q����L5��L>7yw�vIBH�h9q0ۭ�Q̆�h�QM�nb!���[��]	y�]^
�fB3�'�k��q��V��P�ر*��q���r�7���e�lޢ�M�qM{�XwS�uh |țY��	+�/�{���SY=��������T�����r� s/.��<��5E.��ƛ3j�W$w��Ƽ79M3`4Gsʗ���W0�Z")2��_�q 2�b�."b�Bz��k����f!h}U�C��҇ݙ-����-n�����L*�/����?�/޲gyM�1\�.�����	�̖��C��m���Z:�}��RE�4�����"�2^%��Ѭ\����?~X�B���&�yK�4]�K�Q���M.��(�0�Fj Ѥ,~� Է��n8VP9�1��@������;��9˱6�s	z3.Iv����TQ/&�T�=��R~������K��A�Ъ��E���}�\/�b'q.H�p�§��bs�#�s��]7�'��0����lv7��1໡�3]2���sG�̬�Rvf2X����l{��m�dTI���Q����ˈ�?���u�H٤<�v0s����+�Ł�ި"!��\���-�����;���*����&��L5�ț���WǑ��[�~K'��y=0[�9$�B3�4V?+#0��BZ�^Y��
�8w,!��0����ZV;AfZ ��Oژ��=�)�ϭ����8�|7�\�� ��V�q�<��RSgA%/��ޣs�zx�����I���{Q89vLo�i����$D���'���3�}$�m��E떯^(�P�Vn�:�wwK�C��A`�0���e��Uh֪��=Gs�c�<�&�~���y��<�Zz+�r�ú�&�E�Q��M��*va�#��������0��f���y��Rm/�dX�z��Dr�-0���.��t�/�m� h��=�i�F\���̜���i�@�U�f��4���.;3I�t�ί�?<I���(�b��u:K܁W��R�3sgف�g�����>A�2Ts�(�\.�!�Z���JE-�����o�w:�ͦ��YW�S��N�w~'@e����We�A�q��zӲ�b��̽K�>�k3`͂��[]	�ނ�I3��_ z�Z�pf\>��-�rx��P��ԑmf ��i��墉W����R�Ȍ�:gQ���kWy2�k�p�9LY��s��K�E��d�F��7v$���p���Lu�;!Qij�'��A���Ys˩��R�l3<�\VM����<mv6��u���N?�k2E������^���"�[ؾa�r�F}���Y�N^�u��"ҼP\�"�G�%� qޅ����mf2��XH_[CP&#�/
J_E����,H��H�tȶ���w��w~�U"�0~k��Ic�\�
j��0vy|^>���4}�7�%��*�%���k�s
w+#d�$��HD��a�"�� 2_�������'���d�U7�,����m9r�5 �qE�FΔ�~��4[v�A��v��h�.�E[1����%r�#��`vG�Ǖj�Zq0�g�` �=�w%�'���[�E��e�򀳓�/(Юߐ#�2�����`Wΐ� �Щ���o�hK�;kI� k��n쑵�eJy���U��3�d���$�v7P�$�Ѣ��JB1�;ghĕ��]ԕ���'�^E>GTs��ߟDc��
[9�/vw��s�	�M�6#����^Pe�-�>�+i�b�P����۽�>!�O�,�[1�e�gR��{��Q&7��5SEH�nΣf���	��s�O8J��ˇ��X������	)��^%�dX3����7�A;&�6	���e��kL�� k�2��j���[�Fd��)�6aG>�'o63!�1�7���?�#�AD4�c�O�����Ƭ���V���ɲ�$y�Q��Y�)�O��h��G�}=X�PG%+3�����>�G�������-w��ȓ��J�2<��Q|F�mwf��٪k�+y����G�i�o3��,��Y>�"�B��-Fe��Н{��[,2h7֚n�9��Ư�z)T�Z�sM�Yc��Âֻ�O>�ך[�z�ۼ�ͣ��6e<�p��P�Eb���)���<K����b�SMP\y�R�w@���Zx8C���l��6���J���#��5�a��^��8��!���H�w�~�/�Q������m��w�֏	�� �տD�p�j6%���Lu���ҵ,�i�rc`�8��cb끃�F�D��oy3h�Pv�������8����|�<0Y.�H%ܣr
���w�%xJ���d��S3�P_ �D1�nzRx�������܎Q�bV���	7��F-R�gI�.�Ȧ��[��HKBΣ��B������f�j����r_�&ʝ)�U�V� �c��[��[2�9�A�3��0\!�t�3As�5��D�t�ogDF��PK[��0ah�|5_��rX��/��衔���t8�
j��Ś�XR�\/���I
~7�6��E5ī�.0���|��D��H�T��k���MD�S�R����r��9��	�v�ѽ��a3��򫞗�[��?����T0K�W���RV3g����[��V���3����PU���a.��u,�nE�v���\Oi�k�������	�I����N 1"�ξ��NA�cĻ;9-wB��3�x'��7��.辻︺|�����|�u2b0��l>=�(�'Y�A>���P�.�;�]�}��	N�����p��&o�`�߮}
\����/ ��J���e�b�����������*]t��WW=5r�5���F�Sޒ�1���������e�`ɃV�:�$E�/h�t4Ok�6����o�@5����~��V�d��34��ө�sQZLڐ������x�P�&��[����� �J��X��N���j���T��5�hM??��kx�+1=JF��9��bݖU�7��y#��X >�L���>KP��t�Bc���� �U��K�!q��H��˺l!��!.��da"���i**!��W�G��R�X̯�@���Qĭ����y;�s=%vw"������i��X�v�(&6O-zLF������tBH[��E��{Р��l1�0�ʜ/���b�Sct�|t7s=Y���^.�J��ͲB�����%��pY��l3U�B��M�fZ����W�H(+4�:��Ź�Fme�>X m�Y���~�|:����e��8L(P���1\ܶ��T"��A�\��ȕ�M�����Ą|.ͽq��ɒ����]��\�]���x���4\7�T�l=��"����'�qN���Q������;�w\W�\
�����"�/+q��$ ����A������*�E�ɥ	&pqc�B>>�,#��av�c��m\��M�xw�R9�C"�ƨ3�v]�����8pE=��Y�Dy���OO <��W�8���UB"��F�d8������8U%��|1�I�l��afnD��s��x�7ޟ�c�h;���u��VN�~�x�6���͊���d�U�,61y��CX �+{�@>e���{\.mt(�v	��*! �hL�k�.��M��_��&,,����Kx��~�"��	��JB}k��Ż<�Ja7����=���S
��| �H)ރ7*��	Y�F͑��q��,��캱5�iN�(f�:��@*��L�=�<�@�h��>;]l��x5�~�}�ϣ�v�]h�[<�n˳��*�~:w�L����|�|�n��Z�������E��8*��}�L�sOX�������4�w����z��&��=�Z�t�u��T�ܒ	ۥ����L�4�n�GC�U߁�7��$��J��P�5���()sW���gI>g����{�d�B&=9S�w������/�AHV�$����U�.u�(�$��Pk�j�#�>� �":�?]p�3?6Xܲ���Rt��_r�h1�Z�m��Q���R�W-��D��>X�N�y�Z�����u�VeQdɟLO:��S.�wn!}��໎����f5˝p�ܫ��]�C�c[�͜�,�@[rw̟��	�
�,6�:.L�mx�:�(,�[F�3R�_�����x��&Q�^[g�P: �V՗}�D2�k7�U0����,��N��f1AꖅB���h�:eO��T�H�1�k�+�]�u�a�&"cN͗<�����y�q^����Ɇ��L��Tv�'�З�U�h[/TjO�6�n�5Wۗ�������]�]��P���^��0��;�qm�,�rS<]�p?�n�*0W�Y8c� �<�H!?�mH�h}B>�}G����,�F!�W�����cN}@�����6(΢`�b����O�AʤSc^>�5�Zsw��g��C��������l�B�?�*Htg:�7��. ��da�$����m�tƥ˶%Sٿ��^�b!���g[��@Sl�KS����)F�껖�9�?�V�DL+N�)��T`����z�V�����^W�\��o�OS��9t����#��B�~�|4,�x�Z;�+7@�Ѱ\�z_�(ʳ��%�o�/	c�vI��b��@�F�J)��TuaWf���\�ν�T�Sv�S}p��#"�{�a�3��M�`���p��k)j%7:�3������I��]�Q�@(+�Q3;�}����Uc�fpOk��j����h;���6#���/(^OH%����{te3�C}H �����ڻ����k*M#���T���9M^�xi�N�7,�M�/�*�-?�?�)�ѢA��W�����C��$�����	�jYa�K␖z0�A�s��0?&.�e��]�ǽ����1��[:����O�Q��9掣�œ�1�L��a������7�y�M��r�PN�5�1ג�t���·� ���g����źw�m��#s2��V������/�������}�r0L
��p�
�3�����$W5��J��m��2���R����񙊡�UV���nﶺ��G
\я��7U��x���Ή	K�Z�dS%���1>B��E�4��m�P6{�"�l�h��R��b��qp�]h��vI3P�!�<dg���3wBW�)� n�K�Djl;�����C��X��h� �0%�p#U�?�W�%��A�p��"㗟k�O�i���>�ϙ2ς�u�ʥO��u�+L�gvF�R��/�o�Q�nP�W�8�w2
�U�ә�l|��v���D.��1R`��܄)���O��y6�EoB)�܆ٞTO|PwR6�T_I�����d��E]$����:��;�Oׯ�q�������t��կ}���a�f�juU�<�~��r$[����/O<�w��Dggʁ�7�>So^>��7s��� ��abJ��Px��pl(� ;��+�d�Kɇh��~}�vĤ;�- '�	�gJQ	������
��C���"zv\�y�D�SIy�c-(?�e�N<Cq��r�l�(%ubi��?��d֡�p�p�|�|m� )Qsi�������f1�0�O=���^ǈ�m{�ySm~PY�i{koqk����<��^P�%����/·��_O<������Qk��O(�+Vj���V C�POaN�/�[CWu�X}X���ײ�h��^�f���V��'��lE��yI�}w���d�*���*���J5ly�M`�1�^�%�I`�� ݘp��2P����q�M%
P|�y9k��^�c�� ��f�M�b[��]�u�[f�����N��>��2�&��J;64���2Qw`%�k�������l�nZ�����S�	�F�!$�5��b�¿v8�i�:�BO}�&�`|�):�Q<o����f�;¼���t��CR,֌ס���:TϺ�m|e��`��4^Kc�����A�$�FM��a��#/�9�$��}��b~�q�E���s#{����d�]Z+���X4�Z����vEu8~8�-)�� Hct��Υ�8���p�b-=R�7r�Z�?�M{n��9ŒC.P�}W��~D|S�|�H�yO��*w�'	 ��{�m�?�R��(5���H�)�S�(%Rk���qs�?���ܤ��^���'��]����58ޭ]�k�Z)O��%��2���W��q��o3!����2:�u��(ه�)���l����C�o��<��S�$���2�Hj���_w�<��Pܻu��
��:��X6�Se1߫y�ঊ��+Z�RF��)?���_�kפyF`U�M'�v�N�!#r����Q��
1,����6�pMY@V�4��k�R�y��K5�~#�u"aᒓ���.َD{W�Ч��vPU%��#�;Ԗ��~�ka�I�uM5�E��ͮ��+�����;0��I?���&W\�o��'bG�P��Y�@�c��y���ᄅ|y�`:�T!J��+O`�̙���4�~�C4��ė���fg�:�������$vЋ��{���I7H�8�E������l�G4X�Cx�����Ңk4XS��O]�9mì�<1���@��k�cnb���ֲ��s|���h��N���5�NZ�	��"�CG�u�S�k���U�?�Fc6�������/c0�C!Yģ�R�p�ao��Q�*�k�eDj��f.]���H��K��J�^���\v��»5>��c�F����4��Y���pŝ�|�'M�WG�3��{t ��-�h.`zV��9�s�;W2%�_x�r3�A!_�vɗ��$���7����?u,n:�w������Gwh#��.�S����oX��N 3?��*�HޢH�|�2��'�A����J;���I�W�s*�b6��Olh�Rԉ��W��E�Ey޿P���R؄�PB��Ȥ���D��cJ�3�e
��)�e�=������fu����L������'�In���u�Zt�(v�zV�L��� �\5~��na����x1�b\�;m��[N]�'U�9�B��j }m�g��j�Cu@�NkcaP �}��Y(��o�b�����Vi�YD��/���*���Y�1��،v�ۯV=��6z�q����|���j��kb��dZʗ��	ߓ��*vL7G��5����X!�[�J�Q�"�5�}ķHE_%�S��$��t����B�a�#��i*"n���L�0��@���7��O6��B��G�v��.�
=SQt���q}�Z�a����:�s�Ó)���t�ݵ����� �f�ܵ��ܳ��L�����m��qqD��Ky��`�n�����,M߹��&�"����Ms$G��|n��z�gHA��\$�=?����j��mgI�i�$#� o���|U{�$���`.�'(2[�G-�Bl�1`��f�A�5X.n��[n���7�$������X�����_����hpS9!��k�(�/�;�5Oq	F����?�[̐D� ����mx,\WUa�o"��J����7_r��2x�4!SMv/�D=�����HJ1��D�)�~>L�D������=���>n!��T�E�\N-�a���v�'Bh�$1��[˷�Z��#�]2L��f_޵�O��b�U����ǥ�ܸ�ߧ��5�H���Uj�u&�����dAW9B��%Y���I�������
�O/|��d,)��f*$�lp�Tᕭ2��N�.z}hw�0�O�B��p����#jzb��h��FD!iO�s(�{}�����G�qV�m�J�V��r|0H��/�T�soZysd�	qj�5����=�0��H ���4���/��[lݛ�ɒ~�*�o5����ݫ����ﷰ�t_/�e1�x>��Ο�3�{ap5��Bn�,��g�RϧA�d�kHS���L��vf�j$f�r�#���y;2W��\�%���O{��v�=���s}e��]x���<��!U���b��zzК/��0i�/^�G(IB�GZ����J��u�H;!��ѽ�<�iO�/��c�;-���KN�b��vm��ޞ͈�}�ؗZ�֝!��Eѷ�����f� �p�aGEO�ǀ��+�q	�Ź#bW�)"g�`�~8iF����pn�v�΀���)/�X�e[<�1�f����Τr�a����5�Zh	[2a����b	�(���l��ԫ�ĠK/y�q���E��Ɵ�����8�Ct��}��-h����Y��ޭ���v(_���F�aƂ����	8ur�Ƭ�cT�������\��Joȟ���\ڰA���?.Ѱ�5wT'��	�yg� �o;cn2v�M���YEݤ��>orKH�;1�}��y�0��t�y��(���#埐wf&Х�=�K�f;�-6�ZiH�P�O�@�c�k͒	ֿ������R�0-{��M¬]*׼�B����oUh��s�a����s6�x�h��[�ܜ��'&�m�m�J>�{���b��!�;�(��r�`/��II���*ԉ�z�5�+��4�R6e�f:xi\/@ȏ�ylc 3Y/@���}��*�\�>	��8(��0�/}�bVL�K8��U)�2V�9uC�e QDg��6N���7?���J�X�����R]��>�L�E�R� ҿ��h�?dtʷ�Ŋ��5*�B��>j��)C����|�h��@�O�&�"�Y4%�$)}�Ou�U����e���}`�2FPEu��#&[;��嫹��X5&+O��Ƨ3�GJ���O���W��'8'k]�&����E�$���P��r�Ym�s[�xWܓ�_��&
�f|+ٟ�t�;J_��YUeֆz��<lB �0�0�XR�ؙ%̓���+{�u��g4�A��1r�QZ����;�E�8՝NhQ�b��/@��G�obǸ[2᝞z�e$� ~8�핊VăK�Ow����8������T�����Tzn�be�
�NI{
�ބ.�]h9�]PZ8U�����-�d=��_l����E4�TX���_�p�:l3�y���6�b9':����c�~�ۅ74�������/"]�R&�q4o�XRi�}-=��i��
&ؘ��b��ɒ��J���u�yn�Kה'i��ԶC=��<ʃ�8kɖ'�|��X^�H{�(E%�L��r8�.y(��i}A>P����?�E&�==���d�+�.����T�
d�^��>D|M�+�b��R���x�ga<�?��?�7�o��R�Xˣ1�O��%~��*�S�Dz0P8&U>/%c댑`/%6FFdPVZ(��vdgZ���m�'���=��v�A���ܱ�����&aD�f$W�֔�^���Hy�G�2���N�&�e��V����jĚݤ�'�����������D�ݨk/�
��_5ud���'6����a�4vb13�2g�R<�&[��Xڪv�%��"Y�ۨ��f݌ЗڄF��&�Qq���t�!�t�R�"��B��1oa����k�����N��K<FR?�n�7�V��Q�JJ���<o��^���i��#D:"�D%(�Og�)���a�@��ϟ��>
?Z��\m+���$j;uZs��8�+U�&���u�1�3�oڜKՃ{kO�\�jO:���L>(���c�-�w'�FG5^{Vh�Բ'���pC�dM	�0�W�(Mt7�>2�R{���0�B��A�׷p�8�t�<�vF9w}콏22�bG����^��0$&�}�Nqr2��}�T�Y��r�2�/lI��X�=/��v�|���&�"��^OD�[��[1OB1�� ���g���}	��W9dm}Ȑ��(�w��\"C���w�ϩ�t�]�	`s/�?��*/���� ���ԂEn�Q+�D���A���&�Խ��|�?V簃�{� =ȶ��D��ZQa�?C��̟���_��Ng�V�:�i�,�C�^-�<-�x*h����i@�����?s���<c�
��ʢ�y���YJu��Ů���;dNˑ*��=[9-�05дH�r��Y��S��ʔ���{F^�sp����
�����y�E5:��yOT�c�YJc�.]���B��o��(�SOT���d�q��ֆ�O�8t9Q���ul5y���R&�c�Z�-?X�r�3�#Tީ�.�����!N�W>��r���w!��q�]=�Y�V��t�
׉�<���&��wE���s� ��"r�s�'x
�+)�	Š��Z�����^l�ey�d^��|�\��}���C�X����:5s��/|�޷�C�Q�N9e�_�J�9��a���pe�8a�b����>z5tq���(����	�{��]��z�;69*	1��\�IZ}�?$9�:	����DT��%����>bV�p����i�(���`���I�7"�씥ˉ
�4�kc�yB6�P���L��l��*H�X
G���f�v�m2
�ro^sEg�N46�p�\��%�=�X�Q��hA /�� 07�4}D��ʗ�l$�Ywm��%�b
�����!�3�P��+���<f��x׊�gFr}�X��V�%U>F��N�H�f��6��	#�l>�������Q3�f>[�):/�d3��g�5	��)�4�#����eޓJ�M��D
6��%���RS2�{�v����M �X˙[$m6������yNٟ bh�be�NGyl7��5k/G%�7�θHN�t4n$N�ɭ/4��[$)Ԡ��v�`t��1b�!Ϭ���,���X�a�L���K�8h�l�dh�Vu�謾�w���a�-�]��9�u�[�l\�l�ܷ���)2P�
W�ǰ�o���VbjP��C3���:E��\y��ܰ?��/�	z�]��T��Xo�K�$�7�Y�HrIo�����e�V��|t؛4��q�( �?_����d:�3���M���|-�C�w�_!lP�6�y�QKd�SVn��]�D1��.��_�)'dY�9>��x&B�����+`󟕿��9t:s��js� `I�o�֘�D�q?Xq�Q�����m����wx�yD�� ��H_R����'��LN�M��X��Z��7�<
gW��8�Z�u�Z >9�hȘۦ��D9��P�0�p9����*��D��
l�WR8�I�[�k)R�`p�1��]N��Y5{v�.�w�k���m���Mh��7�&��&y�Ш�E>i��䶝t�3��[,2%�@��9�m���e2����i�A�!���1�hL�υ"�a���������F��� �@긚9�~�|��?���L�5ގMqrߔ�����g.)�%�߅�߃Guq��j�7 Ս����2?�#X�㢈�	�N'}\9;(I��4�>C�Dэ{�N�n9`��_ܝ�j�x�	�m�P�΂��9�+Ղ�t���$���Q1�I�ZtGD�l�s!����79h��x�\����r���C�{m�^8?��9�q��A���d��Y_tc57
X@ߎ�T�S���v�ެ�T\dFT��۟�Ԭ���e��Z��	�x�.����T�j3+���y.���}�X�ѱ��a��3�#�=�4����j�y?UD1���tG[	�{�yh������W�c���>����'�3n	����#�Z"�ٮ����xC���x&�4���(A���2�$<`�#+5W
���5.O�P��ڔc��GBA�Cv��Z�d����EqSp��h��ˏv��n���^��n�/K湈e/�&J��V��J�q�)�Z�i��r�0���uo"�,������+�@2SqO@�ڦ�Eb��NH2*|�Aɇ��	�:�?�L�н�\b�ƕ������,IQC�A������*Ѥ�׃��Vyf�G���t�A��D�z_�֐�G�t����}�b�U�Cm��I��u;3�����tӨP�F<4<o��j�6��%tE �o/�O�/W��ND.�CU�w݉�Zl�^�e�ݹ�`s�<B��14&x���-.�.��'��%D�{َUf�����a�Q>NTV=+�$�폝��!�X_����H�R �Ml���x#ÇU��]u�?~1�ab��~[��4?��������THra�l�4�3a����ֳ�VaOyP������bJO��V?��+�9ri���'b8�?e�܅/�d��=���A6��~�1
�6��1I���KJ���֩���,�i5�����D�����=�|�bCV���%�L�L��>�Q�u1S��t*>�&�m���h/�/�T�X�x<���6;K��QS`*T��j�N��rk�ݗ����e']�,��L��~�p��y��(���k�>ѕ�ѳ���J��U=e��#=��|]Q�"��[p":\99ͯ>~s���4���h��l��U��@b���5@���TG��{T�����0��A���i6U��l����H�0�߽�}#��H�����%�q� 5-h{fl���3��P��G�^y<�A_��{A?
��'m�����=
�;?a(�{y2ͱ���k���mu�U�H�ꛟ��?{dB��5���ZO�~��)���P�z�T���:���=S����^�'�D��ŏiT-*�~��!lg��l�}/*E���u|�; �S�z]w�r���:�hEŃ:4[I�Bx����+pG�9��%V��ZF�Ez�? z�E?���W���L��Lȴ�X�ͩ�!�\EOMY5����XUtS,���hje����{��^e�}�Lz�4�<�C�-�ˏ�)����F����e!�Ii������[�f�/b��X��r�/�2� E�5����v�c�|����K��VBH�Ez����5�wG��x57q�o[�6�B\��Ŋ@�JP�X��u��@jC � 2�7���ݓ�(j�i�.`ﻼ�.��sͳm�	��|-��V�~/�V��Uyw��'�,N8��.�i�TB_0e�ɭWߥ�.�H���NN�wT�������V_$�]G�A.����������pm�TuY뭁N����|˚���L�7�l�{������]���������;�T!����ճM	�fr���6e�O8 d��;��Iݼ�I��Uۤ�����zN�O�#��u��7 �Y�ϴ�x�����[��+IĬ��Y��.ӣ(AG4&�-޵0H�Lʣ�t[�\�o�=
r�� ���[�-��a
ę�]���z��WU.ݦa@@�9���j�L;	J0���R�Ť��qcܮ�A�*�Y�5����3q�[�nV�'PyB�D�	D��y���=����=k�8��/Šfjw��|3Y��6��Rp���EEY��V�_�����|�Jmo��[�}��5����T��V����ګ����ek��lo�2˚�O=j�:����!b�B��q���o^i!�j�>���<���ڸȾ
D�����#?E�Y ;Z!P6~.P��0�G�#e�!q��H�,u��m��Ҵ��# ��P4���ʹh�z|][E����H�%�bU�ŚǙ�}�s:ظb�V��Dy�a��x��E����]���-u�����(��(�n�t)����� ���S�bX�_ή�1����z����$�]1���d�1�|��|�M�$[�FmֹTS���Cw*r
R5�)
v8L� u�`�Ww�P��~=�١�0��PX��͎�����/,0rv�jvȎ)CL����!HR3��3Dԯ�p@���J��("I���8���la�jgI�I�q�"V��6X`�<��=�� JSN���QNy��Ӡc���w������Tq�TF^*l�7Q	�<�ff N�_����Lj�ؿ��$l����셟�G�|4�!o��eG|6d��l��0p��F
�0YM�D�KU�;�x�y�S���v{��	�i=jY���Q�A�\-�/����	Gǜm�U����l��v��D����8�g,M�8�mH�p��73az�u�ӗ�\i�N9��r˵��YT���1G)L�s:O\��r"W�"]�ggeWqPo�G#l�Z��J�j���2�)
l���uid�S����S�)�Ά(l$��?�Aፎ�&m�p槸uԚ|�9���n1������A!!�U�E6�6�s�k<����{�[���50v����~��0P�}���k�x;�)��l�bQ4Hl��W2�����9�ʪ�|�	,�XS^n�>���B��+\�Ά(�v@o2T��)�'�yO||�i����%��xz��d �;Y�;}m������m`����f��Cd�����J��>Qf����*oSQ���ʩNw"��$���4�3MT��Bwԑ+J\_���~=WΫ�J� �Y˦��)"	}	�R���`]w�鱴��ؔr������ +LN٢y��d�z��c>^)z�·7w��e����@�9X�HGcȫd���E��b�L����8����څ��{�%Œq�.pF
"j���zv<t�7��-������a��dl���qgrb�3){`��3kD��������P�9��������|�6��� �U��U�~P��>oC�I���X�V��5���k{�~Oƛ��їh�")�n��c�f�8��	7� ��$�;\�39��Y��A33']t�-�x�E�ʱ�/��GÈ	������(�+�ѠP��~����N���c�|+��U �]��P�YuU��6��4{75�7�P@��
���[�q0>]������~O���7�������.��{��H*�!�)� K&��A�p�-L\��Y���Ft��\��펏����\�qN~��0�蠅��@w�#xӫ���􀁇�uY�s�<�1��o���F���t�Fd����q�U�-�i6܀�h�# �E��v}���2wyU�41���YBRix�:t���2��q��$xhLS:~$�~6q�s-�1(��\]T�,O�kY}rS5���n�i�{�&�)/��[#u�d��)ͱ���"Y�=��v���צ�f+*}������ר�c�_fP���|��WasR�!�
�􃲿�%�Za��k���R��������L6��V��g��|���(�o��@��%ejC �]�ԧ���=N4���#n�Ȁ���F��%1mQ����DcoaMLôi̬���C]�đt�\��~'���T=H��8�x�$���o�v���4��בIe=�&[CdP�������<������$�"�[��zr�־s��t)+u�Ќv��=�������u՚��W�*f��7H���^! YRlv�v���_�Y̸
C�5S�Ƒ,��J��v���'��!ƶ�S���O�a�^�
'�R;�����Àa�O��X�}��=�E�ضa�m��~�s�L���"��p��3��l/"+{��G��N\��[��-u/��aM�j�I�#cW}�&4a�2�HO�[�^��5]# {Ԟ��`�m#J��۷Ӧ�C�6���:�۞��tA�����6��H�F��ƶ^J3��m���%�kZX�V��&m�3�B����>�GmI�>�ƚ���eM�d�[�+��ƌ�'��b^��D�ܟ��XPXT�~LMg-V�iX���9@N��z1��?�Zމ���ۢN����3�V���`{��9#ޙ=�`��m���D (�;�,t��NԗY�?Y���K���Zk�ת�H$�����k�������v|r��-��H�b��玓L��R��S<dQ������29�!�|R�9@g�Nt��z����I�������<��Z+�{h��o��D��%�"��	�N�pp�S=AH,���yu��U�S{�=ƨ�T�kab�
���f-_���@�J�����#�~��3���ϔD[��C�t�=��"�a����7�U ��Y;~�F?�ә z�<��&���;�V΢@��\�z�mU�pT���d�*>:2��.�C��r�6*�4G�z��ߌ�A��L�&���39�S�����w�Mf/�겸����֎'0bk^�c�W>�����)RE3��H[���/��U �Z���R�_�>
ʥ~'lZDU'� ����5J�y2��(u��ķ��ȴ�Qc���*��`Q���W�=i�	�Ć�>o !��/���c�L�K/���{Q���j4��2 �PM%�t����!�r��r�'АZ;[��1G��(�y���p�*C��դ��w��ߞ�^��\S����KiAL(�}�JB��Vj�l�{�	��3Z��.ʰ "Cj#a��)�qIg#����Y�V�X�W{��`_ُsi:����؊�qn��%T��zgE�WV��pwZ(�zo��`�i`	w<��R�+���^჆�G��q���9��jC�8�H'8Z��߲=�J�"=J���Փ����ǒ,��ཱུ6b�a �?�\��e�y��*��|��rAq,�X@�2r��Q���7���}�ߦ�.n������1����?�:�i�Jһ��r=�^��¹G*1��0��{�.�,�"��J���+��v�|I<]��Ge���/��cc)��-����q�+(!�뼑<�ꈏۑ,l��i�b�`�%�1 V	U���>���G�jß�P_:���\Q>@>�(��,XgQ!��*��0[�}���^�D��=��4�!v7B|����wٵ�'hE�0k�#S�ޥ�����~�-�r�5s";�Jٍ|B�e��V���?>ߪ~H�Q��,������ ���+�Ԑw�����a9�N�>�����1LAJ��c��ZƐ��Nj��m9��]�:�G�1��l�y��k��6���!F�i��w���q��0Z s}Ȧ����};@��\M)]祵�Ւm1�w�~Qp��hK��/5����Q�{�{{^�39�K�|7?���a1��H�"ȿq��+^�gp�J��g^;�e�IuBO��b�p#���1���r ����ܜk�I\yuz�{��q���u�zr���`!w#��p6�HΖo��=����i�d�wl6fƲlkN�;1]�G�\#���4�F�6�)w�	��3�ˁy��)�rH	s�۩��5��"5ˌB�e%��:wP�Z�z�����*`������x���t��+�V�6U$�j�u⾸�r�Iҡצ�
�f������N�T�n�hP=���6 �K�6���v�����c��o��k�c�c��R���&{�����9~�ۨ���ʣˋ�r�N����ı�*�n�2(.S[JMvf�P��~��O���	L��rM��v^(�J�P���������v�-��ׯb�����ՋYw4��OSCkS��E�"�/����)E��
2hpљ�,do�o�� ���!!�bT��j��{7Ы�R�U�ծ�yh m�����u���+�E:O�ޑ9̮�1���|��9����R��
b����!T�����~�rp��W���wS�O$r�c�+H�G���I���;�b�t�K`{�Xm���A�lȨ1 ���O��fZN�c�W�t���z�t�9�>n]b�	���t,Sh+�mp�OX������>��xT�����跛�[����:��o]������x7T��M���}I��F|�=Deǭ� ]�b�Pǝڍ�.�h���l�h�5U�0�ɿ���Y���4��㰀GQ�]S^ڈaת��{K���3-�q� �}o}� J���:qG!�I�&H��s.7k-f�}e���L+?ʽ�?Hx�
�Y$�\�>���G�����B��%�K���)}��/�$eIqoBo��89�oi&x��M�
^�� �5
F���R��&��jc���B�̀�zVw�o�"�f�����dn�Qg�zc	��o�2�X��w�H����>=1��l4�&�]��g�!�������'�'�_U����~6��ڞ1V��G�i�e>}�S�g+� ��2��=m8���*���^*�$�x��`נx��0��7�G�z��/��2R?�v%q��J#��̧8��ݏ�+�.�
5p~n����k��0�̡6D��ј�>*�)^�X�R��G����2EeS� �- �>}��XK��q��*�y������X�
o*�(�Ԓ�wUl_?p������M�;���:ѕ���.�Y�V$�V�ކ$W�J��j��L'�`NF.K��غ88�Ke���ǡe�h$=�L��H��}�>����C�@���S �$Ր��LJ���Z�1�pd� �%�9y�P�;=��9�3B��V�'����O
����w>��ާ�tb�'.�3i��b�+i��TBQQXS6���=��pI{�0،�nҿo��N�{O+�>�:��E:���s�L���JTY�4!�6�P\'!�Ϻ�mԸ��>��Ƴ~�
g���W}N����ZQaM��X�;&/=��`a�-xX�=𑤀�1TUkƚM���e�G�}��Lc�i���r�@n�;}�cKGW��.׹����v��W�A�٢�ό~e�c��6\�)�]����~6�P����(������h����~*��ˆQ%I�̭�S�+��� `M!��ԇp�����0{��Y���d���)o��}�U�o��[!�z���g�S�n��S���)L��:oԾ�4A��;�L{7�b �<�P�u���/� �b���?�s���V�u�ƴn/WwK�|��5L��4��� �N�]����\_f�%��EG��~��
�L����c�.�5�;�/�(�!<�Z
�ՄC�n��z�s$�R��i`/�.���ĥ��'"���!^��/�p�!�Kظ����K�IRG��x��\�~��0�?�|?~13�r���_�g��* ��r[d���ol�YaPL���8����:�{����JM�|J�؍6 �a��?	
��M�.ɣ)Ў��xf ި��"�l}�AV���Q�7��!������pg�0:/1p�ۢ�W��$]8��A�&��7��\$s8��4^# \�	xUm�iҌqչ��ۨW96.�PP)Wզ��E+��馇{Rۇϓ�B�WV��U��wd6�9ǈ� S�%P�����5��8���~=�j�S{��u:}��_��L���������t��
�\2P�W��"�6�^^�鄜�C]�S��X���Ѱ���k��moy�����B���i��Dm!	�z��.Q�>���w?p�Fi��	}j�?XQ��q��ಪ��`�'���D����Z��Ʀ�s()bW�����I@����Gj�7���Z� m�X.���YeQ��s�x��.����+V�'�ϰׄ�$�Cgf���h.fq(0/�[z�\�<��H��#T�.�S�����缃a�le�^d괘����������#I!�0��R�&���,��B��ʉ3��憒��V ���i�t.��I0	�>����pݓu������nfj��=�Q�Ji����՟�%�-	N�P���OU^��H�R��=Ѭ0�$	u�R㏞��d������8Z�Vӈ![[�S�O����͹>�:E�3I��Ϝ!@(D5ٕ?�� "#�S�.��	��Ё��ukI�(����28"ߣ�W���cu��q��t�:Ω�G�r�z�g�8r���vP
�����G�ʐ��P�"�?�!�l��	����9��^�lu\{N\������&˄N�-�
�Q�aӣ�&���4g!0�
d�p���,�g�O3��?R���beL�MO��oUL��Sp ��
��.�l�e��~h�� �ʧ�k�vIg��7b�$ �R}�2�d�Nj�+� T���}G�SҊ���u�#M��,v�����V�:N��]��ÆD�4kQ䵞�!�6��9T	��bp�$�m��L��)9Jhؼ&9�F0��C�륪�0�!������j�P�ۡxn���A	j��,�� 2KpzX��A�[�Y��hI]�f���8�Z}@���E���_����o�cH��;4�^��n��T��%���%�g��}�g\p��ncI���/��������|)�γ�an�^��jJ����Ա�뮖*�<��iw�'�=a?e*Ҫ����[esYR=XT1P[F��u���9����a���ɂ�:�V��Q����O�bp��\��gI7�WVZ�z-I�$�����s��K��M��${KK��MHoHuK�1���dwq��UMtT�(���({HX(�ɧ�.�H��5u������9�(�>_D#��0MO��u3+��w٦�	��\�I�Y��LL]N�C�"E#��`�JkV���WI�c8'�S7-��E9�	4�c�8E�v���WQ�O��z��:���յ)�R�.9����� ��a��k�g�Ǫ�͢(ǁ� �RN��ݸ �ي��yw��N\(tx�'�)A�2�f��V9��ꐯ�P�>�`�B��%�gw��,%��I3bЃ��+j���WA��SB�l�ķQ6���ڔ�R���]'��IV,�ɚ�i�P9@�C�u^�O��@ 6~
�G9�1	�Wz��ݠ�+�ͽP��o�t~��N9������E��ޖ�C�&�^�8�����>�#-�:"KlQ�+�B����ԲC��|�g�7J{r5{*����V��1���/����	�/�aQ�%��8�X'N'�<������\���#�ABop)�sn���n�QΉ����1!��X��ЌJcA�Lqp�{�
���La�e��cz�c|���$D�eP�����I.g������-� -����bَP�����2�[�~�''�b������cDge ���ᇠ�<ˎ�xp������2Z١�7ŇA����Ug
�!�-IN�a�x��$��!��|+@�!���g�"����T�!���ǖ��1M��C��H�y x��m��-,0[>��B�3H�ch�]p���Gh=X��l޲���qJ�o֨X�����[ԓG\�
9�nڛ�㴗a��{"V���C��$,e��go9 ?��MQ�{S?q�Q	�v?�t���@Z7�n2���W�`(������+/�ډ�GRH����BE��vmS�Ǭ��@p����msG�?X�+y<=�l&؟�<_c�X��-Ѣ0*&{��}*<Y����	��'��sCR�6<̾�,ID-�@ߏ�6��v���K�8ڤ�H�P��X٫L���E�ę�́�_6�{Z�~`8�#Փ��?!�&%K���Ƙ��eP�f�ܻ��� a�Uc������t%�$q��b�"ǳ.�;��l<ԩ*/���L�x��y.Of�����]�ZFx<�����v��Uh?a6��nu�7���*?���7ʮ]��%��Z4_)�`��Y7�GΘ�dqDzC�{��a�|pX��C��=�]�k�<ۉi��c�%�!l� e�I"�<p���V�
  �&���2\��&���Mϰ5N���e)� �3r��J��C���a0�Ϣ��.�{&��Q��y�� �ɻ3^!��f����h�4UO���.Bk|�QH$M#���#"C�Qג^�H��3@�lfЦ[����a��k�a1��U[����i_����	IS�2�s�6��G����SÓ *�;�#�c�u���$�/��h��D�F�F������ݱ �V�Q�f,�`�SN�f3��3N�|Y7�`�E��i9��ګ ���e��s�V�P��Pb��~���L�x�D�� ɡvZ���O̒(�W�@p���, �u[��p��&8���W}��<�K9I�ѧ���P-�$�j�}Ձ��f�Λ.O�N���ۯ{b����r����U���	߳���uG��wf:��95�T�e��%
�d�����V���"d��#;��9�D�)��F��-&�P#ȸz��؛:=߯��Cυ��_U�Q�BDP6����|m��htRV(�I�yt!?��u�,?�[�=J>!8�MC�����|ߪD��b*��	9�	5����i�X6��(vW��IS�|�I�J�r�2�Գ���7*�d5�H��2��oЋ�J�	��$�������j���Y�o��?�4E4��S��x�x�r�Lҿ2^�,�zE����ɫ�e����K����l.}S�2�`+m�Qp���g�q��A'�D��Kxa .�G���� !=U�t�$Ma�_��Z��AԄ5���RoP;��I�Ì4�f�����@�z�[_
")I2��U��ۛ�+���?m�y%�]�*�o������D�p4�R<gI��ؑ����?OIr�x�����OSN],C�b���tC���f�9�Zهx�v+��Q�d7J��Q�Z]�����tڅ����&��
�8�����zDӍt�()o8�n�ݚ���+��C&����Ϡ����n�A�8��[��O���J��0�3�B��S��.n�r.�����b��c��߀Y����s	��S�+��{���O�!��_���ߋ� ��BH� ����ߴ�6y���v�=��tڂ����V\�~�Ϗ�j<�	݋t���L�g3��{%�����56d'A�t�f'`�:"T���=���R��hl/�O�-��5�^��Y��Qσ�Y�G�����8*v2�)ow�iG�
���ł���h�p �>�����_�<[��zf�7�!�|!�S 49�^�|/�J}�F"�m$>�Zx��6�"�"s�Rˑ� 4�<����7?�>U�lN�#nq��È�\%�@J�\J�����M��68>u����`"�-�3⃷����%���e��nԼ%g��kr)��j�F7��k��[l;D�Fː���x� vh<DX}�.'���������%�=І���A�����`��9���DB�?��YHjb����N=IO���P�D{4�L����K��%�-`7ֲ�����&jS4�
�W�󕼼<�P��hfl �wr%S9��1��c�Ul@����.�*�q�r��mc��%�i���#��D��[�2\���n��Z&��q(qv����^�e~C(N�f��
��L�̯�Y-�й���b�Q��Z,�<U1&l����nq��?�d�/}�sޜ�NdӅC���Qf�/�q]��D���~�	�xn�F�*]�S�{��B���J���8#�o)+]o�B�2��|`��X�fy�(a�Y^�۠���^.3�C��>��O�3+�V�c���^RPm��Д�{�	EU�y	�"U������ ���U�}E�O�"z���`"��G�ki���qB7̜��{#���(�
4HjA�%j<�]s��k�*���6���^��T:��p.&��7�1+�dGp|н�o�5ݸ�f�3Z�4�]�x��	�3/?T���2�`3��%��ש�Q+�D��Fp�^b��Xa$�O�H�����Z�(>��)�_!����Q� s~%�׺��3�-���$���Uq���4�gm��&��[|�4'	Q��m�)}A��������sh��KO�H�6H.X':@���d��z��r��N+A0m���\̚|�9��VO�;)��**b��`V�v� ��� �VGvT���	���c�-���9�]D�=!X�wR�����r��cfG�Q-!G�P�7{�l��;n$�+����1�oXq韎��n������..����_S8�<�ۿ-�a�gƍ��m|���[^(�?Bn|������D��_'��YJ���\v�3�?�Y7
���ȍ�v)�Z_3b�
l�2Q�z*��=�s�n��(�K��]f⢦
�%6�����T��B�,�%9��\Ǎ��?��u*��6�RWe��|�]����4gu������b��J�g�& ��s�_�#�bp�[^A��!���l�Sshm����δ����r��,\�.���z�7���Aa��V[i��<nk���O��#��w1�(�i�՘�y�s�4<���O�����KG���7h.N��eJP��m�S=��j�)Jg������ǘ��M��C��\��y�����t�L��~����#�(Ǆ�J�����4C�)����
^Sy�:��̂W�)�O���9�g�/�Cؤ*�Q� U�x��'�� "{o�g+��p>/�N2���%�D�/�Ą�[��W��̄M�Û,_����,eH��p/�j��u~ȑ�BQ�i�C����L9�
�v� 7�{]��̺����*L0S"�ӽ�D!8��	}�3�!v�~�ٽ~�:V2�ٶ��m3f_d\Cw鿻=@��%�B�?�*��!���S�A@�i��B�`� �|=uóB������nt�A��֜)I�[��~`�?��,<a�C�737jA.l_ud%�8�z�{�qOmt`Z	l�H�u���XV+��\�{.Yq�ÂN����÷͋N/�h�V����3W��?���zj{�MӤr��F�݊X-�.9�~��u6J%f�M�h?��?\> ,���U;+'2�� 8s�x��6��5y�}}��ؠ�6���&cvm��� C*4T�l@Qm����I�M�6�4g�Hy����{C����g�i�Z�g����gܦ'k����v��L����Z��͆_�G@�IL�H\��j:�D�z{��kU�� x�
±I������nt�Zf1\������;lΗ���&���!���'6�6 Y`��;S�bj�}q'�@ly�3	���#k]9
�@�Τ]����H��$�b�F���l(J�{��{Z����,���������?!�!�-vQ����u�]^�E�w�U��Hg}>��iTv����b��0�B$��0,s���9��ˌR _��k���<F��|1�sUU9�Q	�k���,k��U����}����y���pJf�m�of+u�6E0�E�Ӎ �#X�����F7W]�1��ԥ�� �G	�~����O���𶨒��3)�"���%�0��
;���j�4>�q`2�`��0���ʗg��I%�ɂ��[֚N1�X07�B5����sa]>W�ś�llb� �&�� ���Ù��lp��xK�7m�D���Sb���q#��6����{��鵤\5�[�*M>44*���ܙ��>uH��86���'~.�0��n�a<�w�I����P�2�$�!�m���|��=�u�rkҘ�y\��Y��`s�
�ܭ)ҍ��b�� f0�]�*�(���F��V/�ՌQ_���H���D�����b�~�y�N�] �(�z1�Wh��F0�v����V뼠�1�!�j�?>U~3�V���o�_��&3jS����E�=5��Q�M�}ڮ �$p/��E������R.ʋł)�����B �LI?��-iʨެ��O��4n�����	�{ !F�V��?PJX���Oj`ؠ���A\N{��=��!��i��$�D�'Rt�<sC|�
Q �g/�]�w:=��)_�&�9�P�bܵ'M\�]J�=f�V�X !QOCp	12}�Fo��,�^`�gh�a�oa���`V��l5ª���9��Ȳ�o����#^��vv���2{t��76�:��^i�i�L�3�~|J�S��Y�F�E9!���i�9��4����4 ��B�X^��\{������-�ܱ}��j�M]P�T)��'7g���$���{�&�6�d����[�I�S�����|��FHi��� ��+��G��oذ�����B ߥ��t���:�td'��j��,�<�����RB�'�k���	��=c�Y+��T7���ů>�BW�������ӓy��� #{o�~�b�����M\Wyb�,�-�����d<j�U�6?�z�-������\QZ��*�Ƒ"
����Ⓚz>hڲh	[�@7,Wږ���n����弓��|f���<�~ �8��T�`l����ՌY{�:7>	;
�ݏ�fcQ�?v!�_HJIBuA��%4x���>��f�ӳO�/5�o�uK{�6ʾ�S p�1r����<Y� �.p�>��#��D<��#F��#���6�ץt[����%dW��M�禌��}�>�0�a����6�P.��v�0�4Ċ��B��J��Y��j~z�X��{U��Ly9�˿(r����K��mu�9
�9�S�SySB@PG���ai8G�����tY���v�qf�2���e�NEL�(Z���Ǽ�ُ�F>;)�L��\��=1uc���=�[솄�p����Pqc/a�IM��n��̓{so�
Puj�!��)'a�]�ː�z�%W�C,��B|���W�9�{XpRk�G98Lȿ��m׶�����V֋����l�@Xg�a��C?�z6�bF��^�C��{��K>_dd-�X7�z��J�j��+���Hʾ�9-@���2���[�j�4�:���Iu������B�[�-�$�`�fak��ĳ�G��6rr�>�cr���V�tn=Mnc%�����8�:�zX^�:����W��ԃf���6j�Q�H�h��$vcL�bn\�>UUc�-i����?�S�5�ЄTX�.F�R�{�%��L���YV�'��p�hd���1�1T;��^:��:���:�7˼�>2�ح�� �,�Ȳ��tlF)?���/ħ5��r$�%Tk���W8gK���F��;��|u��W�x��O����S��h����&"���5��x��Z�T���%��6Lf;��3ȹ����k���h���J2Z��_(tn�����%�ZD��[�?m�VPd�E�fk55b}���oB(aqW7>J�'�NɰTw�
G'��0��:��z���*|��x2��,w!g�٫~o7���YÐ���d�S3�=p5���qz���)�`����r1lmܬ��V.��OKhUy0U�z�W��M�N�,ja <�"����߼0{�h��K������߬��u����/�n�?��B�.��~[�ES���ޜ�,F}�F�Y��U��Ԑ�DRk46�A�,�r�+���Y�1Ns�S�zQS$I���$�s,���	[����Ҥ�/Y��BP��R�K� j�^��
��J�j�yz
Y�td�gy]�6+4k`f̗�Z�l���Z!��h��"���l��9'.^����N��*�9���,��y�g�^l�g&
�0��t�3��b&�ڐ{��m]��p�@J&l����e�oV��~�.'A�Zz׽+�YDݟ���k���/�7��1}4�T6�!�3u�e6�ߑ�|`����^&ՁS�#�Ph}"{WEWϧ�������Д\2���]�B0D��uȦu��� ������b�G����աV�p%���z`���U-�m{�E���z	dKVYJ<9�N!����Ǘ����G8��I�	��ɺn�h#Y�ДTg����9�K�)7�M?��.������9�]w5�j�mdgisr{Z���Br
.��j��Gq���-��)�焏X���(���	��$���)V?#�xnY���*t6�]OhW�7׌t���
z������V6ڳuc��Z3;���I��Mr�d\�`6���3j�zq�N7fަ���C��P*�'����0����}R�i����Z�1J{xC�@Z?�-~p&���*���e*��i�ߋ*�%Qޑ�� ���S̨��g^C`<�Wі 1X�������@T;܀rMC�F9Ѿ^v�l�nh��a���a���X(�$I�r��B4e�z2�z<ﱷ�M9{aOۖ�A�wbO�'{Yu*�n]����6s�Ek�����1N��d�����}���-��Yi���Яdj��8}��ug�c��f�$rA�pc!�e�����q�ai0߳�;�t���D(��ɮ0�!���VUj9p��t����j�1 �ρ~�m����΀9|���)�W)�4�LђE,�T���������[���Vd�ߑ���]Y��S��ݐ�,�Bo�梪۶0v��@�<�����F��,)f���<F�COY˩#I\=�W��f�<J�Aبv�S¡��h��W����h�D�q�p|�b�/ ���"o�[RW��jוs��Wm���. �m���w��I��*�Q�LV֞��Qz������xҊْW�{�߿�xW$�~M����p:���f�=m��#�/^�v�Fv�����,�W��h�9I��+���i�y��1J^�gY�@d'��})�����Æ$M�aq=��x��A�TQrJI����&�!���ɉ4K�k<؛`�h�����&Ʃ�SO��^Ⱥ��7U����4BB][�,�i@�ۑ����1��ť��%�׈��K�Y��1z�mҫ���Qp���C5:^@�^L�s�@}���z��АvH�����]i�"���<@��(��H.5j��w��)���&�PX �-�~�����z�H~�|8f�#,
����A?�Q����'�|܅ʍ�9Y�]����S��@�5;q\(�'��X�4����#J�"�'���vn�M�[�r.Ϻ���������¾[���.�d"dy���T-XB�̐1<R�<������i��>�Ƭ�A�^:����Q�Z��B��z��1:���ξ�>
ilb���o��4�p��5�*s[��K��1J����H/�������>���N�L�ˋ���m-K���D
���ۺ�V|?<�{���*w�4�#�#E�6b��dT�Ϡ�_�`�KE��R��3�4�G�K�#㇜� �*��cp:51@���/Vy1�bu�8G@���+���E��ĽMS�,�Y7�\Us�h�g�������Kr�bq��&��m�|Xw.���@f��p/'5=�qCA��� ���3�M�/Z��du�'�@�����L��X-9�&ߴ.�{�G����~�����fu9w���߄��"��|̕���c�Ӓ�ǫ�͘g�z�k���k�2�xY�,k��]�����Nn���ϼ�Re�g��C\h��@&E���dA,�x��0�w�q�]�w��i�	xa3^Z2�$l<΢�"#RӼKP7�U��iG�������.�sb\s;ǜN�!�~O��'�6�P�_��2�]F�4�~�MF�]���s��_�����¥�*�����ョ�fv�zK�(uj���F�o��q�U/g΢�r�<����t�#�+�)SiE��Y7:�;��}� ��!��w�u$��V�튲*sұ��&�Gq$,�p�T �NЍuo�����-�� ��d�9˭߸����*�3�[W��?Ë�+�`X�Ƀ֦�kl�Pl-Gi���t|��v�cԹ�T����(���s�l�w�
��x"����D�*�ߪ�S�	���}Sa�t��*Q2��	�ٳ�΋�wԜh�XS� �k��KW����$�Ow&T3M�s�#[/�8���,����}}�[p��G5���E��\�BX�d�L��!o�昻r%1z���Qf̳���p�hl�U��B������R5-���Y�UI�&G��.�j`��q�����DL��J����>�+ά�A����l��3��g�I"�F�f�PW���a�%��sPd����r���߉��e��g�PR�Y`隝v=�a���{?�fmF��4��{@����)٦���e�n�3�_��5�|]\���z�WkF
!���0Z8*�yVJ�f��)�p����A���Jw�^C�j8��B�K���Y�!��/~��Y��t-O�eH�/�/�7&yԦ���x�J ��7�|(G�e2�9�|,5]U����F�e~E�v�Ȼ�*P>o�>vy�����VF��³�!���G<�����e*`�����b^�˟
H���u��L������Ǭ����7�M��b{A���V�aiѩAC�,���KȒ.�����b�(��;�?�r0�J�Q ���j:o�Ҭ뛵�Y�g�Ima��Pj>¿Λ�l�!�-�=�V���T݌7���k_���Z��1 &r����o-L�ɡ�1�pˢge����	�h9�Q�fq���J
���]ɘK�i������+}3�D�,�����gLDT;�}(f���(I���ҿ`�n�K����WN๓����h����u����;�xSA0o�5\9��B�?̅UO�Wn6_�Q���F�28��#h���$����_�kӬ:ua�	1Oa³"/��C��eZ��$���!_�U8��GD�_����ز#e*��T������=i�������<n[������,����wW	���"��Fz���aw5�>]�� ��nI-�����/[dٻ����6qe/��X�tL{4� {B>S�R���'�����q|R�l�7pk����\�"9��N:H�n-d�xr��x�H>��G�'�~~�]��Q���3���+�;�c<%�Ci��������������pY�J��]����Jd�H�=�C���c�
\u'�����ɑ�1�/�|��A+)�Ы�D��n���ބ������!��~�a���Q�Af�w"��`�1fo��|U8ٝ�y�	�<	�>�D]q��%�ڵI���T�w��Kg1�@��諦��VUL�d��2���/f��N�;��v?Lu#�«�jW�3�#�cl�ڮ�Y9{!�NU���Y�I��&@
�!�d�Qa��n��o�0��fҽ�?Xdθ�_X2#�h~��ð^��o�?!�ARz{b�F=W�͐Ç D7���{�f�=�ؤ��� �7t\�ɑ��y�����>�����߱��prǥc>|iu\w��N	N���B��]e�(�p+�u���a�͝�?��Z���W��Y8�C������I�RTP%]���#O]����m�Q 9���Ș�x�+N��0���TaIo[�֪V�:�)��Z�>�)T�H�\,V�,S�#=
�^��)tcC����Q���'�������h��E��o��#�,�o���^ ��?��-�tk�i�տ�۶j_9N�h�t֙,�A�m�,�g��a������lT�A�:�{�[C���F ��ל�H�b�SNvyIXR���Zy	T�Kc�f�ӱ3A}��Y�Sw9�Ę+N��>4æ��ꐝ*S%�7����@�1�ٱ�Y��.�\(R���H�d�"�\/c��57=cۉm�����Ua�#��;:&�����;��C�}�ݓ?�p��޽T���j�w�#�@� �se����S�z�cz0�-�qM�͗
��4Q�ޏ�]IDt X@M�?(��~I�����o{Yy,�������S��Ɨ,s��6�e_&���[�|����}�E9�-�^l�*�/Qw��}(���>����0�ɳܢ��]�)^�)�57vq�!?`�ۼG?�p+bc���h>9h�0�� y���������X<����2O��\B��9��#�->�3S�BngNL��a�D]��@>�����I�ܵ����Ij?���ر�M�^-��P�X�[nz;5�s3�s�i�ް$�np�g�F@�V�d�3�/8wv?^�#&b��P%����?;����'��{�M�>G��D ���:�TF~3��0�KOM\����IE��%,��*w˚���*ʿ���}��G|�N$���L%w�<���_AbBU��!��B߶�.R���y��O�N�W �����?A��;�>�󟛏��.td,}�	�d.p�;+�'����ǐ�Q�fQ��VQ�v��m�P�ʿ؍���z�K���p2���0+g����X��1Rj�J ^�d/`Izͱ�+�W]��R>K!�|w�.b��;���
ʐh��X//.TY�,ek݄Ф�94��)'f�D�o���t2¯"�8��BB������`9��ﶇA�8;��ԍ��)]�PX8��KV�q>��iyy�c�Ut�P�;f�(a5�<�����
���@'��Y�<~j�k�#�| u(-�򗢽�
k��2U}��-�^��
��������<�?Ì�.� ?���
_���ј������؈Dz���;%z4/��ek��7�0�:���ar�:��I�83��������U�^�tQ�4�Y)�ӹ���7;���asMl�]��׆f�2�?y��Ta�>�3��Nd�W!^�a�?�B1$e �&�}asX���1�-	�Au���¼�I%���R��\ ��]ݦ�p�N�*�>�N=U�43I���NcO5L>N�3��qDvf{=~IC%����P;�&
�E���G;���5���E�)c٘*}{"��^0׊��BX&��!l��:�!�<Hϓ�L����Q6u)V_��51�ez5��?-�y)�l�������k�WcO��Y�j,?�M�����J�OC��b�d����W����pE�<{��|��<\�B;�<޻.��@����=��ҽX��w�j-��SXʺq�k���-��N�[����(eo�YSDЪ���'����Q��ߵ9����=>�k@B�!m�x'Ů�9al!����9>H�v�FV=�����.�����
�b*툵�q�} v���-dۙJ�7y:.S��<��ɱ�t�tC��6�#c�b��#<%{)�{�8�\E_�К%!�o��s���#�pӳ$�鞏��*��"�4��xDӣ���0�P�X�Ɯn�U�}�^�����v��.Ff�WT�S5�}F��en��GJ��B��Ռ_|���ݫ3�m���Ỳ����k�Z�at�G����
t=�$���2U;��u�%lԭ�,�����y.�r�|�9`�U�s�m&��A/?�r���G�i]��,W�_S���k��<P�d��q +��嗴��L�RU�C�g�F"S��M��WN� Y����콾e�TA^}�3;���I�jS��V��Dv�A�a�ҵ��fj�a�ڇ�t�b�QVu*�62~9&6�,���
��2G�\�,�f{Ա�R��z�@�`�N#�+��W��7��k)8�Mpq���Ha�J����~�~��#����&_����	��O'�j+���wv�vۑ�����ﶲ��:�ُ�n�Qf"p=���>��1� �3�4tbY�[��>��ۓ���Z��d���]p4�� ��Y��~SGj<%^��51=fB=������[��
�|}��m��)b�.g�V����5m6:��Ά���7ϳ�8S9`�v�!�:�U��6{�7IY��j��w������=���) TE�}�䛤nZ��$���Xs�?ǁ�zK�/S�w@�8����dVS�m�ރκ�Qڪ�k���oF�	�Q��]^���l�}��2py?�������cĬ�l<,����� ��{��\��>�s���餸�-�w�������[���&?���Y�C�yZN0�Q�w��mi��Evx��6�Zn5�p�\�D�.�7�����ᤴ��oL:�\����j������N.㍟F�U�8����]/\�]N�,p���`�@�)6�)����KT�C�覴X���J��4�чd��[�b�q4Ku�:k�W��tV�uY' 6���d��`��CTQ��s��:���W������̨;4�$��(���5W�տ��2H�%	��i�q�[i�>��/��mx����H��7��Q=�GZ�t���`����*<Ҟ
 ��8%�Ǝ�%Gc�/�|��k�,XH'�u����A4�f�D�}���� %�sׄMk^z(�X�XH�f�[%n�ǿR9J��n��	H꠩�5�'��ݳf����@6�9be��,���j���2�җ|�O.�h����� � دR\޽��LRO�����W�F�O�ӿ,7��Sb�t����3Wx6	�S:��E�5�{�\9�7}���iN�h~��U�pf��ZY�Z[~�J����A\/��w�,�,��Wh:7O݃�
B��o��'/��*T�UQ"˶��v2h$"�L� ����H���]TE�^���L�KπѬO��̎�."�~�h��m�u����p�'ꆟ�1<R�5�H5��%�w0!�9�ZA�}9O�GSa� *;�X^�<
���һ���gv��N2���uvLDYZ�.���I��zs�7�����c�M��A!���
t)��#��C�N�3�]@���Y���&�+���3��e�uH����4���#w����N��6��|(LWF��\��	V<'m3���#�	Y���©���Iw�?�z���D�!G�9�~��f�G�N��-���<zN��U�tܑ�G}��ۅ��3�7�)-��୫��e�p4{^t���Y%a���=`����	��Βo�s%��z���nx\��\i(�f|�%@�0	����/���x]�R�e���.�g�dPd|����j����Z�6+��#�������wE&=��]]5�I��v����e ���1��؈�iT��v��H�~Ɉ-���\��_��,0U�S^B@�>�J�2�n���Ԭ��e�3���+��d�-��U�CCs)��i���ҁH2�]�,xuJ�z
.'*�H� m�!�3�ڕ�I���J�������� ��`i�9���h�f����u�Zyk����9?��(�U����cWks��&�.�],���f_C�+��:�ì�y^�db<�����u��o����I�FQ�qw|�����m�[�㖅��UU�@�f�7w!�e�����(3��IE�1z;�Սm����8]#�[Ig���'�!P�[K<u
�_�ITm��-�����0fw"鑴%e�5v�]���8�h���(���Z��JuY�e3���N���<���ʖ<��P�����m���r�1�Ɛ�1Վ��"�������V��`�J6�x�W���*V���ΐe�Ճ3�� �R`؇�"6<��J@�!�yu\s��1�1�r 	�-���3Z� G�'�
������?	F�J�8$I�7���"�8̼l�#����2��f�5״c�����vc��s�z|�@���]DbF��X�6���Q��7�#?��sp�����!��c�
����!�������[\�m�T)���V�ѷ�A<�߰��&}^����H����m �mj��ٹ� �B�x�(Jp�Q��/���&}���X�:�*2sQƲ��٘��:e�tZ,!W,̱D�����l�z�|����>,I ������:�ܭ���E��̘�_����#�����~w8wr�B�[f�RYڎ�����/�9%���)���GZVJEH/U� ��!�<��j�B���p�#���U%՗	��c~�
3����