��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!���"WYj����i� �N�7A!�@<e�]ң�;��5D�監p�.� ^+��Rk0;Õ\z�7PF���p�e��	��j�kdD/���1M���(���T�e+qr)zD���FWkV��������\���mk�*
`�R���	j�' �� m�cD���9:�DhT]�����۶�����i����ޙ%��d7ܷ��	�:���U��(�����#���wv�pFc�o�m?���<�δ�7P����( ��(�����1���o.O����BE�l�pSX�m����
'j�ߑ?�a\����3!���Dꁖ�0� �a
Ӭ ��W�?Vw�h���!Kn}�g�����׹S&�044�wZt�ܵ�XV�pi��e��n��ZX
�HѡǦ�P��v��>.��l��<��v�M����ws8�Np/�ZS����N�o�jh�C���&l���,F����tm������-wX�Z9ݖ�e�t|Bp0�������NLt" ���;�a���X�7�
�^���ߊhD~�?nM����d��Q�!�rVuz߻m�������28��:��z��Xb�o��_��8�PDA��En�毿�r�~>k=�E��b���P������,�ͣQkW���tFQkQ����i�eF$hw-M�6j'��xqU�@�����%M���nŗ;��X���U"�pH$�p�
l_��B~p�g�O��yY:�,U$U�j7�}+߫���~��8Vbd�� �	���/]ޝ4���؃a��wC��"%lJM�%����:�<�{5�L~�/+�{�x�v�ݪt��=��3�E�{�v3��%�ﯔ�E�����{~�^ ���0^����NQ
���qA_%^�|�/�����<%��x�U"���k5m��Q5�6/>��e�M���X���iX�'N��'|��z3�לx�mSP���0�{Y����y; z
����[�J��f��b�.�z�a�5ַ@x^�c�c�(Ƣ|�X!?��~�U�-��^``8go#9h[y�#�¹�v��y�q�'��|8<��؍u�t�������q,���m��$�~�^�q�\���(�I�KQ����4��8#��Z�jM%@-��\ m��P�0�V;��8$��0Zh�w�_�*�����_�9�k��C��X~�j�Ӽ�Yj���F,��T������F���&�$c�ǘXfo�4�^��iD�彨wg��$����D�94�8�*�՜&DЏ�3}
��2�`5�6��1��4�Tdǭ�-�d�}�r�d+��S(�x��Ğ)�.d�w�o(��ޭ|��]��|�&���?$'V�O�\���^�D��]M�����&�a��}	�|��"㭀 K�M���0
5���/�/�vu?��o��:8=T?obhD���h,��K
��{�5�� �CLJ��F���^�d}0�\nu,m�.���,�?�l�ڐ�D�5/���g�smX�%�a\��~�J�E�͈ڵ�֖ ކ�ݡ��A�bHL�B�J�@?u�2���@O�sK�JO�oM��2�C���q+ �IҳUJ�b�s!12�s:H\ElA��*����-��ZQ ��Br�,�-� `}֒�E���GK�6�"P�$������]�d�ʟ���s�hpl�+��w�"c���;�s���e͐�ף�M���n0����$���轍n�?��|�����v8��\���Kܪ^�zլ缾��7�p��6#������/9N��ѷ�Cw�/��U7X����e�:���\ޏ��j�L'�#�����MZ��?��2��D��3K���z�ᣜ�)���9�ZR��Gz_\���Ȑ&��Ф'\p!�
��2��٢��Ѐl�v{�K�&`6��9�>H����)�K�z���R�%o�^�Օǔ�|�JM�#Ųz�1�����,��i�3J�󬽩�������R��]��{l�?�C�)塚<7�J��5����5��mb�s�t� 9l�d�_%(81G��3����yX�O�x�Q�ZC:m���-\%f�R��#��̞�������2��n��P�[�jɶ�n�����w�}M�VT�Mi�H�e+���
��4�֥����d@���6lc6%<,�����~��u	��*I��*|/�uܺ��6��,M�yD@�����+-�6�dԪ�S��f�I��N�~<�f,$�<KiÃŀGr7�5��fЕ����A�7=yt�l����]�z�*u��}Y6��N�BtA~����`��c[����,�3�Ly����(D6���� 5T�K�I�� �P/@�m#��#��1��A���:�2M&�������7ӕ���Sݓ�)��*GA^���ޡp�aX��eN�%1�|n�r����f����;��nD��S0F����}�U�>4�<���g4�X#�$:J<'oV��qƵ��s�����σ��X��]�����r��Ht9W�(�OU�<^j�ǲ�3|���T��]-�ueFN7���X��;�6Eo�Hv�%F\�Μ�
 ���b�u�I;�J�i�Q?Z�F`(:�ܝ�/�.'���C�جD�����֦
�#�j�c��u��&\$g�j��mwS�EU�>�4�ކ*T�󤜋񫷸y�����F��φ�x�m9�r���3mi��KٞF|e�.�Ɯ
�r=�z�����8P+���q�vT�R��Z�[׹!�3�_"3�b���FE�]S�*����Ձ&�	��d=$bei$&󜾦 ���p�0���E����
Y�z�fJ���n�D�[�$yK����ef�xL9,߰h��?uσVw(@�
"(�FTf�g����xB�0�5�_���.e��w��L ��Ғ��G��Ȁ?K���W_;�>x� 7�'C�-�H.���dzZ�Zp)?�2n���~�AMڔF;:B��zy���?�Z��� #��&'���>M��c��5� [Iq`ԾD��Ν�iaSPO�8<��yf��S�)ZxW��H��c�� f��WpS|gdΥx8�c��B���<��S��D	���]��������6V\`�� �-j�ή��,�F����]�/J� ����U�o�� �d��B��{��D4�={;ո�-k��Kn�P�����A�<&���YҞ&�3#9�f ��ʌ��L�Y��MWs�L�Ƙo�+��d,�_"ۙ6ʨ��tT����&��Tr�.ܽF��-@���Uq� ��m��Hf��|�����iwC5���U�iS�r�Yx$����-n]�7�߈���?�e2����8+؄��!'�n[9�hz���	���Rm�� ����ĵn���I�>�sm�4rs�v�8�_=����l%GY��jt��:���1��X��W8�3?-�
F17=�ݨ �T��L���H�^�=�4�yM�9o�������^%���j]��v]!�&��M�nV���Q%��<�P]�o�*OA^��~#�Jc�0h�sn�dA�Ad�8�z�8C�k�͟Q�L�q�я�::�ú[�E���q�g�����%�I���^"�����w Q{��fV�\J��@*v��&V~1= ]YѦ��Ru~�2]�
��-VxŘ�9�B���8̊�����+�o��_�jq7�j=�k"�!�3���ܾB�)��S<�#������E}O�V��ucݰـ�L�������P�"���H-��w 0�
/j$��!Ѩ��~�s,�2_įo����|'���	��*;etx��~cͨl�ɞ�7}��?K!����ӷ���99;[HeE�ؐ��K��7Y���\8�bd#��Kk��qM���:y�PV�-� �������"XƟP���R"ڙ:՝�__������l$�O�@
eJ��ڝV1�T�Σ�2�=��$���@���mR�).��� ���P�ƫ��nd�$�\+-�h��R�����,�v�����������g3�r�+`�!x��]8��@��i�W��]-�s�iN���j������GQ�!�kvMo��������9�;�.|V.v�)OX�
9X6m�{z�+u���w5��8���=�ܮ�+�E@���N<���+�ۋC�]<�����}�d{�b��Œ�N���Q�I�>j�R�ݻ<�R�����)�?���eQ��A����P�*6�7q��o���1�d3s��``����>�{xb<�٤���(��&(L���#PY��5uà�9.���$HXwQ�̧���\k'�tI���4:Z�w�C^��W(kT[�}Cq~����t-������2���-љ�XiXh�֔�5Z�����\�;��fT4�n�G��5�� �)&l8�����.�Dy����ӣ�q��	#��� �����()K)�-A#`�*���V�"�@l�%hz�s��bJ��Oe�g��u^̣1��Ntt��/<'T�
l���/Z��%���`)�������~�kҸD,���i�8bJT�B[�MD_�o�����=kP66bh)�R2�XV��IxJ
�@.�v��-&��E]@��� ��f�!����ŀ�j��$������4�QDq�K$�l)ɀ���~��f�)�ŵL�h�<2i�i,ߟ㌎�b&�,�B?L�5N�k�-���)����{��֐a�F�:�a4���Ր�ah7�A��qJ�t���@K-�g?������퐆�w�R������1� /���yU/E����'���?=ݝa��!P��x�l�
=���o�;���{:dE�����|[`BU�&h��9�[O�7�E���ٳ�,�������:Ο�Y�X�M1�B$�^�퐌��.��|)���Z��W��s���
^痺��7��p@L�<�'$��{��WX�j�e�P6�8S!Jjl0R�0=���d�X�Mp��������!"9>ޢ�>Ѓ�@ �q�FSγPi�O���6��9e�IGU(TZ���vH��O�S��Ǉ�-����w�Pq�!�����YU���~��WW�{�h�v	QbI��
����.�:p��U�d�7�AB>(tJJG��&~��0�U��Ek'5Xs�b�.@%�P&��s���7�NN;U�=���d^z���`�:� 6V�Ir��(���B�Զ�&!\n.�c��o��ڸ��lw?�8�M�0=��^F�<TR�]M� �{��@A��}������&n����5��wC|�J-:�"VN�\�	����h�<�!�k�d���Csp��<8���`J�/������R��S���agr+�l;|X�e��L���3w����Mj��N�HLn�zw	�T6�=߇D����ǂ2�?s�l��Y�A�b���jv&� ��6�8�I��b���	�������4�㼥�UU?���*��î��ض�5m�i��H��x�c$0F!�j']���z��a	j���nQ"�]�]E|*�֐�tj��:�E��Q.��\��l�C�/��ݴ;�JE�N=Uݞ	�5�3�ps�Y���M��^�,ؑ��~�p�N�A�q������~�zc�$�YP�@bpZ� ���6�D��/eH��8)��ru�����1i����c~ |���&h�z&k�~�v���-�7�R�������$l�Ӽ���u+��[(���"|�xxI�D較��G¦:gUL�#ϝ�0 �����m�W}����*!@5��p����נ��L�L3W��)���BW[�*
��Q���,�d^ߠ'����##�Xp�3�6��D-�F�f�m�İ�5+n�eO[�e�����9m G�<-e�3̒�┅A����Ac��d�{�ox��F�u��#��G���Un��6Cb���u�)�O��.�L��O�h�u������"�qw�$t���N4��h�b�9�o�:�/�Vo8���lcd|*О���mO��ۼ|[`�$ǣ=3d�Q�c&=�=#.LM������4��Zg�j�@���oTZE^�$�{c��|�e�;��ghs!��t�����������(����є!��؅T�}{��:y��W���	��7�D �s	U���>�x�(��ɵo��c����5y�3V�>���Z�f`���J�@�����X�$Am�!9w�iAj�%�p����ރ�4��;6���2�j�|GW� �F#��^��0��o���;o]7����YT,z"�Ԭ]��ܕKn���W���k��W�@z
�i���K�x0?�*������"��SZ�R������i
��v�{�65'�N����2�j��uIi�g���M �]� �����0���K��TFz���Qw]�
&P%���������Ӳ󏇟��rc�M��& ��J霚� �<@攱��@��ץ�]]!D0�=V�(�����񕛡�q2U�U{J�j��r��	�yr�H��苄hgj�k��X}g �Ҝ��6������H4�h�ѠGc�g��� �ׅ�9�j��x?�tAP�{��;D����E\�y�@(��/���o��`�~T�_O"��b����w�kM��'����N$��[H/μ8�����1j�v0"$d_�p ��d�m`0$�W�rg<.���a/5�_�O����|(�⧚�0!\���B�2��vSD��1�r������rt���k3n� ���b8��@��s�0�-�s��Y_b�����,�<�0��\�S�C��kK`�5jo 1���KV�r�NV�M�\����]+G�[�{�n%x�qpϲ�����rC,�&)����I���wb�&�E��F�B;��7J�
Âcd?`�Q�U�"��p�0�3	r�"��{��o��`ǜoc�xw�3�P�*�}�~�x}��W��W�����5�[SΎ�(p!�r͙��C<Վ����|���R�����;�BU�&l�b2�mY�tj��w�}S�L�5�����(����t֌�[Ż�*�z}"��k�g�A!�̖&Ml�*3i���'l�ss�"�?\a`o� ����&�O���4�w[�a�v�;���bn�C	P�y��>��HPs��x�@Y(�\��M,$-[;s��?,[�E�-�)U�-�����,0���@^ԏ�r߄k�~�U�[n~�Yk5���')ƭ���$xme��K
�3��S���O]���˄s�8l��hjv�׹��6����6��ّF�m��
���B�g�?��,����\�Q�\�[*N8?����W����(�x[�2�n�̃�:w�a.:TQ�4o/��Zd�����5�X~�E��ߠ��	8{w���G,!Tv��T�����T�A�dwM��*��A��rwU8`<���n
,�v>p�8橉��&5����zW�w�QF�р|�w\"̲���M�f����N~EFG)��z:ᕇ���ؐ7'8���}�pl�d�N�38.u�{}a�*��z�N���G�����h� ����5*�[cB�8�1�@(��c����%YLhF��b�s ����#�Y������xsv5��e���n����#Q�n9�Z��?�io��4�P&ի�P�$g�d�����01�������T������Ǟ��b���EV�y�� Վ��xer+��3�|?Y�9�խz�fR����/����#Y�%_�G#A߯����c���>'q�Țǽ���أpC���٧tTL,>�����nO5]���k�+%�T�ܑ��;/J%�ሽ��;������I��`؝&��G��>������}Ͳ�$T
��ċi�-�����D;�R��uL�o�`KnV8��:��#]�T:��ЄP[��<e,P��R�G� K!��.`��CjK[:��y#N#�npǃb4F������T��V��Q�Q�o��5�f�NY��F�w�M��b������f��,e�0:?���M��֦���
�92�j/;c_qd636���g���Ꮂ���	T8X�;&3�ti�D����6~&�"��hr2E|!Q��̚��&!+E�i|S����/���2oq�}��33�7��X8}�n��9��?xkn��4�޸jd]eq_%�7�N��)*?n��e����"I�;ͻ���-�9��pOy�B]TՅ������TӥƱ+��?Y���0;����	0�\Ѵ���(�;br<|y��s%�D�:�JKT�}�Y��}�å��<RRbw���X��6�g �8A� �Yx���6��D�yȱ4,�����͚6��B?�EN���'�7��wc�{s_�],0��'��{'ϧe+:�a� �E������'���W�G.6֪H���Q���(�/kty���2iLU��$C�X�Bڰb��JE�����<ȺE�Q��^���7)��%j�L�D�T��Ϙ�y�~x��c��[v#�"g����-m ��g#��c��_�ȿ�s����hнiC���������K=�mrF��� 	��� !�f%�Mz|D����-<� ͜ff�B����`�M(J�Nޔ�XN�����W5�a4;�a�6ӥ��8_�=��T�,��(����ڄXd��Q����M���Nj���"�e\{7/��H2�=d����?�` '��>ʅl�_%\��|i[�t����K�/o�SP��3�Yعh̫�K���q�lf|:�Ș)o9��Ay*����-����5�&���7Wu�Uc���]��:�v��=�ߋ����6*�B�Vm|}:.Ǹ\�N���=�<�ա)B0�s0E��ϘlHok��G��s��S�������%�Y&�N�&�Ә�RX�l���'�;ǵ2�W���j���
�6]% ���媈��-ܝ���ko�#ET![���˥�P�<?�'0��@˫�$쵟#�����7���t����D�Ir�ŝ�œ�~SV''m@�������B��L�	lf&	d:����7��z�@���"���]٢tWFub�ߢ�OV�r��3]yH"̧�6���>���_�n�sOHV�Z�����A5��|�NG�0aI������\k��^����iڌ�������c�1��q9bY1�L%�����Y����w�=t�"���f᯿�NH�1�A�C�~��[�yTOn������%��$s���h��Qp��^꽚�!�W�1ŏ�b��{K�ܛu�N��J�c�$x��Z�Z�ez�#����7gN8�񪉇5�T��ai�U_��C����G1��_������e֦_��%��|@�ȦKN���{OF��+GX��~Eak7���J�L�i%�t�xD<���-���~;�����`l{��e���d�C&�%���1�\��7Gx<�_k�e4��%��Ϫ��1��ʅ�I���(�k�[h�&�EG�N@�]`���飗���3V�}Fu_�"��DP�?�cxs�6)���.�A���Q.^B��NT7}dK��"������ ����{U�$z5]-,�՟Og4>Q8)�0�
A�{I���9��R뜚��l�i�/����6�;<.�K��ǅc��Gu��Y��!�i0�^�/#!�<�dɐ�9��oQ����9��x�⾣����-A��e�t��F���� \M��*��?��$�\'��J؂��S^�QK��b3�l�O����ue(���qn-͞��Q^�F��w��`��U�q��/���2)��jj�1�cʿ��0�Vaʖ��苖�_�Dݣ�'���C�N����Qo�d�n��*H�#C�h
�];�u��/F���}N���r˓K���b$!�2�Ͻ_H(.���S�p��\]x��Pb�/��i/�!�.Yk,Eè�#g��'_�6x��-7p���8L�k�=�c|��ߐF��
�q�M���씧s�^�$�ؠ��������_ב+�r	�'��b{R//�M��<�Rˁ<K{���V�A��ޫ�ZU�塍����,��Rh��\�:�CT���Lç8+}��cw�;;<f�ߎ�s�I#П�F#Ҥg*�;��߲���CJ�����쒸o�v��u�CE���h���_�	��b��+j&��PH�l���$e����^d�}8��4���I��*�f�s�0���!��t���k
�3%"ד]�=��Q.]?���M����yY��Q������!��m�T�I�hAt�[�1n�k���æ�0�3��e���~��2G�����ԩ�'�4u+i��*,�bT��ukC�,���Q�H��x��rB����q��m[���#��m�,���w�ZY$i9����0o�Ai�"�{:+r�N�_�3*!ca""��`���S֘x]y��:-�$��v\�*�����$� �hnC��K���ݸ]�ںWwD�rOߴܾ^�m��n��B�� 	 g�~"董b"��L�KO��-ܩ��
����2LV�A�F��y���A�w�f�`Q��ҍ%�)�������f1s���:F/l>u^�h�)~�(2���#^!La$��Q|ؙ���cY�|���FT>�������B/��ތ<���IF�ۻX c���3��7�hw�@"��ю=�,�@�
=�J�5'�
�p�� 녃h��S�y��>냅'�8m}��U ��3?W0Ȇ�x
9�tb��yY�u�G�����Y�{�\.sa�~��#� "8fXcO��w�Z]���"y�M�W	\K2�bm�IЄRp�����/��B�ɸL�+�Gr�Aփ:�.�Ē�Z�e�8*��	�`�i������ O�$��)2aj5�Cyl�X�ܵ���J/J��y<͊0-l6�Z�}T��U,P����6�L�@���cw�)��'�Zn�����Ã���Ѓ�_wA�{.3S�JD�?���d�.�/¦�+<��|�SM�[n�p������4}�p#Ƈf��EL������7>�*�cB����0	YT��Fk��%1��Lo&��||"�K����#@������櫚��-X\�c�f䷌��Y�""_�+nI"=� U"�<��`m|2���:u�5w�q����u^|�E���S:�����ß�J��8X̲�����]1K�?��	\����,�������}S�k[=��U�9�">�1�s�J���F�!�}���T�K��#0�*%��8���zӭ}�pnrp�̄�nC�pQu��Xe��Tlbu?�ߝX����)�ȹQ'�M�gm���M4�ZQ��i�����#;��b���Fr��k������Ñu����/���0m:l�^Ʊ�Y�þq�Ӷ,��f�tD���\Q�.s����=ۃ��W�Y.���}�ͮ�J�8yQzp��2�X�;���u��d	�N漱f1�J�7���I��g)ԫ�g� }c�U5$X�ZB�h�y���a�O8O�~7�Uo���F�iЁ� ��-ĂY�E��N�}Nb�T$��'�J�&4�vB��6�L*8#*P���jZE�$��ۚ�����x�h����_IQw��<�At���6��~N('!/�l�]���|�F�IM�j@� �����,��H�w�\�FH~|iC��F�	�u���.|]J{��F��K��ޅ����J�0pv�>���]L�� vc����˕��ӗ�`u�;���`,�3����-�$Y��_��X�+�W:B'$�=A���z�a�:=Ӂ��%@3t����{!X���JT�edbsW��*Kt���K���q���"�D�f,9�KL�;��U�5
?���E'Ã3��V�1TN4U�u|��8|Γ���l�c�7wKo�IE�]�8�D��,��vd�e	sѻ���m���tA���^�Q��~w�����9��2ڕ��C�p5Ʀ#�/d�ҩ+���8\35G+�:H�:�
�U0$�\ADMO�sl���?s*.z�q �N!� ���K�`�Ao>�F߻u_Q��8HU�IK�Y�c�XN�P��}yc������D����?.�KIQ���ѽ��Y�4/C}@�.�aܾ�b�44�fG� �qð�x��(�ŀ�"�1!�:^@�B�T]�p�Ŏ(�MG��n�~~s��E��k( H;����B��~\�xX#H�kCz�R_����FD2�!���k�4Vs��Up5���z}��%Xu)�ZE��P�%��DɈ�Έo�"j���ΊP.nQ�x[a�]Ȼ%�3���E��N��K��xL�P��=a� Ȱ�{]MUρ��蘷͆�ಓ�f[zq�����O45��`�_\%�j�	�yP����m9Zó�ڵ��a�����5{�Ozl V'(��Q(���T���;\��y�β.�j����]��w����	�.΂��oaD9	(s�dY <�O�*�FX�h�銥zn$d����&V_�����L���4�7�+z���k�F@����C\F�Ɇ�e���L�x��3�b���c,��A�����Z~̵b��mW@D�����@������z�vg<��,>�%�C����q�j�5��[��r�B���iXSf(�$�:%��7��.����:� ~�m =#R�~���^_�cE[���Nv��*lF���
�����c贼+���
#ox�S�+7>���,-bQԱ]K�%��@��&�lԞ�Wf�,T�+�B�>�&�U։��d�(���$3KR�&����qk
��%6�2P�TW�Hlw]ܸŀ.|�2E`9�W��r��l¦�\t��[�V�uKPꐌ/U� 3:,:VV����b�#B�5Y�p�:t�'F���k܀��-z�'�*p�E~7:F�Al��{{���cq?,K�:�/Y��9�:q����2���ٌ�T�=�Q�m�c��Z�S�%D�q�#�����iY<^D�"���@��_Ɍ���rZ�G�{��;����I�30�7��vO����Ti�i�*3�]_(�����+cɉxS�5�K`k����$�C�h��"T<H)�?Ʀ`��hmU�k��_f)-��?f��������ʹy�! ?�X ���j��{;�
�W>��1�}��B��Uo(f�Ge�
��K�^tA�u�:���`�	�-�?�z��W�N�P^ɲ��vęs���@M�8���Hc�rN��T�l���>��+7
���Ǘ��]_�<�{��n� 2��i��#���P�k	T<�;�.I�i�)�il�ĭũ��1�l�����\op;�Uj({<�A�����ɪɐ<-��!�u1��,9�G���XY0�|�߆���\����+y��Ii�Ř�^�o0R��z�������Bkr���2�)m	�����|hn#���n�3y�/��C��q�2P�@�K�5���E<[�Z�F�[C1׺Ƙ1���;�h��A�a�U�e�>�5���kj!r��)��L��3k��/o��Ұ�����֟qr��a���
{�:�-V�Z�;��3�0E�т�U��Ӆ�Dh�ĵc�;5y7�����K���+c������A�"�{�a���NƜO�z�%��ꆱ�x�����N�}�^�)�S�@vWK#W�F�����/��G�.��k6����OL\�Od����p*�s�ɝ4��4�ssV�낏_	�6.D;9�QK��j���u�	�*���-�G_Jƨ��Ð�ޕm��;�#�裐D|��k`�� ����-D"sC/�V�C�|qN�p�e&���mF#Z4\�L3��:���[ 佸 |�l-y�tވ��=W� kµ\�)��o;1Fyۍv����xI'�n[\��n,�3��`#��v3��Lkӿe'X!{�@s�8��J�h2D\���EtQ���x}��3��5#�JU�y���ryu��o����]"�0�vES�0���U(�UA ��=�Ma9�\,c�z2ٛ��tdy�v�b�ӛR�K��ϒ�aZ�͵������Ms�'p9��V{
j"HQ�鱊�v���0�؟���P��4�N�fz������*U$켹f��.is��E����XJ�dqm?��w�IO)d�0LFz�2���.A�z���&�������{�9��f�k��T��[�޹*�*�Ӆr[5��
ĹN�?|�j���Κf��7/� �U�� G�= �N��+]o�b�e�0���V�Y��z����;�����`4]Ȍs�V�jX���^�"�z�Թ��-x��(y.�gb��qz�2�$Z���r+���d���D�&�|��a~ў�,�J�f~���l�=K�NY��[�+���Q��#=ѠS5�f�T��\�������<��4�O&���Gh7�-=�F��ϥ���Nuj�?��g��_��%+@j�<�bt�h��vքMT#�����!̠q4?�x>2��Pf�BRc��W�z��{����1\��8��z�z������b�`�H�:�V�0�����=��GRA�%��k͵�A\<�m�k����"Y%��
�O��u�"�{�%�58x��@BI�-�\P�	R���T��`H�h׵�)!�(.}���\WL�&UeK��Xn�xïr��R�{͇ M���[Y��z�(ި�Ic2LW�[����s�t����Sؔ4��3�	�\��t�R^���'��\���x ��V��2Xk���D�j����ɛ"��I4Vm� �k����WV'�M%��홚7l_t�W�.�|�7�D�fH���筀�24
U���L�T&�����N?���V��܋E�(J�yD���\�&Lh������>Q�.xwg��#ڋ�&�Ɇ����u�N�F������NH>VbVܽ1$)���o���]�ƻ�x�k��R����?q�7���c�dv9H8�D�J-:�4�.��V�1B��S���N>Ǝ-$�����[���.]Q\V̏��6$W��1OIDC^�����װ�b��aS~}2���<n�vy���@9�맱6���M�g�zE�|���s~=ۃr����o8�01�wێrnZF����h󇋓���M�2T��& ���>��>L�-
R.Z��d d���a�a�	7-K
�3�"�Y��Rj3J���(L��*����d��B 	����>��))>�A��f�f*~'��YП?�v_���gK�f�I��%V{�n�z|��I���e��g��1����{ ^��=�5�elh+A��T��bCCG�v���gi���֓t�?'l)O>p��� $�����1��R��_�.�+�~Ztj��j>y��u��gafS�[�aLX�Z�9�5�䞀@O�ʴ5��ƞ�s);�:�yʈT`҈�WF3������Qh8r��R�w�!?*�PG?�=���7]WC���3�4y���������]���XN�bg��T�q�q�ݟ���y5�e/���2ͅi��Q�A5,V�Af�k)�Ϻ�2R��2%ä<�7s�(X��I
>_i��(m ��&B��W;G~�Ē��j�i�"��L�	���p�IOU�j	�G3��z����һ����4'fށG�[5��dVMZ��f�a��� ��W���!�26�z|tq�㠧�B ����ZƂ[��B�m �����X��udR��#�?��z �~::��=�0��s$)�jT�E{�����3@,KC�܈���u���`K��V>��|<8�Z���|�A,b`cB&l�OX�=��JP)��˃Z��Ǫ؈�Ղ}gZ�ˤ��p"�:�S�Y�����;�L���&�]����N~�[=_�6��K�]6`U���,����`~}��SQ�q,��đ�:���R������Q�GA;�eyLm�|��B4��T1%��QTc�V(��I$hT��B!]����)'��'��'� �	n^R�e8�8�v,��M!��8Q�[��<���L�$�ZX[F� �����x*/(
�i*��]0��?D_�M'!,��!���&+�/�޷�W��b���ڐy��sNN�Q����W���DҢ����w��2��Mg�&j�H�fҧ�$��eE�Z?�Z�	�j�vE:��l^ �{+D�Xvk��s#�ԯ�YF�x�����cy<��~n���h�`��;2����&~�BC��F�uk٤!��|��U�p���]j����*�4�s]ޞ*�Q���Oǩ~����u�/�F��0��YU�nm^�
�͈i������b֥^�|�z�?f�s�"��&jK���.�ǔf_sol�z�eH%!��`�H}�������i����98���� �깥h��! ��8�C{.TB$k��ٮ��}wf�~q�x��#B5�}�k}pp?��Qԧd�Fܾc�{/ڥ;J���"D?oȆ��|��~P�9{�_��_��2�&�n3����a����KAc)���!��ñ�:�*|V�]D΍��*�Ea��t�6��['����aܸ�'I�<��r]���^�0yzI���Z��b; �E�*{{(6d$`5pX� �ܥ�$�/��ҬI;juj Z����m�M������EH����fVc��'��Wr!E5�|��C3*�JC(Z�� D��!�${T�\�v��>�:sFi���AD߲�D�W&t%Shw;ϊ��%�3� S�lY��&�����*R�wT �����l(��J�Txʾ����\q$jahȽm����h���>��,���;�;���[�u3)��n�Z�'NTe�7P<d��ztH�f ��Ȇ���ow�D�;@{��]���h��(�Ł��X�\����!Q����,:��G᤼���=����0R��{$��r���CܕCp�߉��$F�%XxL�X������,I����:�_
����ޝH���03�4�+O�?�:N����p>g�/0w����K?��k�Ly0��[vf���"L�R*N�ޔ�F����F�!��f��d� �pXH�+Z.$�W&�z(+��j��׈���[�6�1�"�L%*DrJ�����X`���H���O!���ԏ�:�������I	�j4w�\��>v��[,v5;��1s����'��F���Ԃ��2_�5m&��Sg�|��j�z_��s��[L=<,Z,�5��{G�$���~��ַ��$��2B�`�\�������v�V����o"���Q���k����7�
9�w�nҥ©a.j�sO��__��w咇G@]6_�C8R���%�ME��3�#�y�Y�k؃��跍�)����iF��o��.+.�Cw�,F�Mɺ������u�lܿw��!�^�E�ʿ�1-*#W�j(b��3˩���&�Qz$��e�p? ָ����w�A�w���]�^���M��
>d��wŨ]?��Sl��p%�����\������Rn���z��zrj�~�O��il�לH+���>v�����֐_S#٩��z��y=��ד�9�PO��Q������u�	Ƽ�7�𲖕K7�R=�>��1$D�3y�X�(~N0�	;y��jԕ�~MDФ;�ַU��U(w?��������^�xw�����8=��.;��Ǥ2b�	��i�����$\��!0{Amd΁�qtCˀb�
o4��v]���(
�cy�GQ���0���8I�3ˡ^M�LΊk��N������}�D_y�>��g]�Sv��p��5I�Is�~�Ϙ,\�D�*��ۄ9��
�����62jo*�i8���I �_E�y�v��vfz� �q�X4�c�?�;m���6����!�ZK\�L�C%#\-�����i�سYO`�@�r���ޚ�L~��+䒪
X.=r�L�� �R��v��N��f�T�k ��-�:�������^U��*y��~�]u!�Y��K�#�Q�\y�Q��&B����,%�@�����������;�B1G�RI�ɍ/�^J]x��J �H�Re��+�C��o��#���#nCu)�T�,�=��8��-~HAO�\_Or���r�� ;@4׋�� }�h�x�����+J:`K t�r
����y��	=�6���c���>�D/��Q�k���*M/�-�ړ3�& �?[=�O�TWS��i�!�S��א��c�W�7?ϒ��-Rg��b�r|2AM���Q}�5�t�M���`�xa�~��އnv��t?6l;��v�=��Fk�����'*�����p��C+�=Lݠ+�	،gIh���Aӎq��� 9/m����İ �i�Ǘ��r�Y��V���ы��<6D"�1��%5,Z�`��m���n7��~w����奻����ӗ}��!�AO���4_rZb�=�\��[��Vg8��酺A�����{/�I�K�=L>�c��%��D$���QuC��Q��޻ݪ]w�~j֛\?�ă�E�4�|�e��Men��W�װ���L:����+�x؎�q읭� 	fi� �nf*�Y#��T�>v�6��� �U�8s �����LA��o��������
���T=E˸�#ld��g�+l1� ���͑K�10���������EZ��6�
�7�`@��v;�J�Xw�7�uGl���s��6��e��rК���w��Ď�8���1�;��e����\�7� s�&w��U=����4��|��� ���R��g����(-y�[4���v�w��Vp^��E�v�qFA���H�WO�˭�oI��٣��/�5����4h��!bE%�	�Z���VC�W�P�� �|7
H�Q8�` ������k�UB4hm���!��Hp�:�w� "�&;IW�ơ��㙣�X��e�CV�Al�˔`T6"�k9� X�����Lṿ�喬����i_<,���RzW��Q�f���y�{�PX�5~��W��x�<����� �8=�<G�D��5�.�Y�^|=φ⣸�A�k���L�B�]�Zh#g̥Q�o
S[�q��Q�u�;E-ĩ��ނ���I�����PuUp���/)��j�w����7�f�����L���z"�(@�:&���z��3`T]с�%�R�^g ���Z��i1X�{d�q3��H8F�	녿-���2^VMRǬYN}�{JGS-\i��솫�<K�P +3Ϙ����
x��n����������bο>��X{���n��/�k����B�i>���#��"m��*�&���*!F�8t��QK�AaVճ勦ts���:�Q]�?)-4ZnX�CkrX��V����H1�C�ܖ�y�{'x7�rPX�k}u��<���p��0A��ٜS�|���D��7�[a;,5�u��f�\��ޮ����ҦK��B�R���i��!���H^{ч����m	ٿ�^R��Q� i�����F��6�Q�x��d��u<�V�V74��:B����,���o�!E-|�*��L��!��o���T�5Z�a^$DS�Ͳ��g���?NR�fQj^5�N�q�Gh5��/6��Ro���bo����Ͼ0�Ua�@�F�q=L;M�؇�������Շ��E)��-]j�@���Cf���b*r.�b�l�(���RlF�B��qA��ſ���/x8!��;Ȩ>\�T�d�|�zG{�'����ޓ��-���~���gO�:�9�b����D4�*L�En�;:u%�b�M�rZK7�v��[?#=[_�>��*#5���X0al��;"R:uh�'�>k����HYvd�FR0m�彗�;f�e��W�������ӤC5�j�U�U>��Ut�ت�`��~aoÜ�V���t�)5۞�3&R�k���?��eo�AD���X�o8JX��
��� ����0�Xd U��!�1���QO�@[�:�g�`��G���m�ˀ�@��̶��D!i�2`"���p��]"M2��"&��0O`�H�3��W�n!�tn��X��nO�Fe6�XX#�J�ã�������4q�*��� ��*�H���5w7>["�#s9ܦ[�­�$6�����9$T��w:`*��c�^Z��Z�5��������#��ݞI����i3�[Vv��S��`(�ϝ ?���&b5�w���{'��$�
�(-���	%B_K���5\�e�Aק
^�7���t��@��(�?59��1�')��찯87c#�X���V��b��QE��9���&�4%��<e�wú;3w>��O�e/��#B��D�̽g���Uq��T�p��uS/��!��h�W�֟әާL����?�J쀦��!��8�&ؐwR�˪��X�%�w�,4'y5_�A������;�l�B��g�+u@oz�:�|�=U��N(TDMB|�r�Y�$A=d&f9Yf==K<�v�U��L�N�e��g��E��VV�b#�v�"j���e���6]�4�a���m����&�7a��v��p^
'�lo�I�Z�,�o�s�ԋF�=9����t�6��'�����I��=\��kौ�F�͗��.�
#�$j�-F�B���pNI@s�F���:>�?ؖ�5�����﹩Ӭܗ��Wި�h�v�F��5�9 Ld����G/mY_��(�g��N,�i��c)^�M��h�x3l����M煨�?�k��W�%�,�wTS�1\�p�����O6<����|�y�pBAz��==�o����]�
��]��*`�Հ�F���TU�?L{��_�X�{��8��@��O�_�������\&����y�!o���,�q�ː)��X�jO�Am~a�!�F�DGL�eˈ�b�?m���۲���6V�i�}?�h�GL�+������i�@
]:
N�;��i��Kk�t����F|k�����LۡD�/���j������m�߈�_3sq��>��(f���D�cr�0��Q�9��A�b�X�UA }q�(�|�<���<���Z�g�m���¨�z5�n����Yg�>�䢋F��[�6�25Nٝ�J��M
8��䖶��G�_.�x�$� ����[��2ӂq�