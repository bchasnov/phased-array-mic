��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\����q�?��e�I8�b�Ǽ$��"����ׯ1�V0���ϱ ���u��fi�I� �o���kwk[;�3��l�z��}WԌ���������Vp=~�.|d�h�ύ�i��b%[��l/6�@m�(�}l^���LkA�$�(��-K�@J(HɃ�.4��,UN\��Lnm�/�r�9l=!ߘ�+���[V�)��j� >A tc��V"�4&sf�z
��a��Wz�^3FgL�w�Pb�-,C��צDR"��~x%]���D�Z��i�~6�҄�QH��! '�-��T�gt��.$a�Zp7)➹�W�F�뷅B֝D{��^�9<AdNW�:p�o�A�;���X�5V�<4J�ű��������Nտ	�T���Bb�d�i�p��SZg�i�J�����Lq�q��"�n��+��p��z�!��K ���@�� ��X��� T�M�8�i��lة�GP	����?�QEGn��
W���/�wCmyR.n����#3 o`vⱅ��\x�O�����tHCȱΌ��ȸ�S�����L�Nǉ�5xl`��
ұr�a�s�$�'�m �{�X��{�0�%;��eR?�;�Gj�(�
'p�܌ǅ��1��ȥ+�VШz
/eڟ�z���<`��	r
�U�Ը;��c��f.�ܱ�c5�bg?7="Vcp�I0�5�2)MW�ا�feA��h�����#��L�C�Q!*��6��N�N�B��|���c����o���W��?���Ҫ�mtZ��2!�Ģ�p��6*�&�B�P�R�k@x3Ib2L��L/�iI�/R��N"��ug���̿
	�]��A��q��ß<ή˦n+��pg��؍` %���dtR�G�,т���+J�p�=��O1�-ݙ��p:���gH��Nf�/(�k��v�Y\�D{����a��L�O0>������INj4�W��T�P�c	���_�O����\��i	�FF��od��5=��7��8a�j��Ɲ��SL"��h��r)65��|ɥ3�h���1�-���JY�B��c�K*��I�dOu5�F�|$m(n�gH�}���Ι�"�l��?>�[_W�I�D��HҀ����>P��sd�k���"vp��{?���E�	�d0F�	Gt�Āf�'>%����i9��` y�w�戴�y�#M�8�`�hv��(�R��o����I#vp
B���4�^���A�fU0�vU�Բ6��/|f��ƒx���u��)F9���*�N��kM��l�r����h�)� k�a,�A������o]�g5�m�0'���Py2p9�ىh���x:l7���l|4���as���8��d�}C�Z\�b��2Y6��צ�At��j:!���>J�8� �b�bm*
��wh0W��Mm������=9�q�9H�\�'C�˲�T�k`�	��[e���͠*��X*~�.��f]�x�T�*`-kz-hč�F�6�~;F�]���AK���I���Dmp������IY����O�)�ܒ��Eŵ�i�逧-���چ��bCnE���I=���������0�!\��_ީu?y3@6�ފ����/�=%�-A�H��Ҟ�,D�����78Os�µ��ȸ�L
:tR�cLFLF�:�b>m(L��c��=lsw������Dj��V��Z����TZ:���w�`򼌝vxL�� _a3���˓�Xx�&z���~3�R8���~�?�E���k����p|mK��� �2Y�[��p��\��Z��f�{�d/�I'��\�u���3����3�2Z����-�r���H�Qpuy,���U�b"��C�u���R��D�%\O8�~���8RM=�Q�"=Ǻ�4������L���>\_I c�&�^��@a�g�v��$?�5"p|,n=F�& ��ߧ�1S%�Ez��zб�%�s�/��wᡳ@����F1�P 1��*��zS�Jފ�`X���!LԫR�w���?�

!n�{�ö=��;o���&��Ԩ�(9\�,���֊��gfH2V�����!KTj�m\\�͟y��W\�,f�jT�B���_���EWE���M E�8IH�J��Ec��$���H����""�z�D�H�!˺��?`yB��$k�?�?�v���|[�.ZW?71�T,��`���/L���f^p�H4���Jay�:�b8�=����D~�9E����͌PnL�`�1��x��g�N�x����3�N+�v��u�?��Ea��Z�<�����%�I�f�����e2���D�|/���	�Lb������ NGj��#y�/�!��M�EA��X�b�g�q�W>"� �$�.��}%��Eݘ&V�r�Q���MC�%U2�����*LI���u 1��QV�"���e��!Sy�dp��;��U���G*VJ�S����h�7?�F��ő|C2��
�KlՉ�1��f�0.|������a|p���{u�vXo&?�Q5�(�Z
�RV�t��"_�f�ח:�H�>��F��S��r'T�}4lp�?�/��v^ܗO ���l2a�g��©cyQ�4Lǔ*������TiYxV���D��`']��"��ӎ3�"w+�׺����§�{��V4']= R?�)��1Q�?��f�aW��4
����\�^�6p���]�!�G����2:�xm�����/�KU���{B7���Y�7
�f���$&������u�/�xѽ����83p<��n��×�D�B�Zs�O)3���L�Y�����/d�9��8�x?�I3A�MB-EY���Z��(rdl���e�����h��P� zHva6H93ƪ-=�1���8~���^q��j�$����^-�ҁ:����Z�u�N[2�im���R\�ir9v;���� t�y9����.z�����:7���)%7~��=�㇓� ��֟�]VM˧�H�X&�5M���;5��Q��1a�1`�l���򡹦���K�t�/*)��A�Ê>��R8��"�a�k�Ƙ4Y�ˋ��$S����V��� ׇ�=V�F[1���B
�k�>�K1��GKA�4"�Ɛ��؛Ѷ=�Ep����l�A�m�3-i��w1aq�p���ڻJ��˜Abjfh!�V���׮�Մ�,���L��|�bB�V9��(��<M`�2�iM�^���=��&�
sk�)�do���~�7jm�ra=��V{�����X�{��<�t]��{&��EFOS퍨��[2g���yK�j�5#��&�%�ŵ��=��2.����s0����8l���������{��T��b�jQM����O�B^[7Uo*��P`���	!vI�A@)�"�ؚK���~f�9�b�R��JWh��Z)ʢ5� ���?��R]��e�]��  �LR���[+�y<�V��f����2ֳ��I��ʒ#;Am��2ƙ�+v͙��z�Z�@Sb$�-m�P��a1 F�"�y��z�+����r�2{=-�,����|me�@���t*_0w�RP4�E��	̸�"�nd�؂O�"�Q-���:!��ۗ(W]��7BmZ���eRlS�K�J�I$���b ���Na����^���( 2��w����O��q ��u��Mo�;��@Ճ����I'��<��L[:�5^暷�yb�c��!̕/��]g�]�2V0���� �����I{~�)�VjKYM�ƾ��^N��f��ȳ�i�@���7j���?�����T��s������3����x�U�~(��m���5(��a%�h��<t�J�Zwg��3���${C����1�q�0e��K��5U��JGEk��e?�ԑ��
����3fH�&��)�){��êL���0�n��w�'5���U�?+z�e�#ۭ[dJh \z.�;�n�)!#�Z�sn!��l�!��%��\H�����I�.߅Gl�pG����a�qbnyc|1`����>���,�8�ZW��� �DQ� ���w� 
޻��U����1;)�|$L��XS2-�\�dq>�_.���ej(8V�A��Z�k��8 ����o�d���?=Pe�c}RMhf~������.8�di��䰊-xP��#]�X�8�|�\��V�B �K[9[�ݞC�7#3�JR����36�Jk� �I#�b���q�>.Q����=[�3�_���		��u�4}	D� �ɱ�y`N<����2�Z�m�9����~��@�� ̠����%���4A^[��!�����4��)�RF����JpQ[IB^9����7�g�3?�9gհ��x��"A�9.�"I���R&�C�7׬(��a�:5m3|C������D�˰h�@���� {�� I�H��A��*��9)	�i�|t��8���1r��F�d���=�)��cw6���B��!!G�E�C�gŹh��͉$yO1��L�dg��RIV_8{oG��w�x<S��M��J݀Ji��[K�����m �3$S@P�kwRHJNfAI+ᡄ+��<M�RG�?�ۙ��B��47Sc!S[(3c�̣J�TCRlӝ�5��]S����{40$��5���C�I���2��GΑG�#�,�d&.��<(�k�꾙�E�	�)�Ca�@��F}�IQLmn��J�(�6���Z��z�9;y��d׵�)���I�ݳ�*���{'��M���Fh��g~p#<�1D"a@�Z/����Ex��]��P���(#�!��]��T]q�� �W,���4��k�3�n��(9�K���	U&*�֙��:5��;�j�H؍hKOg�R]2�[.yn��\g�DѺ������nJ���Ǳ�G5�!���&p���58O��?����8�V�5�	��۶%S�;���ƕ�)� -�$��=�j�\Y�{�EY� !ܪ�4�5m�S�-\̞`�.����Y�W-$��z��
�����8���T�1�#����L�5<�_���Ec�H>p(C0߳��ܩ�f:�E������(�	Lv�C4D�~.��z�W_��iG�D��M���B�MD����B^��6���G��+PJ61�v?��wj�\�X��C�?>m6��~���',�L���ظ� H}}�L�:V^AT�l�������� ��v�e2=�Rٚl�Om΁#��ƻ"��ȥ�C��4�9�Uc���Q�~ٕ�d��ф Y�$Z��葆�VFX�?�c)��x����H S�>PƓ�o��|[o����R��~��~L\�������o�;��/bա��n��m��k��7�����{r⠭`%����Mb�.����%�?t�ā�&t���.?��S;��
�e�bt�']���y�uA���@�K)����i��=���e/�x�,v���k7��H����i������5n(���?�`>�f57<]�$����v���i��(�<�3���?Ƅ���o>�s3�A��5@�-����������̮�C����gi��s�\�k�E��fب��硵� [ht������G"���M�qGx˄��빵�U���/ ��ĩ�����
��vS�y��]��6w)}x���|��gI���'@Zu3j�
���H��j�X��)ˡ��:���oW@��mEM����NU�[vo$>:%V�bi�W��|0Ie-�t]X��*�r��4��`�F'����[g��ko'u}����ߏW�>/�����N�)f?Ɩ��V�o��U%^��P����HD�JjCP�y�%��Lc>q1��}N(��3 �U$S�To�}+��7)�!8���6;M����v��&�%�Ь�$AʳhioGM���loZ*@����M39�[�|$A�jގ�=�7D�z%�9�t���W�t�H�"�_��V,Y��T�w��dZ~υ��zH]�L�u���:ho��m�����b�M�5������4Ӈ!{�H0�[L8�����3Бv-=V�G]���%�E\�E�-�0X�,b���m<tR}r3��~�ƴ'��N�����Ӑ���:q/1x�+����7,�}P�`�LW�r,����At@��P���Y�ܟ�4+��:9�9�������c��1ѓ���0�qb2��%5,�E~m�7]؄:����*usı��h�$���\l#j�;f.r�r�6o�+J��Is��� �\�(?w��:Φ�����4�/}�Όg ��zА]�d�q��`z�y��2��ħ�@	�07^���ϳ�	����|����K�Ϊ�'��We��"?y��=�-���P�av(ec��6y�AԔ5�s���A1���
߀�^�3�vF刲�[�؄���@��N�����RÊ��8��P���n�:(j{��%���2%x�s���Rk1��V��Y(h���pK(Z�q>Y�P��d��U�]&��]�4�I"�ۄ~uI���[����GS\�}v�F�������3#��o�9O�z��	ܿ�qק�Ǘ�c������q�l�Q��[��qX���j�;$I磧���K�ʜnlC�l�^ywc_ޑ``#]Y"�$߰(������	;�l� 	�|�b�C��	a;L��T���l0���hb���X�:�EZ`'���Ds2Y��ؤ�1���HFL��h���i�E�e����
E���~F�Xq��<���O��d�������7в y2_�=�R%d�ez.��q
��� ɠ	�\����q]\Q@d��Ms?���REW�M�JX>�_��Z)�KXdˆWU��,��L��Y7!���O��D�!2�#^��^�O���̊]�c%��y5���Z����G��0��Ves�@��:Z�ԄL�h�d��b�4�B���})HT����ô��J�������g,��Ἐf�v���"�ݭO�
�叉��o��)���;	lk8$&�[ �1�㈮|����P��S�%m��T`��t�t�O��x�M��9����C�4SVK7�������Kڹ�	�����6���ZN���<S+B��{�Q#�]�B3yC=Ӿ_}[`���j�a^��7�6s�tF?�d����q���Iջ�ٶ9���/��& �!(��T��1Fjً�48��]nm�"2�����ڃ$�4�];��}�j#s޸w��0��ݟ�T�M�(�,2�_����i��{�tZ��������|��N�����ٴ�]�ʴ�uD#� ���N�:M��-P%�Dki0I��WI:��9-��[��	`M��',�y~X��ߘLAO5�ɩ��|��T�N[�� u���)C$��'��%��B�aR�6|Lܳf����#�vb1/$z�_��Y��L�b��x�Td�!��o�� Q�q�L��KG	�͡6��E|���ߓA���8�f��[��-��Fy��wh����Dx��gՎ�'��+�H���l蓝{��T/������ �.je-�*q�0�9�S]A_riWGi,EI߰s�>R�dW����`3���%u���ؑoq��XC$��]_E���ɋ����9���U-1z݇i�}��a�Zҿ7<5B��F�$�Vm�`Z��(J�,:Y�O�\]!,~Dnɑn�.$#�J�L�|�6w���'dD��n����E+Xj�*]�-�Z�Ɗ���ܑ���,|�����x{ ���x�����ܑc�}���u�?�x��-9Pk�]������A@B���>Ģ�>+n�(dm����������_\��n�i[0�˞�N4S��im��/�'�M��. RP9p0)�$z���H2�{8.w�c/.��sG���6�h "ܗN��3l������ǦD�-yz���B�c�=�����orv�o����inT�#�_��L�.�RS`mQ�����a�%���m�tH��F��\�ؘdZ,�	��^9���@�z��8q{��*\�}� ��3�r#+��,��� SD[$h;��>}Ln>h������:�À�.�^�+G=%��+b�o�.տ��e\��Wl�N8H��Tk�Xz��)�c�ħ�1ݽ��O����VC-Oۑn�7k�]��`N�u������^uy�/*��3�������T*��SGt���pl���V�����'���X�G�Wv��N%;�|l���2GU�\����#�����K��F�p�+6����|$�f�y)�7*M�M>:˓�O�����8!@ڡj'&�\B�t��/�һh�~sQGƷ�4������{���.���.�.�e��\��=,X'_OI����KA?��,����Z�
�V]���~qE�`s��*2�t���k�d��?:�"K�����潕bS��+fw � �����	���>�[/XeC[@��?D�H��S�[�V�4�`���t߆n�č� ]==���t����E�N��{�u��������n�b���,�m��#z�}.�b%�%ܟ���D�ω��p���eu[��[�F�<�B*e���z�e�{�
k�rZ*�W�,�	.yA�����,��#8�5ug�Xk��;��O����H@trC�ι&����ݢ;��KC3HK�Ȁ4?I����0~4i���@/̅���!�.�i���PW�}g!'�<i�P�fht:jC�X��)X�''��?JE�̑a�����&� m�=�M���@��o�uLR3����b3�fh�c[<6Kx|��2�oe�6d���u��ӐA�q��ryC��x�mA��e}�O�c�T1z7�<X:����2Ru�Ŝk⸣ZH>E��'��R:�Z���1w 'i�2"��	��]��S��G������/����׳`���u~IK��d�'��#]��s ͞��-�����P��{x�r��>Z�57���������I��P�w�v}�<���̨�x�L(�N�}G�[���23�>��$t���ߠ���a&~����{�*g5s���V���ؙטcտ:ωr<#8F�5���w�m�u&R���%��co�n�c�[[��&��I�Z�t��=�U_gY:�GYV&����L �����t�� �}�@�ƿd�bQ8��?f�0 �8R�&� �V>	�r�혒!��f�}K0���	�?�3j$S�/Q "���Y�9�-���xg&��*���;�#r���z�Oڂ�T�3ƥF�PÍ'�l`>�o��)D(23�7cmQ�}(�f�OPx/FUF�;Q���9�NNމ���%P���l�2�0>ex.j��ِ-��*y"�����A*����8����<��z�с`$_;�'L�.(���A� ��Y�@ )���e�{Q��I&)	@�ZJq|V�c���cg��b^���P�Fcxj��|�DJƂ{�D��*�f�q����Qv��L����Ϣ����S5 ��eF=mԛÏ��7�y�����`���:'��m��ǽ�f"�ʕ�(RP���m6ΗM��&���:z&g�"v�34U�n���sfl��$幼q�}y�^�
������r�J�Gw �\�B����Q�8��\�l�����:�������t���UA�Նs�?x�Cc�U�؂�k�l��af�ohS�8��1IE%��d�̉1�΅]h��O"$N\0Wms���v`��O`:T)і,�X)��ԕңc������õ��/X������8�s�"
QR���ɭ��r�-���5��q��ɷ��
�>�&�V6�ƀrY��;��~���P�*`�3��۪�')/�x�^���o�	�x�X$/	���h]DT�B��L~5��[��߿y��S�~���D
�j����|VX�9d2���Xv���4�X��[-+T�x�}��_�;��	��p��OPx�:B���{}h�+�[3nZ����]Ҡ9?6��g#�S�7Fɟ;ǩ>�O�bJ�8�-ťx���m��I�Z��leඨ��qG�]U��L�ҍ�w�-�sS��,��K��=?<8��A�]��-Ic�U��4�����er�-��pl��% I�eiw#� �C�i�L��H}/�B���i��GSdy:�ow�l�S�YĐN��w��/�G�X�/��t�`Pgq+���$u&�x��Jɗ�=G�!���N�>d����ӄ�=`H��*ϻ��������#������W�R	��VhE�(R�w��@��Z�*�Л�5v�ɗ�%V