��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\����q�?��e�I8�b�Ǽ$��"����ׯ1�V0���wR<�o�Ȏ���U5�:W����td,�&]"�,���;T��Q�^��	��ܶʰ^�6�]f���\���v���/1�NIZ��P�k(ET��
$;��(^g.�� )#ٛuK���e�ZT���7(�V8�b�,���O��H���e�2�Ϣ4�ob���(��Jnt��<�-�	��r?;��;.���99�gdw$i'c��MC(�GL���`�C_�&3v�v2�������`&��	��K�����$�n]���$ұ2'���{K��0�􆽂����w{�DG<��.Y�j^���"bٙm.J��G�È��=��0�R@F�|�ip�F���0>����7���i�N,�v�鹹�`VAnb��sx(�c b���%#ipm�S�l�#䚥��R�q���>��5bY�zN�H��e���/�}A��[��#\���(��R�OY��x2�����l6%R�,���i�.�jV�W'a����"Ҫ��MU"�Ԭn1d��c$%u?p��\�Vh+���&�c����t�z�A-�����{'��	`CUӪ���MoXR�Ǯ����(Q��0��ͭ=ZWSu&���c��càv��#T#"�*1�׭�����/��f��&X�</�r�l7��h��A�����[b3���pfz%��<x6���6[�d����Et��8mgAR]�A�2&��GE�P��ü�L$*]�~����8ǭ�_H���qA�Һ��d#�///!���9��Vj��M���#�s�/�����w;n��zq�؁����vH5�+�hvf���a��=Q�F����a�]Ɗ�F�S~�`�B�Bͽ�MP��4��<Ւ��#�H�MO�6ԓV���P�b�_��Hc�@v,0��1��;]�8��}pA�7Ѧ=ck.
|���9�ɷ��]U^���D4�s�@ā����
h����j漂mZ�����������1��F0i�Y���B��lW��%�� nBXK��e��``���z\5(��k[�᫆`�fvշW[���s����M1&��޳\���X,V�� ]˾3U�Q�@�j�X�Q�5{����a��ӽ46_��7p��el΁y<qM�U�W<�ݒ���n2(�������&��ݦ�X�)��Ђ�ԙ�'#D�(��M"����ت�%��({5�b �d��S̭�"y�����R(I~˰�9�#1��l؄���AQD.�w��d���?�Z��D��~��*H	�KQ���}r�\Ri��	9t߃Ge�O���ɸ1��#��Ί�
$���&��$Y5��va`�M$#(��D0F<�,vY�֍��
v�d����ʱ��<+H6�(��>D.�͌�κ��\t㢵�O>[�m+1筙q:X_f���{�����Յ�k_hfdR���^<~���K�?����b�kK���D{R����#Ǎ�&��%q�v���j@�9�����?��Ia��l=@�*������C=�*���=8�ȥ��(w�8�s䳳��Zۇ����~L����Z�|	Ry~�����p"�z
��
1q�� Ԑk9u�a-���i��ҲjH��.�t�q�0��lGI|i��^��#n�C�-yH�1�mw�;,	�J��%:�-!�H`�hu��E���C���c�!ϙU&�DHF]�ދ0z�0���K���"�I��vh������Y#�Vb���S�H$�<��{c>���V�B��V5HJ��R7�]Xh3��Ku��<����-�Z��g��Ǡ��i>���VRg���۠[`4y珄�n��B�:��Q,����)�U^���e�&:��u\�*J��
a���*��~J���e�F�K1��|�_�\hU�l��s� ��&��!)�Ի�2w7TQ"lp ��hw���6����PgeyA�{5��y��w�:ń�;�r�y�V�x!�f�:a���Uk����� *�*�Idd�,H��+ݟ�B:ԦYy\Ju�IKZ^��`&.h�� =�85%ڌ�0�a��>H\���-z���S��u�9(:�ɲ�)XE�H�b�`��MY�xY�V�0I�a����Xa9�J�+[q�g�[p��&%"^�E ����ʩ�9���G�������k�Ds�V��1
�sv�8�]ĪꔃY#-`�%��S4�"��uJ�&�A�E�T�3��M��i�G���<�."X�;c�h��XR��'�T��l�����P|�y�?'���K'�z;@�����ܐR�H����o���4�����&ҳDE���-��Z���=�W*e�V`�Z�^���/R�`��)�q\���P�������I#l���˵��;��r�>4T��9��A����s��@���5�LC��5��,h;@p����c0�X]9R�chb7���c�H����a#�O,4\�n���tT�p�U�n�ͅ���+�P��(GKȷ){�)����:=L�z��]?5m�Rp���D���e.�	,5��bj5S����Ѓ8e�>���y��W�5�Ȕ�v�ltMT��l�ɞ9 ���sW�.���1�?��]],,����������[�U=T��2�����"���T����qS:�鐱ksTʞ����3��&��g����N�aZ-]N���fAs�7%�N���E����q)����Ki�݄����N�7[�[���A�*�+inz2!�Jnh2F[t��D�2zFQ'����g@F8�Cv�L��T�e����%ϯ1I�r�Ǻ/��s����L���HA��gg�<�ki�{/-ʝiBP����\<79ڻ>�оu`_�����{Px=�R86�赱��ݛdRg(@ɈJu]�h�%�-4�8�����I��}�Z
��!o����U�Z6(�R��w�A�셺��;�TzZ��e=�ʣj͐8-aEH������"V�⽀�?�,
ɲ�:t��^���h2���<ܪB�j�e_�8�����x���� �R�)M-�	��d����Ӡ��0�t<;z���S&mh�I�s�}�)ˉ.��j:V���<�PD
�����:�戉U�ΤU�mM�i�O�U�$f�A�D�{�= D$�LY�BS�c�:d���Us���n���S�@BY��k��6E�8��Ub����H2����*�8�L�΍A��hZb��U�ʂ��E�&?��YSG@I�۽s���:R&~�ߨ �w_�t�9��EMvA�hK�l��:n�~�ts���!+�v�W����A�.����� n#"��X8���2>xk0&8�IM��=�����?�G���`F��M��DW]'���QѴ~]����Q���L��}qfjy�R�f'z��P�a(	[��k����YSk}F�����|R������޿���w��&5��U��X4�3H �F�8���dd��W�����d6	���Cf@�zЉ�SQ����3��B�->_�c��f"��mډШ���#8��#���ĸB�h�߭c�u'��3֙\�MB�R����`���G�SG�l��y������ �v�����A�q<������Š{��.za�i��1��z<��2(2k��8����#u6����@�K�S��$��#��&q���J
��u��[٥�c��A�Lg\����Q�&r���iS�,JZ��Ya����i���u����H}�&���\�̙��K�+P�~t�4���L���OCF����c'LX�)'�|�0Q6�Ɠ.���h��6�_���L��Q�h�����,!��flsJ��ԲI�,+�����b�c����h�́O�S	+��!쀒�l�O���d�,������=o��+�"D%�S��'�ɦ9�d�in��2a��0��}��6"����.�^�*�� ���!;���6�=N7�\��@�{W�/��N1�H~(�w��S���F�(��y���0v({�eXݷéb�
(D%����e�yG�������S�)��U��!~����e�\Fe�]	��M|��U��sO���$�U��C��F�
s�.�1�v���Er�o�
Y��=I����+��,r]4�m�?�_gTLn������l� �X�"1+`;�Ӊ��n�po��G8/����ME�,YrY�l|vq@R��7H��X�Z͆k*Z}.��~f�4z4ݧA�nev�Y
�r�����țĒ��k�ë��"�	�	7m&}.��`1
�(�t��*B,D������O^$�Ӳ�N"�ўB-Oކ } ���I�7�x\;�����u�n�j�WX[�-̖��f�'=W-\���T��!#AIB��y�X���߈�Ǔ��*L�'&V�,��ч!�P��x�|(�ڻ�hF�?]�G��� ����w�j�<rl��d���'O9 e��8�R�����mB��e��L#厨�mO�y�Կ^�������C��/�q��h��7mڲ\�����-�s�X��#Ώu�gx(Q�}C�<��^��"cp5R����緓q�':���v��
����3^d����]��������v$�ѫ��⸼o�,���o��jD�3����F1QGx�cO�w����i���C�O�3��h�=D��fh0���O�������8t0�6B0�:?t4�L��`�i��q3bAkb[�W�%�Ӄ������k*i������x�Tq��.|�
�Hr���x�Ԝ:��b�{a˭��E�B<AP��f���a���Z����Uùړ{Ӛḫq���=�}.r]�utY�3Ł3����.���������"�P�53^w�����&A+��Y�����6�rk�20�t��nѧ�v7R�Qz�r�Z�ּ�YN(�����U�ԞCI7__E��k.L�q�l�`�[��?�lb9������|\m�p@	U���H�y{���TE������̴��� )��L��To�͹n��7@NA_:�\&��;��x�1��ڗ8�ǉ�G��;Pg&L�<9mϚ�\��_	[H��K��6u�g�xE�i���E*2�AGj5|���5L��hh�1f��A<�$Y�T�G�;��ׇ��{`�^�0`������8�B
s8����Qo���3W�}SP�i&-����B4p8�� sqg��'˂H_���V�lƦ�Obիs���e���h��~ArM�����e���q��=�ੰ�w�`���-$�.��t����8�3�A�..S�$$Â����WG��fb�o}W��
Bx�:zb6̡�5',1'vU��>`a���:Deo@�ί(KL>�.��&;;,��h3�@q� x
���yX!����M���AE�}�[����r�^�Z�_9IPL�P#��3�I5Ĥ�
�����y��&��ۮ��۝=Ɲ�7qt4]w�e�0��by��Ѱf] �:0N���!��;Ac�f�1<h�B����z�#B�.P�<��q�@n65�Th�z�G&�NL�&�/��Y��4��z��T�.N�+��C�X�7�i-\_y����	v�6uJ��QFWI�۰0�|f������C�+���V,�7ivo
��)Xq#2Ԗ������q+�dU0�>R���Dэ�v��6���^A�භ�j��eZ
_�ùA��Vڏo(�K��4c3e(�Dg��=�	ǯZ��:p�X���=��NV4%���KcaZ�Q�A&�=1�e��ǿ�~�_�M#�~#@���X�{%�u���V����x�{��jVb�����L����̰Wnq[��C��h$Ig�\�a� ����vЀ��ށxA�bUf��~-��>1����=*�eʆ,�(Y��2b"�bm��FcZpx��D  ʝ�	���e��S��+�tN%l�HT��(�̃砥O�Wf��^�1T���La������]��tf^z)jP�C��+}T}{�ic��~u��ײ��݂���4������Ut���Ѹ���M��������h_����k�NBF��(a�$|�����5��A����!�F�ݠ�L�6p��g蘛�BZ�#�2浶�`���$_bu�yV3��`C�ʧ)3��&�)��%���Ù�Lf�r�n��+im5��@�Е;��ךΉ0Q!�2�K�K�8�V���E\�@���47��K68�?0%� I��'[S2+(P�
�%;�f>��1�%�K�VG)�wK��E��	��6ɑ��ۡv���վ8T����!iZQ�)�������^e�!@��V�Wp�8r�(@�
k�dE�(U��Lm��L ��<��Q�kb�h�\Yy�����q�}.��I^v��R�7V�dޤh�־A�!����ϑ�<K!^���Nz�}��2�`����W�	�Fx�ˬ��>V���A��<	���Q�g��L!ϊN`�ZAp|��җ��I�VY5؟�T����~��/��{�$20<M�=L~��'jyծ�U=�BgK�j��~>��,�XFj�%H�&�;׈F�{�X�y�[�,13��0�)�8�I����p�v*U�D�g/�N��|!�4������r���#6Y=+L�*0�������C��(���my"Fp.ԛ��Ul
�9p�$j�#��R�z�C|ѓ��P%�]A��:�!��rG9���Ѿg7�aQp��H[2ku�R���K@��Қmn^v���aCR+@�'0LT��r�h%#Q��������w�C��ǉ�����AkUV_�魛��-�_�X	~7i��͘�^�e�'�0�5��1�Z0���ɉ&�G��Q�9��P����f�B$�ك�0�拕�.w}�NZ	!4�/�&���)=�FO��B�;���4��h�n)�;���T!��Km�B>�t�(H��	]��1�u���?���`����7u�xl_�Zą�]��-L�;��"$���%��(�m����`T$�y�)�϶B����h�a����x��m�V�N��\09�Jt"�u3����@Pn��-���9��s}��[�ݥ�o�j���&N����/��nB�z�A�p�E�/� %3J����0'�Q_�	 ��{�V�"�e3�8�>���,�%��W�sWv���U6�\�zR���񠘷����s�L�<$����W�{9�[�{��u?%�E=<v*���BS�j�i�O8�ჭu5L��ގ��Ɏ��Y��/Ð���k�� �IbSf���@}�=��00u�6D����:��=&b�E�D;Q�O*ڞ_X̯7�ۖ�.�tr�B=�n�ǅ�	�d�_0�i)��M����Ͱ���wo���.����}�nl-��h� 6_�t1L5���ԡ_��	��LD���!����{�dwDbԋ��'E�++M�M;wd}^Q�DF�#�S�[Qp����o$]��8��s� &�� 0��	e,�^;��l 43*`��e�o�q �"���j�E1*�4~�-��E��z�������]��/�p�*�+��aL N�f����sTfq�ʾ�N�%5K�龺a���� �M�/\��\�3  �p\/��}S#"�֪�h&z�m�ef��
���xj���r�^�yn�ЌŤ�^�z\�`W�'}$�,`�2PyE��b�jD�;�CM.���KsK�j�>����\/bk�$k����n���d���~B@��Ĉ���ڞ`L /�n�G�7��R�&�TN@����^��
����������,-�ߟ^���haf�s��܅��� �)<2CM��í/q�k�j �S0�_]طf�ng���p�q/����׽�,��J0[��zI2t�3ǌ�D;7��4�`g�II%<uѯ\mY���ɀl�b}{+�hK����g��$n�ef�P�7|���ꊿ��{�d�FU�a(�>n�����eH�ښ~�j���i�6å1���x�9�����1-o>�*1?�嘷��඾êV��Pܬ���$�'�h� ��W��р�9KF.���'�%s�ȥ���ҩr�.n,Q�
3H�g<��.^_�~�1D�n�D�c�0�m�b��|��A��{���.�'7D][���K3��#4�cǹ���E����R�3)�z���,Cܳ�i�GN�>�K�.UAg�ܠ#��'�� r���6�x��1���t�bk�� B�D#3֤�^_�/�[��rۗ�OY�{
V/i����r;qE8��}��&;o��Sl��f8�ʖ$IԞ�,�kZ��Yi�Ԑ���gQ��{S7߽̌�;^�L��ڪ��0뫬�177��� �G"�$�Ҁ�ѝ�a�0ι���E�A�ue2$"���Ig=�ɋf��s��_H�zK�-k8w9c�q�ƿ��Ȳ�y��AMн1n��xD���ݛa<��-�;2Q�Lؾ����H�Vk�!&/[�L��;��I�xj�q���?�u��Hybo����D�����Yǻ�J9dII,�>OtA�Vb����>�X^����
��>�t#cr�PrJ���r�Na�Ĺ��R���qw�dl�úR�W���5"�O�6���e<&�f�9J���gK�9H`��z1�c�~D@�����@Ke��_,�`{s~i8��F���gD����7� ����v��1������a������#���H�-�`�F~ZSn �G jH�ڙh	�5���U��ϣ,=��@�� ��}8U�=TPC�q �㆜u�@g���ev��,��lx�Z����茁b���)�d`�à�2a�����4���s:�:p�	-���R��h&ZE@�+�}����8�z�%UY0V���c��ck�S<���� u/�]���z ��N�TP�B�W�'�qYj�c���nI��s��L's)�#1�g�fa��o��v���Eo�#����Ok��;U_�!Đ�_@L�v�aN�;$bS�¦A���Tڛ�n�A�7ջ����F����+��ΐ�a8�=����#��2�.Q�+���R�������G�vX^f����#��C6�P�>h1Rȏv��(�����V�аn���|���!�DZ������W].�Dba.1;�n6v��[sKȍ���8����a����+g��$�lڍ��]D���^�3h�.���d���-MD�1��ibF眕ءx�����wz�fTp{�o��Ԁ��(G�:�>������Z�iS�l��6�@q�U�ذI�p���D[}q{i~���Y��u�-W�p5��t�ݶ�����]AR�q�*h��W��B����|&,��i}����ԭ�-Z(�� ��O|�-�m"q�H%�$��#�A��)�X�ѣɌ-��2�fW�/�����qrE���A��O6��ٺY����F'֖	x�"v��� �ۯ^�2�1�\��Ȼ>�P�L5�ZN��O���I�ɦS��L����=���E[�b��Sl||�J�����p��������T�D�d����X����5��"i`so�.i��̙�W�y�YB���D���c,Ů$g�E2[���t=k�[*3�B�� ޒ�<��k0�⸜��o<�dl��x�J1�~/��9}�P�b�Kt��*��e����O��8Q�����Tn���~��E���w7fgW�X�ej�3�����)�54�~g� r�~��(���F������@�m?�6�&�ىˋ��R��z( ����mܻ��G.x�Ta�J��a�1aUۄ��1 � ��V��TV�"��(vQ`t@}y��	��S���;���0���)o=	(��,��� ѱ��[��ӕ6�����ݰ���6K_n�1M��W*m�rj��������O��W��p���Z��Zrp����R��#��/� �c3Oc�m�/tA�y�׆es�$�� �)d���6���Ǳ�s�3�V��ks��?��#wU�F�Y���g�-2�y���<)
�Z�����cnxqbR�Z��߂��}Z�T:��Yc�f�c��1��l�߫톍�G��xeo�
��A�b�F��0�/�j�4���@�~�jh?�}��R�5n�E@[����
	:�b��t��@���4s�\"���;1Q?"F���@����C�K�H`�+��X�Hq%�e_�D�i�W�<���pn��?�)�6	\3i,��J
�e$,bU�CLz�` vɖ���5���؝yb�}����q�=,���sV<T� ���/ʲv���4¿��+�q�,�SL��:r�r��0B�$!�`&�"����ʎ�O�FE��	����@��!�ZȢ�/:�YH[|����-Dٚ���ԅ����ĈĶkf���d�\6@�܎���g�]���b��[h�����TS:�%N�'�����J��h/KyZ�U���z�Q�����}D��q�k$�J0�"�������U��g��$�6hڟ&�TV���f�el�O��-v������Y������@�.\s�L�2����ho�W��h��4��t�l#����ߍ腀�Ό)�K��]����q�%]����-uK⽶��z��;O3Vw���z�����X�6Yf�� /'��j�m4� t��އ,"�<{3W2��X���ק΀�:}rF"n�Z(��d�j�UM�ny\ß�[`/�b��J��z�X�X����)46��J�k<��5J���Kƪ����c��G����hg=T����Ŀ
d	�cc��ŦdF��(;~������]��d�Ei$����C��r&Q�5���O:Q�)��;��y�3���VnM����T��&7
�r��������}s�Ϗr�ֳeH I8��^q�b?c�U;yO�8`�ԟ�`󻶾c�2$�˜�C��!U����;y
���!�$����������.�j�#2��ǆ�t=���;�7��.�D�����bm
�=��ё���Ш�T��9:�t�w)J�(�G<ܗ:N���
w(�''o{�@�H=�o�]ө�@T8�p�Lo�����1~Y"��a���������