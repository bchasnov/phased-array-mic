��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|۶��-�E����0/HE���ψ)"!J8n�t���,��0�*��W�T���-��ب`�Aolk�AT�$���Z��VgWC��U-%���W�ep�8�"�fkUS��c΂62Ȼ2������hq����Y�m�<=�����u�4�G�?��K�읒�(K�潀��tQ�34Ϗ����=��Ǚ�\{ζb�x���}�` ���%�!eg7���#�no�/q��҈�g^X��P�윅􀗽�fG��"=h�G� _]���7���]�胉]Y�#\7|��V�����^ohT����b6�厢�����Q~0�¤�����f���#Bq<��R�����p��!�J{���89��<���P��x}VUQS9hfe]�"����^�m/<{����1~+`�Ws�"	��+%��v���kC�s!��.�Z5vvM�� �|xM�=�?L{��ߋH�>�$�n�HR����Mt�#& �P� 2*�`3]������7aʂ^q���|͟�wJ鼘��K���`KR� E�F�Tќf�������$��Y@���H���"�o�hg��]�l�?v]]z��7�|���i�~?��BT~&�����;3�f�t~������5)8�,K�@f��XV�B�栭�	���ad���������yP�?��F`+��� q�-r���J���Ő뤃{���L� �1E6�&��)#�n4$���JT�d =�YpW���9�8�!=�%|$�7ؙ�Z�Y2�h�����i%�
���_w;�5�ݪ��)]*�����0�9ݴ���m���x�S�l��x�[w�
]����MN�z���&��)v�/C�7�:>��R%UCML�يm�v|����3Yr��E��h�<ps!�;�U|=�B���|9'䈙��M���|\~s��+q�$�Ŵޥ�@�r�o���p��9{�)����?�,�J�A���F�sf��a3����D�(j�fPD�ر���}f��\N�~ˋ�`��QL��^�t����:ѧ�������h%?W�o<�ݗ�xx�O���Ħ�+��(��������m��e(|��ǀ\I\�+��݈62�9��(V����n	Z�E�����]<��~����L�+���^�r���E.�Ȱ��7|��Ibd󊵛	�ӌ��BG(`��URÜ�a��]�� P��ǯ2nD���O
]˗�Q�VΛ53B�0G��a��ѽ��ܢ
1V'�B��$X��[<�99��@�>Y��u��V�g��خ�)�G*�৞�O~�2:eY�* ��ui���ޯ^���^�3���<L$��"l7KU#���K��v�^<�QJ~[9��?�6������ *vǤ���A�$�)T��]���-Lk���vH���LN�O~u����fj�И�%�F�'�8JRա�!Rﭥq[���%1s����F��(5���1�������K�!]��yxm�\�!Ǿj�F����U���o���d� (<R�o����Q��j�u����k-t P�\�o�2[�}��L��tc8��
����6h��s�ن���}�����6@=كԏ���f��=*�Q����q>�?���A�C����b����){a0RqU�>c��ÍQ2�k�[(��?��v�E~��/y�[��  ���D��Q B���@r(f׎�/�h�B�N�@<I��xZ��y�8�HB�>��[����K�k���ޡ�=�%�zF�j��PÆ�҈�d�9��FA�k|���4R�G�(����|��V4m���2'�_���J<�S}_Ri+���%^���j�ҵ�W�Q����������U����'�lwqƿ�G�����~]��6��̉@m����;I�D5�R�����T�-�����4�M�r�����ș��s�e3d�vU���2�抽#���y�F���
RV���sD�1~�~��Z�A^��¦�eН��U���
v�I��Iͱ>�dE���W7 ?����'h�]�ý�C����;{����%\�`�s���f/	�s�[U��1��T�-�ˡ�)U��n֨؋���|��B_z�}��^]j�x�6�����,�^F�Ph�H�����sq�q=���fA������\1��k�H)*0*F��%"���j�d��QҚ}�ݱ�A;�zEk�Щ��F P�_��A�j�Ѐ��2��#�������ƣ�?�IkQ4�]�y��s���Z��m�W�mq~�7�.��f���2@@boN�~�>���"�j�y��R�m¬�..�M%)25�N��>��Am[����Z.�u>��	M�f��C������A�:9��鬷}�ػ�s�T?����V���b�M4��v�J�{���{�5�rL=&���˟�R�Ɩu�����r43��#�iCء�̍��>����O�;k�m�3l�ʬ7���9��9enA|t�'D�ͱ@��M:8�C�6�8�`��Y�4f��a�-�Y�q��7%��2��Rw ϖ��E�J ��)�b��`8;�����	L��ؘ�Vm
mE����U�"#M��G(��r�WlD��~�s�eu~�@c�l\��_�
���':v�xv�ȮcdN,���W������p������1O��� q�/���[^1��x%�A+�Ve�p��|l��'���nR�军�#ֱ��ф���8)�B��}Hң��B�ۭ-��o��@�P�x�O���N�s���.4�S�́7�1�c���Q��[�t ԛ�?v���3�1h��P���?�d��Ȱ!�`�IO��~ac��b���e ���ow�{�(/�vڽ�gQ��o��.��7u
դ����[C��������]?����hd���̜�>��9��h]47���ه�2�u�
'3��8�q��4��m�[pRI_PL�wF� >���A�|�N+�T�V�L1� �0�?��7B�u��fQo[	)�~_/I{.��t���#@1�mnי%�U���mM;�
��uXDU�}����I#��,��LՀ#M�b�r���idEfW����B5��ja�2}r�_A�?ث�G����A�nf��0�Q�jv��3�[���]$���2E����� %�%܅1̕�1���=R�l��;p��iޒj;�:�#����&�%L�o��p�3s,����1�����o�p��E�H�m���+�9߿�#���J��i��5�q������$�E@JNj���|�j��Ky���=U��O�lu��n�~�$��F؞�_�Ct���j��ڬ�X��i%��cy�~+͖1Yw�)�7���t4�����W[믬^r%Բ�'��Ԁ����.^�����_b])���m.�`[юG���wء[2��0����v�H�� �b��4�3�=:����_n1�-��V$�"s3K^}9r7!�%j�&1U�۔Szۆ���N�O@aC	�������E=����؄�z�=��h�8�s;�'��V��n� {,�F"���J��-�$���L��EK��F�Ƶ����T��d��H�w�i���>w��l˴�8��C�3�W`v�>��3d���ϖ�)>�����oEm�?3Lo�~��s����F8�jM�y�
�"�G�P�e�ҳ(7��UXd���a>.U֮��ئ��en*M���k���q���w㸹Ay%�"ԏ���d��|:��e���G�S/�!�]Z��J�7�M�Z�����pV��m�#��GLx�W�w$۸��u�f��<f�\�tᆿ�:D�K�#U7�6����W�v�r���a��䢕C_� R�kr8�5vͽ|�314�C,x�a�LW��YY"�_��y�2�-�����e�&S@m��g��̦}�A�~�x���mI|:�!<d����iפ�[	���/��l�����d6��d>N�h��wn��O�+v�ƙ_G3n��c ��h
������*�8�+��k*{����q��P���.SM�F�࣑����W0�/����B�H=���a�F,�@[n�f�9�L1յxV��,�DH<4�N�g���BÙƁ�ӝ�²���1iU�����E�1}�7^{~��	f/�>B���c�ǉ<��K�-����S,_�"�d͋eh+0֢+��Ra��V����\�1h����.ٱ���N��-�9�Q�@��T��]5۟���)�Ț�A���Z�!t�ɿ��-ZX]��M�0Ts-����9�8�!3}���v�
n���M1�e�``/2'A	!���L��D����<�Z�j�)��?5�]�'��|r��}�0d��RH�J��!��<�k���NS�\��Tg铊�@熔���[�3��q����>��b�޹S����q�E�;q]h4�oT�l�Lm���L�7�w��� �ۮ��SS��@v�r���_��q�|��kCT�m���GK��ď6u������_��L� $S���bHs	��w'{_b���gE�%H��=7@|/M/��ܑ��,�U��A�`�H�"�����=s!'9�[#/��dve�7h�k��݅��Q���#g��nr�ד��'��_5,��e>(�2o��^^�N'b�rp������8l��M�Eh��:x6"aN:��v��eo�iȗ4Jp���z��#�؎��2at�g5�l�b��|�Ą=g!�T%D�����$���Q�T��JwϹx��)������F��B������b���3LN!^o�7��pn����p���wV��8�(@x�K�$i�4Wx�R��eX#����v8F�a���k�����c����-��*x�4����Qx;'+�!�D0�ʰ6!>rݵ�>Af���e��G4~�A�p����5���ig�U�TD��}$�M����O�Si~�Ũ�I�c��g���M+�B�e �S�,����'�M�+�0ڀ)��
"u,"��=�1)6N���\�X�*vj�V�EեP� "��
_�f��m��4
H��-�D���Ff��8����bz�i`�A9�G׬�x;�}b���Z-Ѩx'�5O!o�e�P��燩��d�sK҈iaBcĻu=P�����lf^� �ɪ��jA���$\�Z�j3$2�`2���a��ҏ��#}�G<ؖE��{0`EZR��Y���Y|�F�B�P1̪ECgK��كa�pA���/�`0�u=��8����nx|�`�� 0Qwjַg�u����N؉��Ddf�W/���i�`�Z;1�X�u��u����)h$���K�w1)�~����R�k�u�/<���?2{�9B���ޑd
5:���c�r���#�/��U+G�I���LG�S�6o*
MC�R^����$)�2��J��Z�����|E����.:)�/9��/vƒ�,KZgO׭l6�>N-�;�A�n�Zw.����kL����J�+?
�AT�G(��۟��تT>�c�b�;8�YUV�b�/�P��U����"��-��/����O	��P	/_����X���[M~X\u��D8%�`�1�-��Or�a%2��CwJC�V�xB��r�ޒ�l��mS�G_*�ɟ8 (_e�Z�?���{I3��L�L���nDxʓ��CŠ9g^�>l�1h-l�?�q-��F����P#�><�Ɣ�^e�(̸I�n:�󫩨y���r���>m܃A�p�.*��\Y���=�7����,U���(n��� b?O�F?�c�C��.A~6�J�[e��M+�o����:4Aġ ���Н6��>�gl�*�uM+�mF��<r��=�����d���C�0Ti�]M:T��;t���h[��ڸѝ��K�kfW٣{��<�JE	���<���S��L�o���Z���bIrbIv�$l���yt����,
���N�v�G�K~P1��**�����ֻ�V�
�p�/�55��izfɦť�zK�,@4%��0���$9/�gw�[
a{qe����_��,��M�U2_b}��l��q6�3Y���1���@���K�@H��3�	���џq��1 3��7 Am��V�	�Q@eɭ����A͕�9j�!�ǉ��a���t�0dqV_?�n�j��b��M��F��U���]���m�I)��%Q�XE�	��o'u�p�i���/�E�Q�v(�9no��t[ؓ����Į��+&+�aԔ�Q|f���w{���blr	Q��U�w��M*��"���7�F�
tD�j�Z�3��S��{�̀�M��F{w6����zJ���f�Ɔd�`oi���!�s�2��V^;.�9f�.I�����?D����ޟ��й�����1z(���:��	2��J�3 z���=���p�;��Q)r9��cT�C[����Q�����oٜh��g��dsh��$K̒W�`�_pꤋ+-D�8|]�*XE��W*9¨�=@�����^Y,��$�Î
�=|����^�]$��C���Ðޯ��5o��XNhoH#T/���D�G���>���bd�����PEuX�>�l%�h��\��Ϊ0%F`1�G8�V�g�t~Ҽx�����P5X�l"�0��a���V1m�j�n� ���UY��-���S	���p��s�ׄ�_,��^ �*�]�p�6!���LQf�q�6Hև|�%�C�V0i��0�m�fRe�� $X��ÕS
�g�r�q��ws-O�.UR&�|�&O9莛��N엑��B���mV�{��݁N��Kh.e�Ya���b<Sg��t����ߪ~��X��L<�y_��9gt���׵ɱ��Z�=Z�S9��(;�in��[1����`�,�x�oG�T�����pf�w�
:�;�-y.d)5*�!��F�eT7�hC^M�g�{�	�p�3{/b��G�v/�۱HR�V�
�f��)1|;�C�s(�\�(˪��>uH]��m��g�i��^�_3���h�:P�\�^#J^�l��ҌSr�{��#a��ս�yr�@f{�	+��=Wt��|b�GV�):/�����	G8�27�%�xK���qT�D9=Y��i��r��ӁZ�:`;op?�{�#y�.!?�K�
�#��&��<ي���I%"[׿����A+�c�aT�7�O*Zw�QkxqHiFr@����[`?#��  �$(b�o*heMG�4���*~��҂��F/�r.�s'�No��9�OH��յ�xgS�x ��u�&q��<xqa~�癙X��Q>w�� Ĳ�C�AoG����1��8v��9>��矒�
0��	���fJ��t�4��a�N��F�A6���7I��>d�.ـ���:_�SYE��S�:0q�z!���B;������0�xu�c�`�b�$��Κ��kd0�L���zV�USuB�Ak�p�ba��\���	��P"-c~��sb�W��* 0���̈qG�����|�C�W��Y�񏔓��!>Z?3.^oOTwU�t�5*Q�����j��Ւ�[�=��v=�
��<����Gf�'Ɠ�|�RIАr��$��@M�UN�Nm���5�����L�S�9YJ'�QCm���"���Y�ᤕ�;i=����l:%|�������HCnz��W:��<~�^b13�ߦ,,l[Z�dx��ث��7ٕ͗���bѼ
D;�!vx_�+�y_(�U�3�[<I�M~A�/֎�$i\����b(%*�e�bD)[�}�P���>�d�w�K���aw�����pyo����v�t1a������qǍi�\u��4^A�G��p@��X,�r��~NQw�ey��i�T ���t�Y�?���� NW?O?̽�j��d��o��ЮAB�i�?��V�UT3�4��!�ւ)J�Il���JA����<�4��tR�%���f��IRJ�O�}��-_�aؼi;
������SQ��^������g�=2B�s	�]f�Gٵ��ំ�����{����sp�/U�hCO/�v��α@�|����
c��wjBi�O�^J)R���mR'V߫���\���3�:wX��R���Z�-�7�B�0b�q��A�;���ܵtP��{1;k}��,:�h�f
V)Y��<=*���r�=��fjU�w��=��q�tTG�Q&&8Mo$���1G�-"�.�0G�T؇>0�K&r:j(B_���%45�,P�$ �.�k5�3�� ]·��ey�8@uuy�uE�5�WiT����m�$C����X}�4iƘ���(�� ^�.h�\�E�
��b���1�/�WP$��%����iO �˯�I���qt7�>��\7�g�{�9~YKg�Uѱ� �oBM�29�!>����o&>U�����je���
I�|X<RIyc�^Cw<�����2M�ʵ��������D�2bZ-�N��-�6뎻�>�Po7��S�0wP�&�t�	cD�͈��ƫ�A�\��#��^+2{Ʌ��-�w�L�ؘ�����S��슴D{i�P]k�'`���Y��M۔���?����'���ƓN����t����;�$s%("�}W����l"�f�(K�S�GƲ�,�w)J����?���
���: �%�uM�d�J��͜@�rH�%/���1�.Z΃^$��fY�i�/5;�b����K����8�7ʹ�q��bRt��Z��HBPmE���y
�G佨����������l��T��������|�ž��/�L+$�`���@[��(ďÞ����^�E}?����1z���W���jb�=g��?�x��<�]Na�t��3,��ɐ�	�s,���~���/�䝼�Y"�]n����Za2zH���pMh�pLc��k�Y�v�������"�l�5H O�� ��U�B�����u���V!��X�"2$�A�H*�2	� )?2ݗ!0?�0��l��s3锰& �f5��Nt����_K|.�=V�=����j���=~$+�Ys�tno�R�'ȇ��+�R�5�b|��6h�_� (��M���g�:�#&OpU��
��S�7�o�v�e��1'l�XZ��я�CjbP$�
�{�pDy������æ�_tè�q�j�M�mo��/E�!@Z����.Ȭ2i�D�Y���R�%+��n��(?��D7ʱ .������.�nI�1�P�d��Z`7=���^L��X=387:*�\��0و�\�j�)4�d� �d���u3�w�x����M��SDe��'=cP���ES�=2��Wˏ2�`�P����q��	M����L���в���H��:�`XT2�fg�@��("G��mC/5*�e��F�l-U�I�&x	�XV�T��M���_c�ZC&L2᧩X�mx%k5T��мM�Uu��jOtá((�a�L2geM�D�+���P�
+k����[F��1#DHn��v>a���~]��,B�{��
��ڛ�,�B�0ns���g�;?&ہ/|1�**�U6����A��$L�m�}��[gl�	��镅�$H�+Q���*ϸ�	� e	��֕���+��Fb]����5�po{ke^��]�
(��U�-6~Ow����P�ٷ�=R����,��EH�пf�%�@U�cFB�Ó/�w��Rrn��Y��r�{5Cz�ɖC� ?�C�ˣ
�4��c&���=�����x��z�m��f�v�;��ݢ/
֗"ܿ�xӰ*��x��Dv��oy��ő�x|�c�"\�7f�Z�>��IW��+�^���q�c}�S�T�r0}� U��8�@�yP-N��p#	�I�Lش��S�9�f��ž��h`�f�z �9�X�f� �Z��u������~7�-gX��J�������>�Rpx v�)Oİ	H��)Ԙ�*|���2�;/��8��h�ؿO ��:�F��i��J�I��R�S�#�r�q�2�����A���9�<p�*��&��i
o��^�7Z��M���F.�����8D���2U�Dg��e)C�6��ms^����9�sL6`�ֻ�~J��VN�Y ?�p�	'w�Q��?���p��ЪX��ID����ڎ����=5x�S�7�Ys��r��3���fzK8Ep'���������W�|L�|T(���]r����Ɇ�8���s��K4�,t`�D{�UE
�樤���'�8[��~��係]���I��"w�_��t8,���>TI�~zC��>��d�\^�c^�W�S��KbR�"���\�ƍ��4u�"�z�'sR�A�|8�|�Wqbh��0.C�Sd*�P_ Q��L����9��۾kh�}��DD��N�;�[�qv����<�el?�sD��^^X~h�`˴H������K�Q�C�Ȫ��@���tP���B��j�)σjw�\���v�rs6���1 (��N��ը��(�0�#aoz1�����X�Q0��IK��5h٢˵^��9�5և�Ae�f�Ե�����	OĨ��A�}z!��UO6Jf�H�1�_�������Vjb�}����h�wf���b���y��~E��H4��3���tr��PK'�o]`Ze�u
����>Wo�q�ց�=#0 O�Vm��En�!�}��=���8��S/C���8���X0�l4�f�Z�B���_���4 �`5�=E<� ���R��5u�*c��;�]�m��-��R/�V�O�����9j]��˪�����%��Z��Q��777��-Ju�-�蝲����l�d�����J�](R�b�&�=8�/����tP�:�d�TJ�Y��g����`�|�+�UA��b�?��gms#�{@�tv�8E�fM�~�_�-r�d���q�Q6c�d�ٸh� �6	ذ�L��f�5s$H[D����\�= Wgk6�&�dX�0�0afȋ��E:���׋Yp���<���	n4?f�Z8�F����1��O`�����&Ƕu�pꕹ��X[v�Tg��ɿ`L�өQ;k�������#'�ĵ�Zٳ���Z�}��P@�3W�܅��F���95[��ʹG����w/���G�E�Z�"��/�d���uf��q�����a�<�&$,L��2�<#q�o��� �i���q��n$+wGѩqGq���b_��Ι7�8�]-_�\Y�+ٹΡ�D3d��&�k�8����>I���YE6\�X����#2��|?7l
�x*Pl��Rk���ز� $��<
w������0Vt\;!���3b��{���qڑ�E<l������}�*PӨ`����1+�0$�r3�߷���U�H�)���\�����u��(Xh+�_�K����D�ugt��|e���� � �9yJ�&^�?����<0}����]&���s�G �Cξr~��!��*l3v���Smn�oGd�$Jh�7�Z��}�r��ʘ`J���p���.�J�vL8N����vQf�������u1\��J����P4��/�9N�#������5Y
�L���\�&��J�����Չ��V��O��d�x#"��#=�^qH�ֶA�0�I��!�]`&���->A�ɶ`b�h�A�Nݯ���=wȚ�-r�
���.;������9a�*�Xl�u�z��G��rN���aw,:�@͏�����̓�F���V4,�O(�X*�E�H���L���p1��q����+d��pX�,I��Ϊ��k�L�j�-�Yymu�>�h�M!�%P7N&�{�UL�����ؕ��ҍ��Dݦ�Xӳ����+�~>�7�&C���=�,�R�4�v�����B�}W�4�%<OSE�!Q�Ai���~!�վ���dC��*��[c��[�;�T1���U����#���i�w� �i�Mb��T� �	",\�0]��\�z�w��;�Hp�cy���򚄸;mI���D��m�]�e��b����8nہv"�䤞p��l�1���N�Ś�V���� �dLԈ���I��@���]����]����A�|Zvw�C��:c¹j+#��P~n}���FZ�'4p�|�����[�5�d�f'e�'�����T��N8g��������ĥ��e����$!c�93��$Ό��CA:b_(3X�3WB�:e������n�;*�����'
���J�;9�x�=�6'�+�uSša��pԔ��!s߉j�GI� V���`���;�۟!�"��V�Xo��L_�_8g�J���|^6������9��©�������f2�w;�S�e��U�y�`��	������;�J�s)��.n�q� G�¨-��A=a�0kJ1�@�cןk�D�E�r$�P�'�[8�1R*�7x��ѻ���mO9�s�^�t�̻�y����Bd��A8k�|][���&����@Ωˢ���Z!�;R�i��x97_M^[5.���)8���U�\e�ϖ�@#Iup�ͻ&U!)q�b����0CEJ��\J�M�fH�z�L�&&�����5�Ys��]�o^�?�{lm�H=�.glo��I]b�kMj�}��ї�	����i�*ڡ�1��OƧͦo�'���&`�f�H��6�2�Qb��^f����!� A���9��3���F�pSuu��/B�@�)+:��0[͊2-9��ba�j�鍯�'�i�c\���m/U�D
lc*_4�<ć��1�<-�P�u�CL���G�Ʀ�an|�,�!�Ȟp*�	%ZB����2�,]H��p�{�ډ[��-�����G��a�*=j�!v[�%����z,�)��k� �%v������3�ٺ�R�Ƿ�-g~ܡ�~C{�������S��	q��E���E�N�^�G�G%ir�����&�OT#�]/���~t*��*C��p�M�9*|!P�	Լ	�*7A��1�����:w;n��g���ȁ�����F��/?�H���+�$T��������vg6||��+*��_�߄t9J#��)&:s�~5?1B#�2M!�Ξ��fj��Zi `Ek|�w��$mn3SD�S�;U����F���-�i!�ܶ�N��X��������Y�����`F�ʺ9��fXm���v�.F���.�>2���ީS���*K�� �5�@��A��yGE���,
i$rP���v~#��d|�b�Qt�ě���fx��� y�+��\+-k(��Y����,8�b^�f��{z4�aP�=��1����{��8�����D��+t�j��|WKȑ���_�%��"_�>l^�2cT8��釶� 5�i�u5Qk�����q���?y�J�*�R��G�����b:+�ɨgD*#g�ʶ_E�`�i��)�A`�)�A�w]�\�d �;���vW<>�t�kkh���L�a�76���M#�=�P�a�Z^S�E�#)A�ys�u$#�V� ����c
��C�+��Cd��]N-<���=s�Q|��^Vݏ� �B�3�0w�R��2D��>ǀ�K�DB�An�x�7�ߡIo,�y�]�����ަ��[��K��؃�?��El����f��[�5TڬUU�:W/s����H%����\��� �H}Q!�	���ޭ�[��q�vb�@$�)X�ˠ�����W[�.w�Iz!x��+��ې��P_X�m�u��3�� �SVv>l�$�;�����3m,L�s�s/R�����Q������ ��֎����Z����ՠ�����
>S8&S7V��w��G$�=�&M�bJ)epc�$�	/䄂n{�c���򄎐#����bb���� $�[u���*����TKUé�������v�P��6�Ö=�3�'�j���k���d�$m�3�r� &�٨�Y���Q�o����S�+}�s��f�iaR�8��h�ƚ��j�Vx��Am�_$J�	�[2;��/�3�)%�������v��#�ci�h������[��A���q���|򐮼��*T\ ��K�c���=��0v`Y�'7�1i��S`��M�z��t�)_D�7��^�8�������b�UɊ.�t�-}i�?��a�);9�S�9�J��ޗ�4�2�xZΧ���¦��|'e`���؇gi[M�Į���ceaqH�Y.W�%�?��@զ,���ƎQ�N�J���/�е��il\���� ��;Q�A�>sM���u7�H�褟�b�A~t�┪�f���EOd:�W�8����-b%D�p�~BP�z '���ob�b�����Ӄh��ՠ^%#ﷅ���efQ���y��Թ�C#�XX� (ǥ��KZ��{�S[��:X�KN a�_<���V�V�p&��0Q��f����g�إ���^��g�X��!o�9�s:Ҝ�PR��Ŋ�ɬT1	���~�B����L>������֫PU
T�&�yyC?eW�Ο]�n,�xE=Q�=�៵���ߺ�||�r��.�G2��z}�%#��>���j�S�y���룮�.w��L���0�M��P����)�A�O�C)�����{n�^�t���#�3.�NZ-��pW��P�h��v��X�RQ�]_��1��0�Ik{N�%#��}Ȗ�#�_�����p�j��	����=����g��E�;��1z)@45� ��Z&�cx��>?as��<�Npn���c���3�����VU^P��DQ�O�����d�xT����� �g:K@�Y��́�i���=�,r�[�i�' #n�vg
KPԥ�g/��ɂ*�����t���P8��7APN۹��\���II\k�l�w)QϜ�خ�lF,%Ƀ�)��~�_����Km�	��Qĸ�Z�t�J硡������a�^�/z@�$O���&};��S= ���T<T��e:
���7�0��k�?��R�?^�,E���e�D�����VN���'��F(2�3�;�2�d;.#9C_-R��q�Y�ųM��;˅`#>��V*���.0ϛ��X��d�>%�(�"��`�s��l)���Bd隍1D`�B�\/�c��Ƨ8�܂��MڔsX�w�i�_K�
���ƍ� ����H?$�Y����\UV��{>֪��T�n�]^mt��'�?��p�0���5*>^�������o����[��M4h{�P�ޡ��ͣ)M���w^˱U��d�T�Gw=A��rk��;��nN�b�f`�K��JcS��dt��=w���;,������?�@���&�S��rZ!��=D�V���9G�X�G�Ψ�����@��ZT�T6C�j�'�{��_v���2�ە���_S�pw|{�E1~��?���0�iB+��� >�_�G��]YV.��i��:/�K��Vk�|ލ�W?S"	?wQ���%eu��0B��ۙ/�V�ܐ�I>b.�-V�}��N�hfۇΉ4h�����kM��tft��v��д�����\��o,b%�5P^�� ����G1�k�@���\��=��ͺ��y�`�Z�!�@���p��z5��'Y��$-�[b� V�9ui�#U��Mwܪ��<�my��f�������9T�3�\f
�phH��u,z��4] jx���̋��O݅�}�B� ���;�*[^g�hIW�i�w{��x ڔ�Gs�c�0�&>>�����%��1&�6�� ��XU��e4�^+!����l�e�`_�V�C�M�RR*�z:f�L�*�����<WQ�����T2r�,�=��5��p`<#�X�w������w��Wg�)V�ʤ�-F,�zЯ��Vk��u�aT!�l�!L-h��i��W���f�x�C`����W}]R���R�*�̥�?�J.���ш���-�c��,�W2�Ř�0���ʇ'�B��4@z��3d���+k�l�eF�D:�1���$�d&��n�Qe"E�EsxK濾[�|:���P�Y��+��^���W��k�o5�\����@���m�����m�Yu�'*'
�uo9�����J�#�c��_�9�/@����8>9�A�u_�1����\�=���:�x�h7H2E)�s��
��c-���5O�_�TP�́U�K'?��U��VjR߂'(s��F�
4@V���\��>l1�gk��N��!>��������
��
x�)É@�."�`l���)�i!�v�.&��^�|�̘]=Q'��oaN��>%��j9�gt�r�~m����|WL�����'��ɕ��s$pz+�h���ӣIV�i�T"`J�j���k�T>E ���#����_0�_�
����������jk��F��Ǝ�f9���I��m�dX���yFE�i�<M���t��\��B��tv�
�I�)G���� @�ŧ;������m	ٿ�_F��P/t�'��HÀ+J��WŬO9)�ܞ-Vү�N��wg��e�'I�=�y=��Z���`��Ͻ�.�4�����Mf�"�
��{���Ǘ5�� �x���\�>	"ST����dv�0���ri��4h�S#zT,��{ľ��3�Rkk�h@��՗�ܚ��x\d�I���I;�.��(2��ޫ���R�V���o�T�����Q!~��jK�!P���"����<��b�R�BK#�x�[K$�؀*��c �a�VopE~C�����{�CSI�������@{�����I��Q�P���f�7�T���н��[�̩	K�w��+M���z�k?K�����_��ᱥ���Jce�����-m��:{�_�J���u�y�U�f��b���uo��7�~�K��F��yN�<���y<<G�tXP�Jf}U>��	��������!
Fg���+=��H��oP�z�ޚ^���8��2��6�g"+�|O�Nĉ�_{�"&SbQԊ�o���>��$�ǟ����o��O�gk��4�%�EgXB��6{k�_��Qq�Ėږ�3#д�8�����0^2#H�L�{�ny,�~����95�Jo���a>���l�\������֒�b2x�l+�Rx�n;��J2G�3Ʈ��8��`����nc�N�`C%�_6� >��ȴRx�Ig� c��G��!��z��(�Ȱ�I��=g8����{.8�N8�T	�_�m?��ɕ&[0=�~u{w$�$���$�u�%ԝ�4�Z=�8�`_�=���ph N��%�2!���Br4�&�ݣ�� ���a�ށ0��q4�_��e�ڐ�n۪�7��>�nZp疍��+�@k��C,d�P�G��`�ż�#Y�$���Er�r�`��D&��*��K���R���w�Ń����7�km�s�N_U��Fv3��8*���'�Þ'Z7)3��k�Җ
�7 ��[�M�	UF0�/��ew1��|�b�{����C,R���7�&�.Z,9�1���8G�V� L����!-X�`�E�b�C��#+�h�49�*�x̫C-�Hf�O���A:!�5�O�.5�x�n����0��骞u�%4%Ƿ��|S�f�#�ŝ%<z.LEpPtl�V�?�z�^o���H{�͙A�H�?��t�8���C�a�A�f�
Mߣ�oӃ������{���������֞�.B!c������d�����o��"�a+0���i��.��v�Z�J�z!�k����Ķ�H-����gAHR��z^->�J0���cq(��Lw�� "�ޔ/a`����`Aɥ������}���fչ�+#�c��;���9���6��;�F^)v�I���Ib ���,�<���f��vL)�{~\��G����p�ĳ��#m2�89N����,;S͸�b*��s�v_�,yp'@�R_y~Qʎ�J�"~�:o� U�r�eXŋ����Y1;�e��>��1�/�-"��������sxe����I�T�?�������@��-��������|�ח!ٵ��@q&�YS���������p�ct@q���XY��졆�h�����J�T������1�ΜVj�Œ�E2!sX!����p:�o��"��͍�rd������kJi �ekn�¾��2�v:��C����bf���������U�/�2�:��Ez fډ��v_ ws[��L<��|�js�s���Na�W���sF�T���3_���C�:�B�1˲R%~���^���MZ�{v�Ac��8^��uɐ����[e�Lƕ�VO��r�0�AA�vD:n�Y��v;��Ӈ�"�݄n��|��r�v ����)X�\������8Υ&��|}�и�ި��HUɚ�'Qg�~���!�DEfU�w�&2��|���E�/�|<���&��D_�HU	l.Bgie��S$C�_,��S��Lך�8��ދ�v���h�o����k�n���B��\1�\���*3�#UG	�,�/-o�)p�H޻+`~j')����*vg�t�����(uE�M^Qפ/���1��!h�un6J1�*�"��Ē,�6�S\��Ԃ��\�T���n���%�[iU�u%`��%��� N�l/����P����|�b	z��* Vf#���ű�x�>�P]�'��r6CЛ_���e1et�KT��s=�}�?�F��bP7���DI%��^�j]JlI�F�m�aN�VB����B�s
�G��8O�HPA�{:d[uu�7OKP��ǂK�P�t���p�:(��1��4�L�Ka&�g���ʈ�[�I'Id��Z�?�"�N���w5�#�
���c�,�pE�f_���L�,7�s,�bw�ޅ˥�isᐽ'4u��&I�!���LS���ܜ����q?��PC`A.��$��v��uCYW��Yny��J�E"fW�6]��f�z`���鑇�(����a�������y?	4ɟ�m/f��3��G�D�A��E��=���X�I}A�^��_4)���xJ���<G�ma��T�U?r�Z鍖�n�	���r�M?��`�F2�.��E�Kv�E���h�d���G�^T/�Q����Yp����x�	�OA/`G̭��.Y�s
��͇
̚z'��3L��=?.�'R��9p��Oh������@���6����;����{sy��	�q̴���I8$̕:b	2��B�`�#R!����K�ߤr/#?3� !$�����5i@�Gͩ�J�aR�7;Fڮ��s���TüsUO��J���ITč�
5
���y�l=��;��J�.��Ad8��l�R�<M݁�q�X��kX�H���ύ�0����"���/vA���F�Kw#�_�0;L��}ǧ������^��d�
�~�9��`˒ӯ�&���>[���,��Ͳ[m��"�lL�7v�@��h��Cj��h��;���/[ӤS��f��Ay^����ԅ�mt�"��V�뮼�=�A�й���V�)`�ؗ�o�ev��`DYhl?�Q�P�$5�v�c�ҕ�>_���xF%thy�� �:B5㛋���0�r�gr2wKz�6w|TG�̖+QӷTb�&�`�e(Ҏ�7��ķtAڙG*b�	�PP���5I��)����߶��z���%��%K���o��Z�@��1�6K���f���6vv�-���>mC��y��V�d������40�}3yA  ��jxP
����?�D$g��V�jPe�f��{p�؅do�s2G[$>��y�L������<��_��Q�-6GkB��;+߳,�#ʟ�Z sΰF�"�⩬n�g���/G ��51�����z�V�I�E����V�]c �3�MvB߽4�Z�Qͤۘ���1"�])�5R���qe�Q�i���
�R)0a���������t�ਝ4!�q��Ǫ���&�X2pb��ך-���@�{kzNG\��~\�ī�����A����G%���d��=mDH�Y � �������-Ul@� ,���lu����P��M�K�G�'9��!�#I��ʛ���4s��b�e�/��k�GZnQ�����q q�) �x$�� �T��ʟ�0��pX��6��B��G����}w��.�(�>Q�T	p1��C���V�=�L�jN�A�'�(7W/�?��ǧ�x[P��#'��mNO�C3��ׄ|�B������y�]��I�>��^�|�O[�x�X�$N&s��8�x�ت��:��zA�#5ͤ��{�j��}�O���9��w#��#!{�yɛ9��?B�J0e��H��$H�&�"=�<�@��Ǐ]�����v�n�[Zօ��Sdw���Nc���wU�R\��Id=4�)��	P`���w6Q��wY���0XD���R�\Y)�&������AV0c\Ղ'���c|�F��1�~/h�Me؏$���k�,坋������U��\@�ci�����Z�B=x�|���ʭ4#*W!0���4 ��V�b�v�FAa�I� ��m��ՔzweZp:���w��i[�Ѷ%��y'4�Fu[CJz�T2��X�T�*�%WJT�D��݆7( �v�E��Q��k��$wg���,���I����?w`Y/�r�@��� �\ƔJj�|3�Z���&U���B����+[W���Ov��a�h��������3�P�������w�n��+K��	q�@a�����Y��g	^ �*/O�6-�WJ�(�Y�^`Q,����=��E��~X]DJż����9��O�' ���o����he�=�)7Uqb��RS>�=^j��Y�,F���d�5�n�����u^�4;E�z]@��Z%7����#]����}�;��#��el�Xi��)��-Paa@��W�Gl%��a�Y��um�j�%	����-z�(�i��u;�u��^�݈HG8�%w{�n�F��z�D"5�}�G�V�6v��v���`�~0y�R ��&y�ъ��)+]{$��X�ؙ��~j;�	�'��^¾}��m�XOmD��K�y)���۵�_|��U�~p�<ժt���a�O�w��"H��xG� �bX�ge��+��~�TS�L*���}ça��Q�v��i�Z*T'&�~����Р���+�:Î�]{o�/}��5&"g�jW�'⨈7�v��G�#ufF*\I�n]�r�vo;u�D��2ndy�@�:F�z�2���:^�N����{�t�Cc1{w�i�,�Ko�pq��_X�'�L��:,A��b+!�6mj�ʟV��֋�Ur6�������s��.�<�2���T���psfd��8"��	}�C�4�B����
�kDV-=�H�މ����p"b�bу�dj��$�1[��h���u0���\�dSF��E�H�Z��C<��s>�~�G�}
���=,Ț����Sh���(�4�ԗQ(p���_Vd�4�ܜ����D|�ci�Q*,���ZA��S��yaq��L6��
P��2�	�\�{p>���,D�Y���3�B����q�7t����a�$jl��d��de���O�y2�,�D��x�ά����������NB����m_;d��e��82��U�M�@�]7�V�G�FԱ~LE�2��B����M���)�q�̐�_2���ȇ����S���ȱ{��F�ELTh�|m�5f|�,I��Ի�=��rg~��M�(��g�l&~�@�r�=h�&��hu���=w{���۹�b6s.o�ӫ�EƗ���:!���@�P̣y0�ɲ����b��4
&��O{�ǋ��i��4�]�97�J\W7��v '��I�ȟ�g)�2��޷P�kݟ��ŏ�
�����л��������m:H�����Y�L�	����⼩xgP��o��2X��ώ�O�h���;�����1��z�L�H�m�dB�o�-����< m
U�Ӫ�gY�l�v�#�x�eG��j߰�ۭ��Z�Ƕ��hc��ݳ�=�����ҹo1�Z�K���K!x�B529�\x��fV]�ÆL�!%O7�����27��/c_[-{�Ҿ���P��Aͫ#��h����p�#wDa��$��ww�&�k���~p�rg��L�E9�g�hHj�f�Fy�9�S�A��5��]������ª�8u�<PMpt�+��,�m�F�}Z�8?�'N�\�A�Rr) �ብU�XQ ��c���85�0�#�^D���i1�N��&ա�޼h+�S��m!�|R���HAbJ��� ���I�ܨ�K79�wvb8���&���΅;B�OV����0��O�����y�wz��`F���6����ȋ���哮U�����;��@�]T1��bib�)
T�c��0|�m�!XQ�a�A'��#�ڣ��D����tl��,�F��%ev��/T;���#����Պ��'"	��l��e�� �W�س���VW���%4�W|��,_eG���Pb`�de���"�܀�}�O�#h��,�t�<K./�cf���[�=�C���3��Q\���?��1�\�	��=�V3�K�*B6��6ҋ�r�\$.$�ȉ������(����&F_�c�����OnnJ_�n�:$T����x�e�=%`k~�?:\3��T9���v��e-�7U��N��@yc	�<���0�f�5C�=�L�賃xXY4���%�O OG�C���	7�-d������l�cI�0V�M���Ll������Z���IUp,��q ����lK�R�o�i�����K��lc��t�w#�Y�&��i��x��A� npi H�0��4�
�5D����:h]#8:�*[_�X�7����ϲF��fo`oH�b��:�h��7��0]La5�E�����6Lܔ�q���¥_���.�
}R�s�־YΛ�@����36�tE[~6���2��_���e�Fx��ƻɲ3�?6�;�e�5-��>8⺧c)���$�RVw05����eĈ�k�r&���q̐ )Q��lUMP/�wy��6��JE6\�Yg���]��O�8	����L�PN�����a����3�\N���h��VJ/�7.���sl�M.ruQ�4 <$A.#���~UT(7~�����Ҝh£c���y3G�(�LePp�Σ� �S^v9�UiD;�}Kׯ��� B�H�)d�XHL0��~"TɃAn!�?��^'���!=l�!OZ��|��U=k�Mt��X哝�HȅS-�'�ݝ�g��c����`?_`Ж�q8�yuڃ<�����6Қ@�ThM��_����Oq9Lt�] h����N7�ڄE$���|��r\�З����f���b�l�u >�qg���,�<Hv9�>�A�vY�e�l�$�M�Z�9�ϰ�ѧ $t�,�M<y�崪CbG͍=G�UH�#P���0�3���@�lo�Z)S'���d.�u��>S���$��m�%�T�Ju��ot��&my�	�3)lDK�Z�Q��ؐW&�� MZ(��q� ��9V.�l�5IJo4�0�!;��Qy��� ��v
ے���|�)����G�=R��^*���ͳ�SF�0�_�6�ɜNy�n�Ϟe���L�v&��H}�Q�F�L���~�M/��e��3ME|������Ռ*�t�4�O#pB�@��m�J�'<�ƚ����cZ���a�>h������Fr&���~�@7bۉ�[*������u{�kG�>L���La*$a_ٖ��jgB��a_-�K�@��y��C�AVz�X/�x�	�j�����,�g�[q��:���ꊱ�}�K�d3�/@�҂�@�o9 I�xq޼8Oє/�$ѪK��ۮ��U]���G&ߞ���� `���+a��T#~���C�6� �3(��T�G_n��� �?`{��_��w�3����a"i�n����gL݇��~����|*�;Oe���u��,J��Uضv�A�P6���x� ��{��<� �^��+�-�J1R�B͚YZ&xG
c�����`�W��z8<�ѽ��t�������������W�*���JZid����O�%7?�] E��Kg	*s��>��s	��χ��F������a(Pfu�c6����=J���rJ���X���7L�t�˹�P�eV�[/n�%sΑ�4�_�
׹�}O��ej�Y):�ʎ�,��9]��ȑk��ʐ��]�e�
#.���j�Nq;��ז���>;f�i�I�Қ6&ƴ�o19=?��~p�]���l�<V�.F�O�t,������b⟬��c}���Q?�b�ʈ_���X�?���=�p�xJ���C������	]q���gc��.�?�/K��A�S3mi?�'�����A����p��z@�]k ��?��Ś=�
O�TP�#Ye���.֦��K����b��׀W�%}����[���z����G��m�;H��fw��b����0��orT ��_N�(I������4�xE"�HlpɊw��\�SF��(�˺�f��g�ç#�TITD�����3�����*�;'�!���bpJd,N���Q�i�74��mVr�"eE�OZ�W�)ҟ�v�N��m��Aζo͊φ�ҷѨ��@���/�-h��ђ��ݛ�)I���}bl>(\P �&��A��g��@��!�h|���FF�i��$�K��*4��&���+�������JH�L#�i�'�w��w��/�Q�OȤh�|hWщ��(v�ڳJ܋�ȃ|�[RF"�r�h蒜��h|}���&]CX�:����ܵ D���_G8�ժ�dx���gR�if���9�@�Q�q�*�R��P;>X����]!�hD��na%��,�A��Re�u��1���uťi��P�!�d���`���-)��+D�Į2D
����"}l5���No�n������'�P�ѷZ�*�:�z[#�
Y&J"��J��Y�t��Q%J�Y�giV)���2�<.�Џ(�DZC�V�K*5/���g�������z],nz=:���A(�z�/�����d`��5G����N�-��nZ��Z�� ��β���a��K�s��UT	O���q��jka�ӄ3�5�DOd�E��Tڥ�R����d�}���)-,�&N ���=�+:J�I��}��у�*c�i���D�L�
"Ր�"�I����t�wb\!�y��3�WMCA֜wyT[0�m�x���8��x��fI�P�����!e��U^^�L@m�߽y�.�?6��$�-	�fG�f'ڇ%�(O�ۊ�-]��ß������+��?�QNw�,����)��y��$c��_L�����l8�ޏ��C������A�䣻(�C�]�F0=\��(D�H��`��EO�
u[;�E4G���)�|�M_�� �k\�Q1�����^�8w������%���G0�}j��L�H�ػ炌��&O1��)-�&�%n�\"�����J�̌٭�G��G�?a�d��@��nM��>(�I�y̩�ɢq�䋥� ��e�*��1�x'�l|�3:^sCq\���.�Ls�<�F������׿�4u���62ŋ���cyb���_8)��"�)t��Y�w\��\@۳:�+0�tΖO8��C�#�!5��$72���g�N����{ò��PG��ǅ�Vr�Ϝ6��;Ve�����3��	� �BB�_g���x��dmQ����k�L�=ܲ�)��v �vh�����6����( ���b#"�n6Ҽ
߰��!�)�/KC\;��<��,�|+^0j��?�Ф�DÑ�q�R�]��m-&���h9�o����E�m~�k!�w;-(J�N[�  X�U��VKj<�c}������\�&}5C`�Fq��ƭ���{�;)A��o�~^�$�_���^�s�[������ǉ� )����\��3Pu���FU��,�6���Ehe&�%�O�M�{ٸ��f�~�ŝN�8���h��Tf#��(_kE��~\Q볠�+�zG4s;5tE������W�x\zK�m���$�ZBy��<{�y!`����p|:�^_�?���f��;����uu��B��#Cm��D̪�aI��z��1�����<,��6Qu.x@�rQ��>����R�U��tmNhq&��L�J���J���Y<Y�����9���j�%Ss���֒o�� &�A�>�T�����2��t����ۉ*N(i���	{�.�=�������+��_5PH�hK��=���ke 8׳b�0a�[�J�>x�U߿d�b� w�y`Gi)**Wq���E�Vw��?]����e&������`�^�,�L��Bj؎��~x9��4���s�ҧ�$T=H�� �ޅ8> g�_<Q��ͫ�ESOT,�r��Zf��Ğ�2��srޠG�/�ty�V�Z���?�h:/���O#�lf3�)#QCA^����+�\�.�A����bq�aIO傝�D��8�-�C�������1W
��}����?�Y�*$�M�֕��i/<U�'ڂ3|m%V�?=�(󲝪v��K��n�d�LR���d;�nq��x��1
'�IL�J+�&�� 耫/�eU�IXN_�}��K�BHʾ�s�7b�`aG���腴�u��?Θ'�t�6��86{3] ^�[�f�[����{et��J�x�9�=���2�h�{�Zy�FJ�=-:
��5�{}�&P�ʾ��1�<a�-n�+�]�y�P}dn���9H��̓�g�Q��@r����rɯ�pE�����5���}�[�Fx4G�?%S�0gCځ©�*h��0��w�Ǩe�V���M�Q�H�j�8�v�k���Ҏe���2�	���}��*ȗE-TP;��� ���p��=Kt����)P9g��i2�+�~�@)���o���]�d��l|&�ߦ3��U�?S�W�r���+u��9�;(�n�މ��-�!������D��a����~"��31�2�·�-�_��0��`K����.WFo%y�k�i�bn�hڶ��{0L.��s*l��5�$��z�Ƕ:;��ag�Zd(�~�&&y��7!�����w�'�c�/�Wf�� �֭��;��B
� 9��;�X�*�lNQ9�(��g���$����CԬ�테��I�6��JpգS���0����7��(���t�������R݇��©h^M �
�I�U���@'�H�#�ᥖ�OUϊ��j����'q�!�H����0�YKC�x�13y!��Y�w��}��}ԇ�K65�5�1��+��n�$ a����(=��٦gu�V�.�A�����p-Θv㚤(Jp)H�)ܨq���
�E��u�����)�r I1[��7��}��|�ǂA1��^'��>+	9����"�5�6J�cX�:f���17��L�jb��2²B~^��iRjG�qw�y(�$�+Rm� �y�=�6��*�
|%xb��,�m,H�Y����V��!�%#"^�^�0@l��	��(--��n�m]�@�9�5�]�a��/��m~�O��!\M����D�胛O䡬W��XM�̐���b�45�P�������C��Ϸ����� ����0��7�5-*d$�+q�GU�Xz�k p��K��beC�-6���v��\�b�܂��H�?v nta�!�l������Q2;7̟AX=�L�f4P��q��t�k�q�x$կ�f�)�s�>Uca�{��}����2�н�dc�c:�_7�jڷ�0�ʚ�@~q<6N=�η�&9Woh���^�Q�>��U���ʷ��,O~�1�`�;�#�?E�B��ր�~@���ӾI�D�
�1��h 	R�T�1.y8�#���H�Jwݼ�x�;o@V���O��{�j�_ f��҂�#�ML�CuC�im�|ĺh���BA���q�-:�X�"q�TT��ED�=��&�mn/\��tڶ�-�s`��,���'��z˺�_&�;�y,~[�Y<dDk{Q$w/�,]܅��]���%��902!Q�aFw\a4 �\y�ޙ��b�P��c���A��Br�İ;�>���}�>CS��R1��ЖY8�:'�økf̘9!��KW�aWEuN/P������ (cF��o���.N�-�G_Ll\l�*�����~p�G���_�Q]���g217��c��mi�%T�-�0���#�ye.�X%���F��tH��-��"�R4T�4<�(7f"ц�<cr��'�e�p*� /�	䟴(�>�H��PcmZdƄ|k�1�K�x�c������ Z�eO&{�#6�`��a��J.8�<V^q�%P���p�B��ta��q���56t�ͪd��]xg�υ����V@n�<8��Us���ӭD���D�C���Z�&i�(_�D?���a�,&�"��F!���Z�P�(�j;��s��(n����*��ĵ�2��55:{J���!nX�I����$`'%���%��XH���l���'��z%ib"�(��Uٟ��)�fe����8 �g��!��_�����V�E]��|-ȹ����-��޽�������^g��ղAF���>m7"��>��,�W��J~C͇V��b��k�4(!���E�����O�|b�{��|��k�s�zZQ����>�;6)Ӻz�;�:u޾�V�{�S�
��]p�����J���Uq���ڋÿݎS�b"����N��|(�J).%�9(�E=G*�z+�}N(�kMq���S��E�'�3T��6��z��A93F���j~ߤ�1�jܤ8LR%�DS�ȣ�u��j���hCDN�m��@� �~sB�)��4���Ƹ�h����h`.��I�.�I��2Q�i�jJ��r-gI֢Gr�KӁ�U�?b�J��tK&|���%��z����f��N���='MY�ذn�NYShO&�ھ,��$7o��%'�b�2�1�&>����8�b���U�G�k�6���9�"���֍-�����%f�2^v;9@��I*�������Hʝ�N��d��b�H
L�I��]y��D�ғ��u/����w�_�G?۶'ÄeI�&������ꊯ�L�@u*�{?�O1�M�v_~'W���-�l���rP��>�N�*�
�YBg�x�7����v"���8Ԙ�� �O�[0`��3-��U�%��yw��7ҷ�@��=�<��`����;�W:��:�Y�&�P�Ӑ_���W��R�,I��8������n���Ey0
VjP*���qa?Zږ�.?<,�ٽ���鄊fP�1��B��H��
<Դ���W��A����$3U�aG܍,œͺ W%n�Ei�c���z�B�A�]%α������E_|*(~-�ss�r�݁��,���ALq}��Bb&h�b#ɚ�����k�* O%w;A�U�t�\��ц_ >�<��]R%��]���T[&I�N��:4�L�?} E�ḑ�{�qܖEt-� ������&Ba�����k�ueC�z7�mWg^��
��Fvgw~v��)�.Ǳ�7�.�'}�e��T_@Dz�#�bq"����d=&̘���*�4��C�*��&+qPl��C�fh*K�%&%w�𭞄��="�k�!/Sӳx�N/"qB�>��(�N��p����A�$/���4����O9�<;�Ŗ��4��(�0̗���Չ�*���z�ݦP��e�Vo�U�/��X�΃�u�ŧ�a\Z�u��r6DX�F`	�v�	�H#�$�_�{�'��\]z(���Qs恇�&/�5C��S::Q���F9��#�&m��Q?FiU��X�/�N�ʱ�������&�8Xj�3�]��U��6��R-�-T�òG~�r��[���^w�|3�[kW	O��_�=Dq��-MG�	f�k,4�δ�- K礍�F�]0(�N����R������MA�/t��g�;��	��������vdt�����_�G��g�L��jr�.�g�c�~\��}jI�*t巌�\=dQAU��F^���xt��&��Iy���\ �t�$I^�E6�
��qQ�ߤ�mC�q5ͳ��Ѫ�/J�����c�� 	�mM�Z�?ѵ�&�@�᳥��r[�Ll7:Ru�S��N_��w,��V�޿����cNH��1�Hr�*�ʒ��S}�bO�D�Z�.�����xUG,�[�?��#�A_BF������&�٤ ���a��h�rv�<��`#�V��mˤ���mu|��0IV�Qe�D�7+Qt��賵����;^�������t� }xnD��H�m�hؓi(�4a�rce�(G2�t)u�T�����ڲ~�~�*�o��r��O)uM� 1�Pt-'[�D���VjfSt��;ɻ[�����ñK8�ѱL�z�.'����0\ܖ�/�D��߾�hͤF��<d��M�94��Wv�����'����J�,~*�S�%tqht�yc�흧������+�sb31���?�w��w��J�D�>�,��%�ǰ�� ����\�����������]G!�Oۛ��4t9�AdE� �ϡ�[�LJ��g��]R\㩋0���r�;��O��|�%+��؄��	�F��?�*��F�Y�>�ݏF��p���A�zm�Y`�n~��k��T���{t�"o���It`r	nE�y"�Y�{���MJ��JZ�ߢl�X��
���H��8��Ֆ�
��+\�q[ȯE���&qv��;m�a��;;=�z�]Е�]�W�����L__t���tc�a�{I�[�c��EW�}#{"!�A_{�,�$�-d��B�l��tMl4���Q�un%��t�I��<Um�U�Ԣ�rك��7�x��Q�a��o��03�ߐ���Qʟ�!4����|�l]+��]�=(�Rp����Sk��ebnOZ0�<ٕ�׸/�ufpc�ܺ��$=z���Է��e	h���w���~��ԩ��%�n�n�38�wٕy![]�l����� �U��ί��#�B��[��^³����=<�^"�l��;�x'C����I�RfQ{:�D�U��2�4�
�{*/6�*�u2��SO�S�%���?�������ࣾ���@E�A/+�x2x/�<m���^ݜ�5��d�|���z�ܻN��J����F�m#7� l҂��r_��{kˁ(H0c�}|�׉��ݿ<>�A-��Li�L�����CB��H�Rw���4e�"�����4Y��q����Uu��O�+�ħ�H�$��g��a�ʑ�n�s�*�`d��+����^�31�ZD�Ɩ9��:Q/�_�3�wjt�e�Z�2���;)Gγ���Wd6 ��-8*��¨����<�ō"��V!�44�m��<������qǘ1sWV#�: h��6_o��h����}E59����\@�ٟ��y\U�|Ԉ ���&=Ũo��#l��c��mSa���L��#3xC���$�	'���M{�6A$� 08�~#[*���$�3:�Bمs@`ʘ���v��	0*QP'uA�G�)C���yv�!��/����Rה���-���6��z���a9z�K=�w]����̜�2	.�N�BO]x` �jI�hp����9���6ջQ�)9&%C��4���,-2+#�v���y��)�A����v߾�K���j���i�����م��#:�Wt�kG��G��i箰��ϵo�'�����r����=�f�q�ix�*45�3q��P�n�Yjm�d�����3��M��X�!(,�ϥ5���˥j�o���)��D��p2R���c��猆�q���K�}_u����[%~4FD9�.��>l�xqH�:�M>&hлƺ!�+�ovH��{�KG�yĨ9����a�|j�h�X8"{q�_	$2��qe�oF$!�uZ�	)[�5�o�F^�a�󪧩���!���b\Y�S��5H��n �Y���ʺ��qFQ�B�ڗ�e~'w?v;�OU�����o�w̡!�տ�zꕗ�RM,1��2[���Дi��w(8���#��w�Ho�R��,�"����_xO�V5J]�Y[{�.��E�@a���7���(N ������#
�ғX�ݣbT֠}�#�鲦Qߖ	���t~,�d���pur ��q��]�y�Zl@�
�^pl+Y�T�aB��iKW��|8*�N�Y-M�K�����7M����3�/`���wq��
��p�
��ñi�=�|�p���f��UV^�Ν��q��=��]��[肌R�h��$9�����8�=ˌ�K.��$zq�}��\�,n 鷰��b	����8PO��
�]���2Xx#�J��i���ʼs�����*�7.z`˜
��XO��0�[T8�	Y�Y���.j�5��ܸ~4�p����9�@�{��.Y��#0$1s���=NƋ�v�^-\�@��������[��	�q�����K�w�[n���v1={;��g����l.za�	O���di�uѠ��U�S5�cl��JU@kI���T\T\���������=�w��v��ڴb];ceh�l@i_X���-Y��w�[����#�;��� r�c"��F�I�cM���W�CX0m��a���b��K#m���i�5ll�pYp[Wrc��F]Sꓫw�z=�0lU��۶@^[�W�2�K�{�u��g�m�=P�����6��D����\ɣ�[ȝ/�%]a�C���06O9C�o�6X��������,����\n!�1�?q ݧ(=��b|��⩏���輅�$'g(w���c��j��6[n��Ӳ^(�A�q�㹕����5E�|.D{	In����.u�����H�c�w���m�:(�eX(*�^"��w�r
����_۩ڄ�y��8q��Ր2Dm�
�Ô�G� �Y%���zY���z+��!эbtH�*�ЩUx�zǂ�! 9dsDBA���ъ�R������I�8�\�(��J�Z2	�X��#�~�z����y�&���[��s&������ˀw�7��6��X_���;�XR�k<��},=�\,9�r��=围� �d�o1� ��Hf8�2�,�$Q�����f6 ə�{,�CKg:��'7ⷐ*�FIY�O���$�%h�AiAі��d$��=�%`=P�:��c��E��5���K-��Ӓ����ԇ�"x�k�d�7U�z9A��L�Ϡn�������C('�S.!0�"U�'�'?"wcoUK,3��C7���C<#��zQx�����ٴy􅔔˸��sc �"��9nk���f�����^"]�m��S���~HT�N���{��̼�^��
T�i��i
갣�KM 4EW��="�`�q.�2z��["�ę�%�ʀGbcv�qs"9�ϗNo�-����p��F���x)���6uDi#���X�^ץ�o�76����������^�x��p�.���I4�HP��
zT?(�%8*ZV]�/�;�ǁ�=y�� ���=M+W����x�FL{t1�nGl�*��|Pd���M\1��+�K��D�Q]K���>�	mo�5���ub1���-�u\q�@F����
mCH=P�N�|�RlF��������M�"u��`!@��ћ
ҔԒ`l;����8	����;i"ZQ�C��9)���֬��u��&g����fRsWZA�ʨ�ih7V0��`?�wnp��Ge ,�(�
&���A�!"�G�����{`i)��eʩ%d���2}���J�W�aـ�����r�Δ�a'�l)(s`�&�EX�W��ǂN���_�tGA~b�D^��iz�=���
��ͿT��p�$�`_�D͓��x&����j\�0�̹>M��)ɟ���B�O4�,�q~h��᥉s��X��ҏ�=�,��_��M�e�(z)�+ϛqI7��[����]�}y��s�š���wC&p�1�,��X�+���̻$�)�?�=s��Z���5���
T����������_ 47_���ɎO+�lU&�<�.���.o�,7�}rOj]ث��hޜ:���v�.��d�M��uӈ.��bZ� �X~?��alD�_p�%-���D5�he��yq��*�b���e;�ʫ�)�c�l���$KE39R���o�vݲ ��=pbJ�qT��A�`�:Ճ��>�P�M�b�?���5�AB�ذQ
�*z�=uW8�K��p���%�z�_��&Ek{?��ʎ�oLc�T� �Ru/�x{�(�����ΟpI�9?�%L%�<��DP��&�6ԭ�8ޞ��pY��Z!,�,-�����m٩��̲�4��W�zq,���b+�w�P�6��Q�z
ч��	�=R�q�msRr�/@��;Ѹ"C�)6�2ն�>�ll�}�.���kՐAj �o$V��:�S�WS*A
Se�)��p��>��XF��4�Y ���$ot��Ro�p�)�1�����{{=�צ�L�h�#�D�j�p��
��3��8�|q�{滄F��ZG�C�����.)#��5�9�L�$��|f���&I(���ښY1Ԗ�x�	��g�B�������^�{�9�|�Z�-��I0 yU�NJ�g��T�z����cC�2��������2M}�7�[%Vmݍ�BP�%A���q��x���K�clY�����7

�f[k<�T�V�1۞��R��Lu�EI4Ji��I'`~ݚAػ=a���F�ڝ��x��Ӆ.���kw�J�Gt����U���7%�@�uʹ�ÂI�d=���j���'�:BGu�������Zvp�/���=C$�(�[~H}��'~��_D���$Ҹ��`8[��\���#�Hs*��xѭf����lH��gܽ�/��m�oB7R����k��Զ[�JX-���"�  I�ho�dP�;OUG�!=�����6�)l�#�+_ Y�}�{z´ 
׳��S��������x���,P�=�>�t�FuA��aMk��a�8�͂���wRu*���+:�c��	�Ñ�W��!��|�5lw5PF�'�~M��_^��qp�a�z"�s5�%��xa۸�C����bh�_�������^庲���x��Ӗ	����ɸ��6��nfE5eq�쾳v�C���8���P�X(���X�9JWl��-j�8G���[�cUV�y�y/�:�zF'�[r������sF!�劃��4��*?���2~�0��s�l����f�ߗF�i!q�7@2�ȴ��tL�[�XU�3`����W��t� q��;�ٻ�beu&4_���Qx�v�,~fs����
�L�yg����P�������f��b{߫��)���rU��R�۟��~�@�i2�bԡcQ0/#J4��XJ����L�]��E���-�~��@��tu��f����pz�tKV��Q�U�)��a�$�E�rP��E��<ȕ <G���W���w!�iINƣx�/
@]?f�HXMJ?�PmTq"n
*�7x4��~|�*Z�(dP��`�6hze\�����b�d��]ʈ+M��M�B��gٝ�~��^FiD|[BXie��I��U׻�S�q�_a�dS!|���X��=�m����\�M�k-d�e�����$P�Ą�	T�����с������u�����@f��A	9�a����l#��8v��m\>�8��2��3�bǓ�/%x���K3P�
�(w��HD��  ���A{l,���Cr�ΕG3�bF�"�}���K`��Ą"�`�Ǉl��p����\kU�t�~�#)P͎m&���7+��'�|��n�z��O�-O¬��}��FZ���Lfㅳ��߉���f��DqK����ogM�p��'�F�K��c+,
�wg��$|�����91��I2� �.^�\�O$
��Wt��oe���[ ?��].Kb_{�[.0)��`��0�J�fb��5]u..�Оl��z?r�[��y+b��$��V�� JD�c*ێ�<����|#�C-0���+�?6���ϔ|�P+�{����||{T�D� �x�G�m�n�n��YШ�^R�k$
U�����K�Kx�+���^���ώ�6�0q����e�ڌ�N$��p��O���L����c1pC�7p��;D~@ui1J�-��TJ�(Y�޵I����K��1<�(�w���Z�E�yc'p��N��Z�l��O��-��YV^@�9a
�NH�H	{R������R�����W0H������Į�!/�c�3N�>�b)/�֒�ݛ�L�ԭ�jNL^Y`FM;M" z�D�i,�)�F%�[r�|��oŷ+	:I��������]�*�7.#}�c۠[+�����a쩽�=;�v��ѥaP����L:�g���c6/�Ajݴ\kܮjնĳ�C ��X5Wh�T��E��L;ک
F7����'��NM�A?�r^f�g�
$�&��w ��5n;�a�2�$ҩ�Y"�-�)�CB�d�����*M�|Sv#��� �����A�:Uթ�
h���x׊�g(�~�'�*����x�l�):�����
.A4́�޹��#���:p!�+1���jN�'�Z������C����r���@��'L�������pJ:�<�e��{m�'�V]��4�7�}%�3]�����f#�i �oV�}�{����^b� y~�6l�B��P
icv���x���8��P�i҇��%륪,
�]�������Y��y��%���v���l��������?&����ΖU�->�A�N��J$�u���f������v)y���G��Jug�f*f��^!��陿���o.08�o�%(����l�n,���jPmv@�F��(-D�u22X�.�y�4��z|����D� �,�'D�9�E�h@%J	4r��1��䏮�1��0���/{���n���^�[�R����S4z�H�՝�Ѕ��󺯉ch���i�;�a�P�HU��P�z�M3�DJ��
����SVtN�dX"����e��\:���닼��H3���/R��a�ƥU��D�d�G M�c�/'[=H�V������e<1ۄ�,�m����ַ� &�=���P�C��9�:���ˬ��7Z�,U�GsJ���ҷ��|^�����1�JX��-3���:��sM4�A��_8�|��)���� K�t�>XD�T	�ߗ��`�����,lAR��c�X��-i�,����eڕ(����3n�@�-���\�v�<�[��n*h��2���[c �`
d�&R2̰�
I��z����,���<12p4ثY�ۓ�Rd>p�-�E6�,�i�:Ŵ�̠:y.�3-��)�>1/�8���,�)�/<9��$��r�6'���*n]9��|���=	6���a�չ\@�j��Q]||�4�����b������W	~�cު9���GQh8�.��������;NL@[�-�;�W��sFz�D17)9��i�#<e5�G78�#�s;-����	MPgU2�<���ܞA�u�D���y�:�N�
��/��i�Ќ�,���p�l��Vn�ǿ���8�V�H�1����n��n��N�[u��
�E��X�%�3��]}�4�MNc{K�}>�[_ň
�4.f����-e�����Ρ}x"S�����G�j����p��%���^��P����m`]JS[Jr���_�*�	��^�����@���5xA�����0�kK��~m�nn7��P:B*0E;D5��2��/���X A�+m�o�z�6��'G��Wk�����U5����-��� ��4�7�D�*v��ä��gO[�L�J�|�8�9�40�]8qȭuc^���5s�us��e�������m���5�K���E|�n�����Ȧ�֞�ī;rj���i����4O��ݚ�[�ZHZ�0k�ӎ��A��8fT�2iFv�#�C�!�;zq������p.�}JZ�t[
�	
���֝l#ɺ,�z�]Rd$ >��͆�]�g^��G��Ǯ��<� 초Λ��}�흻B�V#uL���t��F�[$	��j��Y:��"�Ɓ+;s�b�~��Ct��v���������Y����_u�F�6I��kL54b�1w>z�?��$J��t�z�����A�ϰ#^Ш���)�$���;�ڭ��-�L�db��]���^�/����\�()HǷU�4�B��B�5*��TV�F�Rw撙�.�2�f��SW05�MF\�@�%aה�	�������r=�6��m�USͯǠ�q� ��׸�54'�ϲ�bEJ\��BtI�j�/�1W���L�D6��mں���r1��C���^��F�I��<�q �ui�#�)B:.�e�P��( sm��A|�H���*��A���"��mQ������mR,��N#�	�9_i���ǟ���k��dդ��/C�� �n��3fSdOr	��|�����1e��Dռ��Ǣ���E(�ʡѶ��Å�U������e��gz���z�t�%FIt8����+0r�p���ql71��e���|v���U�5O�.��
ӻ��z��2=�K��s`�b�b�:�q�6<����:�����I���$�)N����|���R9�[�<o�Q���ͮ�e#e���r���BI��If'���RC?2���4��}P�F-w=�+}�,k�F�m�P��L#�7�SOE"f��0.Pz߰���x?��t�x^La���ˣ��*�x{��|_K`-����v���shJ�ߞ/X�T>\��k�UK����#��/Y��T��)�����uŤ���>Y'��'��{gv2Y���2��z=�(����$�e�:�O�Qk������/���r���p?] �t��M{�"�6�@�5x�YnC^��|��&X-�}�ߜʿV	R��p!��qi|���	�1]-�I��z�m�/6½t�cz����c�p5���=7ȅ��L�à����Fz�S���T�v�8�+z�3^�kا�����vj�rX:��R(�o�]&�?�Y�J�t�)���έB�� %��ڙa�)��Yo��B<-�;^\`����7(����޷���.���$����j=��ĕ́Dƥ�0v���[�Pe�⦈&Ν�v��`��U�-2��?�rz(Q�{yi�է�����ﵟ ���蘵�;�(���p5���+���Ā����� ��X�1/���vfd���;���ʢ�B�����Iҩ����׿&|�Ӗ�F�͝��i �؁F��z��~!r6��G*O��b�'ف�Ax���d�:��2�TbD��x/�PoG]g�awI k[���~��_j	�k��.�:��pP_�j�����`E;��f��auB�F��$��f��On��i<P��؜�l�{���
���sT//��X����lZ�fk�QNן�/�V�m�FGVN�Sf�]ft�ʭ�4$~>��l��[�9�-����q��c]*qҹf���ɫ־�#�(u�]`������rS��������&��m&���iK��
X�����*y'� 獗o�Q�'�-F?n4<h��f F,��ð!
����&��%�f�-P
���"2S�Ur�y��YohA��a�׹;M1�M�5��j;�u�LP����L)-�"�y�r��hJ`��Qj�υ�6�!E�N`�)^zs���`#%���w gͦ1�N7��< �)��43�Zx�nfp#a%�Qw��ET����#<�������H�������y,���y�>���S�l>��h�|���~�+ܼ$X *^�?���->PP�9�^���x/���^k�wѴ��Q�S��YzX\��Z7�Sto�a	B�_� ��Cr��^0M9��@s�cD?��|ٚ�R��\�DAmN��6������mxt�LQ����w�Ca����(�0��n��S�PT�}�W�KI=�%��*K�`�lg�ɹ�Pƃx`�	OV��l8��[3�O���!B���u���?��C���zh�Qo�\��;+Z�ϹG�z%S�t�v����ߓm3�����\v,�����y�+L�O[�j�yڽE�&��w�W��ו�#T��kz�x�긜l 󾝀��S9!AjZ�ޝ{��}<�B����VI��Y�wl&N�K;^Z-.�mF