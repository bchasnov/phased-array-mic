��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ��5���5dδ���KdXyݕ�2�j����B�}��AlU=w��m�C�}�S�[U ���c��6��u�������K���ֵZ$�<���?�ޒO 	��ȿk�Ƽ�o���n� �����4D�������;����l�{6d�0
�Z�^�^�2�;�D�
�UjR!�1�2>��Lb�`�D�l�W�?��9�J�ס�Y�u�kK$�ɓ�#�NA��Y�o�~8g�!'Q�Qd���1��+j�i��|Dσ:���x4����j���g��6��� n�벙s���c� v�f�GMcˎ�����0���6�R��$́r���E�^vq8g�O�jl\	��ч9ݢ���/�p-Zo;i�c�at��zb��M�պ@
�G{���CM��0Gm��w3���Q��ɛr�v�^7�<��cq��Z{ۙ��]l���gw��Eh��v|ۻ��&�xN�I��X�eъ�_�PB ��'%xRWh���e}��w��X�ə*J�Q7�j+#�1Q"���E/n3L�r�~��(>�,^�"O <r�b�?��cN2}�8��[�sA����+k2��\�8�YҐ	��~��@�D@�|��u	T�IU���|L��Ms���<��ˊ��U��F�5КkvП=5Ǩ���-�a���ow���I�@нr���\��.C��JxNV��IO�,�{�F�\��kR�[$t�c[��ܘ:^�� ߐ5��nV��m�H�p�m�:��y!o�k*y��P����P��U
���܂��BQ���,�O�/a������2B��1�f��oĜe7�拙���{� &���"�G1����E0Ja�>��񻺼�\�z�aA�=a��2Oq��VG��6�H���c�1��`^��uKr��Q�p�Fj>�ZJ.�~�:�4F�eV7�^�q��M�K�u�� FK�J�={��T�~�+��jΈ�
��u��P�k������}dY)G�'B ���$��J�jF��ke��O�p'��~Ѱ��U �&�h<`%0M��C"W�Ubj��Z��F��;z���Tf�.� �k�7�S��>��#0a��hѹ;����e|�c��ҫT�b��P.'���=��{I�������@�R�#i���l�Ť��zKB%^S�����M��� '��ؾQ�o�(��[{[zThQYۚ?jB��mS�|����R�?d?l� D��>�¬n8u�����]̬��#��B�|'�"�H�.e� 1[h��e���V�
��7�<���z�E�w]�Pedn�k'	��w]��0R�ҌN&@Wg���B���.���9�[.��������FSvS�xz�W�4�}���^��7)
���d��|���}�J1�I
���g{4�}p5���n=!�p�?��1�#�|� v	���P�!2w�8C�8�Y ɓ�h�⠂����!kQ|�AF@�
�$���L̚i�H����S��Db��h���[�u�/Gulc)_�`��"��F*��V_<�����S�d����/H��
(�d�l̥��3�s�����	�9>3/�O,(#j��sҚw:X#��Z�TG���ؙh�����A(v���N��哿$$ �%d9j�ST�凲wjӌ�T�gl�\�93۸S.:��9��B�Pa\��bc�~��ί�J�/�X��C��}�)�ŕ���VB�,k=
+7A�CI�ť��H��h�A�-��!���z���J����7��I���[4�UڜG\yM��+vW��k��t)���XKڴK��4���=�m��|��,��
^����d�t�Ǌ�����	N�੶'�X�	�h%*��;?2�-Ш��ޔz� �$K���R��ϧ8�<�>x���?���FIZ��y�(;�	�?|*=H&�m�]��(��E�w�T�9�h���Q�6���p����#�P�i0�ld(q#� �]{�">����P��WV#�ә������Wb��E��3U���^m��#8A[�<=�$�\
	����tCH!e��~��u����=[�&DJ?VDK�e�V��jJ��ւ}9��7/�	���ү@rz��dP������-����cq����-��Z����z�K'�?E��[[�A�<�$����7�p��DW{�6k�ĤC�.4�����D�=g��n<��'����&5$CW�� �Ѳ��n�^-���������FV'M�~�	��vy���E��W�8�;���P��+����������=����a<mwԗ�m�8h8��c�Ƿ��v���s�.�kB�ķ��ig�"���L5-�ɣ���gHTu:�[��`�d��^��A�k<B�һ���VH���y��El)_�@
�ͺ�`I#*��>�:�(�2 4{ �J�Z����?R�����
G�� �P$��>�AHz�m���L��* �fl�{���5oJq��k(u�ه~}�����I��?�Չ@]|̓��!o_�dp�;ٜ����&H?��ʠ�$xD�G��WtO.Lh1���r����t��<��vY�FӈHd	�Q�>�DKR`[�o��f[����%b��6T(���tz������s"��7�=�������W��GR���6!�9�:��W�F]]��Z���W�Vh����}MTm��T���Iq%f�QP�F��O�9p�5od7#B괪~ڠ6|�e�'��E��7ް7K�J��3�|+�ǁ8:��� �\ا�1�:<4��e��s��rW�Ii����&���^�m��_������+qvwq_���C�#��8�	�ry�5/Ľm�`B��+&O��b�y�wQ��]�wzUԸ��U�ˍuM��y�0����{��AB�j��N��cR�@���]�d	�a��p�D����������K�>�������M�>����o����&[�/���Rq�{r�$���9���9�n�ƅ�fR:M��� t)_�E7C��O�y��-�[�gw��11��FӍ�\�S
KZB�]1͔U