��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|ḱ	I*�ɤ�i>W�WrƬ��/���>��|���e�Ν*�,��<����߆4���;NF�.֟q�G��s:e+����I���2X� ܓ�e	A(�o�W8ٰ�����}?ҷk탹V��5�Q�����|;���>���l).�!�IQ_�C�)?�?n.�;D�a�IA}j�*�>Th��+���剜s~��:`8m�J�e+%��r�4��C4v�����&��:fr�=��l�ܝ���K�3��Or;�x0�|gNt;��Aѫ���%엿j���뾚7����5�=�5 ��m7�Aƨ8�)sM�ڔ8����iRlZ�B�B��_�y��<kJAz$+�2���e��	�F�:XmBb@S�h+m��Ǜ7?9�ax�/W��jn����y���嬌)N�/�{t��{:ǽa��x�
�Ѯ ��X���)үJ���kt�H����@����7�y<I-���u�f� V~�2�����[���%�������jd��(�CC�P�Y�m��*[� V��Bm�C���.�\��f�T.�x��u�J�	���܌��P�_�#Ԡ)?��L���S\�i�u�DPя1S��<����<v(ȍOKc�>E4P,��Qw@s�u��*�3G�GBT���
�L��;o�JN��ݯ��$X����Nd�[o���Þ�Y�A���.3�d^q��"�mD�����M=���GQ�"�_âe� Z�B2���u8�� G, #��̳d���_�g��S�����"�Ж('I@)�:L4Uy!��p�ǘ����>�~��Z�9�ۀ��E��7fy(7����f�i	��5�`&P����bJ��P�'|��|m���E4؁h	A�>"�;a�MPS���>�>��G���go�
�i�}M����μO�&�`Zނ��jbA�h*.,Rm�(rs&�浖��I&�	��m�$l-��6;M��m�1��^nc�'�`���f̩����/���Tj����j�v3D�l�_��Ƨ����P��/���Z��j1Y8%�Nw�j*��z�U:���|b�ٙn��avθ9
"�$C�Cr�~�:j�o�F�+ui2Ց/����5jėz�L8iy��Y�iW?�K�ԨKv��7�&`2�W�`���P����R�u�{�<�i�@5��'4��R�ӫO����^�bh9io�~��}�4H����qUSS���.���!gR/�E���1, �]ףs�ЄH����גOlB�+��O'kP:b�Ua�[&S���|��'/�缂G35�zM�~H���h��E���2�H�
%���ڍ?S����ꞙ�ɇC��)�6������sj�	��\"��^�w��FW�}�P�D�9퇫_w��� :L6��ٱזR��"�(�����c��]=���82�X��MǠ�� �<�)}v����4�\�a0(/��b�]_����'$��D�w������}�d_���ԁb_'٦(aY����%��`i�b�يyv2a�������F��{�cT>����7����bm��dw��_���$+�����r��u�J�V�@1������`(4�x4td�/��%ua�-��(N!�D��f�����饜nP*�o�ԅoA�p��%C% �k�}�<I��8�+�{$�j��":᪢{�h�3ϩ�u�3�{�{�$���8�=��&��gS��ȭ��<��sѷ�1Wn[Ć��G�#&��.�[�"$ӓN8A�TyEGA���,�\O��j���]r�-F�2��4��}��qA"a���Qx��g��LAx�D����dT��/O�
�[���F�$�Q0l�a[Hٵ�-��L�QQ�d Ϡ�{A���'�`�T|4�X��֕D⧆Yl=���,�M�*1A�>��)o�<A�Fy�ʧ�vڥsx��ɕ����	��&��ٗ1E�= �\��%s;זWy��~)�X�}�y]��[�� W�]�\�{	J���d���~�X�8���������v�|�
^]��� �yb�$9����g�.�~�3<p�V�C���r���9M�GG��� S�<Q))�àƻڎl���p�<Z��'��|m�I�_#�J�0�k?f��oP�������;�Ǉ�ع��.ᩝ�xfjQ!���_k����l��.�ņ]¾�M:S|ѳ#��Vu
2�+��F��Nbt��o�cwZ��.O�2w���,d �y4;֏L�+|&o�ƊY71ü�4]�WH��� ���$4�Yz�&%�KQ��. i.q��"Ѽ��v�^d����K�ǐ�y�}'˜�W���3�WX�AK-�ҍn������Ҕ��0�C��1�:�ymw�m�C�p�i�`�+J�O�U��#������9rh�e@va'A�:�qg��?%ڐdL�3�����)Nj�$��խsCwݽvU�� S�n_��$f�zN�?�hl|J�C�y�0�/�N9�!#�U@:�J�m%V��!�?V�٪�]�=�t&{ι�a�}��kE#���F�+�3����%S8$�<�RF	����m,��,jl�b��O"��fx5�/32��TP!�}��#ĵ+��9ʹ����@���!�s�]hßF�����z=�6�+N�oo���z
�����	�#ړ�v�J�	��'�%P�aҕg�l��N�GnT�bL����\����p
���F���JV�[���o��K ��~�����UI��-t��3B���}f�W`�te��?������Ԙp��>�.�+NJDݔMrs�����t�_3�9y|�Zt��)�25>����WP.�!��;mvX �	ث��8]<�1�m�9ި��
#ײ�H��33�S�|U�K��z�k���H��㤒ņv,m������qtT�>�5�(V1,pY��콹W�1���Y�"�/����l��;"띆t��u�:pm�w2��7���>���&Kl�0��O�P�%�sk��;O����ʥ6�g.&|����3��L�J����b�Oo9�-h��q&�8�&Uc����
�O��q�R7�
#c�CF�%�k�f}�;wQ�D��#-��a
�J��6ӟ��1�޴��ˡ��:�AWw=	g�6K<���{��B�,��w�� ��R�������f�ݖeB}��P���d�c�zJa-_
�5�������f�qPX��#E%�"N��,�AX���h�;�*�>,���BfP�߇��=��0!A����V��i�4��9X�
�_+q)��Fk�	J�"V���(��W*�l�TD!~��9p�����-�:�W��@��b��N��2�snu�x���A�RWOJ�A��*�pc��n�{ģ��vaV��@үߞhi;ZP�L藟p�^��:�/��xA�Q?).<u���2�*u�,�R�I��Ӏ<뷌jySq�q#U�2ͬ�:��[�l��N8*/ӎ��w�O �kC��<R���"Zn)��d�4�6S ���i6M	���s�
Cc��!���&��	!��A;�<��D���&`xDV�[~� f��0h������va�y�����m���Z�P4Q�;Ks�x��Lkp+�i��I2����֟��Kj�`%�?�zi�U|*��1�1�C8՟��=8�6��_6��)��܋�FB�N����D�T�qtqX��h<�����8��(������z_$>o.=�7�`#��%�Ni��X zQ�W$Bi2]�B���`��y:�]uv��K]+J"��!�Yp���ҜK,�\{� 9�ލ��ƈ�@�S,���"f/��a�Aՙ�������q<3�;5;>��)}o�S,���s�J��G���v�n��� ���H�c�NNq+$<��e�Gq��O=���m��e+T(cf ��������zsg��,���Sk�ך�X�]�)��7 ����1� ���p�`/w,mHn�_��
5������Dg �1:V��8i�_~g�� �)��VdRK�z �3�g�@�
��aC|�c����=%�� ���VAPR�e߳�dQ���]��s;���}��l�'�
W7�-���<�]�y7n����pݾsb�@������(�^�����6��q�L�T�	�{9Ce��T5=�g��bw�>�-iS�ѫo0=�_�w��8@���n��ˊ�`V�҆���gڏ+q�MS�z��yiie��5ίrt#�������5��L�8�G?������m3"�j�)��Q�J�`��ZlTZ�-��ǡ�T��u�	�}�B�O"r�*=�bYtk<0��X�\�+f@���l���fEP2��� ��������oJ��g����v]��hi�?�F�̈́	�8�3�-���rb�K�_'Җ*��sJ�J[mJ�j��[��`������p����OP�����:�D�G�k�
�)���-t��(���W�{xϨK(���DG�B�
{`�mz� ��«��f\t����x�m�0���4���e��gk�"�lF���l���ڔ�慏CAWR:%�js�X}��v�P��ʞ��|~��I�z���r����=-\�.�]9��4��ꌳ����~i��N�%7��F&��z�S�"�)�ɵ*u*���@��NP������CֱT�~�#v�&�ק�e��N	�ȐJ`���rJ��an�`o�n)N<E�-��D��z�|�ˮ�Ɗ�b�x����u�jLM�Ѷ�
�ZJ&?�:>d�nw��ߜ�2N�2F��Ԕ���i����xa��q�� rx)°��5�<�Gcc��o�)������R��3X�v��aOxNr /Sln�׊�I�iZ��dU({=��H%���ݙ !�F���l���L��E2d��T�
Lې|��H�{��F'E��U�DNc���'̻�'<�?��p`b��'�����Tu.4�$�|�t��-��a��[&c=��6�_�-+PwXh�PiA$8��������t�E6��h��'#����S��vV1���w�7��8lDT)-��	  :r�>���"���np��������^�4�E���5^&�����l���O���0Z���n�$ч�/Z�J��H�.8��p�kնK�֤���0�����L0��b�Z!�dW5���h7�r-�$,D�����d����r����������w4�1���FK8�Ğ��R����Ǌ���s$^$�VS9ƞ���W��%��{�;/�����q)�or_�Y���0��q�Z1����sB�gP��A/m8]Ǣ�1C'�Z��7�n
)�1��"a<��D��# =B�#���$�+{a��η`��|�Z����x�.0[�b	����I�������A����Q4MF �2�������Z����.W��9��8�X\cG����[o6�_���e�����p�e�
	��?&[��jQ�4җ!x��	�{ �i�~C��QJ�K���Jx[����z.��%š��'�O*�?q�a�P�:?@���cRX���ZI�ހ�<��]Ͷ����3�g91.�$>��k+V="7~xOC�����]¾��m�eh6r�����8��߉��y;¾�D?K�n�C��e&�������Īi�^Yɵj!����c"r��(��W�4���eϨ8��u?gh�b=DS3=����w��78�VT��/���*.U�6%D�{)�
���7�k��(5 ��x6v�%�%Ӱ��L��� eɆ�u҄���ug5���)JMwɝL*������d ~�?"o �Hq��oa[[�obU>
�}-�?d���q�\�h�t�n����U�呏�h*��CP��>��R1֎���z���G��}��ǰ��D����R~Z��h��=�Z��.ϫK�t�ʽ����_��/U{m�������Y��������$�@y�Ą��R~���I때����B�ض���:+ �"�&ƺ�����=#�/��/���^���P�5��'M��v&�w'����,�Hh���U�7n��{�܋�ۼ82�����w�F��g H�����
Pe�ܼX��^I�q�|j��sĪ�]t�17��#��n[,SV�7���uED+�w����t�܉*+�*�Mg/�Ӛ����6h�e�-j��ٌ��������9�q��A��-]U;���QF�C�&X���(�X��]�W�9�)h��
K@��xd����]���]���ѧ��D��%����`Mo�L���K��'�x�J�JT!@���&�k%1a���y�G�Fÿ!�ѥ��3��0��MѮw'���y"=��Z@`���;Ns��6���3�iEo1�lk�*��AI1�|y�f$0lY�]�t���~�f%<��͸��DhkKrZ˧d����=�E�j�RM�|��-�Y:�	ܔ�Ğ&9k�ؐ�{�eJA�`a@����|��aV�
���U#�/{���3J��ɿu�ϥs�1��(�)�)^%����^1o�ق��x�4��|h�\��i[�O�}�Q��Lns�JG����r���s��	6k]�@���}E1���@�:��腻,0���=_\{�_��M�E��o�is�4�&>yي"o�0/#�R�u>�9Y/�YE�<~^�#�>zuӆ�t�\��Q*���"����<��Z�U��jS�Y��C��N���F=n�B|��l�1g���V���e�.��]��-�g�	#��tn`��l1�'3��{/�n�]����1t�o�td����W��rp�U!���ܦɚ��Z��{bЊ��#`]jo��3��hD�N��c��=���E�� �c	�X�}���" ypR䎊��܆�V��Bފ�A�+�??�7gا��d����]���$s��A���h.���/ƃ�2��Ǽ���P�~�y��W�2Hw�JB՜���>��!��%�<F�?�D�=���쥧��EI4�\�e�����m���%޲�	���2�V'��OAm�;l�� ��+��ĚdqMO_�
nV�-"�b'�v%~Fy��R�L�]r���r��̑�A"\��p"|38�lի�4}qR*�u�y��V�&M��a�%�/�	���h��̎K�Dȼ���i_Ӫ�� _���O�S^p���?R�Mba�Ṽ)%W%�h� g�*�	��3ָ[8:��x����}��l�G��!pv��17OA�n)��&�{��ϐX� ��@���e$b��� D����(�Rf ���+�� ~�����H���G�)3�Q�WW#�%��+u��O'��x�x��K����׳�}USueeO]���������8��vA���f!���b������Q����-]w��P�
�iVy]�Q@�7SH���^�cp�9!�}���A�������:�������|Y=�L���Z��C���{��[.*��<CO<M5�k��T�-�;�k��x���7�tΟ%��0�s�
	ۛ՟��!I+'7���G��ܵ+�M�>�S���8d���Y������V�-�k:܌?��^�[]/���c�9��?�V����E�.��K�h�CF
\�aގR�B��(1���Z��վ��Q���^��D7(����w��R"��t�i�������Š�p2��^�P5�X�B��=�'na����vhd
�!��?[ܝ�5/�,
�m�6�e��w?.�ײG�4��e#*����S�y�E<�r\��8 �[K�W!Hl�O&4�X�햺S����%�x�}ꬻ~�;LM���`[��f<�ͣ�q��Q�����!�v�3�,��v�K���`���&ߔ��o�2�I�q�o��R�0b�L;)1��!)�+w�Wl�}��j��X�(���Mf�-3�$�3�n����'\��JGV�'��ƨ~!b<M$��Uk��O��� 
O�ܑ�xK���M~܁�SD���	�}`�S U'j���j*T��Q�|�n2�𰺓2h9�֐l��OI���߱>�?�A�2b�B/E`���QqdB׈h����nb~��%�{� ��Е�3�)���[�6��x��IS�5H�D�~�ԝ��Jb��@;u���]���6|A�]Ti1M�ԣ�`V)���z��Ǘ�yU�?1v�FcXY��y �d���R��{	LY�H���L�̮]��pM�&���-��)5&.~�)%Ljs����-���qp�?�1���c>�^[��� ��H#h�o>;�/�~5$�b4N��	Ʌ�C0Y��$Px�P���O���/�K8��X�K�SE(^�Sk�<�l�i}�q1А�ed�[7����~��D$�{G
0���6-z$ݎ���?���W����'[J�R�^i̊���Qy���߷�0��L>�̑	 �;M�
�%	��taF��腽�Oqt�q�f���2��ּ��h��f_����u�FX
ǳ_��1���d�t�*:�]o��~��&�As͢��� b\�MNzBJ0��
�F~i"إ�i���=�������{�xۛ �����8H�w��T���j2��O��nY�R�/����5�/UZ��Wi����'Y��(���ڣ�C��~(̹��m�� �K�u�s.5ם8ѽ��Dݻ�C�:rT�T�:�L]����x��IV*���;�]�����"��>��l��@p~�<_pU��^li5�Qa�6���@}��~��j�����)�j&^���~Y�I������M�j�T�+$*�Z^��[J�ې��E�d8��4T*n�J=2qh)�^�l�����4Է[��p��/	�H�MS}P�/�{�'�8�1��"�*��P80;�x��n�F��$w�{�IV�>�Y�t�2�;���Uϧu*�J9� #�r�Ӹ��s2�jV:�K��(��T�%�"1����p~hF�~V�5ۭS��h��VK}��C���:E�3�ɒ.#M�IB1��
�!���g(�9���G��{a+棚�U�JR2���ʳ+��e�Ǐ6,Y9
n��LL�	p�-m�U>ht���b 95�^!Ű���mx�}���n&Q���xut�ǡ��:��<Z�Q��7�!55{��������]!16��k4,j0Y��,J�V�J��V�SKm��Y4����2o�)qo��F��_K=[�2���Wwu�d�i߻�;�g�ӓ6�r����*�b@6m��xܺ��oY� &��R��%�)�I��]5�xc7
��U�!��*kz}�.�f�x}�_�R+����Wy�v^����'�����:ΔAj1Ư�K�GP������4�(�B�2��y����Xh�~5���gu���KΔ�E�*��T���3X�V˻I�l���sb�;d�z1��Y�!�o��"�&�9����<��C�a!v�W@�a|p�[:��1O}S9Y;=_4�5�T��C�
��^�/��^7T���=Ih WO�4�cT/�+(	��\����_Լ?�� W��镧�=Z�P�~k��~5�<C�@����(W��!�d12#j�FH�u�2[&O��1X��lbw�@z�?`�͗#+&���f�	I~Y�n��2��Qˁ֬��'P��U^�G=.�U���pՔwOj:�4,Z%'�'����#IZ� J_�HrwL����p{Ф�Y�w��u2���M�ś����)W}��eHJ<���qV�yK����,�E�=�d�
;�u�\�������!��3���n�>�@��vp��	CO��3]��4*U�b� O�������mɂ(4�`M�zv��z8���6�)�Ƣ}�B��d.�!�\�6�f
V����s#<����KI����
Y��P����M�B4�o<ʩ)7�)�G��U���0����-q������v4�?�Ee�1q���מW*�X1ԛ����'�p�K6K��T7�����\T-����?'k���g�;k�]�7=�/�0�����c��pc�>9i���A��)�+�!ib�h�}	�7�z*���Z��V���{��K�Q�&��;��?":���j^��8�tcI��9�?>D~�����4޳���\չz9*a$2���{�7zLVrBޯ	���nO�	���9 r�8�dH���ľ���/ ��"�	]���F"I�_���*78�9��s��g$�4Y �1a���:�+J�g,�S��l�	���l���>���a�#'ȥy�2�����Dږz�M��r�-n{��GzO��Z��+j�2���<0
j�l ��X{�EQ����(�ۭ���-u&Y��d"u�V ��d3~I���H�_��q�U׉�u�&�׭�#
0��~j>����+0���U��󞼍����U8Pm^����Hv�%�� {����M�f��a�^W➏䆼P�6��;�M}@}�����L/i(��t�O��(���aCAM�A�>��)ûPܲg1���J�<�]�${��O�����bɩ�n��2�1����k��P��r��F���%/�Q
@?�%?�ͱ��Ӛ�S1��:*g�lB�F��y����hP��`�G��P-����@d�=���~�M�ǹp��z;Mz�������҅���T����&~R��f���G63���1!@�UU���A��^8�{bߋUyS�M9)Q�7�G��T,�b��J�BbJYSK"k��ʊ�-�$O�_N�%>�S��~�7�tK3p���p$Y�dא�{:>�ʏ%#�sʦ���:��'�� :*|ț�X'7y����($:.V"��0��D��m�?I��<��-Mf)��̐]~EW9_����$�����Q�[�<�#���B��<�N���Fʃ����3Ǜ��}��#��FV�Qeì#.��长[���v:U�p�
v�&X��<cK�J3,�����G�����[�y�O���7�(�f��{Y�|zHK��	x��ܔH�!�eA&d�ϱ7����y�6� �`�� �@�ز2b	k�9�ê�j2d80���0�j�Og��=�T�Bm�)q�Ș��Q��E�x����Un���7�LwƔi�l�N}}�4Ӣ9�> �Q��H���Ӻ2�?6���< t�>F��;m�y�ʭ�����s-�����Ɇ�MV�y<3��W��}F�j�d�,F��$��4AL.����q%�g1��b�.�����sBc�
[i�"Sp|MWzR�W�2���M�d5�g\U?�6���I_b���;Ɯ���^-	���T�r6ڱv4��#Ӿ��}���Ԥ�&���P��j?��y�c_i�������3�ǣ�����˝��oH��M�]�U�<�l�Ɩ�'����?���Ak��d,���Z�\��Bk+t�n�����`����������A���qK�i#d���#
0y�=w�<�*��?й�DBk3rk+�Qk\K(6�VEI�j<|С��� l�����i�ۂ�z�h4�i7A:R3��6޷����N`����L� �]����w!�@�AK_sZ�9�&��T*�3��"C�.�{��N�d�Yq���[�G�W�IŲS���b�Y��'©!��`fY'��^�E#2����D���.����g�#eY�p�<qG���`��J���h�Rޫ�X�Ap�$�[m@>�&0����7�TZ5����ڒl-�p�cxmy3%���CY����yֲ�p�MH�3�w����:�]{,t���P�Β���K�X�?��IvR��fg��U��C辏��iO%�D����/�J�O���wz�+�ϩ��Zp��Y(}�[h �������١�{F܆��Wj��	�`Z-�\��.����3�"M*��6���y/��y�OG�"g%����J�|+�BĚҤwA�VO"}m{$8<|F�yf^E�.#�ی�q��V /�6'�ڱ���?t�I�[\�٦��S���_]K@����8Bf<J�����4��x�s����_�M����F�+��x'k}nU���f�Om��Yk.E�2@:�9�q$ű�٭���>�{�Z�8���i0���7:?m�`�+��@/������[y�����|T�⮈r�N]S�K�C����/�Y�o�V��m���dxK
q$W?�dI)͔�X��u��sw�ח�� �����⾤|kl����Ϝ��5�����ȆҚ�Y�p+S5"�$�o�3g���+�bu�pi���A�&1w݂냛c��Ve2�B�A�	� `/�7S7���AS�}�$���� �"����Hw�ڤq��p=j�5R�t2����%?�k�i�RQ���������e%���f��%0<�A��}�T�Ӗd���݉#�4'��K%��gπ�9��%Էh���E`�7,���P\�[gf$� ���!�
F�ӟ����¦��׳��v����`����:.����j��T����E�(�Fa]�l���t);�#C#��Ei��]�ӡ���!�.�x��>��=�h�&ls��������N~U�%@R����H�`�0cL��u�c�A��xJ$.0׷8p�kX�$��D�M֮^GL���0|��^;C�P�U�-�3pԪ�|
�B�����/l�Js+ĿE"'d�|��mj�Lg+��8�@+|���V	��^�4q���cPs��L�o�!r� ����m ޜ(r�$DU���-��
B���$1Ϊ6��*�f�����r�J�8_�U��B��Msu��ʲʩX��6�-��>=���5I�۩�0ӣ�z����Ɍw��vƑ�p�zV�
G	a����A-�L���;Lo�P���4֯Y9m,xKX�4������A�(Zc5�u���C��w#�P�t7���z&��ܪ�y��GN�n�?ix�C�mG��C}���M,]�'k+�-WvU�x�R�F���!K1?��������2��5o�l%�l����^M� ��G��ҽ����1E��w�+�B�hƲj몟4��/~9 |X�IM�R��s��^��~͝�����$���U�W�����w����-H�B��P���'��˻'V��O�!(�c�Pg�b�GH ��&���-z�PcBٌ�䑁�vBn�_�K��C�N�iϒ���ƣ�%E�Y��/?;�.��ZD�RVj���fS���tz*�>΅�C�P8=`�ۆ�IK��4��M�;�5;�y��_�T�	ַ��CIwgL�����w���0����ֿ�CV~��%����(s�Q	i��2��&�5��G	��n�{��ŇL)��j����s�e���2
4	����ꒃ��/~y�Xԩ� � ��2t�Ne����3�k�H���E�����C�!x�kA+�bsy�2V��	-���p��m.�ҫ3��d�<B����K�f������SR|��(��!ɒ�oAs~���}�u��i��'���)�������#�ɋ��"��zv��҉Hן��݇l�Y�JͷE9r�]���+(��==���FKƌ'��4�""��9�	�zG�K���x��y�E���B�Z���/� �O���wWH�����X(����kAA��������ĝl\��ۘ����fɝl�|Μ�����>݉kvȆ��_$�>�f���ˌ���P�0��a;#�I`���y�i�	�v�$1ȵE/"mu�	�@�g��*B/�Y�#���� u8�rz��rrV��D������A<��-b�
<G~���g��t�	7�a/�WI�`?U*n%���zI�$obWR��
��R�V�Y��k����zrV�f@L�
�&zl��q�-�0��JV��s�Pc�R�$1O �J����I�"�3�	y�6���)�k]��x,	弭�f�����y���6���|���*1E�3����L���=�J>�h����Icg0g	H-"d��5�W�� |��8��Q;��8R�������v�mj��䱩�93H6-J{tsVk��;K&�f�}��ڿM������ϰێHH.�cE�(B��]K��"Ӵ�8�^�K���9ZN=?( -B���zJ'Cۜo��+�����n�u~��X��^	�8��8/h�n�� ��[���Y*����2],�����VK�1��+�@�g�~�QvR�iF�L@����	�S�a��5�A�%S@S�4Rz*�+0�����_��h�(����Cz�"�,�|>��;�I7	�ˤtf�����͹.�Ya���⛥�;Le�/ۊx��a�"���=���қ�c%�A���tY"�#.���,���8&N���%6mtB�s
�%�m��m���h�R�o8A��6��y2'q?�'��$	��~$u�����B{�t�40EN����M�� � W��G��P֏!��cX��_�S
���i�]�J9��^`���� b@*Je��&3K�Ϝ���t�a��� b(/�j�;Ap�'�g߻M �Ɛ�_i"=�YSb��vְ�G5�2Mϼ��"��>��!�3�l��<݋ڼ���1�Ϸ�؎U�Mۄ��#Y��1�,3��J���2A�[[���g��j�����"�Q�Ф���T޹�q�fr���FK��%V�����Ae^���<���6���:FG�,{IYԢo2��댐g��b$-a_f]7;�>�<mǪh��L��l�4��*��j�d�e+�U�
�
�DD��Ioҙ�+:�aJ���������pѪ��<ϻ��u$+��_U�>�JH_#�|��\�:�1t,7���O��g"L��gWK�J�?���1T��&Eb�q�H�cO_�Pn+ݕi$���\��I7q��3�_�5N��+�]�.�x>�x��d�z�d �"�� �K����B�E>V,F��o5�Km�#�W6$�u�RxiY�Ѕ�������1)���[~�Ds�JSG�[0v�r�s�m:9N�A�ֺc
#�Uʺ��1�#��`b�#6��P��סޛ��Tx���,s���'R.�kiU�j k���S���<��Sf��p��BiX8��u_rY'9�}��%S
�/���qkM:�P^��/���'xG}�)i+�Ɩ7BD�܂���H�PZ�Qw �eX5	���<*�����Y��[eZ�A�&�|��Y�z�=-���a����E��ވ0��՗{s+��X�s� ���B��e��6�?�cot>4�.�w����SCD	�C����7�Γ�1)~�d��$�C�R���b^Wy���5?}h��&��І�u��mr-�Dd)����)��\�;����=7�q;��GD�-�q}��j��c�_��R���]+�C6Q��_��F�U�f;טۨ95��ru,1S�ch��J�g-5#'N*�uw�f�t&ч�ھ�r��3~�^0�_P���P���a�O����
���,�5�&]֮���0u�K���Ŵ�� #S8���,��0m/#>� �.ʧ��s�L��a��܈��L�-�Z?M��[(\�Q&�*g�b��e�E�{�S�"���z'�.��ei���yH���	l���
�Q^2�ux�hwhJ�\��l�ؐu*��J��T��VZ�!`���6���T��V�:�ک���u�(kRL*��CC��@�Xd��}�k

�	~�g����q�g8��z)&����8�*�VV\c�U\��;��$�B˙ �� t2��3���PJi	L�V�.@|��G��w0>����<���R�O���R��·���N��]<�I����b�p����J�M��tP�]���dI�/b�T�v*%�c���*�|Zg�F�[o���'���r�V��N��0f`�*H\p�E�T��`ǃ|��~�$��)�5p���jb�J�RX6t�f`���t@?��B/ת�Y9�&�J�tK�C�x�h�}��e8j���5R�ʲZ)��W�gxv�i\޼U��5ᛣ��Q�JV\<J���4,�w��p�w�X��F�\���h�C	�����S��byw��}�M�Պd�d�)_e���֒E� �߸pK*5�$p͆�1��xV�"��%P�6�M�V\}�?g�_�徽���WP���g�%�
��	[�M���}�l��=�m�;��xK��"��@5�x%��V�0'k��Oa�W�;��Wx�Y=�PD\���^�=eND!�l�7�+���y�,�i�B&0�/"����V���n��4��B}�ɇb�N��hA�-08�u�
�� Ѹ;q�eh��R�rdߩ��j�kQ̏�#��q�J��M�wq�gne�t��X��|��W�.h���t_d˱�Li�^���f�J�r�1��c�$��� \���X���b�A���]��}����x~���L~gdz(5n�^2Uq	H[m����c���G��#�eţ�<q���s����%�Oz+�x����ҙ52�ˏ���+XYWl9u��
��^�t�� U&b5r��H{F�,���H�^F{�u�j��S2�ui$A.�D��a��m9g(H`��tQ��\!���ݳC��92���&o�,�"�_)q�`��R�:/�,=[�sr6�!�}�0g��g��Ņ�,�^s��8�JΖ�����=�q��w]O��zc]ܹU�O23@,Bf�V8��7�x<`�i/7�A���6�^��%C1Qh>�O�~�_�� ���=_������[]V��S+� 8ҏۛ���t�T#�6{�#�����9���E*�1)&C���� q�y�����?�μ�G4D���ϫZmF�8LT;��a��*Z�)}^蕜����dJ���ө���d��ܱ��ڝ�"y�% ���
�63��'���i�m}�1n}����;λ����Ӵ�F�����HD=�Y�}�i3R2���/H%̇���j�:�Gs{g}�Jʘ���	!侫#s�ܨ�I�Ď�#�%����R��$Ծ�q-�.?Һ�_Y�]8i}�R)I��.1�G��#o�6���]PԬ��Z�	�<��#rg(�7���Qu�	�$p��@�Hst;*�����E��E]�9Ţz$".���^������o�u���l!��,�%�!/cF��5Y6ȷ����Ww�:�*f!%��Dy�7�}eKf��y�W���8�U�.q��	�������o��J�,-AS�����x�!A���$���ܐ\A�5��ӊxz�-wa:Sú�U$&�V8�h�<B��/0��LP��U�5���k��N[
w�9�h��m��W����r�S����fvΊ�e���))]%]����'I���� *������=�8�W-W|ǋ��v�'�UC�J�YU_�J��'d�+��!�k��W7}_��'�?�+�Sn�O�x�7f9
$:
�9�����	�����^)dT7�һ�6�ጝ��T���A�jrO(���5�UZ,�h���c�;��������;�(W��?_�X�8.�Ɨ~ז�[�1�yti&8�f�E�R>�����	@� �8���{c�Za�!�޳����1E]�7��_�>2���6WX@�����V�nx�&wO
�y��Y�g?��٨�,�˜4����lٿ�>������M�|l�o�mߍo��L�ڲ�� Z�Lz��r��b�x����xnT� ���pԿD��*^�JP�3�����)Jn#n*��r������8�%�_Q.�o0��oǣ]�z��x|�O4�����uh.����A2�w�� ��n��/4%�q�}Oe�|u�(��з����!Œ�ʦC	���(Tf����ԇ�L�} %�W�wQb
�lZ���GZvOgE�{���G�B7y�{���Q2W���J����������F�XP�$ƧHƃ?�.��%@1��,_⪛�J8h�	�ʺ�Gϩ���|I��<8k��'�N�o���ux���"����g68���1z|Yj�0��~��L���a�5��U��+��0�\�}��Q�3�@��Q���Y����R���z0rF�Ҷ�]�j�i=?��OFS�I�,_р�c��q�h{jN��ِ��-���!e�Cy Kv�U��J��U��ˊ��IӒ*�ؓ����)-��i���D��1���O&򶾷�6׬:��I�+LfM�lԜzr��J���	�v��<�wX�,ge�%��.�\w�>S��``s=4�]S����?��	��Q)����׃�t;�`���R��X�L'sX�<�VOqA�ruC���1�{%��Qw�`n�B�O�·�$o+���Y�f�x�M�^�1���Q�\!����$/�:*�eR���˔W�&\��u1���Ԗc��y&�\�l5�.,L��-k�g2d�7z9O,ӊ�X9��c�)13K�~��Ơ��Z��h:�� �1�T�
��X���\5�v�m�ᙏR)zɩf2�\�p�v$����6��;�@<���HQ�y{�z��W� �j�n��4���{'ջ��>%<�V�]����U����^�����-u)��i�+V۳�^1�c��y��y�#����8��da��'�L�\Eg?��{�P�����'(aXdKAĜ~`G��ڔ�����F}��t
�Nz�r��mgDU�~��/���e�5}�^Tp:���J���̄_j��P��6U4���ns�'71�J+/&B�9w?&YY6�VG�Ի�}aQ�0!>Kk����U�G�ĭ�8��kH�Od�?L�8%e+y6�gs0~��8���E#�u^*�͹;;	�PL~���!�%p��8LLQ?�C�4����%�;m��r�<�{^̌{��\L�<��o[�ȍ��~�V�'�9�C�zC������b�@�x�.{��zk�u���r^r�}m�B������3�nV �
oj5��FMk,o
;y��vrw��I�<6�� ��(	'��ׁ٪�-?�?k�:�g������Gb;�q6�l��p�^x�� �����R�Y�|��Y��K�G����1�F��ҫ>��JN��6���Nb�>�N��N����c�Jl,Gx/�j���T�l�f�/��.%����W�!����Z-�g�9�4E��t�����kK̫�C5'l^�D5��47/��Ĉzjfr��d����ā�H�S���H�q�Io��^A}fE������5�����'��r�!�<��&�
	T� �������a����=�W�7[�t��g'�y��ֆt�J�R�	"p�Yj��6�8�U@O��Y��b],r]
�7��열b��n��y+\brƦ�t��,1CC6�*hC8�C��ߥ�e!��m����5��WO��r�P�J�E�h�&5��P����G�36�Nf��_\	�.*��Y�7܆�P�.b�+d(���t�$�9Uک��;�!��愹wi������X�\��	�r����!��3y�c�+�@�E��tXh�u.߳~NB'��T~�.0mg���n�g�2����]+�#fWi������hp�6�4l�+�����}�W��gMQV�^���2βϩo>�z,�nz�z<'�(ϰ�^(��T�GE��~͈���N��"q׻ȷf��d� �~�hJ��q�6������f�ø�s *c���#[F׈u
�0�	�i��|�۪�;G-�@y:�#QQ�L�U�'��%h݌����&�����L���9����ԏ�A��w���d��9~��RPBm_-5{�0�	�Rx�όމ�jlt�v�"Z��{�uJE��t�~�,ٛ�NJ$-K�5n))P;�S�������r*�X{�ܥ�����zrS�K���� .�a:��H.�*�i�0���I�c^Y��v��oS7���CPLlFh����F����y0���y��u ��@P�m�������I������2��ۖ���=��^��	�fb(���.~���.sB�
�ߡ!�ګk������&���<�a�Th�	������)���*~tJ5�8���\�PfPrY5#6�
�"d�l.}<��Cm�|r��86�^]�tv��CH��@f-�j���N4��t���R?�Aƌ��������	ȱ�p�9���i-g��3,ãj������L0y����V$FG9~:M��"_�D�� �iK+pj���^&��!� �>�Y3AghO�({�t6�	b�9Ok��մ��WBA6�%�\F���_@��
�Q��>�Sp��
�gY�⠝�m;��� H�"�����ŋ�5����զ����}�#�$`$u��k�%�Jm�LPP$M,���1�lY���$#��\h���P%�Sȸ��"=ȕ�^�\G���C��������$����ˠ�|*>��vN(~;_ǵ��ш0nD�/�L5�.1e~T���F�_�䕄�DXVXt5�I��Ւ�!�L7���"�L6= >?�;T�����?^�$0�N��x�t���bV��xe^�̺�9�%Ǻ�;2�Ŀ�â�����&5s��J��z?�K�+%�w�ԑ�?��KW��_����3�"ޏ{���\�pXc;O�Z�A���e����H�,]����<�O���mG�9��2�J����t*T�X&����z ���F���9�6� ��hG�Af���o!�E��[Pˏ^Y��-J�cO쩼#���C��,R�1�~X�{c�(w��g��%G�c��/�Q�*I!�Ԭ d�p_:�J�'���x-ͱ�S=Ks4H"�žn*j���[�g[ih=�8,�[�`-ɶjEi)UzÕ>�)�E������r��y���1�Ү�ujF��ڠ�`�����J���l���Ί�vִ���1��bA2�
t�ݏ:B�ټ&�0E
����!���hۨ��;B��7��G !�x��Ct��:G���'F�d���%{��ed�<���P�*��2����!��M�&v�sؠP���e7hS��i��/����R)'MD� �P�z'$y�zs;QB�o�k�|������/��9[���ո]	�=���`��D;7��U&��1�qxÆ��;����D�%3�RZ�Io�:Yy�%޿������/�2)5&~�� �Ӻ�H�6\�j����C`�������l����7��岚:2'3�GX�%���^3�[8�g4�2�����0�0����X$>�T�.� vK2����P�₿�H�!��u ��l�oﶃk>ZS��ಱeYn�/���L�[�{�'�F�o�yf����g���&Eض�<�W+�0��'����/y����zX�u�r��p�JD�,L�����W3}��:O
����Ķ�ܷUY5h�Ũ�+k�g�tJ�:��n�$��="�8�JגJ$&�]>��A�N� �V�|��	��6� !a��x%7彃�~�
X�Y���P�^#E>�K!��m����黣qzCX��Z�3o��f;랇A����T��9�{��QMb4�M�DMף~p����6�c��"�T{���-Ӱ���=a"ɵ�t����K���gqߴ�7b�`o�4��SYi�,~lW��i�(��&��L�ዣ�A@۝�p��yH��]�i/�0 ix�[��L����o?9�I�+d�K��A&�����m�����Z[�9��_��[��|׎,`������d��2jo�k_�|���,�uLý��x���x��vh���M^�D�
�$(�wpCj�S�>L�����g��{����� =Q�5.�9D��*�ǷÙ����M?��y�'꓎m�
!���A�(w$|w*����vX�]Y��4�/��d6�t�x��"�ɍ��$>�{3"�_������a�����j�"����o��E"�3��s���R$�}�8�I)cf��7o�3�����UI��1�� n���%E�~]l��+Y7��#��9!��~ױT�W�Ҍ��G�V����{2_	�pu�=�K�pD/3Y��B�]���z��u�m��Փ���Q�7���6�X19B֥��U�<�4Xo�ؼ�mh�`j�G����Y��߂��7�3��39L�T����~2%1 ���~]41����nUv��U���u���AtN�����#�v�:1�H�8����ٺ�����3���+�e0K�S6Uy,��h�}�r�̞"�Йk�CN��+8���hd"z4_I�����nCUIT��*˧��c��9�:�Ҟ�e�xc�Z�pГ0��S��;s-�M�@V�t�a�{��lk]�-��W_	3V)M�%g�"�I�����
g{@j^ڙuL&h�BƂ�T��>SR��%='�`��4���(%��p-b��C����l��#�hѯ�
 ��*&�R>B>4ru�