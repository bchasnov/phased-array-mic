��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,G��U�	�oJZ�@�z�����>*Q�p��~!}8~��m��sDmN��3\��\�A,��y��,�y'Zs9|�v�G��Z��J;����`��"��t�������UnRt��8WP�Z#+ϙ���\���~��/M���jы�IFA�	�]B�6_���Ʌ����&8����9���
��n.��ii�����$jx5����q�\&��x�"�UhU��	�8U�^|Y^oQC�g�]�Zl��7�Du�te;�|���(+�R�g6h�Lo��1��t-�f&b��1wKF����iKE5��[�T-l��Z�>��%�6�8��ƒ�Xp�rB6��?�3�J��
_!������C��Bnӂ�!6�2��z//�!!
h��i���JBK��@S�z�%�O]��íJQ>�,��n�����$�e��z�zO	�sp4��8�d�(Ր=y��{�^�	�4�]���q�T�)�P��W�@ֺg���Rz�n��47˭���������q5��U����0����7^S�a��4��#��_m��x/���������%J!E^S
Dl/���xÌ���1�AIV_"��H�C(4߯Uz$�Wma�;�2�y�#��C�~ߺ�Y�1q7�gd��ʈpz �%�3�Pړh+�Q�n�Yp�S����ϳ:�
�&S� ��[�J��X��ң*a�G������>���"��,,K��<�̌���A>�}�O���B�F5��8 l� ���K�Y���s�9c��_���Υ,��׊&�"������]27���O��_$�L�rJ�<"B�]��D 0���9�+,�yq^�>[�ex��h���/��f�1�z4�9��5����5Y��N� d��g�7�������>/ׯUz�.�Jy�J��GU��7�Kb{�e"w�σ��re�d�c�4Js惲��o���Wم1b��J�~'岔����)9a�a���v�#�L��/���Z��j}u*�����q]M*an����w'+_����Qa�a���4?�xy7�џ�i��c��奨Z����a��2�\��M�U`pd9W=n�9'��<_!ʾU�"�3�|��0�z�o����.�G0t\p���q��	���2G��׫c��I�/���)��C���f�j�C���H 
C�S�*���I7�0����_^��?��bl��K��ϑˆ{�ԓN���mGխń�	P{l��� GN*�$T��%�,��#��j��G�6�3�ס�|Нu؂��H������2C�$�������Zx�{#flpAe?��,<�����X�@TL�]˔a��6�k�7&��R˕=d"> ���5`Z�ioش�#��������IaS��(W��0x����.���C.���Wf��E�v��d7ő�8`?���1,��l��,��KJ���Ux7kYGo�֥����T|2@�f�v_��6�柴�cB�K�Sn��g����R~�AϿQ� ��3�h�;~#^��GG��y�NS�~z�.��V(q�Y�T�#]��.�aL�l�6�Jz�̇�{�|z36n]�`!QF��v��(?=!��t�_��b0"�L�����g�g!P���S,����RQ��z(��.Qy��m#S{�A<���r�p`7�T2j��J`�;ζ�(�Q�q�B�c������)C��GHj��{���LH��T��E�x\�Ѿ[��#H?����`f���8U)x�z2�Xw6�M���B��g�Dc�}�&��t:�,,��R.X+�zm�F��whp��9�l*�x�*@�\��R��-��Jc�dTv��X��i�����������A)M t.�ˋj��F�~,J��ܱ�
/��<�ג[Q��'�<��P��F��p��-�H9�
�Hu�	 s��5���Ǌ|�|ޥ#Ji���=������0r1%�6�0p�H�������*lCo�oˉ2�0�]2�P7^�[������
�\X�GA��$�h��  ��ƪ33ck��J�g�E��$菠�x]�(/D�»9��X������s����L��P!���H#V5�N��"W�l�[Izwԑ���c��Ӹp�y�@а�j|���AMx��#v�AT߸���^i p�4�E4�=B+U,c(���n}����L�b��G�Z	�(���*o�uN=�t�*�cT�nx�Aݺ�`X�t�8'DM����@��*G�ڇ�x#?�@,fz�uzb�u1���朏؎~����2�{��/�Dl[}J튫��E����`������tI#���bĳ�F�o�q�l�yR@P$���VF�ǀ�Z9o_�=U%���Κ� ��w�3[Ve�ɖ ����x�o�i�}���FC�؉`e�m��ط�/!RCk���7��#��XL��:��c�=.�q�6����p9N�T2����*�O<��I���S�Vl��#�B?�{Z���?���跨�}�^���y�i��,�◃��0$FD�.����<Oոbc�fs�6��ld2ˣ�)F��0��l��	�0�դ�V-�9�J���H.y�r����N�R4�ݕY��3��\z݂�N�6�����A��L`�]s�q�?����ܹFT��^��@,"�ɺ�mB�IH�_,����f�.��؟��Y9C�1�3�:�Ձ�V��ī�eZ����J�����c��vgTy����i�R�hK�
��kc��/"��j��P�� �`GG �Qh/HRZR�!�z�M�����h�[��2�v.��Lts���au82���[�����Dݿay(Ew*y�.6�O:��c�0�-۶R��[u�v��6t�N�ۧ|�Y����hEM�Ԑpl�u�` �/�-��V���RWcU�������#�g������*[��(V�R���Z��|5\ڋ��GW��L��I��-v���U�q�{�˞j3��;oe͗I��K�w�O��x�j�-���b���y�{*f���"���ݞDRlKcI��y���9N؎A�郋d�\�����:���SBY���nB�Ϋ
�M>���K�2��	Su�Gd1?y�G����1&�U�i*]n�'F�\���C�t:��ZV�G��<��Y�$*�0�^�K����P�'����eA����J����K��{��o+k'��S�O�h�|9�|煐�� ��]�w*K'��'���pg��i���_ ��0C�f~wD��Ey�.l"M2�:6��U
.�.�FƼ7Z�����7��G�;�"�%5�uS� C�3�RPg�B�X��D	���h�~i)��>5��)oM���jA�e)�p+�3X\�Rq$G�� �#N����[g�Ѫ��%B�j^������49��B%�X�vU����S�sV�%qɄĖpdI�Z"!Iڡ�t�D�|��x����#7תQa�ܛ \�L�-��{���zSQq�[T9�!:ek������kq]*� ���NV8����Rc�dM~����b�/<g~��kcB齚!<Z�gGr�$�4����v&���1�-|��w�@`P�1 ����$ɤ����:�܋�oK���$��l�e�#�;u��$�9��ŭöw�>&�, .wh�9v���g�b�e�\@�
0���RzW$e�T����y�r�1nFQ}�2�ېyR��CuL9M��Se��skD�<�ke.OSz�`�ր�3o�>~n��G�#{���|��Q�%�9�b�� ���m��>D5��t����2c�=��$P�)���ס͉9�2UV���v�H�h+;�0NAt��Ʒ�TB����B&���w�t �C��V�'] ��ҟ�4������0��yc�+N�6 o:�@1tM]���g����T��������x	���ôY����:�u*��s��SH#�|��N� �cP���ֹ-�}��yx�ȧ<�����aY��\�th���}������m+�p�ף��?��{U��kn��d�k�4�{�(R�*�}j�� |�R�v���	��C�@�K��������zb��f�V�_F��	)�����n7K!��_
����,��U�� ��}��k}�ȉz�D�B���3LdRa�F�-� ����Xu��c����1|�6e��O���Q(�ʄ���p�Z���5�]�h���;.�&0���6��!M��/
'�u���g�"�[���~��l��L�n5�~(�N:����kNw�Vky��Z��Y�����Վ�׍�6����|�����S^F�!����R���	 � ߶�-�_��> *w���h�nV:�);�;�y�q6L�jB�F��U�$�e�p�8�DIe�޹���[9�?���G��ɭ�赚����VӮ/�0i�k3}YsL�@fD� gʅiƴtt������>��6�'�\���)�Ԃ}�y8\ ��5��&�k�e�xMP�:�&�xv1w�� c0�;i�Yt���W&���8R�35 b@�=4Je�縬?���4_��w����V�͡��t�����]��@�c��o��KUt97�K�R^��t�^��P�C��AwgBw��Fޮ���1,G����~Tq�?�T�В�ڻ���4(��C)�v�C������鬓��ʻ����)�D�ݗ�Ǧ�cP�o�������~�g�J�~2�o���N��͉n����RJ�Ķ�,��B�p���Ĵ��E�GK�
���*́����_w��+!ݧ)��Ђ��6�_�q�$Ƒ�L�0���T��2�5H6r�e������A�	�,1��P��-�E��L�:�;j�H�� nԺm2�~/$�|��K" �撋�8�������s,�:<���<={ڕ���Mw�q0��`
H)���H?���/��T\4�wdo������3�5�Ƶ�~�;�Yk��G"p���
���/E�#}�a!O>��[G��Kʀ��:�}��~��%���A!��I�7����8=���rL�1��O�q�B���0�� eⲋ�<?���d5��PTk��~�"�Y-�B�6��'v_��!6^_&`�C��c���i%M��A]�G'�����2��N�RW���x*����cL�<�O��e�##j� 5/�����F�ys]��$���	s.)G*��S��	�������zR2ب.��]��Q!V����*㧆X�� �#�qS�pf��[ր��y�"�׊����\1�GCG�t���|���҂XSm�|1
V��c鴤)
CG���!��\ǆF�h|���zڷ�e�O���;x7�� Pj��D�j"W�i�5-� ʏ�Z��!�Y��]g�:���dH���m0L��Ur3��(��l�U�m¤�{!�q
m�Ʉ$�$~)���?�_��cko�S��{�_�� ��m:�+��V�lB��<���J<P^�����n����dH]j�����BI �� ��#
������'��џ��q�����[Ɗ5�h��&-��xD��Ò;���f���כ�����%Z�lPٵCp�7�
�Dp��9��UQ���W�� ������dy�i��|^5<=��(��00�}���(�u����8�-J�O� �T��4������hrq,2��!U
G�b��}����c��>���qI�ʙ3�2S%f>ו����B	^"�P.+���K�R���Z�n.D�!n�hG��}�߀c�6�/���(�B�g�_dAf{�Y��q/?��F��(^��q�d�|IP�V�U���94=P���9��.f9�<5-i�ЇѰF���β�n���YF���iE�{�����!+�$	���SP��\�3��$��L���.C��}$��ǨG�H{����<����a��`ΐ�G{�OP�&�ki`f�q��З?	G�%5�QW*��l0/xS�q�_2-�*.�9�~�)�ֈ�jm�?IX�s=�rX�-�=ۂ]��9�?ǰ��Փ�d��t/X�4Iv|̙�d�8�D���q芾�8�l�����r��"���s��~���OG��C(5�u���~��3�u�z}3���H�t��/D"?���"Ԛ�/l?B�Ù�T2�[�8Z(W�\t�]�x(sV���u������ᘔ��+>�a����|��0��bcI������B�Z���g�ז����ť�pJ�����t�