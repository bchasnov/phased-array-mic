��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\����q�?��e�I8�b�Ǽ$��"����ׯ1�V0���9��";/s��pp>�z�AQ�:6��-4��IzgPi� ���*�������Mj)���Pg�r���=DXi��]v����%��5�h��g��Î�,��/����[��8�z�jf�~/��I�e��φ L����1ȉF�N�F�Ä���qx쬼�*���$���Hs#/)ܛ1��B��]��AJ֪��̟�a�+��śl��;[,.�I�3%֝�VU~�����N~(�����|g��s}�����n���1 �o� DG�{<E5Q#��� j��ͨKw�x�l�ďa<H��{Ӹa�}�	�v�}'S,�f6M�ǎ`�����Ǘ��`>�}�l%A*������(����BU����
�ㄻHy,gQ�<���0Ց�_�������vs�����^x�C�ܤ���f�҆�e��^�mH��_�H`�-��f8j��X��,Pq���c/����pY�:�Z���\pR���\�~%�9R7�1ZB�|�%P+�ɋ��¾�վ�=���4�Z^f��t�n�0;C;��x��ƥS�b��O�4y��
x?�.�Wk�P��xhC��ޣ��Np��K���H�y�N��Q�������e�܀�O,���gnZ�OLSs�.9����[B������~=����V�T�| ���x����@,p�Y����� �?W�u1�%h�h�E%���%�E|�
�- �l>�<�4��R�P �cp��Dt,�l|��q�ZV� y�(*�I����R�2��4�})ߗ�$�.�!W*��w�HH�Ze�HұD�攰�.��p�&�|V������~�po���<�+�#��;����·û��D�A�{�����aj�ؖ-T��_�rB�z���,������������3��u������ֶ!��tH�W�������<�_���˘�'I��<>�Ʈe��^�|p�M@?���������PܱI�d���ȱ��7��+��.ӫ����Nv�H��,q-BmƆy�����_��*�%�4���v�|�teSk*���l��@�&�=-����t��C#��g��3&�I�Fb�p=� �G�,��ˍҚ#���./�m����I9Dx@��$&���b��ܯ������Rh60d'�s6�YJ;0͝vb^�|w��ے"G}ߦh`}�:i��}�.�����S81�mN��t=Q�=&�ZJ���
gJ���$&��Sf1@w�{������NECYOr�+U��`��1����HP��kt������P�M�����#�2�y-Y��9��rs�~��\�҂���f�j�JPG4�f����5J(�꼟j�ɑ��
�­��ΡF�����_e-gW��!a�L�߂��Ec��1��Q"J>ZٰN�J��Vh*�|�*����69꺵H�SMy�8��Z����8LQ��c,�@��|oV���?��<l�8�g}p`��2�cũ�<�*X�`�W��!/|�m�cO�[�����5����/�}Ἓ�,��<����v������Fx)ԟ W"�C�:tI͖��ڐ4���'�4Ǎ�I�f�ݻLP�ƾ3Nr�]o��g�G����=gx���)D1K�[�LgÒ���x�38�2GQ3]�p�S��,NNX��m�>��|�[� ���%����i���]�M����o(#�1&Q�5��.1�`��l�Q��!����+����5Hf��|�7��Nw��؜FU��+�����_b(qL��h==�����!{�sy֨�y��Z	��7!^ae��\��YH_�@{��;�4�1 >���J�w��.k�pC��</�U�6i��O2��\�8���c]%�"G{"��D���_�\����m�I-n���.�6������W���ǁ�D��/�$�6:�_E8@	�]
���>��.�_)a�p�.*��(-1�h��wn��n1��4vj�	�,~v��2ׁ���{ͯ����3�(&
�85j��O} :P��ΨI�t���� }S�62�9�h>Nc}�t�֑G���TxQ�_
��6�|������:�M��8�YF�+���B`KX���7*;���~]/�i_K�:ԕ1�r��d��e�4�&>�2b6�*��D��,���c�v�R�C��@x&^^I�1Pn�a7�E�[��kb��������Աj�c��*���8s�_	���>$���t�r@.��>/GVO��F�=pƽ�6������
�Y�5�B��r��Q�J�~�$��b�t`�����y�L��V�=��-��Z�	k�W6� �ɦtw��D^K�G�$V��Hn���X�M��1�x�d<��$b�;"&�j銕e�	���hs��=ζ��5���0����70=�?-���k F>�ͻ2��i�ϒҖ��gV4�(��P�W�O�ε�/�fg4y���`�M�p��{�1��В�ȏg̢�%�@�^���VK�9�����:+���E&����6:��*�;�͋C�bY�ִ�i}?%O&TB�����)��4w��)Nn����ը��7m�K�=m�$�.���ރfB��vu�����d��U�"��iO�q-�Țx3tL#�NBf=��h����<�I+�C�_h�W࿃ ���f�R��5ۉ5���N�v�ym���ڐ릮8����8�8��--m�M}�*�|p�}�^��+e���3br�q`G��[v�@�s�n��Г�����h�5~9���*F 5e���m���JNMFM�"`�QKb�o�ٲb�eN ���F���R(��{Mނ�	@)�D���S�B���zW�,�Ǽ3��j���̟6�4���
^fk��ᡏ�,׻�&"�<�)~��I�j4Ag����&ߐld���RB�L���h�St;��!�U�a?��7���C��SN�v�cEp��fi��F*�	a;̣�W1�PLplP����F����j�ގr����F�9��!�I8H{&cE�R��z/&���t���� �� ���s^��oŻ���Var���-i�&&s �P�}��	�"ⓨ���M��+/w.4����I}��|���~t�@3�e����wTD��r浗�o{���mg���9�]��C3���fw�#��^p��ٚj!�+bq���ѭ5�T6�9����̑;�*��LnU� v��
��-0��	���� [�/���yᖟ��0�k.H~���B��
PɻPЯ޲Y�[�G���%�F4���_�?T9�� ��|G�ŷ"ט����
wb������6ؓb�'6E�=�!>;���j��T�!��a��
K'e��u��^[��F�3�7�&��x�3,n..��58]�x�X9v��q���C�ӯ�G��F���^k 3j������fP��P�(u�b�c���{7K�:�\Y��Y�Y����������H�Y���a��Z�����T�O��F:("��.��=f����Ӣ��2~�bӰ*�jgCp�৸P|�V"���X�c֮/TU�����s�W�����Ű�۷�N�֤ۥ$��c=y��j�@0���sʢ��.�f�N�H���FU���9�}�e.��`kY�u<�[������r���F��~��y��e��dA󻯱�>�Y�����Bb�d���
,)
����ӭ�i M*���P�ޚ��-�����/��X\��:_�Y�k�|�gs�j6��N���K�(M<w�TOM��-UӖ�lז�C��
��Jn�|j6mݼAP�h��&7zM^Oޟ=ˌ����UEu���ќ��
���⋇���,T%5:��&�8i����u�IU���e��ۥZŐ�� ��*F�ԊK}x*bxHX��4����F̳�]:n�x���.�vJ���/*w�h�rجBY	���絊hT���_�ʟ�YWʢHu�Iup��y�LB�A�2�2ɸ}�^�o����{���w�m���r�mT�̅z�TcK��ap!H8k�O^QM�CT���d
�����3��?���)��u�<$b]_���|2���{�
��`�	�s��
0��+�On),��\U�����㚠�)iHE���V�oK�0N�_x��>L�iƏ�נzt��w�U��T^!��'�Ck�؜�����B��0��&[<������β��v`�{��O��>a�U�ڬF/HuGt����Q��
�8%K���H�ǙϜrTO�GE�D#7�m(^����#>1�ߩ�2�Ȝ�
����&Й�/���lҳ��"���n��ӎc�b9�x����ɩt�����<�
�!F���Ο���ר�9���G�|�N�i$	�N�S�C|���|.q6V��K�j�k�A�K���;���c�V�BH^�3	F�YF	�@8�KG+�g�SX#�	� �(�J����&������'���	�yZ����>��X.ɉI���Þ��J�����Āl�r-0�S�9���3���pFX\���x3c"��W4׫�(a�s�����l[d�����d	L�e/\{�~���H2O���:�N��T1T�W;��KS��u,yw&GX&��H�>��I�'��hi�.����$�ߛV����24d]�gz`q���Z�A���<������ٽ��������w�����ɥ�w�����ב�A�D�ҩrҮ��{L�'�lc���r���h"�h8��<�3&���\�,���i ��1���7��욥#�RtuN�R�.)T0Axq�����䜼E�a���AS�U�/��#͑�ξ��%xU��<�yWTl���O�1qq��+uT	�e����s���b�})��砏]�5�,ڪ��	,�lA_�d�B"���\��a��Q���X�����Y����p�v�N\w0����[�R�w�::*�xy����\�j�90%w�;�-��%ϟW�X�Ug���l{�t�Ӝk��٠��9+�u�1�J��P��A�J��Vߦ^�O��X٢<��OO)X\���t��uF�b<.�JG��xؘ�6j ��o�d��!0����꣖<h��v,U��A$��de�F���J��Q�(��y�� �$��ԉi�|��	��� ���9�ē�B,9�����T�d�W��F�]s���9aD��.)�.S�t\~�cx��)��_���c���݃�r��BJd-�]ȼ������զ6��u�� KdR��/�*��@��t���_�٭xQ��r�������wB�JX�Xsւ����(M޲�w�$��M��ϯ�U�/�!I����^ǔ�b�y�(������P��Jע��@m��;=a�u�]�=����b<�h�sFA�y�,(�Q#"��)������$��Cj`~���o��?$>��rY��F0w��'�鲩��B+Q�?5���h{%��S~����Cg��"��T���b��=���X&:�$DͶ�|�2��$.�E淭%nƧ$
��bn�ￋ�%���.��lD"���Nw	lWk��Y]��\a{rB�m�︳7Y�[jv��K(	�-^���C���Џ+�p��yUY��؈���sLޟ��R��_t�s%t��'�kP���D����ID��y(��H�2�����]�ފ�ճ4�i�G��P��ȴ2��c��^��>�N4�J�J-o$�L��I��c���J����`ؼp�zd\'�w��Q9Pc���.��U.歺-kZ�2w�ڗ��~�K���皖R��Gﰙ
���JB�R�j�t�|CH�؏��u��#���4��k�d�щ𕗀��ꛗ��`�߁�g�MZ׈�BJ�sz�㞧��y����>q��:�8}=n�����\�F2�nB��K�}��)g�p�I��@Y�WO9L��R�j��k���ڵ>#	��KV�����@5j3�s���<����a���x���˹��6���ʟ2�����Y���R�5�Kz'���z������qb<)������y�9w��-ԗ�� "����y�nY��'3	��2'7��=���9M�Ι�����ȟ���9����[=:��<&W��~�m=�ǉ"�n�P^MJ"E;��p�<�`e�Cڳ���"G
�CgF����������0eU�ֱ�F�=`��(�b����W�����P'�u��1��
L�g���[T�#�3+�@@u? ��a�.����>���=����R��-U���i&��nYƭJ��ba�T4J]��1��uk?a8F�f�'ʭBD��"��G�~��k���2*MG�1BY�?�$�9�U!���° �����|W�q�U{��������}��P�w=Ơ�z�v*Q�ę���懸����DO<=��i$�VH�ui3�F��-$~I�ft����=��&��0z����Q��A�xj`�cR2F?��5ʔ����� �nH{�p�7�h��!��K�a�݇U2��pʀ9��[����ޫ�c�/j������u�$�8�F^��H	u^�A+&Uu&���^"�¤еӂu���{�x��9�2VF���vF���iAB��t߹Nz_�uA���C�.�Y��L����8�w��M\�/Z�^�����p���y�3H�Z߾���N΢����T�1wT�!��R���/�գN�t�{d�>N�|_Z����8ݵ�Mü�+4�JyՎ��9�f&ɀ+QU�2����!F�~W.�pF;ŧl�lx?_�B�&{,��:��Ɖ$F��˫j�4��vK���@�J�)�<x�t��n�ӏr,�h�R�d����iz�����?�ՈI��X&|�K�ԝ�Q�j#��<�0K�BH��OAk��t�?�R2b�y��$б]7�MА�7��_���ʟ�tV���Jճ@�
�?.556<�ݟ�Ƴ�Ʈ5�0���k�p��	Zd��gdlP$ȫW�I�
�����/+�����u�N	dӷ[&&��@��\c(���oj/YW�p�C"|X�בQ=�̧�zƿ����6��~�C��%ef�Y3$�'�ޜG�:�,?f^ga}���I��L-+�	�x���zxY�#����0�����;r��1dB9]�|��n�b�R	�'��z�	y��[�PR�=��z�: �	��)�����_(hq/c04Vh�}�ŗ�����f�f�����j	4h�D�7zV�D9p��Z�
���H��Qc '{��MoX���,�P=�j"��b;i�eK�!7�}���->ɔ�ɕ(f�Y�;ԁ��8uQV�Tz`�"�]�]u�l�:5hc:o"e��S�>�h1YW�%`��+�V��qU���gex W��A����؛�D�|h��4A4��Zc1���f*�藀�B蠾���M�olb��dJ�~�;����"��K$��J�
������N>}G5 ����ۼ�X�1���P��U·B U�	�.| ���~�;
>(��`/���ʓ�d�X�Act.J�����B�-�KDR�����H��m���f�Š��Λ���=��u  ;v����m��`o��;���#�E�{l0�ѺB8���Ә��^z��^��2uha�B_�0��V��d�����D�N}��[߰�e���^����r6�^̜�U���O���w���-MIr|�PD"|��r�z����?1�]�|��_�i3�ϲ�3��"�G�<��(�_����RhZ��ȗ/��k�]ᰜ:�9�1���C�A#��տ��B,�G)m��&��Զ���]4�����<�ca��X����lly!t`ֻP��]!@�H���ʘǿ����m�0�d�'��8��'���V�VW����,��b�ܲ�O,�Q��F5���)ǃm�(-����_
����nD��3xV,9��x>�����*�؛/�x-��i���S;{�5� 0��n�5@(� ��u���Lw�������P5ΏI�ֽi�At��]`������ڝw���"U�VJ8"s l�zau�&������~����Y�BFhY�e�?�9�)j�]��P����t�˸m��ܲ�{v�H�m}���{0:�3�J(	<��xۋyWW��*��C+R�\���1Af���T���nܷ�ӣ�:Ƶ�!*��
y�jXV!�1b�fE�-e��� ��@�8��
�jDU?��ʷ-X��&Z�� �gG�b�Kc�l�������"@�(�;N$�&�q6�S}���s