��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf\�|Vv �|�
����:C�q{����B��\�e�w�s�v�����ē��ZzkTqk��A>��4n�pt�3�AƓ��F���$:g���2��.%�G�[�P��U��B�/Kݠ�os�ΐpBOd2߻���G�)I����~y]N�53���y�����pnGpj�Z�cF����/Ѿ���� ��\�E��7��Z�E�΃��~F٥��������Y������c� `T���$4��^�y���oF���{�vn�@��y������S,L����	�BÎ�H��[�I�O�,ͱ1�Q�b�:h�\��"����K,��rp�g
�����)��;�/�[9hqIya��XnFʯC�)cɛ�:o�J���H�m���tĖ�vp����	f�)��pc��F�}�瞐n�Ƕ�݈[f?����-�l^�@a7�q��. 1�=@Ț�ٗH1��b�rGl�bX�k�d��]��z,4�� �7P(����:��i����V��x����4�M�"��	�'�_�E#9��j��y��������+My][?��r�-~7\�gFbJ�G�I\��u�������@�`��vXBK
�$�M�!z��C���TF,/�͙�d���|â�Z���5�җ5�G8�n_�د����\yѳK�^��7U@�#1�U�`n���׍�RU��~d��bdv�y37y1h�g�N9�앩oݸ�Z�V�]r�}(��]́T<mÁxf�������c�|����H@�!��B[1�"�S�<��x��]�1_'P�8У��?1k�+T���|�z�}�W0F����d��#�o㸮����#a����y3�!a(�}�Y�p�=�B9��I�6�;g���x�_R�"C�ӊ�'��C�<b�$癄���6_�7~��k�྿ #F�
�Ĩ��	��^P��r�S��R&�_���3!��ȑR0�5Ll�v؅y�����ѽ�}�}7J΍YR/䳂 f��T���4�>���D�j!��$�Qc?�rn�sMw�R����z��/�<�Ԗ\�����3��JqC�O7&I�Ρ��lXEf^	��
hE�����]�����{�����y�c�oL�B���e�]�#���Ƚ�}�����<�ǌFv�?N�&[ȑM9�F�b���z;"���c�Y�&)���r��]��}���x��&9�J8@�UG9c!ϛP����ә͆��N�2�Y���S���3R�:���߬_z�wnɘ���F���-\�҉}~���>�&�Ȉ�ws몺{��n�&7�r'�%�4��r�tdMh;/�)�0Ĝvٺ�UZ4'�VK��u/
����epm�Ҏ�
��j��.Я����_�-�^�P^�����%y�ǆ��ud��`�m�q�]�7�{i�Lki��������C���j����a��_S�>;a%�{�k��Ő�U��Y@CV��TKK|z��2ѣ�Һ��xcշ�Mߝ��f����R�U[:`A�a+=���!��̺�O3{=�K�T<�k����fN��(Y����J�>��/I�ߤ��z
x�C]t@��h	�H�S$�8t�K�{�<k.B^�
���Z�|]���H$�q>�l]�"���!)�q�H�©�>e�5��Ĩ�Xu��/��
��� ~�4�@A��*D8䆭�V�k�L��B�Ŷ �msĦ�]�ܼ����u�d�x��4�V�	�6ne�`.�ݘ�6�;O���:؇фe��1�J���5iMq�`���z�)��Wb5�Z��_#wZ_8ҧ����,9@WI��:Ͽ�m�}�_Sp��I��S6,?�0|�ǫ�����I������6�Zcai��{I3<d,e�.k��·�A��-����.��:r����ϬA:t�rQ�ji�*�@
�9��$;,W]MN�G
d����@H*n=qp]��>�S[���<a���JIܻa�~��<V��Yo�aP}z���=�� �HߥBJ��OtbG>y�����٪���k��E7����* ^oCI�Y�p)�Z���U�y:����ξ��� "��uM��� ڵ/��e�.�!�)�&5鯚<�4*�y�����X7�ل\�pxΣR��rʟ�ςTS&m=z��F�x=����_0v�]F�o�%��'��JΡMP(��$LoD�C\�N����S���O"��L�F_�s|M�x�z
���0�`�t$M�W���@����7��I���B�6$I��y"��νGY�=�Wfu�i�f�������J�yEt��U�5G��A�g7�����˭N1aǢ�"��j�'�1��2��e�f��u� �v_q�Ijq�x�j�Pb�l����)WD��a#=_��ɏ��u�DE>�.���Zu��{6��X=����w���:���4MN�ʂ��b߰6����ѵ�AWL�4y�5-P�����jD�9.�5���B}���C�hֿoU簺��3�Y��&�_?C+�/ZἌ�Xtvn-�wH�>�SY��%_�vK*�]�G<����P���4����F'k*�����W��Rȃ����ɤ~�0��Eq*:��̼h�έ�rN�+��A.�4�E��A����x��ծ�p)��3�DB��������9ۤ�%���?Ԗ�h���f�A��1�W'������D���i�,޸����Y�:$7�֫:N�+�{�U�$�m�s��!���P�<b�$[_?��Z˜SI�h2�GX}4�dm��v.���ƥ4��?��>��Q�Xq�t{����'j+j\=T�-:l�9�*H=��q��˱��s� 4
������Rj��~�j�����R���ট��l�\ٞ�3�L4á{���L�$��M��R��+�u|���+�O�̣�P��r��� �z��v�@j7Y�D4�FW����HM�P��꽽�Nʐm��J��%�t��hq��}�9>O#^���p��=XQ!�gO�����^�qӑ
�����>��t���}���-J9�R[��ր.i��!�N���3��b-)Π��r��_gZ���>���>ь	�잜�Sf:1�֐ZƲ(�؊�ݠ�O����Z�`��'�s�J���b ��]��>�I�/�(�u�5\]�n W0s/[��������:��*�J�݅j@�/@Uz��o�	%��F�d�W��~� ��.�@�]����S��^��fW���o7�O ·+���`��	f۩B�C���t����C��qۍ(�o	0fGv�Y1���!|Q����插��0[:6�S���״k~'�
�3/DqsB00\�-BL����dN������Js��,�v�j�EB�6\ee����i;�n�j(�ߘ�8L���?� K����i�S��5���G����v�{��dv��~�%)5�;���jv	Q�4 ��8z7oT-꒼��5����&o$-}DJ8��zN+f����V;�)���fP��g�3����"{y���`��{�1I8�#�bn�c4���dv�h�=�j���\ŦC�
Ai��ފ��r��	xTr��b��<������T�:�>�$�(D�`��Fc�-9�:����W�tn������L��{�Z8���=��[�v��6��cj�_T=���J��b8�>�J󽏶o��j�J
��b�n�ZSꉌ��D�1Ԏ�/�:��
�h��V�:f���6����/�U���H�Kb9��M�� �Q:���у����~" ���6��1�!�����n���S�:ʈ,g)�E~�'��7�nR�V>bQ��5��b��lS*�B�-7�y��9��uh;o�5?�fD����g-�j�����
��=����"d T��Cח�S��-Þ0EI~�+�;&0w�H1�Zx �A�UZ�LB�~x!�(�Ӡ��lܕ:�)PGé6X8��:�}��s�H��ɜ�Ɩ���::dK�R=�m����ꏶt��EO�m��K�L�)K4�,o�Uʗ��{��#yb��y��3t<p�r^w��5�17����b��m�$�UZ�	�-�>�k�$������xL�.�˭J�^�f퉕�1:��N�y�Z�P��!¬t4���
K�d�܆����[�ac��3P3*}�}y�ŵ
����?�d�A_t	]B�����2�ە��`����<�R��'kv��Zr��_�|y��������ɧ�4`��xԇ�\%���I���� ��-��d��z:�����1ؔj�D�~Z ��0�*���{"ujފ���q1B�-R��;^A~����	J�c���A�3g���-�����/�!=R�J>!˦��*n֡\�mW�$B�Q���[����c�{��Z)�T�/�Q� �l1s�R�ɭ�"~TH�i��#t�G�mM�]��v�q�����q�_J�@Wsd@��7��1ԪՂ�a�UN�䣾u)�՚�w9��ڏpޫ�a��Ov�xMU���^"�s3}�|��E���b�ד�vw;�� 3c�,l3��N�\�tMZ��r\J�.�`S�Dx�&�,�C�V��P���5+G P���2G��1��!��%�8H��ެ����Y�A.�s�m>�9!��V9��	�d�`T��'�O��䦨����R��9lySkf+�e>O�5[{3���Bk���B�ZF�ѭ�jwŢ
�,Ef��������/"	��0�%��uQR���<���.᣸2�
tV�'7��ip�'�8����(x'{%�{� ;R2��m�B��LF@��?�H �!�i��V�!�P�)���5fUS��h��>>7����9��Y�1�jk��a �?z�/�K;��U́4����<�]T�02��F��.YO^~T��]ԍ��Al,�_��yYg�i	�!�"Wg�NG�d��ȟ Y��z��"�^���]俱�Z�T�([�l9�HB2�*�R��������OL��-�D�����_��ϴ��6'������R�?a#�4;����2���p���`?˰qׯ���a��h�F�3�8ס�&Q?O#%�.���*]+� ��K�8�����%��t�,�Y���:�=q����D�@Z����qg�{�E�ڗ@֛6�UYiMiY��S�)/�B��ϥ�}N�e��$�P"2Zl)�����8�/nTB�o �^��Ȼ�~:���`���1%�x��X�k�sk��8�'�酗��oQF�mp4������N0U�lLsZBN�e�#,aK�aDZ椅ްe�')�<�Ω0���c*��i��~偀�/�Ҝ�Z?�8Q�TZ��� ������$�I�r�?�`
8�#�j�Zvt �#G%{%�4
�c@u�y~f#�0W�v/���l�"�v����9Qu5Z��;�1>x6��b���%t^��n��
����M���6���G�}�^
��+��%�H�8(�D�}������Ɛ�}U�,כ��9S�3Qݡ'_����+1�4�ҹ�PK�JdbJ��Z����W�a�ˤ�k=Mg��Cz�D�C�J��0V׈'V�_�Nn5�@�˖����j+X)3G\ɫ��Ri�UV�;Z?���r��Q���2n���L�����Ƃ ���*V��.�\�Sn`޽Z-��:�Re�
O4M��y�l5K�߉fK_���vv�S����i�����#�-�����ʄy���FC�m���6ۄ�Sꡐ����V��y(B���T�}z�9e�����m�4��/��#��qZ4A)D�3�-IR A&[�I�t�1z5��h��A)K%Y[�r�<��R����+�澃i"���2,��(����v$�1i*��!�8�$_�����ǚ<�t�ɛ�^����4���W�c(�TAM���L�u��L��3ǵ�-Ra���IuS�2��l�c�9�X(� ?^,�d`����I�η�u4Wƣ����r���
Dc�)��4����"Z��N�`pPRJc��$J�������Y)���C���V�h����WR%��z��f�]�(��:���7b�B�U�u��o�P�y���<��G����f�˯�_�t��#i�e\!�s}M1�O׵�~�aRI�{Z� �� ��^8W��'V��f��p�������ν����A�Џ/�����J�<=5�V��;@oeDWq�Z7�֣Ƀ���6�#Q�&���Q6���
V�8S�Ho���iMS�K�$���n��e�|Yo�[�u�r�x����~�b���^�(%�$iu1cj��Gщc�A��>����׌п���ϯ~ɏ��r(��TXjr\O���0�2V1U��CI�e�n��}�'��l�{$�=�r&���	Pf[L�wS�_�#󢰛0����E�׉#�o`uF�������Ԟ��e r����x`�����%'���0iӸyюM�y�� �%aAf�|�RD�_K[���v�+Q���0eUEt���/yZ
_K���F�!�b����e;p��t��~F�,�X�M����^HQ2���v��֣iν����M�
�p%��+��r�':G@+%�2�X����޽�|�P�>֢���<G�k
ߗ��><�%Ffd���A���.� {���fc���S~�bCnw	S�n� �.���x��X�k!�����q��qr%��	��z��|2-!����~��N}�,bY<x IY?�	�z����{��h�
��ڀ�\-�7l�&��ڒ��)�o'Wh��n��x�նI9�g�a�Z��V�p�$5�u�R��zM^�0�:�>�밪0-�u�})>߷���ty��/�s�:q' >���X��5V��gvv���ufhi���Th�N��,nٍ@�i}��:�m�W!�e7���OD��a���1�����|�ך��5���?4aT$ܪ��?Bx�\)U��t���g�-s��	������TGW뎤�~S��J:��,7 �mn���)ь7R]��|yude��3@���t���o��| T[`�M�hto
uvr5��)��thuCS�����e�K����ꈚp��mq������#�B�V0!Q�� h� E\f���g"��/f�M��h�� ��Ťn-XI�[�p���6�K)��N�����`s�w�:|��3�Ea�L���LP��V������hZ}F@��]�V��@���}����y�����0.��!�RK��}4��o�!�i�v��2U��A�]%a��;��r�Q��"��J1č�e/���RD�𧨋�d6�#���"�v�x:�A�m��cm����B���S���(켂�H���~�����c�p��JB_
>"�Bx�8�$6�`�`�޷�W������ �t�(ϗ��2:�ُҗ|���<�kU��D�@Ik׏o���_GIff7�4y�<��'��=[�Ҽ!�LN�̮�/�o���!U˥�rԈ�^'�$l�o��Ԃ�����<jU��p�)Q����$��I����y��A����#<b�;d>��),��@z�����}��`NF�-�א��"J�䱣��g��+ )^��±���{��'$$~i|d�%�����f��w"�٬�o�����z5D��[IӅA�ԙ^�ﴣ��Cr~��a[I���̏��'�%FP֫{r̉�>�ttKN��2}f��4U (l5Ki���Nݥ9ݥ$�J4ԒB������(S	��Z��x��nM��m�E�>�˞H�!����U�V98�ě�y�ؐ�>�J�c�^s����]�T+C ��Zu?S���z������*tZk<��Y˰��c~mG�Ȯ+�d?���U�F��a��0R�{����'Ppu{���m�_������R�;��'����32����Zh�N�۝�ۨ��t�μ̵nZw>�tZu�y_��p W>D��Ė�5��am��=��99�푄A\ ��[ k��2�ڟ�
h����^�`��t���לo���2_���&���_��X��y��D/��1_1u�^�����m ^�V��'���[� �Qh.wsi*�Q9���`tq=��!HII�a�c�����K��C��`Db �����M#�L&�`����N��~|�Tu�[��/�/�D�[���o
�,UVQ��xݮ^F�Q4��A���>� ������)U��_�)[��5�ٸ�]����E�W�SU�;��0N�����uAO��'��?[�ˡu�=Y*�.p�	"��c��L	�m渽�#�6oh�o���i֬���8��Ԉ�{��N��E�"T1?��`ef�\Y2zf#a�X�����N��Y��=��M��$�پ�4��bn٭�2��d��S2�~g���3�)9j+�_���JqB�C���&5��Ů�ǹ���<�!�PeƩ�i�Q%-�%JM����vY�ےqK)�6菉�%�����?��n;} '���Ȝ����-�d�������E��z���o�8��uDP_ǘ;�oX����N���7��T.��(��pJ	Ct�����Vw��ߨ		~d��c2��Ԕ`T�[*�d���n�}f��0�YwN�$�0�gQ�-�)�%�*}���svԎ#S��o܎d�WM^�	ũ��}���宱��P�&���V���g�A�\
(��)VTL�H�����Ja,���y���y6O�D�0����������$3y��޴n��B3�L(�j8~��z�������0,\�<���A�Kq44@�ƕ�*�K��Le�~L�_3�ޒiS���z�p�I>�R���9�WUR��^����M��ӊ�������OIH���5�>c .C¦KR����UV)�u26M����g�?%_&EfÀ�n���w�Myh&x�,Z����"��O��(x��nT��`JG ���z�L�R0s��s>i��Vtw�� x�
�,E�)��ac�x���j�a���׽8�V	o+=w5uKG�`E�����v�on�Q[r!^
�5U[ec�P�r?b�����
+���&J�Ɠ���a���o��o8{�/�@č�*��[i�a(mk��@C��V1T�,�4'�Wl���k�bu�:͓�{M���cs�لVyCթz"�\2��v�������#C��Y�%�0&�HZW�*a��}��=�hq�~L2�]�WK���.��|(�Z%��|��Ev[�t-��Tl������1� ��*Ae .�02�LO}:�An<T�V)��/�\!���ܽv'R.��T�l��'�q%�
{YT�|�"�3�)=s{K&YS��U����Hp�Zd�@ʜ�Mgv��6o=����u�;��*�h��u v�F��r�Ύ�B7�W�@��'��@ P���q�����>`�dM��XF1<;�P^��e��Jk}��Zo�����D�ߢ�g݉j�mS�T}%�����������lS{����Z�c)[�t�ċ�#��n@!�q�	�(�M���#Uɩ��s�W��nr���Ө=I؄~W�b�n���)THZ�e��8�����6�H�
��#��«�4��3|���~��и	�b�S
�PEm��s$z3\u�2�CdovJ�I�]͏��͢��.��ۍ=�� �D�rt�(�\�6c�^q�(����s���Æ�V��2~,�:KH�Z�j[��׫��\�ԨH�PzuI�t7��YIG/��h+���urG�S�9+�ҏ�I�6|�����W ZY�<������W8f��+�9K1x){Q@��$!q��f<D}��Ȥ��`�V�c�ŊK�SD��Yc��XNa�P����P35��B�δ�@�᛽Mۥ$'��CP��'��@ j�f<}Dۼ��Ѫ��)�d��aK�3�9R�y�����4	4���4=����<�預jUϱY!��h�6۟5�*��2�伫#BaN�j�%
�މX�шy��O��
^a��~g��WM��� ��cV��v�ͬ�N*�@��1y/��.��:N���9��!�f_'�O<����9���� '�ip]_����% a������f�����"��� e`�,�0P!�j��/��Q7�MC�q��X�.u!����0��i�3�F�����M�g�� �7C
�Mm�t}�P''�]�+J��",�2�1ņ`@��rw���<��1ry�զ����������4��%����������e����M<\v�BF�d�UOZ*�Ɂ6��/�b�B�q'^	gU�x\��l_yr��9� >�p˙����6>]]Q`�����e��������{������/���ԓ��y �<,��ԇp�MSS��U+t�Gw�vG �� �v�m��b���
��j���'��fTA�m���fy�'�߷�k���2c�ߴr;��t�j��᭄_����������%��gܜ�jI�����\Do�VY$�}���߱~��4\T�8�rsKݮ��}N�(�d\v��\��_�-��5O�Yr̈́�;Y9��n�WR:1i�eA�>�'��s;��6��5�I�}�a�Jغ\#�<�����8o�f����V���L%+�O�[�wl��s�f�T1C$1_�u>~�G^�b}4�= ��'�� ��:����&J�h���<ʲ�B,�
���k}�	��v̹��bTA�B�<���!m��H6�b�=2!P�؆�4I6s9�XWWx=7������ޞ�����+��F]��I��7#��Wv9��&�7̷f�L"i�{���3�w��� .�w5��I(́:qO��L��I(���t5��KZ�U�e�@��`껅����P�=�	v�ňB|���z;�E�D�&J۾;@o}�s����E�falz|�����'���p�j(��[�h�Yd �f�}�#�-'���a���$�0S
Y�ߗ��ܧPK�8�eSf��U��fefi�A���c3 B�\�]��$��sQ3˸�g�s��� �~En+mޙ&m��=ݣN��1Jϲ���@�e�;����ܲ(�g�xk�kA�b���ӏ5�xv�W��!ѱ�ml��h��D�=H�2�ڔ.�)%��2�*�DPA�q9�c��)B�.#䮤_=�ȵ���=�8�5��k��IZ��x���z�+ҕ�<\ʅoLߨ�jиeT�t�N�mغ�)��i"�4��@\�%Z���hn�VihlTۆ�����B�Ӂ�H�v�M�?�v����+�"����s����6��W��J�T�Q{�^vŊ�
�)Pu��֢J�c�m��3.����:�T@��LU���L��-p�,}���/��UC�X+�lUu$��YH@�$���t`��v.�2ừ0��d'h3��f�և�-�Td�}�8�#%M�%��W�=�Do�y�h����5���[mT��һ��l!r�-s����y����e����ss�ew����y�Sd 4��.�\	�`AA	�~�|/���P%D,�����)�~��JG�k��RҼ&4�r�0�Yء�yHP�k� �O�V�8��1-���7-��r-MQ�3UW�I�{j��.Hl=2��0n��5��I�F[�DH��/��n���6�5��� a�0��ʝ��]�(l�Y�*��c�.���b�! �����_��cR�8�T1_�F0�p�bEdT�7�-;��{��I�R��,�c��vQh���o7zT��szEin;C���8�ǐ�S��ۧ^)+���ů}�%��ޣ��@����&�	[$��KD� ����Õ �Ka�Ji��b`W���� ;@���0�
ou|�(`s���"�� ��M G{.H���`�p��v0���{�
EK�%�n�D��:;�`%��֔;�1����{G�W��c�!K\\�H �B:���<�ɚ?nX4Lӓ~�L��]��+�M�Ӕր$��r�Y�n��� I1�>D1]�Ѳ���w2�������%����տ��pQTU����H��rc�h3�f��(T�Gm�z:ɰǸGJt_qM,%�g�n�n�/v��	9
�Y�J�I�5	F���J>k�7���S	�gc�Ձ>o�$V3HQ��C�`�#N!D���q��W+�VR�{H�����G�n�-�19 �悝-q���� ��#x"����a'OX�A��,���K؂�a5'ԁ��v�������oh!��^��� �ʲ�,M�7��sSd_�|����cU�]7i�U~�^T�5}��>{�;)=k�t��H���y���8��}��5��<��\�2P �u�Ww�ގ�ᾃ�0�o��ae��N�KԪ���X�uH�>����&^�Y����B�I<�A̻!���)�KQ���X39�͗��!M��?x�j��)�d��I�EfҴ��yA�ܑ�f��ѱL<��a�g\��&֟m�7@_k��THї�ZJ��S��p�"f>+��슪�V������������:���V��́�JW���7�����B`��lR�R�M���\����!���'Q��Q��8�&;��_�Z�����@|�+z��]JcG�1ːY����޽ݫ����:���іυ����#|�8=]H�����*r^mQ�^S�n�O�6HU��-��|Hg�&t�� ���စ��W�3>ֽ��рq	$/iW�P��>9sX��`���%�]>1\� teJ��U��5�15%�I"@� ̗�?K}hk1Y�]6�#U�u:<΁��ơ����^��զ�M����-HC��$��u4�9���ގM�(�B�<UP��tz�h�T>���*�LU�w�N!ʎY~�TZ���;�N�D>������ׄ�z����*@����[�'`қ�lh�+󿟯!ҖU�\�]+i�Gc���(�(YaE�y��O��Y������:�1 >�bۖ��k�{s;��z��2��(ߜ�yJ(�1Ƃ�G��b�1m��ʥ��0��4����r}��̱�K�AB�Fo��8B�V�k�_H�Q�|��9�N����G)$Y��Kb�.d_�/%l�j2ʻ�yZ�ݍ�m�=�0����:�Ւ�FJ�ā>]�T~�.��y$����K�v��Z��T�n�04 9H�A��JE��'��,/��+��&2��顝��]����R��L�%������8;Um7��B�:j��}agzo���ށSK�uS���k��@�%i\<	�K����f�f��$T{��=X���aFl�*j�Y𡡝=D�M�6�3�(7m���VY�HƏ����G>�$J�x���W��i~����?�P�}ѡg5��!V�ȭi�{L+]�=^f�c��.��MK͢.|�uj��R	��4V��B�1KL$ �S;2���J��iF�;Rz���	��ʴ��Y����8�YY����H�*�D�ޒNt�73f��.2XG Ӥx�~!��z�݀xCxY����e�����D�C{����.n�SRb1}�Ƴ;oF��cW}��Y9\I�%��\G�W��۬PF��l'B� Y������h�r��U ��m����7���H���0�@qJ��.����i�#�� ��]gd��/��H̖�J�@��HV�c�)������4��z+YS=uM;R@���oc�vv�c����G亵2sػ�)NE/��������M���HZy����Q��ۗ�L>���7�W4J�����nh��*�	��kn���<h!�`���0JZ��5ޓ���K��_U�������Qq�ҸG��Qwޤ��֧�B~��ԩ��=�;?����^[����&�'�� "��} ���.>Y�Ɠ������zyM�q�'j �.f���ə܅`O�Ntg#���е��f)��f�f��a|�9�9�$+Vy��M?RI�Q���c����v p����*�!��y����-tF�t��f�̓?ӎ��������HC��GL�-���ӵ������i)6"��D��f�|Č#�U�1�U	L9W�ju��:��ћ�(l�<Q�X��]�&]xy�Z4���g�)^���%.<m��m�*��8�vI�m�χYv���J;Ѩ�/pi$�J� ��1��Ň��3l��Lrj�Kb�1R;���}���G��P�K	����m�	�r��}�� �����:��N�����v��94	�X��y15g'�ȳq���2�M�#B�l����-Bv#6���� 9���w/:��!4�(V�?Hwq� ����H��K��x+��0��)��ckT�W���v��B6�k����3�Y��9�C���Q4<;�6���}�����:f\p��֩z��B�ÒN�������凙�h�vp$:.�'�U����1J�*
|���B�AIi:�߸P&�
Y^	>"���h�y���W.{�pǀ���&�Y��jb�O�f���>�j �M�?j�����Q�+u#@wۡ�-0���`�<=��=��g=p���oT�j�_n�@���K-!�;��<ϙ����Ja�{f��#ݹ	���I�	y�Tcw�/dM�F�ߠ��n�#M��c��#o���qqR"��V��J�Tn�|	�_P�m{�<���28�'�����h�
^v�d	�y�桡���ᳲbQT%��|���jGdx���6���_}D{ŝ��������y��0s���Fv�S�`�W�ڼ��5�C�b��MTr�dsC����O6����3�FeG��A��K#Ĭ�PjP��ڴd{f�|ߛ�FZ�_	���Sl�[]��q�g掘��a/�u>X�<I0� O	�B>k꺱���p�j�[J9�{L�!9-|��&ŗT�Q��Q�l���w`֮z뗰[!��E���9G&=��:���iv�#�����*� H���bQޗ^�a�8����p��'�yו0T|��[���1z���Z��>�����w�Y|ҭ�ה�0񀈕e��'���aj/Q嚵�>�30Ԝ�.߁1��Tvۀj�����ݕ���D<k���jp�fh��9���֭���#ӕ*�e��tӋ��8��A+"T�ǭqA�ޘ:TX[H��W�s��Z;�C��"dk�_2cЀS�U��Ȃ���{z��J��)g��mvR(�yxr8��wZ	g6t�m�"�M�����D�S�ʕ L|-p3��p�?�p�?(�|
Sv�~�f�
���/�J;HU�����)�y��#���#���eF+�gl��T�̜瓰���������"+�sS��7DI�֤úL��y�e��Gt�Z�Ş�FE����d���P*��u�������Ai��U�	2��hWW�aKc��������B��C����H�Q�;�[\Օ���_��P�UV�{�܎7����D;�j�
�?i���V�u�����-�7v
�X.��M�cQh�������j��4�!�̞j����
�q=>�{:�'L�LBVی� g� ˶�L�S��8�b���ˑG.���8t2��̞K�+��+�Dq�/郀����x�ډ�lj�Sy&�`�Lw��^+�9�P�����|B�|-��'�"��_�s�~��
�*�mZ����l|i9��x��9`#��]�K2��j8���c�U/��?��D!�RO*&ݴ���b�5�(��2	}'$Ϣ�Z�L6�L<�kv=�~{�k:�]ҸTܻr�`����;�mh7���fh��t-�����n�=¥��ۋ�/ͣ����������i0��X�$q��� ��M�d5�<ƯP�-=�`�ȗ�� �e�����SP
@[��,��Y����N�ӂ�E3@ߨ}X��j�-&�{�	QĂ��#?5�G��NzR��~�{�j��95�j�?��N�.�׍Z;�Ό���=�u��b�i){O�Ş����ͭ+�^c�6(\7|i.	w�D��x�/����~��ސ{��� ��e�<-��s_�M�B��b�ў�r��g��-4���Bt���2P~OV!/��aȽ柃�M���6�7���0E8�Uw�U2��JJ���[({P_=a�f$�7 ߷TVƞT�ݏx1@���P��<i|����v�~^��-!��)D�Qnd�\b���<��e����2A�WVUP��y��Y����s��	��8�o[z@z��A����c��l4�3��w�KݱG�����r:+l��x�G��U�?��äN��vޝ���`0Y��|C�k��)��Iea��q��3�tp���E�d��t*?B�~'�?鳍�nJ�gS��]]����4�l�:gwBdq��6p�^��YFJ~�!\y1�b&8��M����g.Au	'��A�>S�h�;& �*��*m�[�E���Ǘ�q������09������"�C������?�k�K��*��π�P,q����V�֨�I�����Cv�B$�,��q}6�q&�L����j�+����"
���iT댪�*'�bG�;K

�W$g�[T>p��)��`$7�Ld)��Q����FVN�%+up	���Av4f�#1�,d̮4yA����C�\
W?am�9K?�plL����3���cE�H���� G��\�K���u���\���JZ��}�YxT��Ͷ�\��}_�ﾄ?#�J42�n��7�d�ͧ����HC%��
N���,���������&eo+�J�#�څF�?k�F���_�m}_�J�~���qCj*���e��J��S����ԥ��{�r�%�h���/a����T�������][�-�t#w���9jF�sw�xwX� *���f5Eų�c�PֿQ�yO��*p&��M�Af�����|�'2�8�R��6ē�2������������P<U+���}=DRx�c���c���s��8�i��IަY�� �W'��{3��b��-�v��x����V�I��k��9��;�Km�ɌW���l��F��u��H��g��Y����w�G�3�L�LױeC��ɒT��{ .��4Jz�YAd�2�_Ȱ�7�8�\5�Ǿ�����)�̎;��F�8��ҬU��1~9ʽ����VW<���b`�N��Qh�������qD�.��6�'T	=��1�KN� ��P	b���9O,0���]U�
E}�j.�9��*���&t�,��x�Xz����'�(>�K���n�%�Pvw�Q/ jsSx�E~�����z� �ž�Z�{�!nH#H����B旸V�"��YNz�}Ȣc�}�:v��!�v���_�ӆ�(\��JML����
�keMRV�(�M�`�G֛�5H[Vo���w&���!�:������Ҕ���Z�L�D�DR���G�~?׿�eɘ�zxR���ȁ���:�*Z���|��S��J�I�`��n�y�.��+&� 6d��^۔J5\o8Q�Ury(�솴�� �A8�&�>�6�c7�}�0v��#�K�7u�7P4oH������ ��{��R�όSR��Gf�o����
K�p�����3W�>E���)�6e��h��d��>�h����1�X����1��
��eR���Г�6�p�J�����IS��O�zk�K�����W���y��+�s�Z��"W=u@�9�2�WrܑWb����x>�\i��$ӑ�Ӻ�*��'.c�>��	Egn��te����B;�e�87qa ��U�����ۥ����93���k��BY�G�������#�����xW^��`���KW�{��<���B*M^��/��	4�$Z-(�︧�̣$-,���+��z�\��ja�2_׉�6@��U߅\m׶��s����?}�ўs&�Hɤ�X+$y�2�pQx�KM� 8�*))`uMyc����� @p��-x4U�s�S�W܈��� b���~^��8�e0�hLc����ח�4U�-��Mq�!� M��QiL��G*��N��ռ�#�O�E�����U������mQ/2��!o���W��Y3tf�Y�j���j�,
�}q�?�t��8�v�(��·"��TZ���\g���h��	���=ULQȖxN��럘 vj�7Ҕ�AݨLÛ�C�?C/;ʽ�����<2�&�Ƒ,�4�W*���;WP�St����\�q�ʺt��$l*]K�g�W(��CH��v�1��:�l�2 _�wB-��������O�*W� K��q�d��K�lM�P��"u��vU�H��E[��(+����*>N�������R�`�ھ���B�m?� a�N4����-�X�l��)�����WC��`�nQ��"3�|A��d��(�Bb�M�8!��)�f���HC��� BZtfZ����f����xv�C9m�BRQ�\��%�F-.�#Y�v>EF[ͫcw	d�nݞ��Z>��>;�Oǹ2O:#�
K�Gd2��՟�]-�4�$��vIr�����h^�s���}�}���g��n�˳��(���t�L,_2�a0x��X�;�9�Enq�S��2�_���+����d5����>�
L���C�%J��@D~��"�P�Tٷ�h�1n���
k1�Ct�n��ٓ�(R\qR��i����#���2_��f\|��í�D�_�t�pU���Q9������Y��_�)�عS��-6F ������ܲ��d?�\U_d)����}͵�u�%��B����.��z�W�@4�9"�L�6Uk���8��ثS�B� �M]*�B����Ȥ���A����S��� ���3s%W�5�t	CbD�`L�c������/Q�=+=
Mjm֭8l�ݬV\N8��46Vc���Ϊ͂�V��>����{d�K:���26YIy�����)�6޵;��]<2�s'6n���n^�׆��AT��@��O2��v�?����h$�lp�}H��L� ή���g��Ad`E�"��Yz�G��f-		\�TN��~HH,��G"'�����R#��_��R�eH�
L��Ć��\�&1N�]dYb+��欳Cj�o��	�+�a8�7zk��|S�n"���p���!'�0�F-���S�@?�+��F�6�W��v�RV4$Y���A,l7���poPv�/7Rp�?�/7�D����\�<����u�� 7���O�"l�5k �O�Հ�x�=2��o����<33�����2w8��Tbr�ͅ����� ���u���g�t�Q����GX��h՞���\���-7e�wT�nB5m�^��E��p����X�¨�Tn̫���?ףh�e�I}|wyƆEi�0vT�,����@s��@[9І��|^�.J!���K
d]���F��Cib�� 1���K��R�b�/ʝ�r����M�^v�z
�ʷ�q9�5&����NQ d0�#��`ͨJ�S:������@O���`�+�έG����`�H���s1�.�[�a~u�;�A]�p?�]B7U��g��P��	�,TS"aLO��x:�¢{�EK�j"4�磡��q7�Ã?������VsB�1�|�1�`����U� 1O1SE�Xyko<Z>���l�j�B��M܀�����7:�t-���Bk�@�.b�j�v���9�YF����׶���������ꇊՃgV�\{�8��X�����v��t��
=��o~�t��v1+�~F�{=>���&s�,�ŜR��r�L���N���ֵr����"c�Ri��@:�+�&;T�X0�T�Q@�<#a,��i�@���a]�py�i���{�,ͭN�� �^�4O1d,�T8�3x�����i�f��~��_E%�@�F�sia��T�����q�ֈ|g�$�K��d1�K ,��� ��(�HEC�n)����&Hۏ^�Ŋ�[yp��<��.�:^��bG�̱_�I1rt�Έ����!{0b`xƙtD�F���� x�A�y���3�ڮ<ك��� J�;�:�FM��1��m}�k�C^}�+��� ~t�Q����V�	�$��u��ds���R�����=��
���Fd�3�Q�a�m�l�C��d�!�����A6+����+~�,������c��73��I�	u?Q}�	:"��+'����xUksLaw6,�W���}��v���-�f�E@�t;O~�\:@��ʊ�`�9�O�8�ay�),XX�aY����j�+�z���-� |Ķx���L[�J��M�}����u�%�q��pr��o-��F^c^}e}~��D>!j6���w�