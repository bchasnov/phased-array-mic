��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1���e}ʲ��cg�t�ϙ�a�:�KR�%���ݧw���ȼ�$�l��i�� �#�;,�@"��3'��� �� N!5)�G�ˆ<䧶�>F��ð��x�}��Z{����T��@�n��R֔I�m��\���讎#Kr!/����ɀ�Z&2�z�+���f��`���s��Of��N��"jK����sb 4��V���Q��+=̀��s�TZӏ�;�T܎�ت��~'r)�������T���l�L]n�[Z�p�}���mgnf	P%�w�"�\�C@h)tR�lt�����R����T�+,�V���h�8�N�e!��k#�B�z����r��F��G@ɽ��ۦ��Pq�-\s�>i�vS �F��2�$��O�F3��72��>ۭ�DY�;�w׹��p�ɖ*�`RGeVz!�gi�g�4\��i�2�Eڤ�Xd���M��u8u� ^gIR�ON���*1KN��T���婚ӭ�,���"f��P�ao��TMf�\����*G�$�.)E�Ñ�L��+Ì���i��9 ]���k�z���l�2���DZ�zC�`|z�Z�1D��o�E�T�M��-�-�ʂy�����p�VN�ih��L�6��>��k�T�&�?k��f�+v��O>=���e,�=�]J��?����	ȺB$٤�rd����Ǌ1��'<����t1<�	�ݰ��	�'��D�R����Aެ�z"��!ߕ�堼�I�1�U�Qt��=Sp],;�a$��}�V��\���풧 -�����u"���OyfY�%xS�==S7]Y��#��_� K s�0���v�A$V��ǀ�ч�!Zd����&�X����D}@𞰁o��}:z��b*;Y��,rtB��Ȱ��'F�G���D>{(6~7]#z��V�z��=��h�Cn���c�G�癝�HM�f���eт�}��c�f3&��ٞ�b�	�ɑ�7�����]Ey�$ ��.����@�����)���ӎ�d��_�V��������a�9�P
��)�$Vg�5�܊]�iBC�Į��}U�9L5G� 	�I�|X��+�i����	F�0�%A�:MF��T'#�I�S�i�jM]�I���3(�&�H��ӫ�
?�){L�}��[tC{[����W��MPbf�� n*�`��V��+���g	Jm�I�RM���R���Kӵ�h$�>.6KO�4���	��5����m�������l�� y�Z�$�+�8�[x��m[S���gLyQ��6��������=��  ǔ9�*|G�cr��?�B�Z	�s�bc��)Z��c�6��1�h��چ�`��W����
���§�1�Um���]�f�Z1��Ry+�YZP,�V5u� ���<��?��8|4�L�1��`g�7�=�X��U'^+?OZ���2���V)�<���KW�<:�-�#Y��`��eJ����$y����J-\@�w�D�<�l۸��	wQH���pCR�%	9qP0��˞ArQ��I��߇5�����Ҵ�f������>�AӆQ��V�:s.+m��ɯs�h�(x�}��b�h>%�X��������Ge0a��@����6P,(� ��d����N�;��8Nh4�Z-��~-�->o���r`��k2�i4�Z,��sC�X���5��F@i�8x>]"j���$p;�a��4������w�PQ8;��'Sy�;��D��7<�|ţ29��!Sl���p���l�4�T�h5k��d�n���Iw!�m?W��?PUl$r������)�8f��Ә6�u�.��©�Һ�!`���~+���{��%�))�R�9��D �]�>r��s� �#�9�����*[��E��8ܲ<LF6c#���$pb�������rD_VObY��x!��b�ӈ9��F�;+�&'!r�x1�$�ʏE�BޅF�,��
�@�x�W�G����a3�v$���.5_$�1�e�hW�[O[0�����J�Nn�����k3Ӯ=��� 7J��[�l�d�8?�>q��w����U���	Q��Gc���?/U���zi�:KWsV u��.��9���]��s���uj�A�t��d��9frѳ^Gh�b�siO>����)�����QsQ�(i_����/��|��2W�g��3�P �-���G�{�� �H��GJz@C)"ES��l����*�Iձ�:�6���e��
/s���vZ�(>�C�=�8��TN׼b'����E �s���_6�H0sB��s��Lu3��{��[���{	�:ɓ3�n*�xz	?���g�����MLH4�tJO�7�q>�Ɇ0)��DA�j������g��T����+���&��Rv3E�-�Z8.٪�,<k�6+�#R*;y:�j����l{>�l����G����e�K�Lw���>� p<�=e��|�����c+��O�^�ttv�̏���E5�N�RpM@���ҟx���%�U��;li�x��L+#f�{�����{37##B���pwRO�
�q��yoJ��TLwlB��G�3l)�^���0����f�Lz��E��Rx�XKb=T{��Ԕ)ꃹ:#A�\�7��O������������&Z�&��'Ư*��kr�]�G�����k&i#L�6����8@%��}�E��:W]����J��ڸ�{6C/۩�2�m�2Z�n�+�U��^^ p��v͊�_!jB�2��(� ���xJ�m�-J�b��.ʯ@B�~�y������Q��*\,��ǎh���B-Աpzb|�S ��_ZM�v;߻1�=���E݉��pcX\�� &���	�T�>�!���e*�Oz ?AE_Fmޢ���K�)H}���My+�1��h<��=(�ڪ닦� 慪|�y�({��2��|Ȑ�
@?=O�n��vau�q��B���+���;N�?6f�(�	4I�=[�UW6��.��N�k��'h�u���L*B�$,������$�S�.��X��-9�⡪Q�ٵL�[�Z|��
��J,�k�y6���+͕��3��l�h�A��7*bJ�o-�>����W"@�)6���˼�?Qɑ��M�Ty��W3�+8--@�י}�Q8o�TσA0���g"yރo�F�"z��t�׿�b������l
��.�(f ��<�w���5�ZH���p��A��o��<�8np��2���y�����!����!�deO0�u��̹�ٔ���KH���ՇH���a��%L�k)�?-U7_,tEmt#L��/�~��zv�h�髵l	D�����H"�\ͣ6��铅C"��H�ۀ��pZ�I�����|@�h(�Y銓!*
ʙ�?�Y)򏇔�y$MWL�q��8��V�f~>��Qޑ����:1�J���[������'�l%�ٲ9�
�Ɨ\��I�y� ��%8>�s)�Ա�Vˏ��+sY.��P
���1� ,!��ԋ���#��Yﶖ�6Ӟ�P�LK�I�ϝX��a�`�M����~ڊjYvB�,ͯ�>�}���X�'��1�m�0�l+�R��ǫ�9�2�&���l��=���1�5�T�$��<h�g�F��C��UR�$k�����{X���B�m/�$�kt� ����bnX�_,���{~�|xX�rd�wXu�@�}(b��nky�I�Ӛ�߼��З]g���glC�x��V��$P�~�]��2�1"�h�!�����])����W�%����Yu0��=h�c`Λ��H�$��c2ցW2G�����A�����4�Z�ij�4��������oD��+�0h�8��\�ɷ�BO��?�ڛ�0�B���@i��r�,����~p�Tw�.�6}f?���rn�V�ޯg�s�����r|b�g
&����9�2T��/E� �@�"9a0�7l^��^�Y�Fc�u��+:h�eё���l���Fv�Uo��̲/�c	��uE�V����LlFǂ/񖈸E��#��)������җ�.�����P���h��~��^ �,�T�[��.)+��Zh5~b�%��>}� =��_�2#��m�����+�[y�1i�U� �*��צ��U2��d��37��UH�R�&�Lt�܅Dߨ7y��G<&�W�5��	����5u!#-:�����]�0���~5���hl�CH؄Z������\�����x���{O�q;_}��mZ��/�Yy��� �� �	.ݻ����u�-�T��2p�G�7��I�y:��@�����q�-���-��c45���(GX��C����iy�� �⾷E�
�e���_�6V5������0�.��I�;N����d����NJ"���g�q��ؠ���c�Ry�~�̀"ɌC�VE�y6�ۆJ����m�����Y�Ԅ_�I�u�..1!�3ܚs)쐈�Uh&��_㊊�'tzk?T�������Jo��8��]K9d��r���i!*�8�滛���ٖ�g�6Y��8tZ�=��m	;�#�cx���v�Ŗ���7��DU�a������J�_\�
�%���ֳt��y�3S}��+P&���7Ϲ���tkã�ɿ���QZ�+��=c��r���x���^Sbq��%�����S�K0��(a����Z�ȶ��y�h`z�}V�6��@�������Vd䱘��|	%�J�u�+Fʤ*uX߯#�VW�ˊy�iȵ5��g�b�ܞ�h�� YU����I[�ˌg�&~Z�A?� &N{�*G���G��a�?�� �R���`n�X�E��(����5nuvF��5��7ݿ�%��������{��ޯ6�clmVNaΌ�ZW�l�Y���|�\�*xw��}(��ZD�*Kb�
�@�����=19%<�T��a�U	L���/A�y� cP�"������0r�6�F�����H;�]�@��e������]_t�S��\�:���C8��5�B)f�7��m�ͬ�8��U���F���QS���lT�$[5=F�9"J�@�G�DAG�C'd��5L��]V�m,�޽R`�zq�)��"0uc����ٞ��	 ��-����*�1�i*��X�3bR�.�P@��|�cb���g�#R#��{Xjy}�wQ�#����P)��X��wK��`�x�f�W��r)��N}쵀��Y��K��9��fUu��Yw6� +��iB���hԗ�UΪ�`��P����o_V��;+�F��Dx��}H?eE3f��V���A����櫀�ĿY����l�$˜��_lK�rWY��Kz�E�r��j���iF���xvU@RD���° 6*�^�d�G`��P�_��jk��g����yaɑrd���v���\d�L�~Ҳ�lmU���siZ�vO�Y���Тn3<�_%�fna�@�m��5q9�M��߅b�\a�Iu���kв%@w�jTw��J0��A�A��L;�b���&}Z?H#zC����+i57��S�B�(zۚ��0:"P5p?{,�`�wg�N;k�(��8�u:� o�9L��"�/	��Y�`D��ogp�#���&W_A19���ɣ����X�� �T���R8su7<��.64��B�K�`�>{���j�F�\���qsW�e��b��3-�W���0�ێW�X�1h�E.���I���߃]�O`��H��*��H�q'DL|d6o�����F�_j"T)؍���׭��~NZ�7����f��6�8Ba�x��
�3��l�*hjC:���q Z��_$��yZS�/'�5�o��)���,Q�;��Y�J"� q��68<�ث_0�<���8;-�R4�j����m�u8� ��-:Y�}�zSA�&Pr`��mc��ni�z��妕��I~�����LJa@O�l�rlw�,�7M4��iޱ��I�P$D�OZ���J���K�AH|�����(!#����Y߱�i$�.ԛw�t��ؠܐ��Ս����V(H5�˲�`�b���'�*:;"�|mZA;��7�ѣ"r�A�}�S/Z�9T�d�:������@d�M�Z(�Qс�g oE^Ԩ����9+$���9�`��P
�0����w�������}�⻈��è_��Xv���;�т7,���p���c��x��s2�XNv�:�;��+!F#�M=��bi��r��7I�Me��`����c�by:����q�of_�3
��8�jV�2]�'���+ʨ���l��(�
x8�p$D�3H�'Uf[;���M*	�'P�0�q�5�XJ7��V�R��K�9�M�ء�5o��4��ґ���5\^.�R�V��i�#����0������=�pHn��j�('��HvzɺL�,44�J�E��\f��ët��&��3�HE.M�)~O C\����B���n������\��"z1r���ٍW�	~��nq��&��ҝj��EX�0���+&��s̼�"	hOGǐ�� ��:�$ n�� �.1�������̌{�Y?��^1�80IZ��N7#J6��J�Ig9�ͅ�*�2m
~2S!�S<Z#Zԙ/��<K�J���O�-��S��܊~@~��l�Ζ�	ʯ�Y���oY�
��ب[߻C�|Oִ%��������,��dn�����:�G���D6ޒηK���klF㢺���SȊ#w��Ex$0�e��_����O;L�gO��*j���-|Kz7_����ΙoL�0��u)x)Yv��Ў��RxjC���Ν�a�H]zT��aCx?�p�AE$h�%-��vy������2�W��,b�S���f@���]�_e�L�*Y�`�����iO$S�����k��X����d���k�e�r�&@ ��JZ}�Xb��*�?�pW�������N�R�I�@R|f{ռl�_��Lz�����!���O�Efr���J��F2����c,qu��g9���G펋5�?��1��*	͋ ��?�Lɽ�[�ʼ�n?���O��~6'�$��^�i ~J}�o�)�O�)��o��w��`U�Ǥ�K��;�-�(�o��R
�}C��`+ň(M\sGH��cJ*㖸�Ș"-�d�f���5�9CY��`� ���S��V��HV��w5S�z�nx[3rP����#���? pK����S�2���,�A�I�Aއ��WY�SvɊ]f�*�%��km���kL��z���/§�|�Q��RA�'`��Qֻ���z�W,4���0e84#9j����5�5@R\���J�Q�w�D��DP5�p�zfE?�6�j�TU�Ԗ��FĦ90�z���t��4�̔��:`�Lu���r��Nj$�V�+�
��ڢ�%kWy��������i3q�Hu'*�c/�Ͽ?�0oV�� ֠���GJ��`�����G��QT�5��O��O����u�_ү�7AbĪ�i
HqD�����B3�c��7��)����7!)��ȑ�B1xU�[�̹�7۪
�����I�N
�W���ғ��!l8����S��
s,}K���f)u'�n��e�q.���ա�w�R�jIO�5�zA���!�	� �9�m���"��C�$>� \��]��8]���I��*f��L|gw�:'hdU�+�F�o���E�w�@Җ�9OU+�t:v�6Ts�׶�	�L��n*��$��^�14l�y�A��Q���o�_?r�����z�=h���a�0�2�sҤ���N���YQW�X��:�e��'���o��a.�0^s�=��ʑ��3��%WN���"=���D��3�t�Xߖ�p�8�X�Ld*���S�����+��c��H���n��u���Ҥ����ڂ�,��k�M�����w��-���~c�2��<�4�PV���̜�׬Q+h�b|z\��єL�2�+g���3�zZ<Q�oE
�	�H�	�gL�f�3�v����0R t!"�=��3w(�LA��a��˔?迃=C_裋n/mӠ�����ks:z�[a?��'���Ft���bR���G��_ڥ#M6�Lq���6柒ӊ氊+��[�.)�KL<c�i��A��0z�g�97�.��1��a�_v��F+[�I,�چ�*�f�wQ���H눕{�̳i��F�/�� ΐK���O�N
H;/G'prF6L��$������҈4H%l;�/�K6+��[��ڈ[,�7�weŵ<����cS�|L�
���`Z߻W?u1kA�~0��t8[;���1���Ԁv�Ș8�*����է��n�x��,=�د`��J���M
Sq�g򫣝`�ԃ�w`���٥�� �_6_~) 7��9��h�F1HB4>�͉�9�2Ţ;WA�=�$�#s'v��oDѬ��NB�g��.,g��s_�r�[�!��l�[FV�v��L7�lO����.���mq6�n��G��k�xҺ���D�:�<��֔Zof+b��^������캡���dg�1���Do����ciڂ�˵
.�׮���m4__��/r�L��A�_a�U~��S�����͈9�-8YO��HF���>�I4OH^
��70i���'#��b�� (�T�s�nC��j���?Z��ő�gv���%����a>�`�OD���A��P�&��Sب�x�%��'�7��q�5�EX��9q��Nn1æ��b@��~����)G8+��>[%z�|�i�0G;�=��kƩ)�.��|a��wn�B)oR[[��WB�l�.���3tS�s,))�E�3І@��R(l����1���(�d�q�ƿ, ��
�Ih�Yx� ��� �� x�`B�½JϏ���&XZQt��Y��46=I*����A�dqs�8�/,x���Oe�@�:���
��hS��E��y�m�`�]�����X+z�0�e����"�d�*�W{��������Qj��b����J��� �����G����;�lٶː츶HM�jA��=�6�b~Op���䈈G
�;%[�Ь�s?L
Z�@����$�7=6H��*kz���m^�x *�'w+f;�pͫ�(����� x�E����RrܾhZz���UK�`����pC������j����'C���s���3�	�Pt��u�(�\S8M<ϗ�t��@EW���3���T��0�	?�-���|C(��暈8M�4�U�`��ٴ0;��ՔS���y,}����p�bb�y��'��1��o�jcvx�.��Yİl�^-�1�3t�	���ym�*o	lC7�l�� ��5���	R��LeV��4[^���[�����B8�m=�ˋˡ�+{�r�{a�&t]D�����ר��i�*i����ʴ7��������	4�)dx�B&J��#rlaIl��̅nSD���P��Ph�C����y�F \v�`�/�z��ɥD�p�5J��OV�Q��ST�HvkK��#+jy�'�^}2 �R9����(�IuE�v�HZc���"ٖx]1_�$V�u�9�ħ*��ݲ�"s���SBy$�
ԃ�)��HV"�R_�xh$ੳ�|"-*�@�9v�r�6.{N&�E�݉��+�~��k̢�J�ʇ��r���+[�|��/3�1�D�i�%'vy��t�z3�5���`G�K���x��J4�聣2����VM={�M���t��H9E%8���i�����5 	Hh� �\���|5����x��)�&��8�{h��xf*����ͷ�i�B�34|�=[��h<�Е��*�3BM�6�j�5Q���#xY�[o��Z$��7L0�S�kH��s;Z��jM��h�k8�-!93�?5�1�b�ҏ4��Z,e��=���IzPF�M{i3�=4����ev1���)�H�`^v��3�}f ����9�2�_��]��TN�@�W^D[>���Wv�2���PԬ��E{�;�Ӻ��V�l�ߔŻ���~�@�E�H����Rj������"[n喣]���{\^�͉Q����l���P�|�d *�	K�#SQE���
��{�T//�P���E�v$@3�>��W �:�;�� ��a����ĸ	v@��k�F�{�c`EM�]��n�#�͇�Xt�Y���;�l"�Ԇ
�V����GcqR�Y��8�nXj�cSX *(�I@"���Q�.��}Z���JK+r���jLF���
f�\Ԓ�˽�Q�WDG�GI6,�>% �tc�~�Fcg�`��JG��d"u 	��z@?>�u12����&k|�ݴ��#��[;���V��+8���b��J��D`��?;�ƿ���hee��l����#Z��?���#@\��%nrZ��1M����C�מ�?7쎼���3��6l��)�g�qj�Ik��n�m�7*����ޔqʹ��;̽�0Jt|�[~��NE�&8}z����T�'��'��]���gJ�d��X�A`�� }A�2W�q�Q���#7�XL�ڲ.�McF�����Z$�o����}3n(�D���u� ����E����0�wRt���"!��~��J��P�����n5�ߤ�~j�R�5 �CA�R���݌�R��ǕŦ���k�x�e"�k�މ�|��ga�ѽpD�M�k��Fȋ��t%~���7!&�лjN�S_���'�:�&12�gH�,q��T�?JE2�֏�vL��w������i��Ρ8!΄�k�+�����Ƕ��u��w�ߊfW֫�/��I�w{��r�`.���%_U8�L<R������/��6A/v�D�l=���/k)��S���w��?�<�:�������R��v�}ݳ�hݩ(4�Ӡ�=q-��[fh����l�{�r��_d[W5�,q��Z���+����90�S����~xY( t0�H)����T�s	v�&���'Z����jt?j�#W��+A�,�ޥ���8�+�yr�j_�?a'A��LV< u�*��3�=9V�J�L�r?7ڏi4(�[%�X�P�������6J��dY�P1��-�}qGL�4w�c��3�<��N0?DBS|�+5mu�W3�W��5X�y#���{��f�����a�R��?MQ���;�ԡ��������	�͸	�wc���z������?w�yr��?��ٰǬf�e�Yw�������uz��~����������'U��H�]D���L���1W�4|���6X�+���K�O��o$�ٝ ��  �RY)ߡ��(Q �-�6��J�/���sFX��%b���N��{Q�b`��a��⺈��s���_P~�����)����g�{�P�T�3+ulp�<K�Ӹ0��ڈ#0�Ջ��p���3�ĉ7���Es����H8�ӗDL?tn�[+,@cuK����[��/�b�����*n�ڪ!Kb`��n0*�C��GYa�^QI���i��J޴���Ar@+Pځ�	����皡:e����@;Q@.d>��5*ܵ��$yғ��t�߹W�5�g�X�wE�lM���鰋�a�����'��aP}�tV�a��$����$����v�3+�)99]����ˊ�#���io�n�hsӦ*����u��`��d#�r��ať��	����-��%������Km�Yσ���-�+.K~#n�yF"�c֔�$�bi$��(��0��#x.~�>�=Կ��`EY�Eo�e;�����R������y��̀6b�?�6��a�n?�5�&�΅� ��(�+���4�%�cLh|�
3�L�fU!/�N�C�9z�l�rK�N��&� �d?����r�,�6�tYLz�!��u�ѧ�_� 4�x
j	��(g�/X��!~���-�G��P�=�������F��ܧ*����{S3�����y涆+���5m_���W���^W/6����7�AT�������Cl	�xKAϮ�j�74B�6��:??R�IM��8:��v�@��՗�K3;54�x���c0S0`4j6.�u�ɹ���R�:���j��"��6]��f�(q�Jk�#�X���c��UW�������L�
s��0��ňR�_��ai )�p�g]S�ھ�w����ىt��|��o�}��b"<����y�g9��Ir2�,ť?T���XrY���P�lw���B�Fl�ǖݥc�C4��b|7��þ�����	c	@OO�\��&�v��>F���Л!� �Dt(�&j�{���<�0���I��潼��i]6�颫�n���a��˿�;��m�⢯j���nR�]���:�1%X>��r��@�	�z	���w�D)+��;ӣC^�1wVRh�d�
{�\Y�մ��Йȉx*��"�n���Oy���4�?yɤ��D�*�y,��b����u�6��2�n��O%�����oWT�Ǫ�[����L�m�����dg��x��#V*P{W��
5�п_aNA@]#�ڀ����B��Z���8�Qʜ���e�RrD���Y��$g� ��fQ�@�Kx�bc���+�EHm��`����s�Ğq���Z���9Q�J�ޔ�/�����;�:P`�JlI6����N�H�̛�����+��d�c���P�v���A���X]�A����h��+��a�6� R�n��P<�s\���,_$�bQ�\�@.k�����H�dm���ρè:��J��UR�c��훚tn���q89�'+3�nH\���;;���0؉	N�[��e�T+]�݆=u���'Hk.�<Ƭ�ҶJ�@𜝆d��ՒQI�0,�%�Fu!����,�&���.ά_���qM�
�.f��ܩ��&��r+�F�ޮ��c`1,.)�SP����˔u���q{M�bR��U�0��r�������6�6�����	#}9e�nNoL۹��Wl�)�&���U o&m�r����:s�&EvB4JOof��,h��
f������H�E�	� ��G�xuc:x8� z)u��0j᠔ig��*��K�k�N�f�~!0�p&���,E(��_�����#-7ݹ�&ۈ�)��,F��LtȉqD���)^���3��� ;��'Z���TUD0m&�G�Ɯ�:���P#M��ޝy���
,�K���#o��N�q��䁗|��l}��OpFɕM6[�{�(�
��B���r��{,�g�oPS
�����*K��/Z�^B>�f���]���`��w�`!_ �5�+k��.���H�����{��2�3	W����4*q�0^1��	�\%>PD�N�ѡ��	QM&/��!��X����H礋mI�6��!�*u���3a1~�#�����)���'٭�8zzlo���>�W�rZ��E�߷�J�=�V`��;`�t�i�A���qv]����J��a���H㎟��h�:����m�"ǺO8��Ee����#g,bX|7"������Nj��R�%�(�� :~f�\W���Z��n��c���������1~T�������q���;q��yn�9��.�iD��T5٧�	_��O��,��)�b�`����wR<6��"Г��3�2�7`v?~��6K\d���A�ʊJM�.?�b����3�QO�8'��77(�K�?TT#����)�ln��v]H`\�%'Љ§]��J�߽�i��Mr���Y��fb2��(^9��ܞ+��Z]�=5n_�4
ۇ�ː��"�@��H���8L�}|��+,�cK����������
h���)�U|��
61^���s�*pwSk?E��?]��;X�(^�{�x�=��gR�r�>�1[�9�0�9�e��mvJI�G�͘�8A6��B�wY�rݙ*�=�OI��'8�T�pa�W�Ql<�[d�]`����'�7JWp����2!,�V*zY2����#������}w�0F_��	%�)�{�2g)k��?�k�7�%��H��$���p'�R�v�\4/B��FN4�-�xΣ@��{k����r�<�my�!K�a�Ѽ4(/��_�$��d8ٓgs��t��:I~�<�$����7�F�YX�l��g
 
���@l�9���N�qZ7��@u;����#GI�%$i�z<��ACB6����k�����@�0F���T<���
Zy��?�����i�'Sݺ�`u�R�!�jgB�	���}4r+<�Y����u��<�`���E!��M��<�'��iϽ&��I!��`Y_��)����N���US ���b�QҢ`詧p����@�20�FVO�>|�o���%�e��w�O�1<e�Д��k!� ��cd����VUU�?��⯎�[�G��*,�
�9��*e����uK�;$6<QA��)/mKO1���5�>3�������b*/�� ��/��S�X`�-�a��#�G�*�ǂ�5\�o ��̱��X��X�X+Ѽ�"|�c����'^��]x�e
�O�]v�r�|�'��"|���k��n=A�[�gC���ÿ)�q/fpqb\���ӄl��M�	'jlױu%��Y瘫.DkP$Z1\���RUH|���9��(����da�0�`a��~q|�� �ʩ���<���6�s�����E���]O�NK�$��F��.��(��	��HlH�e���޴�(�ּ�Z;\��X1�\�	A�#C32H��SUԤr��?���o� ������.�:<�Ъ����3�q��;�)ǐ5�\�@cVYu�E��B'��,+=ᔊ���f-g�6	e�1�(2Y��`H��U ��+�[
��D_�&�F��h(7��F	�&�<���(�2��������>�I��V^l��&��s�eN4�JS���[��?"/�8'u ��M0^I�za�w�#�x~FĠ�$�����˚��7d�v,�)x��k6� 	�&���cY�7y/���h�0fipnu��D��U]��c1�R��!k�>�Q�}_lz�p�z���}7k�[��!<Cբkæ-��r�F���Gz��@^d�az�|���xL.�q�,���o���=>y�٥�	h E珿�]/n���u��]�9l�Bd�5}g��<��}�2e�!�|`h^H�����<�\��0�1���7iw%u<̽_�K�C�EI���k�r���"�rB����f��/�s�5x�L��EÔ�dY#��%y�T�/��eMWt�g����Y���(4<�'���Cl�%���[������׃`}N�e�|��G��G��@�W7PȄ���7xGx�t�I_���Bt�_�̧!�
B��7��)�V�e8����g�sO m���G�sh�'g(8�1�����jK*M�:��_��J�@,Z7���n��B㹸E��u�D��8T�IR�J�%�U��BrZ���:N��^݄�X.ֺ%��X�2����p�!k�v��eϪvSv��y֓Y���4@r0$�x1\e���Ԏ_�H��&�A,3ئPCIGg�rS�:���N�n�Qо����I�}�XYk�$���%�zaо��R��ɠ��m��%��WL��`��%`(�It�{hD�F�sU��Dca��K����G;�Q��" ��s#��vT|�g��?3�w��@�G���M"I�YAG�Nm���%��7l��l�O�%��.qbD�R�1 ����Ț��o��B0��=����z<�ǖ04짐���]������{�>�Hq��@Xf-���M}����K3��FB,��(q'[<Kʇ#��)�T�=��k�+�7��dV�qx����ʉn�_d~���U|��j��=���<2t�������R|��z�3����9hEX��M��,+㛉1JB��L�/�xO�|�)�Y!�a/A��U�+GM���t�+�ujZ�@�I��J��Q�����)�N��,\��AE/�]h��գ ��*�HU�����o�iZ)��Ԝ6|ɺ68��T`:�K�\�}�[�[?�=��Qa����a�<�P�<��[~�`L*�a���b-�H�h�tѷ���>9�����o��ӭ��AE��s�8���.D�^�)�m��G>|+�.;>���o�1_جJ8�$���c�μ]�; �������h.��u�
�Hs;�w�!m<�%�i�P���f��B�J�K�Ed�9j�l��Y}ߓ����tX�bȌ�����mh&6�A��kͱ�%R�o�&i���h޳v�G��UE�ٜ­�%]�0ƞ��L0��l����u9ۈ3�3u����ߒL�4E���,$:m���r���ª��^ִ�?�\�b�6���T��H�~n�"��6x�5դ��ݏ4`hG�f�^��=��&#�gx����1�{�M�r���Ms�6�b/���v{�g��>e�l��W���+p��I���=Q�L�f ���O�~�._Fj��|/��l=���J�
<Hs������˰6�K���s�J*>m�.�� CmXr3�d{�� �&�3���u��4�߷Y����S� ӳ��k/��\2f����վ��J�X�Oc�}�f�I���We[#h��O� 1ǡ�t������{*�N��e9ɁΩI����cw�Co=���:�)��!���ˋ޷�G�����!0����!p����|���5K3\���\������:��7e'Ţ��&M����W�͕~���hH>���@E*	�4�*nD�� 6B����T-t�7�S.��n���6!AJ�U�5��/lZ�:n|��Hx�C}d��
m����dP<v�St��ʘ��'G�</�w�_��m�P����Pfܻș����g�c���}����6��]�(�k�]�A'�ٱ��s��2"n8�%W:P}��y��)��1iH��Q@�I�~�4�o�Z�����FA\�k�����k�$�9_�W��k�>���T��ʱB�V�[k�nk�?j2��`>��'����EuE�=ъi�j����!��>#=QkP��͠�E��$����4��E��-�K8�x�/쥻��
2n4��,�e2�S���`��$��'�"�Q)�5�v&-��9<;��C �$�4����jq4,Ra�6�|Cf�?�`��WJ��\��.��*�� x����)�./�J�^
4�{Qn����uˠ5�W3�	���r��E��t˿��"�3da�n��%�?i�F�?�`g䶉3�o�0nM��gnǢB��}�����Ȥm���! �B���T�e�v��{;�u���P�"t=�C�5�ʖ��we��ʟl������S�������yb�$�;}7�*6*2��2�3��L��js��6�[�e����]�� U���Dפ� ��Pz�*X,Ňn*��KMnK��w��,��k�w���K~2����&j�N4��-���zEr8h}f�Pm&�]Ny9�
�W)��O�p*�$N6�3��=S��n��������|��߰\W��L��Y�_fd��lԟ!(��:T���R��'ts����J��{�}����Pfp{�Cnq`�V�0�%�g���k(��"&UZ����mZ��.FD	��j������>,{���{>��lIq����+4��˦�"�l��bՍx�M�Rh� 5�q�F�l���UQP��mY�U��n�>S$�G"f��(��ڊK��?����MvloeGI1w,���%�&T��N=�fܳ Uǈ0��ڪ��5~���'!�P����Vfr�kq��k�e��ج��8d_Bx�8�i�D��� /�G��q�}�)iѿ 3=��0e��R\;p����m�f���ɡ���o��� ./�ftm9cq&�(݊�Ł��n ���۝3�7�n�u��Q��O�7�5:�ݑ�����R:`ϕ������\��h�Q��%�Z��K�������!. \S���t��?ibk�"h����ۋ*�F�-xjL�1�]s��"LQ0�����`<�>�
�����V�|tV�8~N�Y
E�Nt��ŋֱ��e/t������P�Ʋ9:%���8��I�\<�Qf�0�y��ͤ�i2�H���B����gŕ�:�TeL�H�2�����+������<1�$��}		0��y��qH$�{4ɵbd�1k|*�J�.�E/�Xޙ|w�e�i�9%4"���9�mG���,#@�X�d:�p�%S�	M���\|@�����>i{�qY�X��Ȉ�Ϯ�hO��-0z�2��YR�6��x��_�_�O��j��|����Ō�X��;�����t��Z�Є��U��m��Aup�<�I��b��[b�y���-f&\	�y\�O �L%�iE~��N %P`����X��e_<{��W@��z��;�]��~jmB��3�&���0�H��n7sX������5]�F5 '���U�B� �0J.�2�>�����/�Wj9=��Ҍ����7D�r�+��,;���+�x��h"i�bٝi����4��F�wG�7uy��1��p�S�7r$����ʩH^�I�ͽN��k�/���~��ԩ��]�x�W踒WOwō���#Gn�}e/��(�WK��Pɱ����{V\ӟ&�d8TvE.��筈��d�-�K�jlA��X>Hs
�����f�"�hFj���f�R�K�0�ע�������ɷ�Q���z��'By��W�媎�\����6%W�JQ���w�����JW��P%;_����]h���9LJ�}N9�:��N$�ݓ��}|D^ȒT	��8w&�O���	�
9RS����*X�;����f/5��1�d˾���p�¦��(5$M�9��"���12e�=��PRۖR轩�ļyQ"�TΫ��H��cMkaq\ɧ@��2{!|��܃\]��:�Dz1+/�ͣ�� �܆i��4.NG��;Om�sv�D9�m�_�:F'���+,�z��ƥ3�Η�e��D�WM6�`\O��?W�t{��(�_P���-<�����&qU��c�) �t3Bw� ,ϲ�Yme�H��]���k��W�
/��f=��@k���K�gU�}NT-���q=G�_;��������
4N����k8�Uj��j�0Y	G�������@�`��s ��e'׿�?t��۹� ,���Y�n�?������
�S3���`�X-��UU�]#-�O�HA�I����]*OW2T�	-u^����f-~�qb��l5z���C�;�����Ĺ:��:k v��/�� o��П$�V>+�hX����# ��N�!-�/l�p�P��{��#W��x���F,��ئ�^=�|��v@��3ӏ���gǶ� *�k������ӦS�[��EM. �Ff�'1�o�������սi��oEoYQ�J��=rTڸpJ�nݐ��W=�X���#�i!��Z���>�_"Tw'G���s�7Un�o_�$R�����F�4E2�����l��h�(���_{@x����rخ[�isAs`}k�ʣW�v��Z.IY#W���7?<��V)
��<�D�Mةm�^q�1�\n��|���R'�7�!;Es埥a~��$cQ?�vR�@�*���^Z�1�s���.��p4��h��T~Y56�A��Ae�Y�%�ˆ�
��(w��^'q�v�=(��] s���%f��ˀ��38,5�-|��ʔJ�җ��.Jq�TJn�<��AO#�M��@1�T3ʔ�-a�@q�f.:6���_\���;����k�,n���@D��P��m8n�A:�T���E�����X�C%6iJB �8�ҝW����jN].U���>J�{�����u/�k�����OaŌ\���j��������\�{hK:t�b�q"���򎵣w��я���54�������[�%�̸�����z۴�J��M�5yS�>�p:V��u%{��U�4[Ԍ����ކ�7Ε$�b;�u�<E�5��bNeŧ.&p�����H�S�U*�6��
��M���W_�fD�Z�W�:���.�Q���,�>h+��=��VL�&��:tOJ�?����i���q7�Z�$�3� �6����m���O��Z�E�P]�zܥ�dHd���h��S�&�-���h]$;�+tx��G�\��� ���g���0�@�@��̞���s�&�S-8�Zv�[e*�J�~O��&/-a\FѪ���ڨcX`�z�w0�Be	��`o�?ED�4h�	�d�������y=���ڤ��LP�{/��;{�qή5�Ou�{7:L��+~�R�dȖc \l��]ܘ��C�̠0af{���6}5�:|	��z{4	�V>2��X�2���1������aJZ����J���?��Jn��F-��b��]_�ۊ>m|������{z����8�~�`T���Q��=?�\�bg�ax ]���h°{�u[��P܎�C��w�s�)��m�a�x��ѷE� j�|P3��M��:����0H>�-�њ�[�&YZ���&�9�*��0��w����W?�����d�>ϟ���8����m�ycI�DA�0n]T��������Y��^�6� /�m˿�p,ók�g!��Y�c�x��kH*6)���)V7��*B�-B��k�j�A��S��)�C3����c^i��!���-��3Rq@6��>G�*�h�� 1x�q	ؼo���;]�'�j~pk�/��.R���ĵ�h�K�A�!0����N��*,ϧ�kԢ�f8��)��d�e�ެ���"a�����+Z��o	��e%��e��O�"M�R��b`�!�9�H�⎢Nz���#0���wd�(����7j�œJ�)j�Rf��Xwiq�Gq��<���U���
��F�-83�r�:9�/g'^����g�[�ݖ���
��l�}�4�Ⳃ��S�.�j]""���4���y������a奺v��e�?�5W�V�gSu�$�>�\�dn+�	���qG���W fI�B��!� �T�D�X�e�_���I��D�P@��_��DA�[��`�F���Wӣ���I�����.6�3t���C9?,�
�1{-edgW��}v���N���Sd彝W�{��C�:\�3��vl[h6��#��Q�f�<l0iXı�*)%?S�%�^&x��D!x�d��N/*i@o�$
����4��7V�^]U ��]w1:Ş�� ]�/'�-4XN{��e=���[�B.Fnq��ܑ�ʃ��:�!���Ć=���	A5<Rz-Yzə���E�!a���":�2UDO�d�$�Z�4LᢿVW.�&���B��?	2����;]%���� {7�f�ҩo�LT:�f���CR�ϗ�=��D"ôޘ�}��s3=��ǯ�)1}��\>��ML9E�>�$��T}��f	C���@L���}�_.~�#5LFf+|j��i"�Ѕ7��	��^�1��$�R"Y$;� �}�q�PB�����H�Z�+��k���D�=Ƃ�l;W��۪^A6:�
BH�z�1"������0���@���I8��؉�h�!=������$�`�9ø�Vp%=q�k��m&;���c#��H~2��m&WY�h�yf2��YW:{7�诎F���gIe�o�ii��W�G���_SR����X�X�Q�{��j {C���e�T��Km�fe�V�����j�|7� �?�)�LT>ne�7nR������vȊ�3��M��|�7�AP%��kM�X5h��3�|JI-Y�+�*�X�ZyM�]r�W��oM��T��u�(�'�wj��2+��@F'���]�^<_<ёJ<荋����=��V&m!��Ż� �w�ѫP���P��L
�J����	��K�DZ]��D�M��{5��׳F��V��;�"|E�9|�Q�A���Y�.Wpo���qI���z!9"��XI�q�b��6_��(���K����t�/�`$�!����x��GA���WB� ��{$����.v�U��q��t�XIL����kEc�V�Ϛz��Hي�
k��%���Ҙ��-�����游o���dH�$�UE5O]J'��y.����@g����y����ƥ�k��D�?��8}��3ʳb^��?���'�k���	�>��Vw����q-o+%���Ҧ+�y�S�wFT��������g�P��>a�?��,L}�<�XO�{����^^91�J.j��pi̯����C��Q<ݗ��T��@#�cX��[��M^r�ݧg����:<��5�K�Wn�R��$�bM��H�f dA�V�����[(�4��a�����:V��:�0���fR+�
�&�gH]#{H��ʅ��P^�|�xܮH������j�8/,�E,�*�3\`��F	�Vlq��YBo�,� ��}Ν,b���
�����1b𓆕��?Ç�M�胥�uE7�ǈ���ܮ�ޏ�����p�>�&�lZ�l(��*�e� x��6��Ҫ*Ga�Y�d��_�^�P|��XH�p�4�g�;X��p�����hʀ_��ǿ�ޚ0|�ߩ�b�TĜ���\����t6��aR"��o3��L� JB�D$x�8\^����x�O[��riN��c���xj��а���`uL�L�w���)ac��S���A�^���Qy�RRn��i����x�v�<�Y�L��T�h���j��	�w�&>��L���ޓ3�$�̫�$��x�zs%�g0�����rX���kt��F�yD�K�zݺJw
���_�0�i�!�Os*�_�nˌt�̶��b|d&���{�R��-�Q����@�妉�g6b*���b|�ߧ�r�<\1Z��:�xG�P�c����L�ֱD��|hey ]9���BxX8�S�>��tn8H�϶�7\:�0I.���A���� �J!=R��i]�G�|���#��ע���T�H�8�9�A�@5x7��|BV��,T��y��\�X�G�\G��7쵹?F��E���'Q)/:���;P"�����ډn���#I`��ۧBv��j�"F1b��ȱYF/8|�s�q[������إރ#��[L���rꆐ�~����	��&�k�B�Ex���θ�@h�񽟲3B��V��X�#���Hҹl�Pۮ�67�`k�/ZiS��0( ��N�RqZ!J"�x.3ٵ?9�;+8��\NJ�[��.<\)Ĥ��p�܎���W�O�D9[R��V�N.�-�j�\d�a���t�[�|�+y��Bj=${|�f�g�G����\8���`�s�vәvЂ�z'"?�
p����|5��;�e���>I{ua+DBT2ȹ�,s!a�Kp�K�+����?�um��$���䷣<�_!�ō���]z�&�N&d�vx
��D�7���($�վ4M�2:�Է[`[�x"�?�T��m+����Eylk�jx�t�ke�bX��#�y�0���0A���q�FR>K�u�Xe��L��]��� �o���/��c��ѳҳ/mc��{yZ�K/P�-�p��?o����eFv�Y5ܷ{5&�6?A�vGoe!.\�!@�Q"�	���&S<�:�SK�:I<�8�~k�c�==$bP�����q��݋��}��_��c�!,%)&�H���ij	V�2Z����	i�q�9ags21}����?7�]>9#�w�Ԫ�9�4l�o|��C�ij����
R[G��B��i�=׋�Ȼ�k�:1\�����
-�ڊM�âH�)U�S�1+m{´o|��#��INE��sK?gFLѮ�C]rk�8݃/jc!�yN�!v�yv��
Kwv�e��T�Ł�F��O�d��,���S�)g���*�ي�5��I.�|��]t+\	Y`�M��G^Aӵ�Xn:�#��xXB.��)ِQ�c8�i.T��p�<=���g����J_�ƐӰc����3Oڃ�.��DU.Bdt
�w$y���u,���}���@�~[�#|��ѯ�b;yx��O�-�C��í��]���{�d=���<*]c@?���e8U�OM2i5�	�YB���c<�g�o/�t���}�D��%��J�l��~nKe�3�f�S<��,�'\�{��lc���j��g������Ů�ʲ�Ȇ�uz�a\<�����מը�=������}�g�����,�'M#�P)��+�r�l4�
�!�Hϫ��?ڀ@��,�D�Vm4�4Cjhw�����;�����u�u�8io����X$)N�z�\e[�K��F���ۈ�����Z��*s��q��d;��-��#{��^LU�Z�y�{.��Eź�����$L�AUD>����!�-{\�̩¤��ݜ�-mL���6
�V��*e�)0�ǏT������]_��8
�]E�٪��P�,}��'����g�5dT~v~��	��hZ0���c�(��h�xy� ��J����P��ɞ�.[���Q�;�Oe7�-]�s���a���p�D��}�0UWQ\����kd0�����X<!�U���g0૞Zd��-
-�6��+G�6wú�\e�5׵W�f��X��l0�.�}}>-3��P3K|d��z�Y���N�g�gQ����W`�x�9���4#���Q����:����A�t�����]��M�$]����L9�5���& ,�I����^Tأ������Ԯw�t�Dj�sv*$_��nz�PX���"&�}@�i���:~��8}#��f.�w�#�Y�<�!�����Ho�$'�>�g�����_�i}$)�e �HZ<8��a�k-5����b�( �}2�x��.ˈ�@�:��'s��W"[`��6f�]3n����
�B�ݯ����p�>!eB�F����;��+�0����6K�L7���V�0(ŭ����	>[�O�Y�_ȫ���b�8r�s2�%���,~,Fp(|dN�$,!$L�<�/`��f~@���y���2���6�6�$`5�.�
��A��f�%���>1�̧�P��W<Ʂ㮧�3�n���/̊����I3�-��AI�� gkcx�):��Y�.DKgm�!F�	,p7�Ȩ7:{eE�6d�(���Ă����m���%��e0�~���+&��
��9.S�|q��O+�p�8"���7c�G�Q��?jn���w��;��=����|����ßwFZ�e6�;��9]��9xN!���U����6��!j~9{�Ɲ^�!b�w�!*��T�猕�43����Ď�}����ф�����b_h:��?�2/��E	�C{5�ju��/������Gpo]�TD��g�w ����C���(��E����fzɢ
�%,�'�rvՓ��т �����NA�Z� �J΅i� �f�-�s�D�8@J6�6$�{3��9�\��f�{�a��'%�:�-ҍ/HrL?�Hl.U�g�P����e"Gj��w8�3� �%�
�Md����<��]r��l�WA[�,��<>���Z�-��# �$�nF-�B�����&=��*��Yh��	iwyW3���� FQ��/�S�)Ir��<���I�԰���Qe��s�XN&�����(���M��;��'1���CKc�ɴ�*���t-��"M!��p=Z�����Xkf)tH�!)��Q�B�(�i�����c7yy.�TL]��[׌j��S����4�4'�1y��U�!�����x8
|�i�]�'#4.f��9q����+�|��a�4T􇭺mĦ3c
����7�� ��Z�(T�g�Ì~��q=�B������^W�鷅�>i��Н��'�Z��ϐ���^��˄
�ի�O��m��y�B5܋�̜ԡbB�8���Pӿ�V�&�e���vX��Z��u]����l�s�yT/�d�<IW[d�)æ�r���<G������.�Dr����Ȓ�;>Q\D�[��_@ى��J}8,����Dc`+� 3f�.��!���T�Y7'�K˻w��%e+�L���o颍/��(�1�?���@O�,�4Nt�.~rE��r�"6�j�c��}pY�&��8fw��O\���
z�mFx��]�g*�:\���*#t��C�Z�@	{�"ԩb�T-]>gTR�79���Kgն`�B��n*���l�	�K�~�ȵ�4���a+���-?R��U)��X)��"��XA`F�5Lь�'\mG��+��KO�t���s�1C2?�wL�lc�E�$�w���M�/[����/���4��pwm�j���0���:w^i�����>��92�i�p5K �����X����;��j���}��j��i��O��R��D�2�^P�
��/fuy��U����������A��i������y�NZBF���>7�粕��L$��&�d�;<�9�b*��i)����>�G_��,�G/�//'B�������buV���2%�t*�"��	�;��a�h�.56����[4{l�.�w,���bh�ԭ��0=R9S�3���$���A�U�cO_g�q���,7�}��J�����Y�8�8o�l��ڇ�k	����
�%�k�Jv/llgBJP@A]�/`�-T�Wy�ΦJ[��ݴ4wyLJ9ds���p$R�؎������Ya����'&� �F�eY�ꊺ�1g��uw6r"��5ԫ}vbm#v�f�c���in���p����\�qA�E��4�z�������M��l�� �p�5��D�I��֙h���j�*�W�w-�E8Fp������*�G{�h[n�H1]���9�y���`��jՔ�	�j�ow-A�(R3P��!����|T#o_wTD3���L��JV*���-��?�¢���7��J�e3��\��yf@��4Za�@�f<쫈H.
V���"��}R�2U*�ZBSN�=�MsF=3�`��u`�Bƥӏ��Kw��Y*R��%�ͦK���^S �owӦ!4@zL_�P����)V������؍J�����4/;L�4Kk��]�X/���Y���@��D�)�i��S���9-`��޾�R�$����G٥{���ź�C�𺠪_}c�&��l��{D�2��>�?`F����H��i!�#��� ;��*os��G4����C**N�FDGb���5 ��SJ�������⡲�6�>>mP�Zxĕ Q�Z���#�:{��ЩZ��r�#F���Dm%�_�xYZ/�����M�"� �`���\i��s���B��z-N?�!�=�$�aK?�ӹ|�E��N��h�p�h���G�2���Zn��h��7�PS���d��mCk��]=�2Cnw2瓋�?��5^�m8$�c� ��JT�
����k�L�#��jYs���}�����0���l9�Q��{�{HͶ�_)H"�^e^�ӇAd��/�D���������D�݁Q壴L8d{���^�pP�f�ftF�Y2�sԎlOJ��3��U:X*H��5��,��9�VJ	�	?�ւ�1D���m��b��։���#t�;�x'�ಁ�ZI��߰''�����|��{?�$Lq�Z�&�M�+��������z6������͙�� �P7���9E�A>|�'�ᙱ�~�J�b�Mۢ;�Z�GĦش�}��	�ј�>�^2p���^Q�pOH�6�VR�w`�=򢶕�� ����aR�mu�Y:���۶����a�������r��^�n	2\�0b�[ͭ�Y�Ģ?Bu��>�X-d�d�G��v?�%��_�,CM��E�$r��\xy��U����D�;d91q���r��V7�H��O��WZ��a�s�����{!�$����MJ��=�R�7;f�.M��= 'qd8��+%�Kuמ:(��՛�q>׷�Q�����}j:�;����Gf�E<��uFHC�z��;s*g�xQ�W�k���oNf��ׇf�5�H&���s���{��,��XI���J"��iY�<k�t��;E���]����)Q~l�-&?����z�Ɠĺ��T��k7[�U����}�mi����'�{�h�++s"A�goK�f
��h1�"ޥ��h��+��F�oF��G��`��g�oz-k=�!���/*��sl �Op�C��(T���-����GG\��H�N9���V��=A;���؇�ȯ��x���\],����gp9��t �s�g1꽚���a�f��
,Ozu�iSD�q*���L�f�@3�W5�2�$F��K��h>:}X�\}h�yuz��E<:gM�� ����,����	 ѹ����(O�����5,�Ar�{GZà��F����:~n!T3���B��ݱɤ��R�z�n���vp$��Ƨ�.ʄH�B9`7�>?�0<�!�6;m}\�p��Qf8m�8�W���$|�At8�%ҽq�M��wөV�[��v��`��~P:��|/�d�ӎ������y���+�M������K���ٱ��)�-9*xc�Z��e���Ck����Z�8����&�A��%�X��>J�Y����)���Ca�������oN:WC��;�\�;�9�g�"��t�)�@A�=��d��(ۍIǴS#K���]6�둯�pXiU}ątl����+�LʔN�a�*z9�~�3Y�#ד�K��Ϊ���[5�s�&M~�O�6i)}��;pL\�m�)���H�0�B|�vY[M���m�=x#fn���P���!�@����>X��&�?V&dwĨ��8�>T��y���T�k1����Kp��<�N� ��U��e��t��R����� ��	7Ug�vj����K�A��/VX1V��o��@�-�����2����k����ƈdwh��iC�-�P�7U�@W��
Ҵ��f޾BFb'Oȩ����s�ܮ���廊p!_y�"����,�p���9g�/�t�pf�9hy���Zm#�%���1���V�Ij/��؊�*�dOo���H�(�R���+�=�C�	�v˟gf���t�~��<�J���l�f'k5�=}�ɽ,� �t��CD2rbW+1�x��j�zx�m�0&L�}Y/�C����`�X;,��jo�܆p�8�����*�j%�P|HD�{����cϭ���o�w�=u��3����G�G��s�PJ�I���\����^A�d�K�e���"��O,������A��D�/�]���J�+c��Ҥ`�)z΀f"�w�n�|�x�I<���X=0ᛙ%T�?�ط��Y�s���+�o&Q�����%�}2�kv�Q;���t!��R�U`��
/��-�5����C�����uBV�
���\�Q�2`����9#��q8�g�c���si����_`D���
�dI�Ǖt�!�R�T�����1/uY�8'�u��5u��"UB����g�ykw�� l̋�Q\EJtW����7�^�1O�\v�)��/��ѦgT��FBwiF�O}���o���mu���Ѵh������W��:�
�3�'�*��� .ni���;gw�ҫ�^�.K�4z>2���
�zɻT�A�a�>���&� +��沏���&��� �d�_ߵ&�f�����a���]�t%4��S���^x	�8ib��1�s���������0����p�|'��}�O��po��E�i�\�6Zt��2���Rw�r�O�#y���*e�/�0&��0@Ŕ|/��q�^�Sı:���%d ��m}M;�����K�=��{�^͆�S?�m1'." <��0Į�\ݙ�F�d���.@X��Tda�&�����T#_.�������8Bق ����D���]�8�myEt�����@H/ SAWp�o;��P��"	HH��F�^`�=�ܬiCj	��c�U&'�Kɍ��!��c:�����a�_ǁP~x��^��$	�����>�)C�ko�"0UĈ�4��/�D�2��M���6�=dH;�M�]�)�Hk	ty�k(���I��()l�u��A�����@d���~���y�w8�e�~;�vEEd���O!�\�v6GR6��\�(�掟PY��\�5y������D�0�'d��+=K_u$�z��cB]���[��9wGf~v�5�\MXk&zS�_7�Sz] ��z�I����u�b���K7e%��B�e-u��5i�ec��%�=4g�?��Q|�f��մU��E{���LUI](�h����m�ќa$6�bӠX��WāB"~�{��Ή�ӏ�~H����X1!r<[��Ϗ��aJ=@Z�-�餢��JqXn��8ಋxW�ԴT���BE����s(��/ϐMMnӀ�+��co��qC�h�5�a�t�� ��Ѽ��S��7����i7�N��G͵�~)�͌���s�U:>��_l�c����F�on�@����^�;�\��T�ek���L�}��N�n� �_�u�[G1{8k6���p�ߏ Ѱ=�Q�ap�ܚbQ��MD?`0�t��*7W�{ ���{~RI8?Ԍj�z���%��->H��6��|���Wm"'� b ��.k?�%���˝�Cm�p&��Ѡur2�0X��1@� �_S����nS��bSm���Vߩ�jmƾr��	�5@/a���[�A����_�U$�@1$�H8������Q@�)�ad�hWKh�$���e1��Yc�)�k���{�$��:x3ި@���w��y^�j�X0_<�9R�)oa�q;G򫝀��SwDa��Jm�[�v�����|	���Tg�/c6�3��7��؇����!!��d�1%��-�
</�z;>Q���ף}	���y	$E��7�b��uϤ�l^3�i_$���b�b7$b�gTK�����%�+\ c�_��;-��.�LF�t?.�����n�pf�"�~����'�F�v(2�J�e���Ԫ2��{�����dS@o)���o���`�9,��<O�*E��8.�4Y��,'���%T���,�u�hE)I#��J�8�!��h�g:辅��4��ή��6���_�ALy���q�e`��~��z�?{��/��[�[u���RҍY�//�e���r3�[��5�ogG�w�ҥ^��Y+<�H��V�ĳ�ȦT5�(@״Bw�VrA!��6��8�E�E�"�c���L�d��3����n�ݗ|i_�._�C*Z9����SbM�7�C��|�%�la�#�V#�=Le7l�l�?r�>���h�?+Y �[�<�w �.A��GC��A|�����5�_����J�=����=��YG~]�n/��YFZb�4�<0j�����f
��OD�_�H�1TS�M�c��~���k�Â�V��e��4U�C������^L�xJo��#�I.����2�W	_�6��%�������&����o��N��,�@7��5�c�T\l\~ύ����̖g	/����c��lD᤬�ޚ��L;��-{������5��f����{�~z�����`���F�՗�3�_������h R��O=��F�Q:�*����'�3�6��e���\��|m5���j��ki.�����,�:�f�r����񗪩א\z#���2�|�e�J		�xY��}�S�sdĨu��j8��<+F�c.�]�H�>�.2�n'S��LJ��F� [�2�
���:�+q��tp����Ѭ�á�����PnV���$�=�}/Sfjit�ޖ���I�,�^T>�
{{�#+&�ʖz���8��U7��="�*7���,C~���]�
 6��7��8�3�M�/<鰿-���I�̜�ࢇAA�&&�@1��J��a�E&. "���.̪�G��֚�ҿ�%���9F2�9Kpt�9s��]�~�@�k!���h��M��y'y�3�!IEp�v!62�κȷ�ax�k�oY��lM-��b�HQ�!��v��SŅTq���|�Yg�s�KR�v" c{�9ak/������Sǈ�b�1v�J��C�΄<�$R4�T��;�6�؅�UY��_��+���+B9��ɐ��k��;Q49�}4�ƿ��<�蕥ٟ�%:�Cv���~�7���2m�1s���F�5?��wug��{&x6��q�Bd�R��V��d��s͟좰e-x��u�.�a88�j忕O�[���ğ�8;���o���[�4zw��������fqǧ��T =:�m��32�"�E��MH���9����rO�;�������Us��ڼ�tJ�{M_�xG���ec�ot"�Ez��x�z��"b^'h�%.$i]x����&�)���&��ł>z7��>��JA���m�K[�s�ӯ���}9b���E�5��6Czin��I(�e	����_�0�*5��=Æ���Sq�<5:=�ߞ'T��Z�W���V8t{�y�^����.G�j��*'w���"J�X#z���%�Ҩ�|��g�V�W���Ȫ�pI&T����IR�5�5\�8O��j���'�I����	��7��F&� �@6�(��>p	���s�a��]>�Cd��3U�N��\8�z����H����A���+S�tU�3۶�c����9<5c&���|>�ɶp�	�w�����S�0o!Eı�N�(1�����\_G�媰�T�1)�]F0� �ߑym�&�!\�~�f$F:&k��{Ed9@�oƑy�rB>��wc�e���U�BD��V&�1�c�$ x�#+ӕ��Gw�CwlmJ/���-5�M �c 6�6�Y�Hڜt�5uf��� ����v'����}½V��ӶpM-�!q.%�z�o�!x��Ͳ��eM�Es���ަ	nx�z������j_<3�(��)g���_l�I��;���aM*���"��X�����UU�]�?��׭7�>��44]�k�ф7i��輇[��\����E�f��e�gևlҎL�s���j��K�?)u����c�(�b+�|��*��V�k��	������1���&gẕ1U����_ՃK�
��6�2�
�k�2��ûֺj?��_|]�*+ogjDlP��G#I�aO�}��A�ش�n��Q���ī�3����C'⼭t�+�N�7�s��4h����L�n$�Δ	%���s��Z/������Q�hR��x^eA�[���q�Q�|٭����֮�O;�"+p4ȯr~\��+6^!@�Z���3�o���O[X��4�Iȹa/I���.p�K������'.�D8`�r���v���Z`�҅�to��QTq;�|Bo����}'~Z���
���n���9�(���ƶ�C���?�OlL��Vkj�^F���V"�3f�/�c�/�1�`]
^~(��1F��VN% �粶�o��Y���<V@r�Zi�za��(~,/P��Jޞ�	�Dm�R��-�w������V�.���a������9	UQ�f*zL5��'QD���k9���1��d�_�op��2xs��������$��E��u K�C��$ۮ��L��}�h3I�L�c��oU�]�'��v�ګXUk����\�"���$Ň�Oh:�I�q��k�p��������������k�0w��w�\7!R�\y��ǎ�՛�e'|j%�K�YO/����	����M�!6�'�0�I���X:�Ae R���$��4�d�j��x,�����퀪7�T�	[��L�ݣ̋�[��<K��M�w�v�A��f�o�����nk3�Uy�5�ȩ��<�C�S����F�Ӎ�M�^��8@�qwG#?����q�X�!=]K�s!�u]�ͺ2�J
r9y��.s��۞�T����I�vw�&�(�@u�oLq��T-��b)B�DX�(+���� �c�Bة�����ǭJ���0 �\��(E��8�tY��݂�R�P-i������j�+�1�Lfi,�d���+}q�L��ۂ�t"��\� ]DZ�E� o�V���xZѠt���՟�YLXT4�|�p/�J�������+��8[B�*_������= ��"̂��� ��L����I��}ٙ	���0��z��M �Ј5A��NO���$	� X3���<�Jo�c�"O���U _3���v��|�F�ؽ۾L�=�X{��d���0�F��'�5۶{GNL�VmęC#-PxK7��>:-h��IW�B�IMceR�4VSrq�����|�V��V���0}KR+���7'���}1o�Ϩ�k(ņ�J�1
Wk�� ��8��1��7Cz�0���>3e�˸�|˅$B ���F�T-(t��}�9�Xn�ɮ(%bՈ������&Z@�1��H� ���b���}M�o��\��=��t���Fs�nh_"oҞY�0*ٛ�G���L,q��('�+_�CD�w [_I	����p;�,���}�T	g3g�_�o]x�ʥ|�I��kD;�W�����ǅI��T-��-�It��Q�*�?X��ׄW�p�%���J���x��+�v�A>��?%r�oKΓ-���T|�O:hᄌ�	W1GM��Q�.+3`1�0	�V�
��r���"�j�!Ud�-�Zv�ǀ�9���N�tWK���ܗ�mw��c�� NR��@9z�l�{�Ο�3cU���;�� 5n�*��rNx�_?pjmp�)���\�͸���!��L��ȩ�탢>I��i �3�2c+F���#M)� �E1��n�'�1��ؐ($Nư*Nˤ��crnSo+���5�-7/9��2*��#Fv1ޠ�$�. @n\]��	VA����~�C��K�6���"��E��'�*4��qxU�Kƴ�����(���T�5�U�WG���e� �t x��led5��j;�S��ᯬb�.�i�(�D�&�K %xhd��k.�U!m V<����`��M	�h-. D��%� խ�TV[D��{T��z��[�x���d�a?����ʚ�ߴT$�7�O���z�
�0�\�����S���ӦJh�=�HM���sXkYw6P(��DW�IY�%_�c�Iߤ8>����r�.�a�ߙL�5@���Qbg'����4#�����(:�;}���xmMm\�gόm�s}ːV�h�/�2�a��[Q�����r��^��C�lHEjaoд����7!Y��ְER�	�6t��MDXJ��@"�{ $�UQJ�-&�3�7+�ÞPR9���,�YՀ��~��3.憗�%v��P,3K0������.2Z\c>�#�.2���������R�*�L�YLۄ�׌s�7tҐkm�p��ȡ���4,$����-p�=��˹�V�$`]U�
A�_>o�\����V�<tѨ�!a����G,4τ��I3o<w�9�ūI��aG��-�jz& }��(U����Lտ��@�^�ڞ
��`��f��-vh[4�fۈ�hN�,��Ň2��jx��?^���hـ�;\c#ގf0�Y��IFz���w��4�j��>�D���ovwq#���e���p1]�H��-�U��	h��5("F�	���Tt5��	R��-�� �?+L�]���ŷ;��F��'���]t�-���������ă�\a�n���af�0:s�A��`�{pr���yB���Z�k��k�"�`X-\KA`�-x;#-QM�^BPBX��\\���2���(�`>��MW:���Ǌ��R&I���� g�)(�㪰i��%_K3u��$�VN�;7O"����	m�ʆ��e1����o�;^ڕ0� ��M�OЫjX��DX�-�ҽ���5�����G�����ʔ����;�Tx�皯7e��UB�!�B�Q�o+�γ=Yxˋ�J�^B���ւ��*�}�
�w�(�[&1O���+_���cJ&Fn>h��
�f1�YO~,�f8���pn������>3�s1���ҁ��ak^j(޵���򚊽�u�O%�	;O��W?=>���H4"q�KR�+͌1�#��"?�@��R�oe-M���mo��;�c
�����4�_/���B۳��ڢ*�X�i��P�	Y�ۈ�C��E���&���ú.F���%d��:A�]	!M�P���^$O=����e�%;�up�(6��`�ROyyT���7�%q(:j���>�}�!�=�]~V$���M�MZO�QHߛ"$�͎�L��8������ȓ=����������ѮnmXyM0�w�9:�B!�F�*~(�ѓx_/N^X��>�XW��qw��"53UN��[,$�ɩ�P�wz�PɌ�Rt�b��IP��ޭ���Z���̿Hv��i/b�=��Z
q��C�ufz)����,�X��PI��`��_�2��V�mާ��x��D
��b>�M<�" t[��u�n�R����j)i�Ѡ"�T2;A�Z&)��b��
��h�����>C�{]��zB�'�Ғ��������d�T*	7��ڙSaP�����5|τ4P$���q�����<���o柸X�� #�gӾ#4����3E�5��G^�jQ�r�t�~#�KMBfA����&O=����f���Zj�ڸRz8�y���E����U��rnΩ(��yW��=�O�ҝ~ ��5�14��4�X>��''Sk�BW�j?e`]$J�����4�k���t��^��q�[S�YP�D�kg�1����~7۫[��>�މ� �"�"������p�ޱ�EN@8�<� �����n�EJ4�wƂ����v�Z(��u��B~}��ō�����V5��n��V�Ň�@:Bnشs���?���X,����m}u?�@[�H�i���ɻpy8L��d�m�A�U���c�`+m¶t\&��f��C�o�F�����#yI�.oF슖.���du��4���$�\h�u�_�%����������Y��B���|�eY��J,���"h,k�l��7���� �3_���f
gk��%�c���k�U��o��#��~$�kw�4,}���}�]X�<{u0!�H�5/sG�[��0 ���(��ep�؃g[WW� y�Q�s��0�
�L����vR�ɬMMb��;e~u�}J��s�V����mp��|ⷷ���A�����7�L1:6�ϡlPR��i���G�A+.����buO�A՗A -:O���%���*c�����y�a���Y���zn��qWn��B�,λ䞮�������u��z�����*��R���8����pq���1��b���d2D��#�n�.,�D�{�?���7��4�jS���@MU=eo9��Alw6��	����Ԯ7�V��!Y$"^
�GG���`�������_�;�W8����ͨ��ބ�����i���
'&7�4Zv����<[Qi! �?��X}���A�K5s�;��$J~�#;b����������f�����DDFr�s�m��"H���~^<}.'Ԕ�
� `�N~cZ�ꒀ�P0Al�8�յ|W Ŀ���6�:d��&|V��r�J��f"k�tsW(WJ(���������>��C���V�8��	b�sE�#��N�5j�J%�F@u�	�\�BB	ґ��������`�:�H�h���h�{̒yɇ�0o�"�t�-�4f?C���NOP墛.�LoU�;k��:���橎��K̲��n-����ӵI_��&�ۏz��(;+��=��v��f���'��;�gP;d(m-k,e�veó��eU�wxD7P"y�\J]ܮh�*a�m�Yp���V���Կ���@����,��*��k���>�Qq2��$9�+�=&a�q����'��ZM��uL7�X�zq���A%�]>�ή06�����Bz��s{Ő�?6�	
r���$ƨײs�.K3�a?Ç�1��]�y���y�[?S]l����Ĳ<�9e՟�D9�.�)��Pz�͂���S�a����i��_��DhU.5og������͔zr9t/_�J^5�t�*/y)�@G��������!AX��<�t�
Em�NHǮr�861��Ib�����޼n�鱅�a��%~�n�4����s�i�v;�c�
�c���(�FSө���5�]�]�	Dkv
��،�>��u�m���؂�?�R�~VDP8r�{�K��d�ǽ��l�G��.C�S��2k$�-N��������s�q�eS�З�=n�(i�l�se�  �m�qð3�:�sHBc�&C���˰�B����O&jb��Ej��H�qq1���6���e�f��_�i�:G��{��8_��º[��_�wŘ�b�6�� �>��`c�6�#E�*�[ę� +VU�7����̊%..M�+�J����"��Y��x��[]q�`�i���3������&�7n^�e��~�ss޽;n0��x|���H�Ӕ̓���+|�Fr<ɨ�)˻���rs��6�����Ѹ�1
�FFd�<w$�b1��obt��ِF5���cQ>���K���3}���jn��`�и���<�"�
�8g�5M��fV\���T��Go��{�Qw�|�L����ܛs%�<����K��%�0ho�p��6)-������X�!y������T<���� ���/���e��W��<�DЁ6�1�Wی)ږ􅆆Q�Ǟ�9���IB�궱G��Ȧ�n#*�Y��&��#Y2哕4i*��3+|73�SkM����%H~��O��%��,���� �ޅ���hl���ddW��B�z�+�$,�2�ӯHg"�³��i3M�\#�9�k�n�R��̀����~���%�8(]���n7�uBE1
&C�!%��ۀ뺷�Z"�z�(�`?Z�`f[��#��6m�`����rmwU:3.��/q�9+�������:g[;�Jw�-�G���<3v�!8:5���B�ܣ�B�ݲM����o�|�Zn�}����
���'�I�92j"V�@�d/ۗ�L��@ke� 5�j�ZV�]�J�b�%���M��4��y[�st;���� ��ўz[�?��;�#��4gD
-��C��������q�A+7p߭�s�ݴ0
h�m]U�e�D2R����-(�`�Lz��D�o�Vmd������#��!�F��4��ny|4���A�����X�p���[�V��)�����Dtl��R��S^e�o˞܁�ez���
@��U�=���Y�6�����k�|�5KQ��RC�}6E/�-y����¸��Z� ��o��Ty��
~�;Q����i�"I�&w��eg��K-�(��t�w���1����΁�*�]  �s�Z�!��`�W�*�N�i��%%��?�GJ��pA	G���Z Z"y��0�B�� ��fS����4Ư�i�dK-LK���?��i��|ϮU��ݞ�E
m��)�����g+�#|q8����ڀ15�L�\������JW���=�r<)CA� +﷞~�Hf���Y>Y�����O�8`���rA�&���HY�5 �~����{1JI�݆
���G�~p!�?��`�Hh{	`�����qL��Dz(-��:!I�)��a�̋v��^=�(3�w�8�Z1��������[{sC1��ܑ��C�z��9����X�O��dB��F_�h�dԅc}0bbH>RQ���c����rn�:5<8O�r,sL�Hl
\��y�\���`ݘ�ksd�����Җu�d9�O�:��"p|C�3���>����?h=C����Ya*��  @�րͶe��b5klKg��j� ��|<2բo�-���1���Q��,�7��Gi�q1(��L�./`�$�0���������W*�u��T���(��j�M���`�k�<az8���1W*���K{5:���I�^cb��ѸG�Oz�A݇�Gq�xmʹ� ,����ACqya+��_�@Z��Jġ%�Qw�ض{�O�ښ�/��
�� �E^avF�<�{ο�8�</�l�6٦M�ϲh+Xԛ��.���D�ji�w�6�@P�i�z�7����[P�9�c�t.�ȤLtƄ~��&�a�R~����|�ɳ�>�6 d� �.i���r�;L��_u���UM��n�'���g;�_P�W���w�z׏5��=����f/�������1�"�NLw�F�w�|5OqzI��es�[@�(�c1��MS�c�j)�g���K�C.#���g�7��̃!Poh��aATtP����Iw�oY��G]�5t��6�G4M�a�<67��[��"f0V;BK���1�<�L�������h�[@�E����|���Z�����I�
j��k x34�T*�E<[�!ip+H�O}m��=u�C�è�2�"~i�塘x-��D!ߟ��{ǅ�Gu�w�B�A_ߨ���f.�%B{�V�b�)>�[AVTrdY[�[20��u�E(�"e����7�{=��95X�9���pT�U�|�0X,V���fN2'r'�h��0�ϝ��8�i]p$��Ȳ�Ɠa�O���.�	lͰxc�A�ڀ'>B%���PڊT<-t��bQ�:Ū� +9I\�>�H������g޲z�Nx��Wäw(�5[Z���]�qn����Tm���y]ם�0p|�[��$�Yfq����J!�:��{"�/�����ԣ��!n�ۭ�� �� �tZ���j$Q��~��/"���A!9�r���OI`�OgN�w��a�7���U����S�Z�n%��6�U�
�$�΂r���h@H�����0�>FuR@�Aj�C���3��"l�ņ�w�װ⇐`d+��.a3�G���<�kO��__�_\����>����
�{&9�%j_�N�2�O��j����q���h�+� s+%�b;�wl$� �E\�CW��^e���&�$~�^f�աF��GD��Hr\;v�0 ߭��������3���_2�G%�]0�Ȯ�!5>�YAgۯ�g�N��q �Iu񧅝�;��J�9���"����*�w��{�N�x����e��z�x�e!��<�PJ�5����y�t�̭�ZI�n̊>�Ƚ���eV#m�3fQ�����n�a�4t�����,���3�{�;�-+,�˝�%�5{X,�d��$�E��^��2ٶ�%�(\�q����3�F�Pz�Qv�S��WVˢ��+��ڕuL� r�$M뛟]� =.[�Թ=t7W�\����2\\���T���lܺ�����[����A�󏙮����ec�)M�hy�ʕo�	�^�vi>�bB��$B^b���9`�(p���p\|�y�Zx���w;�abw�cDb�7�m#w����5=����P,��й�N�8��x�˥���c�|*~:Sl��L�GZ���Q8�_�N���hmRQ��nѴ�xה�Z�l��f��C%Υ��3�w�����C�:��$#6;#zMV�3��]X�P�#�k��Voe�l���&ç�/.F�v>����.���T�Q����8@	ʺ�+����F��C�@�$LCp<+3r?��y`��vK�YV�~��V���B�̀|ݶL�3\ֈU8o]v&�`?jj��dU�e��	�%|OoZV-�i��o�d���h(C�I��#.�X*�ّG�M��������]�?]õ����9���:j�c$['��`͖�ʽ�϶���to"	%g\��yK��[<��C�UN��K�~5>,)e��k���|��|@ŦF2�˭�p�]K,�P��\�[\�K_[��x�b�F�b�$y��ǣR�(��nr���ܚ�~���N�o_ޣ�әU��j�csPdhR蕀a-�?�����Y	0�Ӗ��U~7��������1&�~�w_������ڽa3*(�/�2�`��
8�!���9��ˁ�`� �:�V^�Q���3��������d"��@�X溾�(r���掋�.��j��i�Bk	;�7^>�2pEF�O��  LI�8�Sc�<��^:;�iN�X;��=�"��ޱ
�b�y�J���A�f�a������п=RNcg'�.��ߡ~W2ʌ 58���t��~_#��h�P�2���o��5��� h�KQ\N��F�����i��k�_L���8{r<Ϭs�J��¬pKv�K�Nm+3CCq2I��h�����q�����&R/v:%5��,ш���-��t��$�t�5S����xPh��	u<��f������������a/z��F��ST�YRn��P��'�Kx�;�[x�˲[�p�䮛[mB;�~��\�o�Z4t�x�"�cw�A&!�y�8t��_��u� ��
�eGpK�b_��01�/���W�%L��ʽ��T����-u)���������Q�+K��v ���wSx�/��t ���*�vΠ=�F����U�M T!~���ю �a)�-;�xu(�Ri?PK��f:�n��H����v26���^G�FV�x�q'�5�x�i���&���>U 8�V��H�.~�ߕ����Y#�]�3�qB�"���ƛ*�y��2�Y������4��K�����P]L��Y�g�R3�C�e6C5�\8���F�R�8�Z^��� ͉}�{��T�ܻs%1��h'Lk:�`H�/�� �3�|,͑�q�.�Z6�|��W	I���Q��7el�#������RH�P~�{�貖����A/�h� ����c[��l������ٜ4�	noK�u:sٓ�Kf�w U~Ja��A�ч�,1��d"F�gy��Y�زdL���P��9\{�{�s�]N�?QZ3�#ܪ21+�vĭ���1���}�C<#F\'c�$�J�1rphL���5(��L ���4Wҭl2�2}��jԠ�W������g��û�O�uy�Љ�w�%|�*@���Hx�37@�?�R���h�K\��r��K
�mW��[?��Ԁm
;R�����gDYM�]���^���� ݆��Ț4�%��ʮ�9M� p�t6�����}C�~��(2
����rq*���hǪ��1�}_"�#����L�f��b-b������B�en�����Z�,���J'{�BCh;��lMp��dz}}e�����|�\a��B���o��{�h�noN���wp�ם�K�DTm�hN��/.�Vr��Q�ND�ZP��1�@�l���_,l;^o�����&�{*�:�f*��ƿc������.̏��]	�x���������cn|��8#�;��MlrӄK��F�DTF��8{�����褠W���R��ĩ�N7ޠaw �.c �T[0���j��;C}���N���j'm��yD#���N�[���������G��+ �9f�Yp]@�B"��ݜ��aވg������M-��Z�u���Ȁ;�����8�UIxԈ�u�'e|uw$�����3�a
�xvB02wZ[�ro�댦Uϰo� �J9�7A)�Y�
s���m�?�㉎+c���O�_��Jp�vЍ(S҂xW����;�H��F���w�k��4^�ٴ�\Y݃�RY�\%m�w��D�B��%�3 �� w����Ω�22��$�|�������n��n.��2��Y��s�z�+μ~�5��I
:��`�< �Z�m�zJ>�&�˗@�1f��p��Iב0��/ߌf���|��\���2MAW����
�>y����P�`i�����{�ݣ�	����3ԃΥ���A4��)	�	rĹ������\�#؋j�S
U���Ϭ��f�����Ă$Ҳ
h���:7��:;���b�'�ВQf<�d�N�fu﷥Ң�z��-U��޿�Q#sS��i�p����[�	���:uf�?���7j�28���2��+�6���^v<_���"�.Dt�dFI���ә����޸1��S �ɢC�u�(���k�Ƅ���O �xS-`Pj�v׵�ަ�k��8G�,��@E,g����/9:�зs�gw�VO>�DS�8K�&&6`��((4�����k!|pN���g��$�Fq�b\����r@�o��U�� e��ǫ��|�y����/y�g����S)8l����*� ���O��4;��V3:�ꁍ�܀�X훉A�J��,����d�.ߠ� �r�$���>k���>�L�ظ��B	��ъ�R4�O�o�Km�9G@��p�q���A��A;a�S|M�j�p�٭�fr��٬JMQ�T�eG2� �C�d������^�4�ċ/ZIE�H���j����ՙ�N��w��R�d躡:��J�/�鷺$�z�+=�|��A�#�@���˽y��$%jV@^� ���kCg`�U����ߒI��P#��@;"m.5��7F5�g�$��.t2��U�o�!����`tA���<қ=_Q������8e�����X7��j��B62�t\���K��V=�cK!�GY-$��Qp��;�'�������c��2�Q�o혱��x|�9V�v{�\ ��X/Y@Z�X��V^���'z=x��D�G��Pk|Rm#��s%<f��~x��Ǜ5=g {�Ŵm���s��C8�tB��g�[�*h�,{lE�ա/߷R�Z2X�=��abMjH8P�l�s��D�9��x���^B:��(��+�7��e�؃���Q�=N�.�:E�^怩�W7��0�H�`w٫�Kx`Ky��LO �^[!�
x[pk�2m��Z�ٖ�'�Y�J�L�I�ݒ ��[�����)��촐���(<��$�����É�W^��B�v�~�X�AڇyU�r�dnv�DW�C/��7R~��&s(hu���A���M�����<����+���t��\�X��JӖ�]����^�Uj���\ȅ���4*��Y��[d^��[���+}m��hB�~���E(��Wg Y�o����Btt�����M�&sR�u�pK��L7U��6ig���!8SYiK��2]��2���%>��/�49���pdt0o1s��q�O�2!P1P�Ǫd��tI1�wnlN!Ů��H��Qe�C�L���*�[��p��?PiXr^��K����,�RIT�����;�'g�h��0��;&����dR�.��{����cvn���z��Ǔx��;sX܉^y{4�=�������Vq���)���^��g�3��if�}���H��B(�o,��A�g�}e5�Ej(p�g���k���:�W��ͅm��-�ѐ��V�>�e胊�@�z��-����:y�Σu&�d����;db��^�[2l�g���w�����S��FJ%|��2����#&M��o�ֻB9������J���.RΈ�i�+�
b��ʘ����?`)0_[���	��L�<F�� �(X�	�*�]6ͷ���:a��O
f���ԥ{q�0��D\�Q�����"1f^�J�����ʜB��l�a3���+o�5�I�=Q�~N�/�ɓd�;�-&}��g���Z�f�U���=�~�x->�NUTM)�@��z1�%9@�d����-
���Ni�jX�鿁?y���B0���XFOp)"5V���+iM���u�hW��������4$m�ď����Eq�!⌦�T�B�O�8����&j�Ab���C���#l��� �籽9 +��e>E#�@��~���(����Q�sZ�b����l�N_��\�h�u���~��-�
��y W�÷L��ς5��f������<� �Fo1T�g_d:����7/٦[�T���&V�.��?��h��a	�(!i7�#�h8��$Ap����ؾx��NRAtx4f�eP��l��>JO�rwF0��&��t�CS�E��+�n6�"�"�d�k}|��5b�\39�mȭ��  /jy�u�e�!��LU�z<����-�:��.�bկ�� �j�Np-���z	h�{��Q��9�� �� ��ʪƂ�ϯػ��������K���o>�D��m�Qs��<��hDFo��VĤI�ә�1�i�������\�>L ?uځ�s8�������������H*�<@���7O�FЬ��1B1^���FzB�֨�8!�T�b�;u��_f
l ×GJ��!v���=�h�IOr����Yh#�����b=��eF�qLf*5f� ����>�"�g�|ڈ���l�����Y�*C��������Ʃ�����x�Pu��aC�P�f��4�J|�n��|kb~߽Գ0$HE���9Il&G��c��-\^���C
#�����:̳����os�g.`�<ί���aq���%�ʩo� 
sn�B�<F
�w=��q;������Z�cqg�/	�Ā��I �}�*!4�(�!���K�cP
���#3�GJ��
1�X���XI�O ���s�j���"m�Ȣ��3�SW��P�����_RC�Y��E�/�0���@7��yɤw�;1͘���&�q�]$R���xs\ߜ[�~"+ˍ��'��M���Y��?|��c<�v�2����Y��f�A�j��d�����;�O��c�4�%8|C�%��Q>��>r�a��\@���+f���k��gd��8fڲU���BX���E�A��̿��U��{Hʄ�q;ca֫򯨉�XJH3�T�K	�}=�@�aYi�~�rYV�;q��0nUt-��xY�:Qda|�S����CĹ�9\l��IE������R�
��q���	���&�]&��C. �}OO��z�1�"�-��|8)���.��c�a�	G����U
4*�ӵܚ�Iy�Q�[R���9T'�ܬs�1��-ɪ��J�ߠµ��3'��|+�c-}��́a@��v]��`�.���ߖ�r����v`QT\�MY�c���ؽHh����ǂv�9�ʆb�/�B��G9!�쌏3�f@�`��},K�w�� �8C႒	�]�EX�$�ɏ���vU�P}6��ʔ��������p�y��;a��R�\�b>Y���X^4��l���w�w<+_լ{�8��?����P�~��O&=Ru�FNr��n<1����{�ۅDE�Y�9L�:��_��N�po3�pR��
��f|��	*M|4�q?Յ�!��&I
�z�J��U�c�����v�qnT��J=+)�����D����-N�7�j��o�	�@&����R��罡�%�Z"D}�MGoe���p�*�X�y<P��s�s�ʸ 0�nao%TFp6�\И�p�^m�1��j�Rk����4-����(��.�i2�if�=kW���B�>�����D���g��|��~����Y��^w(��z$#�6���/@�d�rz�|HE  �$r����m�Ƽ���<�^8�Tx,��)_P�1�O��M�D�_�7�=��U�c$�Wo���a|���_Y'V��&���5���Р���i>�$�$J�.�3K��@�T�R��qD�ieD��7\�ǫ�4�j`eO�Iw���X��8�B�*�~�0����v�������ZUf�g�/�RD9&<��W�q��;oh0�������cX��e����joc��x��#r��{�����+�NR�5BJu� �p�@cY)+q����Y��؅sZd�*�k��
�ڲ��~��	9{�ז����8�O�y���`.��gPsL��O}��Q��55�䂟}e1e�)�X= r�?.$ՠn->L�ކ�d�s��<,�fa[C�(�+��ȩX�jg.�̞��{'��"�qE�bUȊ;_\���E�˗�B�Eݡ��*ϭB�2���SO)F&c�t�>iڧuK1��R�HM������m�	}���=b�Z���n��w�P4r��|�����y��ҽ��L���=����Y�H�vh���3BR��S�U�0$�vPMu�FE�L�2 �B�&4�����E�E%LK]����6��]=��;�+�/�LNa��:���	�fKx0Í,�'���2E��Z��Q�<х��Lzʞ ���BA��F w|���G�T����-���0�����=i�����	��Rw����ª�֫�����&��ګ4������Rd=�!(�?]oԹ�(C���o\������;j��>��A���� h� [���=m'�2F�v�kS���F�C��y�A���W�����K$�aΦ��������4+zB���Z��Ѫ�c��;�ҪY��4� �.n[�y��T��s1FH��4�����U?�K���(ȭ}�U��c��-�b��l�^q���p�n[�j�W:��0��)�<�7qNc�z�l7pw���݃�D���78��m�T�>���n���$I�*����Qυ'�-���<�_a��5�k�In�t}Ӝ<�:����%��枏F+h��-��{��*2ik4a���[�;��A�V`N����ÙzM����y�L]�"��;ά�:��s�i����fcɻ3�!��}����o�;fМ0*^t�z��UŘj�Hq���\Q�yķ�Y$�Hڳ�x���_��ܲ���Ow�����] �L%Z�@٘6�b�]=w(�csD?���NK_8�`�r�� ow��������%�;��
��NO�1k��x�+V�_��`�׋.SQ��;�0����	�Q�!���h�X$?o�$���"lc�|�G4���!Qb������T悫��K����cm�-_/�=
U�K���ْ�<Tz��m�
ӇWA���w_�'42��]$��g���

��K0FR��􀔜G�)B��b�e:��xVFܪ���a��%�
ɋ����u?��EC>d�8e<�'�y���]"�:!�	!��P��#�O�{��^�#�+:]L��A�+�_��WZ�'�
��y��+a�T��Dg�_���d�$�9/�{| �s�ҭM'	Ǥ��b5A�ƫ�o���k���,+����$�~mNN�l�S����VD��.S��g743.��"�����s���mٕ��P������JhrA�Mi�d���;����	y��r
ب��>���*
J��k���b����JJ�^9\,*��b�49`9��	�.}�C�MӨ�\�S�t]�
�c� /��Q���U(��{ �:ǋ��N����?�5ֿ#or�
d�u�0٪��I"j��� �8�^0{�,��;�bP�na�^	�<�+ ��l�V)(�<
�8"��k�}?�Y��w��@kv��BL;X4H|&}2�uqs�g�����!�@<��G�43��7%Pt�71� NŅ/{�8�q S��Zi�D���i�`�U��a(���PE-X��9)n5=7V�JS�E�)�Hg�	���qd�EY�񾱍�p�4p��Tf��������5���:f��{�������3�bLp���?<p�v�
&�[��d�,g�M�k2����3V(����h����n���V���4��׮��1��ê��T��
�� }5g�Ϗq$�u�0��hX��-��I^�����"����	_�ҵ���S�݂6��Ѿ�ڰ�.�+�yAyS�X�tb��tG��r*~��' �-L���7NA��g�Ƃӗ�L�e��)�)�An��gY����͗+'�a���<T���A>�$]<6�X]7\㔐N���ݔU��|��E4�����2ImIx���a�4�[�iV�c� fI�sU'��Y+������$���R�w���1g��Eq���8�c�pе��N��jc�3��W�@?�
H�n�|��`�"��n�@��4�.k���_�1�D���[{4�L`�̛�ي"^�BPP���8������������V��dr�C`P� ƥ��)�
�=�A;<��p��m����ע^��AX(΄���ی���ݐ(��Jʊ��%BX䴮��D7�lt�1U;��2'1�1L�<��.�X#V/R퇏ŹF>&1���޷{RJn�VW���{�sL���XͿ)�_�7��v-˩Zgtt���NzL�s�#���W�I�@p+�͸A%�EӉ� <(��ł,$<�������jz�(#�nC���TJ\�<H��.7����.Fu�_���}�C�c�?(�}��v=W\ �qc��T��
t	��<�k�"5b<�R<�Y��������+��J�T�0qXU>�Š���Yj�&��ͪ:�ZA�Nu�d�_��Ǩ v�ER�6(�W�Y�V��_A�]|(�M�S��������eW��6U��Ul��~P$:�P���*�����/���;M*�jq�̎_V���̴m,����`e79Tg5�>#(���?942��5����+�z3�qy�ʄ>�M�Q'�w���[��n���9���Bնr��,<ffL�SȹI�MT��R=+_�`&��I'AHy�S�P�:nٗ�M���,��a�iI�~�WjDgI'A�4��� ���);6�IƢ<���^&���l��M�l!��!�}��	|'I�	�ӹ@��0�w*�)S�њ3w'>�#�Fq��4�yh�0�o3"܇k	/d��\�|?�"S�W\�5� ɷ�V]z�Q�C+�5BA�K@�n�T���i�`x#��YX>�,F���6��/�*��i.�.�{c1RRb)�AڔK�7&��b��` 3(7�?%�@@N���^@${���{[k�u�ыP�Q�D	c��LH��wu<f�7N��a��#�*�k�Qk5���M����{�ok1C2]��wPm�nC��."�g�E���VAx�+�S�㑭k��m{�S�����>�?!�e�8
q��.=$�zT�ݖ[�����Qmm�F���eABnN �E�"�:6���ff^Vǡ!�O�2�%:��2)��C���a3'~����+D�m-�A�0��=���P[�9(0������6����C�)��?�,ȍ����*��	����NFu�_�˃g���|X&�x(��Ym
_�:�:)���?����� ��G��36gv���i��C2�N��t��@AE@k�DlxH5T=#n�1��Yu�{{_(�kg׃�>�t�$���S�IO~n�����K~��� �B����`���k�1�V�+:����v� h.b3�g٧Lj0�&�\�.�VVϥK��C{��vҸ.^
"nX,�|�z78,�f�y(�	?�R�:���q�,"�p�1���'L��,,�v��2pP0����f΄��5c't!�7P���8{2���p%I!j��ٖ�[�+rź-��A�ͯ��Ȝ9g �s�͝�oo�� cs�ls��ǁ�LW�����}e�z���O�W8��F��kr�]��l�P��ǟs9d����)��0�e�sx�	|�j�o5x�x��1n���@7��<K+8%�Ҳ�t#b��$7�Mn ��k09#	+sj��;<(RB�X�6�/7�8�psb���
qg�DQ��7Ɂ&��_��6��'���+�as�wU�ޘ��B��@՜�	���+sQ�~��:����Mߗ@7��1y�����p����U��GK��tp۪B��-��o ���ax]n����Y��2�O3ّ�݋��7,'�<�3�������wn*�m$��9X�v�HQ0R�jl���K��XMQ?%ej�IS4&���P���V�D4L6��m��3o?�vQ�Zd��>�OT��o`y����b�TU⮐粀� ���������#��=@h��i 9g3��0�δ|/��$�u(m��K:�A6�j?��Z��DƩ�P`�T2���͌����˴�gA�t�c�{�i\<��C^��X�2�����r�S���Ò����.��w&�áf�ċld!^��T��k��Y�HC��Z{!"C��!�.��VZ=�Jy�uO3M� ��u}�;h6�kf��+�w6T8����.|�(*�w���,��k�I-�{�Rj�c�X���dk�Ʒ��Ϲ��'p��w-�Ϥ�y}�!7�tK�,���A��l=��Ҫ-���w_��蹙6�2�B5�X0-?�u�絃Ǜ���.��V�@���ܛܯ���wjZqM���$(_^�e�`R�����fu�D���7$���L~��R���Bx�.Ӌ9�-_���S��i��,�]<F��h���^���� P�m-�;�bS��l�,��L�"����ܞh;N��?M�><�N�*WO���mG����2Ï�|���$�B�1�� �R�	F�pz�;N�M?�i(�n��ߠ�(��մ>��)��1'��GƐ���2)�{Y'��%���BW���F_\�t���2�,�?��?�E�N�(�U�z0!�6hl��d��kDZ��J>�&���#u��Ә?����W^s�:m �D��C=��y����/daX>��LO��ĺ�/�;w�6�e�g#����.�� �D �X�b����AS <�9s�^��M�o� 5BD�9���J5o���?�	�sm�A��Ya`��K�K�s�JzDX�2�uۚ�Ů`G��Xܽ���q�ȗ㏳vG�����Շ��cg��T��M�	a�|=��"Kh�3=6	9������4[G���v�)��T�le��?/ A7gb��n�Q�\�=6w��z)\����g:<o���HdJK�+&���"�$�+Q�[���^m��Q���I����85�iI2���{��R&�?������X����-�Gx��8N~?�xb�����]9�����}���A��9���U+rc�٦-�[��l�,��;�y��T^�:�����[��y93�-��wD���ޕ���|�ͺ^�,�+�܁�P0����-�GNg�j\�;`VYD�X4*r:Y�o�9J="L5��C��az�WJ��I�f�p�'B��1j�:jh��[�p��^B�s����C|�`���R�rG}���%1n�
[�;�?�y��JwN�v'�q[R"'���(�!߬x?��EWP��o�˱���/_�����A˿rT_�����Mm0
�.GD*ͩ��f�Hoh�ĩ'G�lf���U�9����V� ����4�� ��D��%�52"��߹��]��P1���vDŗ[��A�
���pÏ���B8K
�M'H��т� y�t�@GS_y �6N�?�r����5�52X��@��*�?�؛Z��'��%�;���#UI�-����lʰ��`\mtOq��d�I�����;_�����eB:��� r<U���&���)__I[x��u�#�n	zB�#�� �|j��iax�D�����R �G�;}��̤RC	�{�jm�jY�N����MƮo)Fx]�?�����sHU9G)4�qJ�׈��بA����7�BQ�%��H���嬧Xk+W�tj�d4���T*������51^t�O�Un+�Dd�+W�aD4��ゕ3�N�OHQH�qY|%���'h���C:��^El�����IJQ��TX�,�tP� ��4�K~±�l�?��6d�J�wP t�uλ�ԇ��u�e��]DL)��4�T�䨫T*&����R��
�d�W�s�eO0�I�G���>}4q��?mبb�vHq�\�@�뛺lѬ���0��gb�^���ܑ�^��B�~�����AK���Nd^F�u���؋���a�:��+�g;���1�kꂿ��"�m���Os_k��@5^��R�Cܩo�}M��@ �A����+YĆ�	�N�0�Fed�X��ڐT�p}���׊�:���)ŷi���錛�t�Rd��Q.�_�R5�c��#:]�q5fPOe��;�o�/w�y�6��Hu��������N�&�Rⴺ�I��6K���4Y�'��R6�:ڭD>)9J1��:R&|�q	u펯6o��b��y�+�\�>݄*5l�x2 4t.�v	~6��NIc'�w�_�|�q�vc?��d���9_��tv��l*P�L��צ��ԃvA�fU�x��n�Fo��#�Q="С�W$��`Վ�~nނ9��:� �Qu�í\o��-D�ʮ���Q�p�#u��VPN���_�e���0{�M�;6�qf�e�'�>K�Y��|b>� g�1)��L�%�k���V��z��zO�nz`�Bk2�p]�%-흾�g������R������Z�K�V�֎�v�C���,R�gԪ��w�����ņ�#܀q:�=�
�R��A�Y�g�TB��|ۨPP*�=��G�B0e��j�6%}�j8$������&M_"���f)�Uy��[j�G�Rvۢ��1Z�,��u�Adɴp�lc�	��kv�F��Q�W���P^��Jf���]�� ٴ��-���( �SK4�z�u��;�^����ښ�FO�-�C��ř�k��߀�:w"D&��H>��nռ? ��Z������Wv���!�MY:�# <�����e^�6��yn4��5�7S>�[��;�	ݒ�S|�!9�t%X�r�����+�Ⱦ/S�����/���2���ƭ�>[�︨lJ(�\7;|DuR��:���ÕDi��O~�9l���׍�oj�ʪ<��D��:�ݐ.C:�&Ҷ�0�	�f��T�w�p2B��yr�|��g�~/C���#�z1}�i��u��5�����khL�4NJI��|�Y�Z��	�>��db~�C2ܔ{֛(�DL�.�X�7���FDJ�4��IMW�E(�藂>��M@�ҳ��	�UD���`�XD!�=:������oF8�i�"(��̱����5�,�*E���C���^bm��S�੘,G@3�#L�J��i�<�O�K)�z�Ԉ< 7�l햻�W���6���L�{��toz���NQX�Iv��峲�-�-�� �~r{'��l��I-)�PK/��7u�xӢ�r��Z����U��D)��ʯ8����8"�˻�Sݶ��+��X���c��5E�w�-e;��%�p���N}���b A��EȆ,=��s��R����\�r'���S��^���P��``e��R�m��x	x�ͭ�!;/�B��D�����?���:R���Uu�'�D7]�:Tug%rG$�z_%�vV��D���.{B��8����UF��5ʃ�w�`���+3X[��Ԋ0�i.�JY����֚Y��C��\�)�l95���w��r�ӄ��,�ϲM�}�DZ��;��Uu=����"���Iy ]��(cY����I�\h��2kgOʎ��R1�\[���V��n<q��c������3RA������X��;{"� 3i���iד�OZ�W�w�5����=��p�˯�W��p`� ]��	�ѿj\��i4:�/��v��JTN�[0G�B/�
�C/�1N�-�m�G���OڹS���������y��Ҏ|p�t�LN�����K�SV�6A��� u�9�-��c��4uC�^C]��pW~��`����Xr�!���=\"�D�5��4���ʖM�+��]Q�����V�m6�L�w�s��Zz�..������կ�']%Θ�ogU���	J���:��8hL[b�A��V��䉆@��$�f�47�]�Q�|�]-�9Y(��&y5�l7f��	i6o�P]�W�L���I�����uJ����.�y|ؤ��"@�U�'|+�<� R��Z�[w��&7�$j�WF��e���9>�Y\a� ����(�f���Uu�x��v�ضd�_�-w)������PI�{9���F�C������.�[�rV����P"4���R��gI���۶ �#�t������TK�l ���D��=d�(*���|�կYP�ja�l�N���3�&�N���V_�w���\�~{r��|�&��0�T}��3KvM�ZK2����*l�HzQ�&�
��tY:�"��^�o�5j�\B��+��*ey�w�x�R(;��r��s'���6�ґB1A��
d������>fָ��M�c�u��SBx��AJ�uD/:Po0��o�nY��w��	�S�b\GZ����{�o=��AViT*��b�KU[*��r!}���������C|g�E��8��:�l �9���Ϲ<\&���Q�`��,]�t��"��c��~�9�'��lVd�{�N/����ݺ�,��劰�o�-�3�-�S�A��`&D ������=��2h�ă`�T�	W�l�u7�R�D�$��y�J-az�n�a/�*�,���Q�f`�i�>#'X��X�2}g��a�iwdҋB�cO�<Z��ZG<9~a:(ln a;T�G\x5K�+O�jO��a唰����ݑ%�maz�-U�=>P*�(�V{�Xѽ�Y@�B�(y�2٤��X]kv� bZ�k��{p0�T]B�Y@�"ɗ5Y�����'��f��4���i�핱�@�t9��0�I0��]�I�q`B�Q</C��?���� m����ヸmi��B�SU͚	��nw�U�l���"��c���|! I��=�zv!܁ջ}�$g�����h]��Hشl����A���._(�+�i�cŭ�)f#Z)7'�ɓ+�� ����,�9˰��8�͔ۡT��y�ے�^�s�q|P�@��?d��AIRA�L;^'�b���hHYe۠NsT�_�Џ�t��VJ���3C���b8������[$j ]5:!���vC�i��I��P�FMm���������������ր�>X���X'��2_Sp2�`���UA��o5�%�C`Cxв�5J�0�u>��op����eD�WgϮf�sw��Q�vR�fI�V�4[<�N�T���>y��$i��Be���{TP8���ғ[���W'�pZ��s��,Δ�1}�#���ⳡ]
��C��!��~az� ����aX	�q̰� ������+�/(���r3o����o���vE����t?ϧ�e/P�Q'�N�ۆ�3M']��7{�L��o/���8J�Ο�ld����T�G'7u\���.�y}^�`	�<3��5�*���iۄ�^�f���Oo)����t��>~~].�
6C-�?�`�p���5�"��JC
V'�yY&���	�,[�D�8�-*�PN�������{�=�\�r��ʖՊ�_VB<����}qpS�fPѼ��dB mP=���!dY���YA"��ݖv�
R��\�!2�Ĭ��1w|�ܱ� r77VK�x�j룁om��Й�.]�$V�:-��ݱ��5~H0������L��&?���ڕm:jmq�d$��Q]�1�K(��ۂK�@�ss^�!.���ܸy.|wWI}���m�����v(^w�|(O"9�|�._6@W֋S��{�Jb2�νV��c��;PR�q'�oŜMO�籠�33�E�F�b�{��Kwuwྕu�)y[+�0}FJ�ELq��w7�lb�������FI'	9���GJ�f���E��^~��R���d��+׎ ^?6^��Ʃ�v�A���QGBZ����mtu�ecx	<f +L)E��P�H:��}&��6��@9���E�:��D�ԯF/@{��b]����~

s����;�y�-Yz	
H`1*��3`��T��Sj��)^�SuPTl��"�C�S�`Q���uuΩ3���騈A��,��AbUL����@=-	��JA�9�%�&G�c,��U��f	c��W�`Q�V�V$=ř��>>/�<";��0{��\�9�~�B��,�%����^�t����\�,p�,��u�?���,��F�y��6_��)yU��O}�ZR���'ټ�h�����/g<Gk��z�}�/��J�G�:�8���i�S��ڙ����G�Ce��@v<q&��1���a�U{��7u\�F�y�����廗�V��j?�)��Lel��r��0u��?����P��R���5�0ۓm�T!/v�sZ�5��</���\��*}^6-�fI�)�8ͪ,�Ԙ2�"8ҭ�\�zB�����8�0�b�^0�k{z��5q)=W���	"�'�u�˔�%_�%dѩ�պh�K9�am�a���&��a+E�3?>�V���ۏg:I�J@ �6 �z4]Wr:j��#P��찇�	d�o��s��rki4�*%��f�,�1��R��M�1�F@k^�D����|+	��t�L��I`P%�.��:�3j�찱��-V�# h��^� |*���m��щ ����\f΁<�<Ć�o?�g@N�F&Ch?�\�s�Fa#���xs�;A�r(��"q���C�LuG�𲯻�\icz��_,~&Q�y�I����_^��Za�������V�8�p)D�!*����%��wRb�op�\�Rp�g�T8�y�1�*'ML�?0$�F$��o�(/Xp��E�E���E&3v�t�ǂ�AE��߄�b�B���/��4ݨ��<}m��ϊD�H�ϵ��ت[)���#P����ԛ�R�d?�������M)�jRٺ�����<���^o��N��=�v�δos]�'�7a�Z�0�^J+AVpy}H�������4�J�q��~�'��q��|#"�ߟ['�[ ]����A5N�p?Md�%�0I��҄T�N�ln����WA�
֑QP��M��q
j!�?8���7	�������ז:> �r������M�Ll͑3&�4ς&PHo��v%H=B�ZC1������c�¥�Oto��[�T���^��W�e�Q���E��b���Bxj�i]9)���=�����Ź-"��}v9����`��M��Ooi�`u����{�+�3g��A�`�qUBzǆ_�:�0Mv��%�M�V!��j���|�y&���J�%,U[�P�1�����/�K }�hB,��YJƋ�|Z�`���Jj���c���/N�	�>R<B�����ѡ���� &B|��9L9	�t�@�����v���j5,����W�aj�Tw�I��m�Ehfl,��u����gg�t[D�޶���ͽ�iMxeGQ��<|).�}u���:9�__���"��.�au��E���J�r�;U�ߥ�b�e�[�@��1���ɺ��x�{Ѱ��d�-&�AE�첉I��(����ņ�^n���9��(;i��l�En"�c��|�?=���Usjk��[=��|���e�_|�}'�*ڽ%;ڬe^�}_e��9+�ꤙ����`К@N�AW�Q��uh��ڑI���m��]�(�k��9�l	7D�fn�z�C��P􍝫��͗1�2�֡F4`b(}�u�.Jɗ͌�XIc+�<ֈ�4�!ߛ?�	��{�zJP�}�}U!�ᗚޑ�鍻G������&���l����h�k������zFlj�N�);�!~8�H'��%��a�H#-�)�)�Ƃ"X��D��/s�2vfq��Nq����x�y�%{(0�
 �jä���G"�'�����	�]D'9P6F؃�{���,h���)	��{]w�"��:L�K�
���;�#�T%e�J5�ZY۽����@15�</t��0� �w	�{B��K3r��a��`
�5`��\r<��$1�<!_�<�k�淼�u-�jT���&�ԛC��|�}r���J"W~=�T�c�$�e�W���F�j��:0a���WEř�ֶ�[���v)�|&'����R��);)x�&�C=�=^F�GQ���kȃ�yS��,��%�����i��r�\����]�>U���F��򦗎�I�h��`$�9�(��$)���]��/��h��$Y��v�@���t/3�!����?��~�P�F�J"?�bqx�O� (e�ʴ���v���!Y�U�	�����h����<��󽅭���zț:QJ���sF{���V���.���r��9kN����P��_b�?�˞�o�����V�R�'|H�_ᜥ�F�A�"�7B��b�$���FO�o�d��G�D��ﻍO��Gx<Vt|j���H^]�f�@΃T̴Z*Vq��ڊ��ɤ5��P�`c��?6ˮF�'��OU��sβcpM7��s3б�g0P�P�٨��w�fk4�-�l�	�������u@��!���oy-�W§V)�-�Q�䖚���%�� Ϟ=c�ݴ|Ϲ�����L��52�ƭpy͂[��G�b1W�E�O�ed�y�Ç;��ܮ�[=�6�=3��-����d�Z�5�EmT�x�UM���WV�e�=�e����j񾛹�aP�V�P�'^/N��ػ�܀��c�I M�H�{��U��4 w��������6v����h�ߠ`�i�u-Q�:CO�6�s�t}��M��cmU�� �2(|[���D�I�f�*e'm���,�d�L���0������H��V��u�`��8�T*;>�e��M���I��������)�����J<�
T��������0 �S �>Wɋ�z���[��H�g.���(��~n���������eJ�� �H����k�����q9��q�d�Y\3/��a$`�R��}�/X�hth#5=��Ӄc�C�0S��z���A�H�q����G���P���ӟ ����z�&�c�45����4�g�7obʩ��k���N1T�lx�i�}�����g��L.�ϝXK����˟�
o廊{�]2Pu���6�F==\�&
�$��1+�*��g���]^s�����"__�ΧU�pq�S�9�#��������r��x��(�ro^L���qړ�Yy���6�<����[��b�!����{{Q�n_�3���OeڽI���.^���rX���vn�F:���KxCJY�1/�M���}��0)j�Or���v�_+0	TCTa���{5?�\:GȀ0�ؚ��t�C󸱡��:��_(��ʽM�cUPZ����~��bŤvv
�`�D13� ��q���SȣD�6qW���.u��p>M)��C���o�>�����*]Ѭ�x>�1��>�b�4X��8�D�Y&!HqI��Pǎb�b���H��z@z���xe��f�Q��
���I��(�{��ihY�)�=�΄nT�5�j�!�j�d����F���E��^R���􁬿;q�H��pEOV��Ǘ�q���
������s�P��*�ƴ>��A0�"6�O��=y8fP����]~�$���h]T��6	�����C f���8ϧʴo	�����'KJ�7�����5��pe��Լl0����͟���x�V���֍��cر.�ἣ��c��A�(X:e��%��GD�J˧��둙P��,	���/�w�����~���4��	�bL��m�[�]��RTyIO����jW���t����wވ�`aX�7���B�}iԴ��a���������h�B2�JӁp���u��2dM��z%�)u��>Nq�]T��hyqN�����x���P{��,�=T#х�;�.m��1�� �8]��ي����6����g�ߣ��F���,GL���ͲR��1�	�2���<�.TB��9kW�pEW0	��{���a?D$�-�@F�BqD�$Y�u��������Ǝ��/+�p ��c�f셹�s�Y�O�����5D{�pT�{y�}�І����_oR��7��In� �^u�EA�f���KR9�s������.l�R����H?�4���/��![�IN�y5`��O5g6�kk�!F)8�����u�hSJ�P������F��b`<	v���c��n�p��5�Oh�+;�-�1�c�z��]X�
@��l� 3�:LR6fK_�ӽ��śϥ`�<���&�e�M67����
Æ�wA���/�م�Xj�[��1W{���}{�N����",�j��n�~~?�������<Y*��?�4C��kp�ML� 6�<���vK�5c̮u���g!����A;���h��8p6�f>��s�5ދ�y%�A��T�7�Hff���fG
)����Ц���nY�F�OO�F�x揤8>�??�I��6�s�M8�H3V�_�\�t��?yDo�����5P{�������0�]�2��0����qS:�)�#�_~��c����۞�#���Y��ç4	����X����r��$�X�-�%�����$AA�n_e��"��zⴔ�k��H���g�Gh�5m쁑őMj�	��D�Cݸ����*���ֽ��/��6ם�J������9i!^��+Z{Or�F�7�5��f���z'	�9�X�Rx�8�6w��5�F�f-��IEF�C��d�%6u~��Y��2'����9�(G��S~Y$2�q�t���.���fR������CE�q��ߧ,�8���2�'���00��0�qW�+�M�Tj5;�+�ڸ��|�ڲ�ڒ2h���Cx0Fk�~.dtY�m�kB�n�Lp�*�5\*8#W- ��'�E�=/K���Nx嗎J�*����P�]YN�KT�|-��i�T�rR���o�2�N-�l�P�K=��F�"�����&1�R-D>��a�P����:)�`Ȃ����͖C�!*��0�c�C���E��]=�쬬� cwyx���o+$I��C��֘1�U��E����,���q/�)����R�.a����?�}O����"ܝ�Z�8�aW����}Aal,�e0�rbIJ��FI4��_O���!��*��`A������(X:��
���ޑ%�Ξ���pdֵ���;kDh\�Ckj��vT�V�׀,����šs�^��W�g橵�T���Z��.c��.ЙH{[��:C�d��PmA�ت���ܢ�ę#.6��$��	��w�u�ji?&�VA��c>Ї��jL�ȥh��|�z��^dop�=yLE�!��|4�C�0���.���x��#/�l�h
�,ۆy:q��Qa��)/�1�|�>�볕SK�0P=Q���P4��;OQ�q+Q������I�&���y�n��zC�b>�!�@8U�p��@��צ���c��LM�D"34@]�Xh�-^t���P�������c��VU�H��ϴж�CK�1�m���U�ƍ��ǀ'��:�����r����Ԇz~�B��=ܺ��U	�v�K�H�\|�aIe��'�X}s�Z>�d���y^#",�A�X����o�{֭�l��s�]঱��F�ߖlZ��&�[u��I���':P�/��\���^�tea�k�<Qˆ�����e3� 8�J:�Mϯ6ӱ��-��1���8��2���C7�iz�d�N�3��	�39y��g=c��3)1-�/4ӏ�e����)���wM��{<m6��IlQN�������a9E÷K �FjE�e�k@�Y��t!��ٸ�4M_j�">���m�#;6q���"!�G�$�{���ǎ$��Z�����8CM��Hm�E"�HE��ȣ��H�`$Ҩ�4%|�ևd	�ۧ�D������'Z��8zC��@9	뢠T�@�������j>>�D��U������S����_�myh���'S��gp���
��I��c��,Ħ&�����Z7*rU��a�(�<�# �;rI�)���w]�r������"Z��6��Dj"f���Sq�x��*\�fh��لE0�A>X��g�@�×��Q��X�$�|��̜
&�v������Нk�g��հ@��r��d*���z��k_.wG��7���(#��lޖ�[o�^z���Rh��ϩ���<m�~���=��H��Vi���P��<A����J"
�|�Js���V<��LZ�bo�Y&J�~R*WX�QkhǱTa���<E��;���(�zJë��߳�P�S.��h̆75=&'��u1�U<���c"zDr0R������q/���bk�#'��O��\���w��D^l�*�&jЋ��	N
�	a�y���<�+�dSZF�4��i��h�ؔX��&\����p�y��c�#j��^YT��YY�ozb��2sZ�~y�Ϡs�����`�����u?��B�A*�SW�|�Q������gl,B�ivtE�A�������;.�i�In\��j�	5�9l�|�K�f~���=��qZY?�w�5e����Jil�Z����1a�)ﻀyR6j����FGA}Q{ �JA�U%]�Ȥ���Y�F2�蘒G�n�g�m�pm}��f5� D�������B�F��7�(��0�74a I��P�Aq� ��̜����&*dB3���;MD�g�;| ���(/�f��"�k�.?����Ih�!{��S�t���J��k�I9���¦�3
K�}p�5\2$��͸�R����u�3�V���߲1��� ���Wo0�7���:��f0� J�4B'lo:���~�49��"v�F��y��
�p�cO�_�ݸ/0D2۰ڔWm�b/pp.^QHŸ�(��\΁�-�k�lK����s�u��Z��t*BHT}��Q�ڃo�� ��-F�;����8�ldrD����ǒ�N�<zb���q���|u��/ �ẚ材F�|��TP(E�"�hE-xY�<�>Zn��K���}{�,O������v���piDf�M���,3
�����RZb��>Y ��=�̐�=
�O��M-8�b�o�F�	n;3�#n<��h`R"���5�x�}h:N�C� mIK�0��W���'P5����Bv��3�X�S���T�n�>r��qXD!����G�#�8��_;��=��"X]�DR��KUyW�����ETP�v����y0ӐbH�!�h�ؘ���0��C~�p
�M���ho�֎�s��r�羾�t^�@��<3�^�����׎���m��d_$�M�Ҫ�h��v�uԽ�萸?q|�>�룂�*�XK��d�ޮ��ʸj �h�$j��fE�n����e��R��;j_�)H������v��l�����@B�90I��+
�%U\��߶Zp��`n�>l݅)����
@)��f�֢��Hy�-�q�Cmh�1�?���O*��$��D_�	��߇�y�ph�?Q�4��QL���#;�i2Ԙ�Je��Q����'4��´4 �2l��B���ۻ�5rXǚ,�+!��T <\�h�ɍ��zɻ�B����&��q�
CDB�]����qn�G{�.��a���Y�K�i��Y�Wi9�h�3�Q����,7��~�|d0fE��+4s��\|tR��DI�0*�3�/y�L��2����>��a�ii��l�֗���*!0�M���1��^~��щ�]dz�M�
�y�c��xE��j��Ē7i`�puv(���n�eS��Hl6�RE*w8\��2�]�SǄ���S3�(K*v����N��'3%�&�\�4&�� �^�����z�WS6�K��L��Q8�N�;����U�.��7�AF��uܲ!���!�1��wS��>F��Q��X��-ĒU�ͪ���X�PT���=����[��]��?��`�2QYWՉK��*0�TM2��h~��%B�~�$�]��y�R3�ت�y�&�D��RB���B��n��a�S�!����|Ċ�H��v��KHkA噠���rWR*}�=QJ/4N��޵>^�^��w����J˗|M�?o�:Ug7%�����ms�g�^�`p*��P�4>�i�K�.��Yb�vf���L�����M��ׅ
�[n?��A�����gI���𭣩Ӽ�]&M�	��8�,$T�b]�!��	2w����]���!�4�)L��  !�A�����,���񩪣��kd�Lyɑ����YP�z6	�߫��Z\��m�njO�I��`T�P�le��I��F'k�X��V�-^��<<C�a�`���t��?T��m�\53��|%�X5A|!vM�����̆]�5���hx��y撍;g�|�>[d��-���R��1��/�ճ��=bvb/�Qt	՟y��Iҏ8͖ߚ�,n������Rv�n��(���{<$J��J0hj5�-�\"���
>�Y��$O����6JKdI��\�I�!�����rd.�z�)��S�7�c����b��;�Stχ��|�A�֭�����E[ť���0I���ZEh�]��E�U,�gq�9\�U�D�b�m*�6��x2��� p^N�}(�r�I)�H&Fu���{8����<n��c�9�A��{��,=`�S�É�܃�`8�ph�	��I��2l��?�3������f43� e���S��F�[��>ޝ{��ґ�*'�)�V6���"��q�o�}�ǵ��2�F�'(u,x�������4�\�o$6��w"�"����Q�G]��|!b�TU����x�!�X�p�ssW)m|���3�Y�Z�
tH�ӏ�B�`C��+5��؅,6�,��;r���I�(��uP�s� ��N�N�;w�Ū��O�l��}����Đ8���Oˣ��T9mAu�b�� l�;Z������$�i��$~�����em���}���,y������;�� 'n�� �����Uh��#��;���C��_��e��\+���W�5tEX��9*1���\TZ��P{�KըJ��l&���hB�S�{ibq��#�]�V M��/}� ������~���:Z�&����Va(-�ʅ�j�������|w�8#S��߳�z� �U���u�p:�{����B�N`o����FN\Q"�i�ltۧQc x\��f{����ﾸ�H�*O�Y5T�SH6�� ۰mx�R����}� T�5�NX>3�+�hd�oS�Ji D�6�vM�<�f�+	k
D�K�a��h��˗��*��GKJ�B�}�9���<�\�sR�Mf��j�g��Nq�����w:��H�{^5��s
`b�O}AJ�����������n�LBv�����xCrL�=/�o8#�W��.(�͆#l�lN%�7���@�}��~^���� ��q���N�3U�#���;Y�n��.���֞l��k����Wt��e�ܽ.�eXC��4��#ȳ�	m�e0,�J��C3��r��K��C��F�O`9_F�w~n{��/��f\0\D�������p%�:���to����w��O�}f��v�|�s3�O9��ոx=I���+���-ho
�a'��3��7�~�uN��ē�W��6�z]�ZĢ�Ř��������E�o(|�n�]T7�c|, �H�	���R��$V?a�j^{�����ۖQ�AO!�k�߆&������3Y /�TzG�X�OJ�^Gb�Byc�'VcU�V�>+�Qt��J��~��'�c�;�h����*T)I$�j
v],tK4=PCz+Ǭ����#�J��-J�v;s� �P�ۮ�=��e��5�A�=K>��sP)���Y�e���4x���:���:D�9����-�M�)5x���@dF�)Мl6�S'�� "��ˍe��4N���^�W!��9�B)��������G�72`Tx�MdfD�I"`uW�`�h��"z�_M�H�;��%^������0�w����m9D�ӊ��J�6b[|B���'��"����S	��q�f���!2��,�oT���uo~_{�9i���h�i��옣��Js����s_<�B$#tu�K�3%��}ٳNXB�+�t/�l�r�ſ�p7!��lǞ�p����3f�[P�%�>D%dXI)ޣ4M)C��ߛ+� ���ij�	�^�Y���e�����n�)��	�ȵ����Tz�-��g�h&C�p���KSc��F�sQVЬ��S6~���k�n�B1i�Y���'G�8-U�Tk��_џ���B(䌴�^SK�m������]�b�WmmT�n�W�N:�bV-ů��A֯�}Ѥ�>]׻;tz�g���3�j$(�l�+M�%ޒ��"���C��/E0{ïI9nh�z'�kN��[�6�pr�K(rOo���C�Z䞱�}Up�"� s�c��1C�j�%������ID���ѡ7�h@�!�뢽�0b��hE��nO/F���YD~1i�=�\$�������Vq�\�����m��j9-�-�f�<7�u._@t�"�CB��e�O��'�Ч#���n�$ާ /�B�|D۾����	m痾�캁�[�Ӫ�\b�_,�0���f_{��0���&)&�U6Fis=1$�� ���K�\�����U�]��\H�F��a�
z����]^�L&i_�����*T�$� ��Rq��}����7�U�H,N�T
��u��CKݤ�.j�$�եc��Wg���c����������1��n��;�e�_C�㉓�q1Li��7>Զ�)��Eގ�ž�yな�����^�]9_��e��4��>y�o��1��18uCjL�Rv�LT�+JZ��V�CMR���q0Ъ��<��A�5�dU�p��ң���>�FK����\��7�KQ!�a���K� �(h�-7\F�#����wh�=⏠���T疁�~b�m�w����x�up��ӛu�4yY�l&Jq��=��-�@�յ�G�v���G}PC=�E��`>r�+WMͭ�bWd�B�$��f��*�����Ӗ͢LBs��ƌ -���XF5L�[�_bu�B�	��?��ӽ��]��7�<���z��I�y�����@'N��9g
�o��7����Ow<������{��KP7�Z�D$M�A���}�A����������Fڶ(m�:;b��kڪQ5@�^�V�i�YyN�Ks9��.��V�@���X�^�{!e���
}iF��1�1����_��� �&��o��	�H��C�A���;?!l>�)��C����K	���y��#����)O�Qv����(�/�RS�Kv8}�6�@�Ť���R�,����S*�6j�:��DVf��a�h� ߭X���SCH��m�<"��F�̤�,E�<`����Ć����{dXUJ�ox=��q�<B�lŬ�����L��
T<���R��Fa�?ZA�Mu����b��M��3؍I���k�\��l#��*U�s+O��}x��:+b���c%�z �I�&�C�`�E��a=0��XBg��l�G�T�<oֶ��r�ZDTK���X�)�XC4v���G^����I
��eh�;�+%��A Z�R�\BK1���O_Hؙ���1wX�[�T:2�2�ٔR�4��1�����7n]�h�FV���- N���	Y�e��̑Mx�݆$��-�$_̠A���3dȯ�vh|��9P6�y�\B�J��W��9J����T��v|��u�{�4� _����Kɠ�URk7�*7+�$����?��8�z��6c����\l�hwbnb��CS`�v�����3J#A_�����oӢz��3�E�����ɶ3\_�QD�8L�&�0���ף�=
�s`�3��Grʈ"��S%��|^��W���L�6D8ފ?=H��lB�q��V������[,��P����!�� �K�o��{����;�ގ���|YŇAg)�5 ��`y�d������D��'�F/�X���$�{NC�Fo�y�[_Y�Hf�A���Z��3���Y�XCg�Ǟ��
�^�[<�Ψ�G�Z����ȸ���1�k��Ql�ATt��jc��o��un���F�5�g�ʾ��Xb��#����k1ak�C�}{�~�%��Bz��Nn�*r$��H��$GBTDM;)�3J-<�	��DLͫ��� ��7jx�-n�o.��nDf:+Xz�K�5�9�Y<���w�G�@oa��.&��OS��
�"�K��|9�����%�&�"�0�x�i���ټ,����I��Z���Δ�`B���lj���!"4�Y��'z|*�K�a��>��S�<�r��%�F{T,xdFJpu>0O�|��:'Vߓ�=�*g�W�����ݦ&��.�l;�Ƅ(c�;�D9�Ҫ���!�K|�]��n�bp���SB?��}7n��=�OR	���@I��_(�i��j�AM������y�+��=�j��gxm���	������u�әB����� �P���-���=21�8�r��}׏��X;<�p*��H�U��Y��ĮcP� 5m�#$,I�hq��8V �Bbr��Do��ge��~m��o���&xK/Q��a��>	�=���Cb�ɻ�2M�w���Z��Q������ލ�^�&��l�o��;TTO\��v��|�[�J	��̖N%L����v:%4������1ڃ�M��P�Qu�%�� ����T4zz_i(�o�[]h3.�a{h;�R�0�y"ݶ#/x���!��e-�{�$���mV�H���K��c#��H�p�z�RG��q�&�`��Ȇ��4L?a��H(��K����2��k��
Ie���f�k_[����]y#�nAzh�����.��C�Nt�t~S��!��0nX�������,�碒�����#:	�/�'Ȝ�m����b	eΓ
�2�O�),#5:v�8�b��l�Ү�X�r��O��'�?���� &�Mn���//
���.YFKTu�.�7��e�D�t,I'�����:�|�T�Ѡ�\�th�Iߦ�J,^o�941��_��8�I��n%=�c�PG<:6�!:�6��;�'?�@�kG��RS��/E�(�
#����|,�e��Ŀ�\{W''�*���`���}�~��N:�pcO5��TUOj����\1b�d9$������m4��� �*���JR��w�l�F�����뿷�=[�e��rd(��O.)K:kP���Ɋ��/�x����l�����Yr���PYyƶ��G��ӒƉm��4@�W�3�u�V�B@dr�RU�b��t`�5�,{��$�z�f�k&�`�����:��0[��Î���[��c�	j��u(��N���_rm�t�,���/����{�P���������,�����[:\�[g�6�|x'����w��7ǀ�2��+�1��DL^��h�t��TE_�ˢ�Uw��h>��!�7�xs��<��m����P��ot�-B���,V�l@ߟi˫b���o��e%@>\�I�h(W���4�v�v�wu���Z�ܰյudO[�H��t�5�G\H0��#\�&�r��� �-	��#]�KLy+r�^� ��~���bR㨆F;]@���S��I����M�I�3i�IzD�A��� /r��NדP��۲ժ��
�k�ex�b�K�J�;C�^��UZ|�ip����E�Xj�o�F��o:rQ�"�=��sb|�0������|7�r��8q�ю��X��<��%�j�T�t��R��߽o�����:X>:�J|��<�g����8w� NU�@.�p�2�����=����/�	�Fh~�� �E�U� Z��t�{Y���ӊ.ק1�#O���$	rs��%��o/I��]��.[�=�4�^�W�����k�|��8�D��*ā,=S�i6}p)L?��H��!s����ȓ��O����K\�{�`��5,z{������{lI<Ҍ��z}KȆ"�_��4JI�g$>*߂���1����"/A�_�D\�qe%6�(q٧�lf�8�V���$�P@�P�w�,�p��%�eQ�����m�ʐ���i(Ac1lX�x&*r�]�n|N�gǍ�0��w�Y���oQ��p�a,��t�����%�؄����ˤE2a�l�-���(��|���n���Ϟv��#��p�F�m�e��*^�sv�\b5ġS����u�|�vrS�hm�
��!ܙ��*C�h~��L��2�����}�ty��ۜT*9��R�'���8�im�[n9��H>W'6�0�h^�>���W��>�I����Y�&���>j[i�a��3A�b�Qj{X�ۥw8Ü?d�a����B�ª�i�a�`���pZ������喙b��t�6��@������)Q��@��mP=%�������U1i�T��X=�,h���_�*���.H�^j���j�a��yPR�D��f���S��p�D]�+���bX�0R!�I-D5�����0ɍ�۲&r#Z���J�u�i�h�����[N|LF�����rs޳[D��T��m�8��&��z�̜�a��#>t��}^�TQ	��pGz���v���v��-��ʗ���	%�,P�L4r��.�H\�ˈ7�ބzW�!1C��@y�Ln�!��>)[�	|R�HdJw��B�OȺ�ނ��(�� �M����2�]CE���QX��8/>5�1����*� wش�����c�ar-��k���v.)�NA(�I��B��Γ'�{jɸk���>�Bk��Z��q>u��-ts������GU����ݍ,�@Gm�$r���C�Gq��`a���d�+NcFO:��_��K���9��\�s���14\�OF�M��Rb-���-��4U�ݙ ��3�Q4�s��E�&A��)���	��L�	����H{L��R��e�L���ZԄ&�ǆ��mP��%M2��/��W��C�u>��m8	@���;"�@��E)�nU;��P��/�̸�W������͓cG��Lqk�� ��L�XjĶn���f39��_�6څ[�w
��);����ˌ�!�}^r�oV`��ض}3�^E���ysb@�{MTn�G#B�Żt�r�,%�4�K��˹��6u%�6]|�c�^<���������ⴂ|a���D�	f�1�ۗ�v1���"�zI�lZ��'�ycBm-�^|��/:a���+�|�k���Ŧ�{��B�l��S��������g�\�c�s�a��K�P-��:g� κ�ֳ�S��I$�bb�[��3���ٟ���;M���s�I��2Q�f6YkMn	8��*����uk�l��x���ˮ�-2��{�RSos�ٵh{g|��<�f���q��x_�zb��_Iii��/�YkJ�_x$�����Kj�P#V�����ˉst㊢�U<<�(��p[�����(W6v�BYP���+�U�y�qT0�?��x7|�� C�M!��ϏX��m{!H��#��YlI����[��x=�y��#'�w�ꛭ�H�����\�;�/� ���J�e�~��ud�}�_0j�p6�����Ɣ{jq ��;����oJ�����<����eK��@��9�*+ �-�W�x�g��� ��6�M]��"���� DB0�|M����f�sv�A��x�����.� �u�������m�xr�`(Sj��j�t���GК��(��]�hjg���+��0�5m��A�s<�V��^���?rj�e$��'���G�Y�=�i��B�k�lv�!�K�;�}�l���ä�/�c[ ��Xr�b� CE�U;��
y�	՘���<?L��[��3�{w����zw��֝�6���C� ��%ь�6��t�y]��k��YS	�.D�`���2�Y�����{y�Pd�[3�T��!�W}E�h�ܞe�*ۤ<.�I�C�crqs�5���<���m�Sׅ�b��G!zW��V\�i���,���qg~�����:��[�ѳ)4)�݆;�a9����6�/��
3�+=�}Q��9���>ǌ���kAr��*8n_���k�q��X��VGF1V�F�EƋP&��e�I ��� �Z~��E�UT�lh�)�q����{&E���Øn�����ѡW�E�ڸ긨��!R�}���b�����f��������B�����~Us�{��D��+ǟ)L���o��������g>��� ɰ>E�,gJ�զC �����K����T����1��β���̝��u�����\w��@��D^"��I��@�H%�7��������w �����m�#�+���c�fy�������q���,x);}��*f�3�c�pli(���egc�P�����5� ��v�	k�v�=�Y�T��r��0�A�E�1�~�e���R��'�".,�0�	�~s@h�������`~�����x��4����t�"���a�����\Mw�������Q���O���Qr���p[��"5����u�+y�)-C��74r��<��M���� ��֜?C�l;�c!��� b{�QC��d�	0�G��ƣ`�U�=l�|>O�j{z�挌l܁l��:�m����=�u�K�6h򤗍���(v�f��.����ǈ�j>�4Uޑ�N��Rp�O)K�rD�b��ٍ�)��uˋ9(]2�:�f@�<kE���^��	��+ଓ-��d�YQ���R���T̈(�����s�T\*�ܻ�@�t�Y�}b�P>��f���`xMK��=˾XN�[�o-�h�n�@�ԒQy���A�o�=�{͑�6	��R��v����܊�Y��^ |���51�S!��܉%XJ���k�@-���͓���5�j��P"o��.�sr�������	~���h����d�ez�
�iDWu׍�h�b��҂���^7bH�7'�Gy�o�j�ko6�C^粐�e=���ɜ�fԗEgT�t��߬蔊����D?/���ȧ^�%p�����B�%g<q�[���;ں�Ӆ���趵#��W�'�����)h��6�[��n�{�HE�gE?�8�I�1�'g3�qI@��G~��D֯;N�C���ē��85r}��g�AH����K\�`��{��F��È�Į�����Wp⽴kQf�B)�����!�Y~� /b���`����e�JW��X�"���OWQ�o�'i�

�P>^b�"@�dp�SK!�=�������q��|�w����}��u%'`�:�P7`[�����'�W2D�;�����v#�٧h�&o��#;���
x��P�S1fZ��& �ܵ�]��%ø`�$�N��[�)Ex8���ah��㲉U����\�E��T��5,����@働�����T�"��7�|�,�.����o�����x�Pty���åj�\���3)a�G�����~��$�:�q��G# ��K岕+<wY�pk#� �Q���.b�+��~�amI*8�D"��Cx2�����ߑ���[u}{�#4����O�br~Ls�$�4����JuD���6H�9ObM_[�'6��������'[��T6��^<���7	�
�9i߾� ���>�d|�T~�W�ٲ��-�k�R�4�Q����,h�f⑁�-���p��	'��,�7�P$����bY�"�ĭ��`�����QP�PY�ތ��A|n�����S�6�
��֬�)�8̢%������w�zgPi�[x�'�k�#E��gz�m ���`HG}��i��z�x���}�$uτ���XmRx�n�AϤf�M��AB� �>?� Q�`��Zbq3v����
sb��|��s�B"0rdu����S��ƥ$��''3>:!3���w��P�m�u���uBݡX��YAr"InFz�Tteq5}t��۰���݌�NZ�O����[��U�:�UZ;:@H�C�Ҋ���@���<k���h28�$�|�����HCM��`�C�D��d�m�B�A���f��Ff7�QR�a+��^V�Y���ԹI����������&�������	����B���GT���;8f2��5�E�[}�X4aw!I�7W��Xܽa?rI;�����Z�l�I��\a�R��+^&oF�	:��.�r��螣|��A˘}=b؍��4�G,o�U-�P��uwo�x�S?@Q"Bcn&
	�C�6�#�Ո;��8�'���@���P�����Y����Ǆ9 ��>�Xd�
�1�f����vߪ��`=��u$��:C���"ׇ��O^��������W��#L�:���W_8�?+{��T�_=����6�A�c/-�2jNR��EXnG3���wJ���.�p�N?Ń���q8X�����ۭ�)k
��&�l^%o�Bb����$.����"�)q�)�&LL�.A4��:�Lt�z\��®���tփeq�&1��*�B�����t���u�mH�/N'�p�U�@��1h�!QZ'��ґ}��*�R��؞:~3�R�}����W)���q17L�sPƦ 9MǮf��L��{�y�~ai�%�~1k�\����'c����z��E�cJ��ň�q�me��
���l�D� �>��i�*_�-�$&^�pA�1"�����\��SmK=}}���ݵk׼u܏��DH�?��Lk��_�
�Ʊ��(2	�c����ÿU_���d3�n���ԡQ��b�a�^��k�kUI*��!�-�:��������ޫU�/ֳd��pXt݀�ՉyeFף}M�߲�k����׎*����g�.A�Y&�Yă�z��6���X��	�9D�"�t�7+�z�v��p���0�)i����i�GF�����^P��e51�=f[��|�XC6t�a�ܠ������X���0���6~�pTN����ޚKz.K��㕭�:�r)9Ӻ��rJ(��]:����E�Q9͇�;% 4L`����ļ�Ђ�"�$���ML��"bAc}�]s�M�TxC
���F���e�Ǐ�����9-[^�~hG�����r1���N���N�1��UԿ2��r\��g�έ�5����e�=8���]�]����c���)��t��WT��K|�E�Ya|3I"{����"�T��3r
��ȶspz%����8Љ�msVt�W��S��9
f�6F�ɊDK*I k/]�A�4�3%�M$��A�E��X�Θ�mL:	�]��2� �Q�y��䂶tq��l��sf��F�e�%>��^�×���V��ͧ���?���Y=>��{Ɩ�}u*���Ri\��W�NX������$#r9�+�t�#�����f�o؜D6��Xn���z:���&R��hBI���/˃��c�"��o�t~�5|[kh��b;�8�!���+�-�I������)�u9�s�P��n�22_@C�����+h�C�NV)�f|�F�"������
Z�M͵��U�B�1�ԡT�Lx���scx#��K1�t���~UJu�����G�d'�V�=M�r��vO���n�����9�&ζmNSh�< �ba�H[���cƐz��n��]���?	�� H�-2>��;�)�y(��4 �)/��
�y�TS��m��}�)�30�`)��d'm\X��;*��rz<�P�XC���g�5�a�!�&d�N��_8�H�V6G� ��9T>!�9��P�[��t!����,�"����3︹�<rc�eX�Tԧ�m��������H(���e��]P���}85ƮƁTB�P��T�����x�J�����cĔ6�Dl>��E]�:�A�pU�S�^f�oH�u�z��V}6�%r&�<�vͳ�/;~� K�6�"���t��z@jf��"���;��[��b����n#�ʅ�mB���W���`Io�s�(r33Q�UB������c�|a
7)D�tS���̉:�@]POF|�x+�T�j*�����9�s9�H��'6������Y������;�<JXZ���>}7M/�Tz=u�,�f�er;˼ߕ74���V=��gT�Ɩ(���`�߅�]�E����V�;q����Gx��_9Kk���3�3�4 uh{u&<J%�lv�s��x�|k�-w� �������*+��[9��Y�0�I��p����G�l%�_Lr~�܆�Wjj�G�#��Z�	��vr"�鎓 ��û�Y��?,���`��R�~�s����ReӵX��k�������:��?��%�����Q��'�u[��$(�Ϣ�]���Rģy�j�U~=(��A��P ?�o�� ��C���n$ï|�?Y��X.e�Z���OH�� w��I"�>K�K`v��ż �ԸШ;�V�$h]�1�!aN'���Av��Ч�A���H{�=#P\���3I��8.Ig�H璟y+S_M�1p���dtq"�؇ �C�$a1�e��:��F!2�xE��kxF^��
��/8k��~r;Ʌ�Y��i)�4��~���͏Iџ9�"mQ%V3�쉖�W0jO����ᄂ2.�@�Rw��a��������~��)7$ZX ��<������B�j����X�1��=Ӯy����8����N�M�iE�� Ƅ�b�Ƣ���o"8�
�Vk���APC� �� �,\0b�l�&<b]�Ļ�/��*b��:aFk� Y�IFԖ�~uV�3q�z�9���W17�a��{eV��=�CM�_ʡ��oPo�!��a'�����I���RO�щ����Q/��?@)�zb�T��-��q-�g69��Y?�{t�aF���� v�V�+��D؝-M��(��q�@�&OCQV�H;y��d�K3�a�t���z��̙Rs���M���D�b�"*hLCfH�W�q����h���<�_`H��[r�n�]���L���A���o�5u&�=k��fYB@��q��g�3�X���+C41�r�ٳ�gkەR�Ǩ��cqT�&��B&�����^����9�Z������7Y@Jt�kJ����cѯ�dWj5?�'v^\#�uIs[�o��Ԇ�P�$	O���V�	L?����,O.������a{�k�EgC����XV-.��HC"������q	�=_�(|�>������XK�1�۠]%��-V�]E�����}fhȡ���n=J\¥v�&m[�����[��+Π��5G��N��mMS
�Ho���KI��,7̦î]	�-+O��&����v�*���㛩��1��=zC�x��Ht'>�'[��9�o��z�����ʪ@��y"2�w���O��w�Pf�ВO7%��k���V�0������)1���,"��a��	HD������+�� �2*�'��v-C�׋Ə-9�f��Lyo�i�,�+B��<�)U? 0E~��s~�Z�"j��R!����]u��zjA}��_�ڠL��u�-�|�A�q�v�yFd�����ζ��Y��� `/�E,�%��Jh�K!Hdq-x��L�لEY,��Ys��>�=e��ޣ��m�S.�1Q�!?�0�=�&	�'��:0.j� <ŏ[�X�o�J�Q1��oQʍ{"pGpg(=��	�g�5�Pi��l0�����{��^Ȓ��&���%겍p������*T!�D?R�s,��4�h�V9�[�CgdS��>k�Sl��Z��;�1^�Ķ�Zv�2��F�Lz�g��<�e]���;6~\���+ �"��e~����BOh@��|[l�!�48$";,��׳��׫N�^!\XM�M+��Ȋ�Y���FM�9g�E'u���Q�%�י�3ݩ�!�b��Q����v��\*��-�\;�{�����H�R鲄�-T),�Ow�Bf���D�b�j�gYN{o�`�e���Ͼ�J���^�sU�kۘw�v�)9�u8��P�����P��_[;d%�\%���Ѷ�3��#�4�j��ʀE}2e_A['��o ϡ��>$ з� ��o�4a���Nǟw���w)=�<�b�j�b}CD�*�TJNoD�������,�ĭ��"�>K�!���	k�7��^�๸j���z�u\��_�S�w�L(0脭u�����2K�c��䱂"�O&�W�k�u{SXy��[܋ R��+�/�ASF�B�,�z�4pQj3��$O��F%�tYfZA�E��2����ߣ?�B������)�dOI&�?�R�}�Ϊ냷�ޙ zg�4ܖu�]T�@��8�+-�4��d��M1����}Ȍ��kJ0�տ�	��V���3�Ln��IK�y)�o?�\ ��*U[|�Kw���i����8��̳�����XR��]�������\����y��/� ����lh��#���|�ɑ�3�K��sΞj�c��@����ui�HAl�C
y���qz�g',I�<P,U�?l���)�f��C,i5_��G�rT�6�Ѥ�MUH�Ӛ��ɉ}:�ݙ���@���ӝ�F*(ԃ��q{³�D�!�%�V�Eɥt}`]�m��C��8��v��ݱ�ꍘ��-�Ԓ�f���[YI�تlF��x������5=��%��� �i�F ��v"��hO (���߽H�{��>fm��qT:f�}�p@��6���e}N#���Z����f!��o.A�z�w=�!Ε(ps�V�����#��T����6��47J�2⶛�������*��ݺh~e�2�&`�_P�$r��!E�C7��W�9�\�3-6*-�����\�"�{d�
?a�]ArDh4^����A�eK�i~�O�N>2N�@����~l����ǵ��p��OH�9IP5o5�p��@��-��q9n�K�U<�����%}R��<��?�[�! n#_�F����;vu1���_�k��4r.�㒤����Qש��9*�f������ DT��á����R#��t�
 �l��F��|��%���T:T�-r.��[�Zz ���j��+�R�\3q�8�0�T�p挥>K�b	J�'�2���Ɉ(Tg�'�д����j��/׾$F�`4#����c�g_��,?^"�9Ͷ�_��<��n��y&I{����-mb��lֱ�VQj��P���@ݎ�E	�@���q�.x��7��EUȝc�h}[��T	r���z�6��R�4H��#b��K��0�6��ʜ�o�$�v��7>��Nv����Fd��v��p>��	
�3���f���q�Z��C�q���r��l�x��U���z����H&K����h��@_�"X� �A�)���>)�v�:�ٿyWy�>���ᾟ��;�yC�B({�@��*Ny0��[ƒ���(��V��I�7 G�0P�^Ȑ����lne��Њ�>E�h#�+�����إ�ņ?�9���:������*��yם0B��-�H�5a�b�M0Ҧ��|�m���
�ۍ�3,�����q�"/�	�@[��ʵ;�c�G]<�u�͢�u�]���#e��El�n�dO�u�����@
vh��m0�:���6U�i7؇Ns�)J���PR@,3k�H	@�0����o�K,e��,K��� ���;��՚v{������@JOdű���An�K���7D�s����"���!V_�5��ݤ��)l�;���஥�1ʈ�+��|��|d)V�r� j9L�:��/+��� �$���2���y\"�-N�~A��Y�Բ|��Ψ;L���l��x�̴̼;�����8|��}6nFݥ�D8AL����mG�h�����#���Z������pm��;V�}�O�#�:�x>i�e�Z�h���p�%� hһKG��v�Yg�}�N�RrW]�:s����5�NEtL^��Ԃ@�H>re������#��bej5/�y��(�y���Щ�/�! _@`�$�4�7{=��$�����0N��
8�,�Td�)"R�bq�ե��S�;rsD�?��di���=0u날�&��=a�B��U�5M���	�����F�UT�=�+b�`و�M\��Qf$ L1�it LD,q�88н
j���
Ǐ^Gun@@�f0/M���AG�R%�����A�T���m���J��t���.C(���gfp:{$L��K�ɶ��CH���e�>�hq]=�Ў�`�7�X m��&Y���npaʄ��a��1����^��:�-ti�8�|+���gp	�T9~�o��W~9}���&�� [\�d-~����)W|�܈܈ZotR��m��B��~��ᮡj2�b?x��#�ϗ���U��ۻ�V���<�����_Eze��35r�Y�{`S��e�Uf���Ě��np�&���L�C���X}��_��̜�H;'0�FH6�Q��J�"�y���.�P���h~D֜���;rS"���I*��R��39y�}�zM�f�3�.������j�u����Y罩H����.�#�
PJ�5Қ<��,:�ʂɪ|��k�C���%�����gM�%sMx���l#�[?�HP�#H�N�"��h\�&=h�����/7�V�	�Kv��i���h��vҌ�N��خ�Ŋ���0�E2�i��of~�an!��>�Hْ\��pd��J.y_H�"���Q��O���s�%����V��&]�M���IWv=r�Bs��Q��O�����#�	�v����ń�i O�~�ɽ�C.�.22
� �-G��3���������g'��Ml3f�>��K;�K>��>1�V#"���ݼ?Ky+�4��w���b�>��n���~Ǐ��|s;c�\�v�r.`
�p�~��S�An���[VA[�%�V�P2N��̛�p�Us��9�h/��~Gg"���:��07x'�����B>6_ 3���ґ�x�v�6��MD�30���j��r=�+��b����7�ϼ�����iPI�"��V�=
�g�?����h�L�0���%T-�Xn��!E�a�w�zAOA�?���6ȫ�~4����&6�ܬ���X�y�\�A�L���6�"l��\�)����t(uą�bUs�;R�w���&	��nh`�e�zKV����-��X�nu����9�Ճ�KhS3+=O�E�8����^j����f�bN�d�f� �Z%m�����m)��(����Y���4��78@�W��"�H�f�_�Eⲅ����2�ykP PH���gr�0,��VA2A壧%0E���ڨ7�]֤����H��ݙv�@qǮ��{`����D�[�t�u}�=b�����r��E[�n�=��Z��,��9>��8h
�I'���(}����ͼ8lc+z
;؟L{݈P���L����Կڵߒ���,�Xcy߻Y<·TFYs�ruhreQrO�e�4�ܕ�h����&`x�}P��k9���0�t>�0]�l��`_ߘ�zހ3�A�j���T0�OQ[��~��2��	���+״�G�9a?RB_A�US�Z����Q��`U�SK���`����hs�_z�IV�y�LMe���E|7��ѵ3�Q��'���V�M۰�y��$���\z��$Ӕ�"�ggϩ���t��n��'gC��y��`��{���eETp�v�7�Z7�1~T)0B�sO[a��9�X�+���H@c�a�sX�lV8�xf�J��VX��9�wl�&�a�@�Q�\s_w�p	)yX���T�D�r���ߵ�أ����ć)�q��P,�u~�Fj��ueĸ����t��kaXR������'�P�X��S�	zL����K�a�;����Kśpn�BDeU�We~�Ǿ/�ßs��8ժ�7lQ���e��D�u$�[(��fv�.����,�:&Ă�{�J�W�~	KA���ŁG\��%����:*�^~�=;>�����f�̻�;b!_�).��01�I��Z�� ���R��2�M��O�QG�Ne���E+��.起�n�
�:��9cY\�څ�)f��ɤE�V���J	���;����c+Zkڤ+	���Yⲏ>����h�ˠ։H�P��F�Z�{ܐ*����񟇝]#�G�ᇌ�c�?�%T��Ts�D�8�2�[cͼ,H}�m�/��\�wHk`�Iԗ��K˥��A�l����SI��3���6���	�k����R�7K��F6��� N/R٥�r�=կ�1(+]�jڔK�gpACw�0�L��"��o[!�)���䞟����.�*�)�6L�`�g���W����~��D��b���ܯ��{�Rg��7�S�R;��l���(����dt���g�*��+yf-/�|�
��@�2!�Ӓ�� ����w���Ud��iS��򊰼���k� z��x�lF����bܖ���ᩄ��59� ٥�()�b�&�/�!O��*_�+(<._㣝頌��Km�w�wI�7�����z1�I�����؏����h��%`NFgs��+����EjA�����$X��+���B���Ʀ�ԜSJx5�޺��&d�̚_	��rwt��i���m��JӲ�����-r�Ar6�=L2���mDT/�d�\��b�z���_�� Py�X���Rm	�t�2bm �R$չ0���!��lc#D�$N���Ѯ�� ��Yh�᩺�K����_R	���c�p�I���L5�&^:J� ��X��_L�~�&�O�HB��T��Ȋ{Wz3n�\�z@��U�M��I�m�w�2�V_C�bb|��|�؏��C�8�5��`�mI3G�	��Lj�����Yq9�\�[�����_k�{��S���)�ȭr�|&Cy����yG����+�y���qWxq2*g����Lt��2җzf���I��9��ru}`B^��z`��W(��������h�t0I�!����FV�;V���0͍)�$A��D�s�@�i������a�@@`\�ؚ��V�MҿOP>���|?��E�k��qgi�Z$�d �#��.}U�(��;
�O��+;?���e��g՘O����M��R��#g*�ttX�� ��"�8��M%�C;��jr��G�dw��CˊPI�1Bә�r;�����Y`��!t8�T�{2v�	D������5�][�Iv�#�S��3t��0!�9>B�[ϧ���;�xn>���P�0�8d���/=�07�	���>��*]�:#��ƣ� �b{DBؼ�p�a.��X�dW (/�ML\���㋼C3�"DM17[��Y��X|N)�b���ض䭂
�!�;����e4�UW��@7=Om�=��
MSy���౜����L�?e^�K��	�O��ǣ*��g�q��n#]}������G�6���A�B����|�����@����,���EàYZ?`i*+����2��^+�-cE�g{��/�E�?��!�Pc���Йn�V��qW�)8G�yv���٘��Õ���qϗ|�B�,�U&�I����D0�������B0���*�m9���C�T�,�a�a���C�:~4|�-x�)��Mw0uJ)�7g�r-5�~�N�6�}���U79䯪e�n��zɀ*�b�?U:�'E-/�wF�ȋ1����U�ek�1����%6U�سTcq�~���f��sQgAЬ�g��ò�जrAQo�M���=��7�w����I<@�@\�?�x��P���͘�L1��ӷ"Ӗ��12�Tʱݟ�,\8�8V�լ#Da2܌�N��Rp�+�L�^т�<<���R�,�s���	��k.���\��8�V�q��/�D�3�qH�3�����, �ю��bfnK_�����ߝ�(�oz\�Ҡ�!4��4C�p��m�͹N!�Ug��j6�6)��,s=¶�/�_w�\��X?�������Vإ=f�ob��;x=���"K����
	�ώoH��sY��,*}J�vl{Yي��|Wg��!�w����
'YUoTr����n��]��6�sd�`�wP�2��-݄s���@�\��� �z�t�����G�2�GC�v� yL<�Ch<؆���xi�X$MȠ�-�QM�_F��$��'b �yh���]��|J+ˈ{��U�N�8fѡL��4�"-,�5<E��[tԍ��ښ�P����o�W��(���\7�Z����K/}hW�'h��k�˨�7\�).:�)�-��.Q��e�6�Y�X`|��}U���$��ok\�����-���P]���ʽYo���8�C�9��ʿx���J�̊�\L�U��ɺ��7���4��˽�ҝ]ۤ�B���	���g,��ll8���rK�q�z�9H~��@4h?��D�P�T�5I'�D��/a�i9#͑�?e�<Ē�&�4��e���SD�q嘵�/��ߝ+_V=��3n.�j����ʑ��:�������wA5R�ĺ[�9CN^�b�:"�q���<9�Nx�n�l �B�����[*���}9~	Mo��T��0_��a�'D������93��% ���1��Z��AQ��٢�~�eKp����j�xJc��-�E�i��N�ςnz� {S� ��WR��s��Uy"1�S1���e�i*Tv�y���n_�&��+��ws%����y�P~�2>o��y�ZF��=��(��u��tP�#��d�a��ܤN���C5�B�o=��Sͺ�C!e��޼�{��聋@&��b��9x >���¤��"/<� �N�L��<j͈�O"w��L�#��%��I��R<�c�MS��R �8�F�+,oώ��=���H�n���>��J��h�lY�͈N�����@�w�zj��Ţ.Z{����t)Z����}��݁���xiz���K���q��}�Y�3D۩�1 1b���8����.p��X��P���`�����V@��4��w���?��(Q��H��gO�����x<U��j�b��O����\	LEC^��"��5ģ.������g��(]�ee�9�ȑ�L>k��03gy7`�0�Yom�k*y@3C��3;q��~5kC@#̜E���̈�:�s*�se�i.E�S�~�n�l�+���N�PW� b;sNS����-�gW܋���?�A�h�P�.-�i)����ҪW��fvb��x��7��/8`����d�6�Q�dc�x��;s�p��ۍD�!�u'`O,�/ ��׺*f��W}jOׁf?�9��FQu�?�+�����Rue�g�,�O]Q���"3�,d�K8д5��#70O�	�۴GW_��e7��2s}4�y�곯��/�C�h�vtw����z����S��HI��i�	�(�_�S`�:b���H@�䋯�y�����}`����V���72�>:�ᘸ_�4�ѹ�0Ô�-�Ĕs- M&I�7n"@����տ�I��S�4)��v�A�^/tj�qRT�Q�<o7�)��ol�cw�6뾊A�
�?�b�K����CK�T�@�~w�i��s�<��0�3��y&^�I.
GA�����u��(��Uׅ�"�BH� _��'�W�]�ʔ�o}��ǿ�2��HNVԋ����ma�R��T���O6�.)�{خ?���#��+.|�A)������}���r?��wF%,��ca#��
;�ZU?V2@�-�)z��F�\PЗ� ��!rb�HK�\��:@�a�g�9��� 1C".-��>e93���n0}��c��mi�'��,�;��}�U�H^���f��zV�Sd��or<�-�xŹ�};(�7zL�X��j��Ѷ��� �S���!�Y�6;��ĵ�j��+�XM��鼽��,��LyXn�%�僎��k0�U:Lg�bw�>�8V-?���oC�J�r��?�k�N�v9�k���߭ �H�k�1�}�$e�x#���k�T���7��X��\?Չ-�9Q�ٍ۷>�U_��fON-���	����G��R�P@��>G�p8d���	�>����[�!�r�@d _F�l��C�q��e=3���;�>Vcy�-'������7}�T$����b�3R��R��}Z����ϡ��hۆ��
9!x+�	��ȍ>��(�W*<[#�h�g��vBNj�� 9�Q8R�5`u�1h``�X;�|�XT�$�Z\�`�c
���z��N�����z�l�p��@
��@?��f����y��u�=��yb$�8�J��#�����쑤�aV_J�>�]��7�ę��%��x6�~"��x�4��,�x���_:�)0�S�2?O���)��~�v��&9����67u�;]8�T��_W+���>�ɠ�ꋽ.��W62Z(J��Eje}<�D��BomP'��s7�rA�	n��hwHx`ǚC�2O�/�^�b����
�n�&�6�m�V5���&a<���H���X�e�5ۺ�]E�g��p5;�Oc[����ޟ��d&WL�)�����BS�zg�!�isȂ�)�b��̛l�)ֈ�${^�H��A���o��_ֽyaݯ"9x�76b�%�ݧ�-w��Pb��a?���OE���썦�1C���i�!4r�%�N��ӫ�N4�'��?ң��`�f�u�LJ�a�S�� �h���S@Hr1�6%΢�)�\��;Z��v^M������0�%*%��~tn
^~\&�dҚ��Q���,բY}9`C	����x��PR��D��; P`J�B�0u���'��DF/��{dj�+57�7�c 8��kB�+u��x`�v7��V��#�g��£��H�����񐭦XS�"��;-�`/��>�Vn���3�r��6Ѱ���.*g��$�� ��h�s���*_��ޗ�	��Ɗ�%�d}���]v.+�_�m�yG���D��_��~]}KU�I��ܔ�K(6�	�=�ڥ0�����$�;�*Zvu��T"�讱Ey��}u/[6s�znB{�%�(�ll�X@�e>�:�w�V0�j����o��q���WP�w/2�e:Fv]�@�YTe�1����	�J�2  V��"�#��V�"�(l3���7�).�����:32tj�:A-c@��Q*I=�x}���NkW�8X)����N�%�����u�W1L�Rq�c�0+>g�Ѿ�
��3yȬ�	�kb&H~�(֮ �j�}�A�!�D	�?��-�Esvڰ�[}��/E�͘��|<�S̩���nPI�-)V������ɪ�0;�9TS/]��r��~F�A��86~�[	>D��U��Q�X@.њg��V��p�㞥��T&�W�q��Htv1~��)���_���;5[��n�|Lz�(	��ÄA=|�v��)5�Q�d���g�&�'TT�Ei`���WuI������8�E�����W�-^ks�&լ)���BC��N��:eV�o�/A����&��u�������O�S������3�J���l�l��#�b�)Ek�RjO}	p�c����U����B%�g.C�ա����yt^x{�x>'̶YJ����(|�iP��Z7AH����Z��(偄�*S��!T��c�M�W�~Bʇ��3��j;�N���
���{���u��� ;���&����:.�W+��#֝֍��(X�Ǧ��5M���nDV��<���kO�M<U�����+���S�5Í��d���s��9@"G�'4��<��j�'O���ғ�UB���j<�����JMqf'��F�3-˺̰u(��UU$C���V��A��6�Z�%d��PZO�f��b��wKwy�H{�b$�a I��Ľܐ�9��K��P8��W�؂���5�gw�fKZDjP�@�9�/���>��	��qB$#9dm������S�޶�P-�r�>�w���U�K�J�+V&���.�����.�vdې��Ovj(������(

Z�@J3Bu�� ۦ�s�9��nZN��ݽ/$���bw��p����3�4���
�o����#`�"����Kw#%�� �,@'��tb������#g1u�Q��r���d�C6�E���> J��@��E��*NM]���?����ymW�=��,.<��I�V^pLFu���]ܓB>���_^�|��_�%Zw�`��Aہ��[�����s�:[��m��\�W��s�>���8���L2��ψ^�f{�/yD����]�}M̀������|*�]��F~���q�'��_@���]��o�D�.a
��G���>�#�Qsj���_�
�O�a�'��� �Ĳ�2�S�g�cS��Ϸ1�2��"b)�Z>�G�x��u��D^�4e؞8X�w8b�5{Tjd��lڢ��{1�Dl,�il�+\��媝��Ң���;Ȳ�z��{n/��@�-��91 �3�0���� aM�WTn�Z��1k��	��	F�E_r�Y�OC�䉢�U�AR�/�PM�9kj���v��
t�o�]ݏ1m~�]�k������d�[�����[M���>qQ�Y/��$ٵ񞦫�����h�D#��@̄$�����u���%it�w{�<g��V���㣶
���'�K@�������?Z�����A�������ZZD-�z�����jӰ�O�˄�z:�k��Wp��n��]��r� B�S��/q�n7��n.�֑7���g>USn#� �E�����>u}x�M��Bf��I9�9؎��1�:s�n�ڵ)2��V�`��eԒ>��2�Z����2��=;�@�6/�f\$G��ݪ�0'G8�G�J�vB�c�JҎ�����bQ3)F$����e��f�f��I�
���'Uo	#�͂?j�x�ǎ�3��?m4�4h��ar�?za�~��ML���%��1�_Ů�]��?��x�iG�L#n��;�o9�}�_���� ��j��ݧI�~*a7�b�" ʂ���g��^��׬ F}za+�b?f�LG$a�<ts�$�pQe�P)��u�f�t��m���]�DeFv���ZƟ����<e�"�X�&i��,��A��7�XW�c�!���R,r���~Μ!�]������wϵ��hy������n8��#��*h&67�1��z��L�(����,JBxtP��W=����� c}��{]�o�(��\h<��צЕ��g��p:�i���٧��:��V�ki�yt���(M�k[A�ؖ�;�ecE�r�4:��R��z�k�$?�L�>���ɗj_�R̼5T���G�,��������v�{�c�e�·�R�U����?;t쩝ͭJNh��<_K���Z>�$%-^�V�,*_+#��BP��˕�
X�2��Q���C��쐿]�q���FD)@������r(�uT&�PN���u'ne��wc k�y��TU�F�"Q!��z�~!�����nI����p���!g�'V�цkaf�v�p%�5���`�}lts  ��k�9y��$����A *5ݦb��O��@�r�;��Г*���oh �D�蹾�0ڛ�����&�&�� �^�#��'��V���rѥ�T#y�]Z-rj���s;���'"1˼�Q&1�Y0N@�-k5��գ��J�Sf­�\ȶ#_SNm���%0�+�o~����c%~�H6��f��6���zR,]�)1�=W��ғ����K\�Xzm�J���i�zy�N�U^Ft�{�G��O��@�|��!���vv�n���`g��u'�H7B���tǉ@u��T�yԱ��t�x��i����<�����J�nc��5֨�砷�f�Ə�����Ӻ��DL�!q��5��o�XH3�-y��W?���<��^�&[�KV��|��i1�N���V]1�Z�%�s`Q�O:�Dg�k� ��e�ٻQ
K�"�C
���Ar�^doD��we�^�7�T<%��W��O2�(r����!�����p�K�ͳS�����a�[x9�7��.�oh��a�� ��n#�J�Ԏ�|��"������j�'qｽ��^�OB�L�0�b�aJ��;���W���=���|�٩8�/�sٹ��3�J^��z/�(��I}8�o1�.�:�28x��t@�Կd-��g!��a�=6ݾ���י=�]�>=����}�.����1^jE��ƒ�Iڇ�nx����O�z����fDL!�JH�40�G74�e�F�<�)�cA�pj^���rs*]��BmG�pxz�GY&e%t��L��e�u���5:3��"���D��̶֗f�kP�fW�`Q޴����Vb�a��@�Lo\#f�:���:��1x7Ŷ��ͺC�����ՈS�3��]�o"聄R�(�K�������r���<�2���IQ�\��#�R�]?�A�}r깩�#"�%3�,�d�I��1�梘?ˏ�d�	��iH��	Ay(4�ń�X@,�b�(�礕�]���G�� ���랰P�cՏ'a�d������Z���R�V�l���rx�u����+2X��7����8)v���L<2>���WO�]p8b�\>�!w��"�F�gA�GO�U�2~�N�m��4{�k�=G�`ʐ�������x$YLU҂���ԥ��!����edeDf�!�.����'��z�LYú��K�/ʉ��8\�$B�w���X_���,h�?L��NܔM��){��=�/ ��_��B�����P�#��2t��Թ6���Q=�xe eZ� i�r"�`�����(֖��+��6~W��|l�G��ɢ�=��]"�F�цpa#���z_]���.�bzzx	o���6Sw���N�la�Uze��$Il}R��۬�ğ�71/�ZD8��VbȲf�Z��T�~Y�RwnV����~ڽ���E����Q�����=э׸Ti��Ϲ�j��U��;�*�zܶu3�Ȩ���zQ�>�o,����oC���V��sݿ�J=�%xnW�o���/3y_���H#��Ei����V���t���_�{�5M�i ��������ݵŜUC�ˋ����_�m�R�@�<C"�3�]�yc�X!�,�k7�b�:K9x�I�A���k˺2RA#�(̀���}|����s��=o��4!M���6��eH�yJ�]��u�c�J��W��m���ۻ�f��n�$�sjƝ��n�a�>�����2����˒�V��%�F�1��wX}�}@��4�O��Xr�ZXTg+u!Y��39��Z�[s�δ6�Ju�L�tl*c	6o�m��?n /A�#+��YI��4۠]l�Ksqֆ�Zd:
�0�	ɂ~�U�>S�^���
��l�.����NrpV(�c�\��|Һ%���&�g���a}���!e��>Ҫ�"�����W�c���_�]G�1O�
 O*b� �����O|rz�@C;�~�#k��U毋��y�)��ϹC��J��ޗ�����s���L�hH|�s�<̛��������Tpv�Dc��?c�I��9Mq�(8��؂�$����Zm?��y��+�Τ���v��C�e�̄9��`�H�ќ	�2���MS�Ɲ#��垧!\5I�h��#��_�G�}�O��̇�ȶے���T4Guzb0gmM��+�@�X�Ж��Q�� |�9s3];�6�����w���f4f����"�,�b�z �tnMmɝǡlb���
���\� I�V�P�g� IM�[���*�pN��0R�^��B��{�;�m*Ŋ����ƨ�gTQ7M ۆ�"%��U���ǐ��iz�t|?��ivG�5�����-���	[/��PI���5���g���^��[⑝��1E��ߒ��X;��i��_R�+�����	�EUgZ�|(��N�?��?�Ӯ�9�����A��~8��Zt�*���W3h����cA7mM���?����]w-�<)-&�*�*{A��:N+��v<�n�ey���Y���H�3b�K�R|���'�*�)U�������F+�9��l!�AkN��`�_2ࠐ�՝���O��_mb9'۵��H��J�i?���,��]Y?k9g� r���,�j���*��'E�b�VI@��m��� _s.rZ'GU�} `�(�H-Y%L,��� �07B�~� �w/�Z��uˈܽ?�h�dv4}5���b�Sf�P��߆�*�,$�Zb����';�-ٹ������ѸS���W��U�6�`v�5�]�ˍʩM��R��U*�����FB<��}�p׷3��g7�P{fL
>�ȓ�wQ %�bg�hg��}�\��t���*�`�xd]��I�]�C��&��8�n��`q�VР�I<Sj3����r��O�	�Z�s�q6�,'4�v2E���氆1ir�*a��}��Ƈ��ġ�at()e���{4�Vm1-� �<�9�XuM��g彿m��P���k'���;�N��<P�׬����fD��7��0����WQ�(� �z�pMP>�~Ơ-���ؾ�eޯ�)o�z<�<�t��Xu:�l����zBP|S�q�5	*�B(2�C\o(�p8��}o uGf�B�.:;�7���D�>2�s�s��!Sr��5�pP��"���nΚ�'j�ow�K
�0H��귎s�CƸ��b1{�llP��c�&+nW	]������r��±���ϚN��H[�E�@y>߻�z��7ݽ4ā�%fhW8P��߁�l��|d'&������9l?��vS`���aɋ)2򧕑x�j@���n/}�d�qgЕ��/�f�_[g�u�ٶ$�b�ל?F�(ܧ^x���ʋTפA����ɩ���lo�V�o�x����:"�����S���P-�a���m�������E;J�R�wEڪ0�Z�-F�n@�*�B�L�KM���[�1D�?ޡJh�Ѧ&�����s-�!�b��.��hF_����� �iv&H>%�k���<�s�)�-ٓ�J��h�֩��7k6��<z��(8�.����ACV퀗��2*��uW΁"�RM�C$R��کY�`�vw�q倅��R���mi���ưJˬkH�u�����V���k���a��w	X�̇�|uj����򪙁\g��f;�B"���P��p�y��a�6��m+@@�ͣ�_�]G�:=Ǽ$w}�^aǐ^� 
^=�L:o�#����Γ��7�6b�%TG��,N$ �^����2$��}�r�U=�{�����!�YO,yOޡ����^g�ח����#~[�c�YŠ��wђ��Z��*XX#�;�0.bo/&������ek���.�&'��F���+��r��Ԅ?:h�Uz��ݟ�x�Ԓ���	HL�ܿ������=ۂG�5\M�Gߙ���Z�	ɑ;��Q��A'���%�/�o�*b�Z�5��N�=�٠_�N��
;�qs�I�])�o���Ӿn����n|����+P�fj�)��ձ��X*��'U���q����7�cj��[�F�2�M�f�ȧ�j��_y�~�O�-:싪�%Ê��Qy�iպ"�˦h�=�T!&Ŧ���L�n�2�\�Ê+��R�&��Tb<L+=J�Ѥ�������w]���J���"�.�JH���ƨu6z��d��upj�s��#�b���vNPTb��7��`zJa�tw�T�
6)�7P��>TgS�F�G��o�$�]��#��e�\�ë^k�*(�
,U@[1:1ɴy�����˵!�lݖ&Y	��QPs�\|��>ħI��s"W�j�|�q������񢼩>d������U�����a�K����j7ʬ� �KeAz�Y���������&��t�a׌����,ɜ�%�4[�`cE����)[�niv��L���l���EMM:��%��c�5�ʏ�B��5���{���vZ�r�6I�K#��Q��تMZ���'[����5����%��yq��U���ϲ��f�����G�����P��M�[m8�-�-evz���F�1�L�,2��#vr�:��|���� +�c�m�
��R"ŭ �@�5��!v�t�1�&\O��i���?��c��3\��f���GN1%�n^ݶ:H�6�W'1-{�I���|���T~��.9��lQC���Hȣ��(���.|�c�MM�L=��_N[r��$A o+������C&�4	�RM^[B�]� (��T��}��D[��$�ĭnj�=�[�S_<���z��q���2�S���{�oξ]�,��I����݂+ʱ2��5�pJMM�����Tcp��E��f����8�H���~S��4����������:dv�kc���IL"�n:���8��oc޼ ��U���|GT��=[,d�����q�5�&�9)��w���AY���D=7�)�Ԇ�Q x�`�l�j�qw X��
+��`�;v�ŏQ�c����W����Gҋ����i���,x7�H���/=vg��&Dt=��2~{8����Iv!_��-)���qH:�Z0j���cx��Y���c}^��$5�=��8��th���zτ_�ur�OD��r��a�1(�	6�9�ڵS�v�rb�7���Кm�
*�9�]^?�-wL�n�I�{��S�HKM����a:y��~����{=�^�����D�� ���Ĕ�������[���۔�� c�")���	c(&L4�B ����Oy���=�_�
5ߵ�;���x ?^���/�z8��Yeؙ��#gArD��$R ���ŋ��p�a�7�x�xެBge���GĶd�H��6��.�sھa�Xt�P�/�$�*��V�c udT��}Y���ZL��@p�A=%ӠV�
Þ����G&�r�����.��mV�*x��|�*s�n{�\>�3�o2�+��t1I��Ph�I��Eo"2 �d�O�)��&�%���P{>�O�k+Xl<LWĘtiJi�!�zg*NOU)��M�6�,F�k�����1#"! �0<?�D��;������2 _(Zjb�P|ƌd�c��u�}���y�*@K��?�A7K�,�w���L��Iu��r�R����VZ��{SϦ�$+��a���Sm��s�xAe�����{�M���M���"�������yx=fY�ϐ�ceaۻ�JȨ�k5���,H�z�6A����Qg�{�$���\[���*�k"���r��|�W�Ս�k�8���s�b��}�'���fq���sB[���0���E���}п������˾�hۚ&�]���؍�4��`��r�]�z�D���%��zS�h����FHLf���<2�=�L+ї���-v�#d�����pP�d.��� �n��K9#��W8Dn�34/6l ��VC�?�5ba��>� W�˸�.G���*Y�����:�'N�e�7�a��+�Q�ѕP�l:���W� cP'd.�xǧ�]���M��8���A��k~%>
*�}�z�e�ǯ�j�~�&kz�4�6ule�f��\�YX4��Ъ���G�RK12��)��ཀ%��aF��Õ骕ӕ���rS�]��E�� �dvd��i��v� -yt�a`�\&�&R�"�E����Z7]�,���ɑf���`����.o����vJK�
�k&�P��k�M��r�G���C#$���s˻.����	���D�� �S�1����[��VE\�G�Q#�o�W�cE/��;sU�9?�N���H"������/��A�{ZF�s�p��K�ʃw���ؘ��B�lc��S�녝�C�yU���M��y��d��O�a�jm�q��[���r�:_������[	�,�h(�=k^v+Ruf)P]6����Ђs"�3���6�3QṀ<R@'O�p߃RΫ�����[��"��z��0.}�NO�]�c.kQ[��heIп�$V}N���"�'��4N��u��P�]s�_�	�Fh�����[+�h\��c��V�FeeǪV�c�MÎ����V�8]��pqm�,W<C6�w(��B`���R�#j�p -�)61*k��Z)��'v\N�.�U�\)DPRHGy�DMn �������yL{Ҍ�U.(k�ǡ����#R}g��4�:b��'���9δ^{���&�-��IRwj�.�XK����wvЗҪ���[��<a�q~�@ݮ|}��	ow~_�qu� �rp�S�`�3�6�FFX�Es�9*w��$O6A�sC�|�Ќ�Rު��_�>T�) K��w��^�?�U���)(w�|��欀䡼���h}TTq(�VmڔkE �0��~5��'d%�8G~�EO��2����Gy�����?Ӿ��r=���9{��H�����I��d���?�D�]��k����3L���L��F���ꈟ�� �́Y��M�5�f���7~���ײ&wV���s>=� �%�|ږ�Aۼ	����j��đ�O�Ò�$i_J)~�Õ����8�̆;�l�G��]]�a*�|�WƟ�䦷:�j���k!�]�q��r#��U�̼�NEI.���}��7p�S�%�_��я�n���������-}p�u^��A�����ȩhKw% ��xH$�Q{���T�I��T��o��;��F��ae4���	��(u~�mp��d���ߒJ��&�Ls��H���m��@�p�B*x���x�8��+�� �&����X��vù��|��0�T�V\�#����w<��
��h.�
��sk7X���}W�Q��0�M:��r,��Z����D��ڮ+-XB�AU�[SĦ��G���܊�)@�"���ە5�V��2��Lwˈ�G�3��9����.(֓�\�!�6����u�����Z5�#*�F�{��,mEdg��!ېD�2�
]�jȉ+� ��h�e��KR��^'��ÛR��t]m���[�vd�\w��E,�gOݎ���πy��VH�V���!�lNT3ZGNc䛜���o����Uv�r��f�^�ϵ<
�%,{�p��j�e2�?��(��#Q�zJK����&�q��Mc�s�_B4F�o���E`�*'p��da���=���5�Z �%���Ԍ������I��+68����I7�?&�û��K�gȣo��nlC��~�U�\Jo:zWԒ��ߔ�XC���,�ij�W��rn;�
����|VЄ( �L΃��}����;�<tK'�,GN�h�7>�O'��v#[��G|�6�4f��Y�,lH��L�)!�|2�L�|,�O���vUӉR8��F
�P٦���ln���*�p�:�q2����j�b>�Q,1,5h,N}[(�����i����A 0	�oخ�/$��$��Oe����3��ɛZ�� N��%B��g
��S"Z7.K�6�8��8��]Qh��
E��I{����+q���u�u�/�CRzCQxq����{��Ưo3�A�yM�A�Ƃ� �ҙ*RӨm�T޾��WXތ��(~�l+���F8�(΅�b���pg[�[1�����`��`P�&Da�"�WDKde�YLV����i�`2�=�Ee�aZM�zل'��+�k� <��3l�����ʳ�:,�U{^�*@÷&���T		���T��)x�?dФ}�6*9��6�5�2�ד>�N�����õ����|�H8a�۟�ǔ]�^�8z�P�����#����
�׽��C�w�u�a�k(.I{��PUt�yh�o.�|U�!l[���i�Cᕭ��N�s&������qÇ�;s�fz#rTZT�<֨N� ���mtn7�΀��ϟج�P��
�����	oJ�s:*8��f�XJ��򐛰���S1�S0�6�`����Tҳ,_F8
�oϳ,&�Ϋ�#[��B��SÚB}I3�!Hb_��N�b��Y�u��"��8�>6�����#��y_i���:[��e���}|���mW��	��4s�\7E͙2�Z�O�Ԅ��V&�1��>am�W��U���F�̗�c���)<�$�v��W�A�I�j1#�әϒt�HNpb8n�W�/:e�c���1S_��Q�mfkO�������À �W��0����ގ��m 5_�r��Y?�V���B�����T%{���($�!�Z�3��)X�	��>�=��j���Q�-�Xea��bf�~���f��n* �����m�`�CB����f�B�}���M�фgh�7�L�+Pʘ|�q���zt�2�=t�^w&.6�Fpa��Fט�.�D��?[�J#�XkUvōwQ��F�	C|���8���f�W�A�J�k(�x�-I�*��j�k"�[Q��p�k	J�>��S� !������`�%�H6����))�+��9�k��>�����"�w�N�(3�����=�z	U�-���+�	 �~��i�%<u�x̓�@��7���f�f����P�@��0�W���4Qڒۘ|}z|/h���)�@�yW�j�{'�B��wMp�;IK�l�ຌ+��VWk����:��t"HH�|�v��@d"�[��o�GWL݅l��p]�땂�'�y
���"x �F�xV�L�:�0�!ʱ�:_�P�w��og�]�ʖ
�	#<�uT��$���%�\,Z�4}��c��.��h�⦊�x��	��
�4'��7� F*}���ps�����**%܏as�����*&���4���9w��������~�6z�^ϩ�]I������Y7U�s��'B�>ђ�����v���K?�1���������}��e&��RIv���y=�-1=�|���g\���y�L��婘�p��.��ʢ]q���j����Pj{��3ߗ'+5�T��b���/����	��U�_�=��6��b8w�E�������} ��A��@۾����ECZy�!�%-��9��Up*ଡ଼�F��q���������tU(Ҧ�]r*p�u��KK�C���<1L#)Dχ}��@����㧘zg�ZP����F�HN�A�2�7���Iƅ�U���R9F�:����o���Jիe6�1X8�3�=�|�j~pbi7\�]� �Ľ1��%��@U�7!r���k�7 ��p
X2��hQ'| ���b�܊�.V�n{G��7��&Wno������-`��?�X�������CCC_.\��\@�pB�Ӵ��?e*o��(�!di�&@��_d�Eynp�x+}'��;�Ucy1a��Ο�ь��~�X0^�4���ʻF�a����mXT�1��x^��؂�Ꙓ�b�c4`��aD�U8��#���3�M��]�Y�Lׄ9S���%,��d���W`�G/z�
���#'m�@88-�i��W5TDm�n	�s>3��q�|)w�7n�u7�(w�����k<���NwI����������L��-���A�"<InrĶ���O;=Ð�M���El�ՠ�|���}y�~e�v��!���m����|;+��&U��wp�"J4�4�R�a6q��3�R�i�����[��i�ܓ/z�>Uș��<�k	^�j�b	\�	KђD[Y]5��!hi�����]�ql ݽ��o�^�!�Qi�q�2,4Rſ��+��s>����L���V:B{G����P�m��c�����Y`����-�� gl�6�>�;����=�J\�_�ꧫZ�\6���ͤ�^�a�����C�	�Jp��r0�����:�ƉDUtݣe>������_��ԙ�
�-ϛ,�C�}sb0IL��l�����K�r9�^��fs�i�=3�F{r� 	JL�J�ۧ(;�2.�uѼa�Xa�>��~$�b�]I�b�_�h́
��d�N0���|&Y)�uu���cRF�V�A�y�x���4�j�N����%j�ǌ�'���˅p����uG�K򾴏���_K�."&�����0k��B�f�r^*If���!����Rm���:`5�l`�n5@������6�Q�"R,����?5��j��� ;%V�OD�OtՓRp��A0��Q����i���ԥ�b7���_�:tz��c��G�j��Y�`?�M�Et���X�����m������e3�I	�7�
�2OtI�A�d�`��K�j�*�H_�Ԃ��^�Q��Z��A#����ȋd�W⧿��u�}���AF��ҰɈ�]l'�
�C�ʃB��#���J�T'#v�霟�ZqW��_w�*B����d�;�H�'X bM#W�%�0�~0@���L��r�%�4"�_ZϽl�#�$��V3�55�W,���J9�Ӹi��|.����$5Ϥ�}Q���6���#�/���zn���֚�����g���ebo�
_������,L�	�UnM��F�����q�$ėT��G�Z����~���k|X������75�V��O��c�!})_5�Dm35̲I�
�E_D�o��z�AWw��pJ�hcmFl+��{�*�EYҚ�؄Uѯ"��z��O��J���5�Bw�p�}8k��Y
	컡� ���A�=�V��6A�5#D�m8�b
NE�}5�uW�PI-d?-�u4�ZI��2��I���N"Q+&���M6�����6*Wg�A�Ha��FQ�]�;��q��Rg��)�\"�ЧL�) ���uY�vh��jo�O�C�J�sZ:�y`��g%�v3�&w*�[X�ʟTt���>�v̚�����q��aP����Q�I����p�����lt��ZI^��ȟ=D�k���F��p*(l�p3ut^aւ=��k��^ ���6��i�!��/��O/�A/�B<���b#i�aA����c٢�J�ܫ���O�J�`\�'(¶>���g,c�wHoԖ{���_O.���\Σ��NNۿ��uH���_�S� ��[��V4�YΜR�S"a�&�8��h����zz@Ox{��t\�ʺz��	���9!~D���=L��i�'���"ܺ�� ]m���8�����kE��N(�w/[���+^Y�8nk��dSA�Q�����{�9��\?@�:Yd���.F!�.��E*�L���IV��8�Q�ͫ�V��8�C� 5ű�^
�3��o�Դ��������74@fml�T'���0���ʲ9����o{>�be�������n����u�sf&�ځ���S��&�(�*Y6����SX�7O#C�[r}���+����B��&G���Q6x�_�ߨ�R	mj"'`i2p���K���߉��q�Pk�e�-z�s
;s~2��=�؊up�I>��|�u3eV��5\�	����#����E��{�E�M�͉�����O�3YH�\���7})�#L�<u٪B@����p��P*�ߎe��i]_z�o��/m3
[-Zi�V7-����C�!u���:a�^b�e\ޥ4����,�Ԙ���f<��?鶚����Ǜ�<Ud�ӵ���6px�{���{�O�����z�w��}�$�[��:��u(�;,�*ɔ�.���m�&[�.T2���e4��Xdl�-�'G�_�5oRaS�U�7�F<<��,�[�[-�;l��Д�/ r1D�G�_(�?��*�hžX�}V��pp�f3G�DǮF��T�}���e��b��;X������En�Rcft`�i��YGᕜ��5�gP2�t-T�p�L���	_�XdT�"����<k�$��X:��!卦:��/���������c�m_�zocjΟHd�{�m��]���?`[g���Z�U���<�?���'|���xlw��,@��N�����"��N)��:<����]�o9��Lg�ʀS��7Q[h�XI�kW�dz mˋ�x�w�x�o׍�䈏{���Q~�)�<�.���ޥ3� =A��XѲЏY�j5���,#Fe�f��C0���e����.���t� �i�I�F6��:xְ	�n2�"s��I�����lI�k! c�\�s~�3��ڳ�8��n�Ii���x��E#��L	=ė������dk��w�ڈ��ɞ�'/rs/(�<�\�$�ct33Pv�r��4*f�fy��>��A�\���pB2׻�Z7 &��^��' !�3U�l�3����)�|┙��ME|�7�iJ��aN��Q���zW*��L�X0ɬc���0�z���)�Cn �}����\�Rb�zD(�i�.��S@@���ٿ@��|���;:�$P��۟�M�,gF��q��9=�&&�]���w���It��Մ���a6�`�<K'0/��Hb��T��Y��y����qOd`h�4����e"�8�l��9���rC
`�.�n�SG׌e�7�V��L���mjT�ū��c�h��/��vd��w��"���=c&g7�Ӭ�BOǐ/�c���V�I��2W8�!��UU�y�Ss~�3W~��
>R�GS,�1�k�~��bc�&)��ڌ�ݎJ��I�u� Ŏ���[$S��P���[��9,G!�R�M| [<0=�S�c��O��*��W����iE���@e-'��ǐK<���R|�ԇ�����̰Ta��~K�̯^c�(H��a�\�U�"���U����`�L���]T_��{� `�� �|by;,�m0Pr+�~_j<��..G~�s�C�%v�bz:���%��)o �<�nVσ=�V̏L��nb���G�F�l"�W��P�Cs=��Ւ [�^4�D��L�G|�y���wrAOiƍ�UrT{,���������"���륁�b���%��(�
����h����zn�{��7�j��q]O\�|e��	hi�qx509��ݐ5-?�԰Q9=?1xƜt�	,1,�;�a�/<��4�����_SMO�@K��	�%���οo���/�D?�1�%v����~՟tŏ>B=tף]WV�$���^ST?q]��&W���른�߃{���i�O�2���p�BHa��2�h �4�/��r�W$�E�ޓs�NFj�Y[Tg>��K|����]��@����ݯ���_��0��~�z��٢,2�+��`q���Ů7+�K��wO#�Gl���t�|�@�22���[]�F6���A��GФa��B�8�]&�d�=����ꕾ|c�>X�sq�|�2��a��"�y��G�g�*N�>�'�2u�$�?`�=��Ziِa-�c���t	�����<POr�M�>?��c:�	?�.�yK::SS�8n�MIζBL��!��0��͊��L?�f��QX3�hQRa~e�~���W��6�/�Z�����k��f��\�5�:ף���r)�+��v�`f,�0ܑ�~n�<�n[�K4���ti�j�DU|�1��J�eS�˝���K�o:\�� �r��Ư���ڌ$:����a�I܆�T?���M+��샬��d	g���6�^�Ig�Mo�)C���F�BǪI`i����6��ea�"����'���	�Ւ�$�hg:��qOKaڛ��|X~�L�/�/�S}Ⱦ1@����9�9�����I��=�W�V������gږ\����K�Q���i�>62]B~[�qz闻'��7lEۤ�
�
�d%ٷ��k	t�૛,��L�M��u���țB A�l���u�.�Ulm����?Ϩ�(�
��h� Y�I��N�����%�AoY,�j&���\8�@����?��@�!���������+iZ�c,~Ÿ4�0�-O�����T����I���E\ M8R����3d�y�bގ���Ȭ�͍�p��`��6\u��<�/��D�
����胇�:�	ի���f��">�4�^���ϸ2>��Bf�e\wja��p�B����P����	�dz��B>��[�����yW9Xi��O�H��˯a�7���|�KcX�8v���ze~���]r��JA����r��EB�{` 5G2��,#?;��~u*03c����=�dA���_�S��b�m�����M?
�CYs��LP�eN@	�xm����)��\m����"1*}3ȿ:��UFy�7`�OԎ�fE_F��+鞙��Q���G!���+�}6>W%g�z�x%���9u9�9�y�I�"�Y��4^�ߪ�ٟ�<�U� �W�3h BO~�z�Ƿr����}�!��wϷ��n:T��L�VcvƋTU��$�ʖ���]��\���<�3�k9�:FF�E�)\�?f����<b�S&�ȕ�e��SLS�6��"�[ؿ�"�Uh4ѽ_Z��Ȩ�ȅmOoh��M���$<_��6��E��r�� [C1�����4��R�Í�JV�ݫ�d㱜B#��;ؒ�L^;?����3�B%Bt�!5I̴WW�t.G�|�7��А4��B�$r��B,��]�y�Z��eHM�x{��� �A��ìz��Qx�3Jem�%'e2?w*���ӈ� � D��0GD���/M(8h��?���M�X���a���LZy���X%h�k�'� ���e����<f�ʱU��ܭFs��&a�Io��*΄Y���H�E�gs$X�*��kaʱ�y���z���Äd����M�],��W�K���b�ݠG��a��2�x��Ʋ�q�st��]g���6ߪ���h�0Қ����p3|\�Z���*�2���������fum<�Nz��E�L@h�U�F���{����	
=�y��>��bup:���t���C5XZs8$�r�I�/ IYS�.|cՎ-�4��!�`0	Z�<����uܹ�eJF����I��$+HP���I�
����V��:�\c��?}[kT����$��1u ,$��XDd
-�F�� ���8[��"@�~��vn�0�����{�Ho��b����{��[Rb��¢�d[��vG�Qʉ�\�{kg�g�a0��osq3Tl���#�����J���+���U��i�����܀{��]�� �l���M�@WR�� %j�L���G�O��+������{�v��K	i��$䯋��ȩ4lJ�E�/����Y���	#�'��͜���Atj��k�pt��;�x=���y��S)t��߆��p}8�V���6_�_�;�����/=��WP}6�^~�(H������铖/�}m��_\%��m���,�"9�4 �eY��z&@].����_�o�y6���0[�d�>��^-б�;oJ�蓗F��DQ�'�	^�V}yG��9��}�+5y��k�ܗȷ�o���X�U�Lx���DWx:�}���M3Nh�͘���B;���<�j�ۇmbI���25tֵHa��ct�N�E;i
�"�w��H����Z�
�BA�n�ܛ5Tv��[��G(1@�z�U~���h5��r�nY��M�>��ɺ!?]�P��5�O	(n�ek�`����������v���oGִ��$!�'�r���~�>>�'DyA�s-�V(�f�R�9L.0�*�)#B�\|>	*�w��#��5K�l?!�i�X��S*;#c�+��(>L��o�Z�ݟ��i>D�2B��-S��r��S�`e�"�V=���K(��h���ﶜ }�\���Kq�˘%��<#�x��8�,3_m�Up�(��%+U6�Ɋ��#c��P.Zq8�5U�܎Ğj���S1�7ȏ�d�v��!5�d����3\��w�0j�����ľ�x�����WB�f��o�@ ����L��Dle�ô��[�#���0��S�-�F@�uU�Q,hv���S6��4����r��F���*��`Ą��#+E�Or�&��9�瓯m�c��g�rz��2��5(�F����#q�/�h�����׷���)P�Fq��,Uw�N�Ɉ��>��{��M��@�\5�x��s���5_��2�Լ��@���<e<yDV$�y6ē��r�,&ϩB��Rk�*�҅n&9�3������.Nb��Ĵ�/�hqq��r��lcTz�/#y���}��E�Y���|�qwX�b�h�@��<o���	����K�9����=V���a6�Ⱥ�3"���I�Mj�Z$�����z�ea�E[=z�g���Zt�aC��N-;k�r����z��7-���T�.�l���#]w����E�HCb����ǐy�;�i�#��XaP��R���������<�ف�,��E�����6�j��8�:e��������7ъ4�CT�=�t��a�ǐ{g����㰋��
$8L
j�.	}��@e+\vr����F�ԼH�$��U��8yz�O@�Ŗ�qp*����Q(������{=�9o#��Yw�8�0
�xԮ�o!�m�eHc��܋�P|��%�ہ�u��~���00b9L�D�h9�<��ڃOS4��@�pe��뮈�i6&\�6@��0D�߲�V]�G�퓘�o��P�f����䡎�������i��]᰹B��'H���P>jP�*���X9��Tyb�����l1�BvS钯������F�c���~���Y�:�#I��"�����%&�s:u�C�9%���1��hC�B�Q�jE��'h`��;%�H�2��d[
�]ޮ=��l�%�Nv��:�T�����̌��z�Y�Tm����L"x4���oy0t���r�Shb�s�A�ƕ]䛁{K���NX?�{�����,a�ޝ����V���A��|���8Rpj/i�̔3˨f%h��Fx��v��(�f;�ck���<[XĆ�<	u�ʝӡј [Z�{
v��@�r$oڕz�)@���3�	�{3O��)$<:v�/�HS�T�� ��.!�¦��X/�,�|W�D��_ʃذ��<�������˿��I%�D���*L�0JZ*�C�����1�H�b2t|�mbB�$f�ܻxX#*eb�� ��V�4��U�6�+�]�J�5L�8ԫ�P��g�0'�0�e5*��,�ܯ ���EI3D��MlK�m�����$�.�?۳��v�E�0~0~[L�!w5%y�x��_0�}�'>:/���&c����-ա��!��O�72&�4�I �66���e}}��6I����c�� ��)�r�R�x"c}Ad8����T^������Wڼ���cjy1�� �

14�� �7*;�t)d�s�g�bH��BY֫�6jt5�����ِA�)Iyd��Qe�(C�2M�I��D�G�4m�>�"�����U,d9�.�Lw�$N���&�\�ˎ_b!jAv���fW�=`���xWv_(~#��2��&��s��C��ː�l��(߇Ue�:��j1��?F/U�["= w+�]�]�ۏ�Y~�=�+Z	�lV�,�_��������tEA��z�ě�֬�(aש��s��*���B��\��vl8/�'��މr����[`P�	S�[���a�#�Ӟ�F`����п��֐�2�T��:H5�L��SOoK���[-�e7���K/(�
Ť�HD�)�\n�Ți k�۾�fD�T~��G7��t?'��e8ˌ���Yƒ-)6��i�����W�V!!�����/��'��^�&��	v��)��Fa�4����u7�՜��v��/�Sz}y��vB�<L2QB�+��μ�8싟�	\z`�U��u��=$�p{iIo���l�6�d@��g�W��~
�Mp�����f�R��U�?�_�2�W�Cr��P9���qkuDbݍ���/o������/��$�L\҄(R�j�-��@[@���iat4uu���r!����1���d��"�R��%P�J���3^)����`��@k��]�y���S����J$��3�#O�+�G��Cpe:f��!d�7�c{�ZTTE+��O����P�K�]����e,��G�Qƈ��Y��6�ϐD�V/Q�f�훡'7t�a�e�ڋ�-�VmM}2�ʽ&������pB��}�����NB���JC�*�I8d�%�����z��ȣ��jU�ɬ�ډ�(��W�ltN8��d-�#B��@�V��!-V��o2�f�s���+{��%3�	Y.�y�֦�mZ(YO�0�>s�}/k�����K�+�_�X��l�>����>�Lh���.�j�V[�!���>��0� �֏��?�7���p��KW0������qZ�ldK��\�:�
���^G�<;���!s����ds�@�����H���bw&��+G#HZ#/\\P7�]��ߒ�Oh�eS��n�ʎ�����'��P�����gW�޶��{)���D��ZK��V��R�؀�F���/?�L e�Y��ﾟNcçþ��\,]]�λu�S�5܈X,�� �Q^��;'��e�(��g��u�6��
J��i8�o|��qdy(ڢ_�����\]����zA��t�WKd�Yh���D��'y�g����Ͽ��Ru�&�r9�3��uR#�E!���D�ކkˏLB̎�� 1͵6�#�FvE$n�M�x�*���k�����\隁í;�D� �A>F�5�o���=n	�ԿF[�h�b���O#c����[D���0+#��a�?�\��p�䳂���!���ػ1��?H� #10ф�<�^aƧzG���2�R�����Wg��w-b2D�Cϊ�V�m�Oc�
)�8d���q;<2� W�Jݦ"
v9�$�k�޼
7���X;[W���#oo�Y���h���˘ �ϙ��D$��QZ��hE?�kE=5��m^�M��E
u��}�>7D��^Oi�%�+WP������͞	K��(k�9�Ŵ���ew�œv]�����:��S����b�=��'�j����7��K:��߾�'s�3�p
� ��zĳK�_|^�W�s����UnQ�$��}ʻ�_�o��[u'������F��W�����j��0>���]���ρz��C�o�pG��˛.��$Ы��5�$K�s����>��`1��x�Z͎��{*�ϴ~�HWkϐ\[~�����о	8&�����{��'�.�Rf�v|N�.��I�m��@r
�� �O:�#��D��<f���O}#��s�9KĞ�J^Y#��������WN*v�L�J讦�N3����ٛ���Im�q�����6��v�gs��<�D��'s
WO�Dw�\u�l�1SB邓h$�r�n��uS'���O�.���vs �Bm�?����_��̝�2����&��rLrf�+�&�럿iGCp��O"-F	6�3�i₴Ӛ��wG� �F��C%r�\F�v9��?M���\u,i�m�Dӗ!�SӢ~�D�Tup�J��ާPLyꩵ��=��a����vW���GN�����09�ϔ;&�F�}n>֘��E����xΪAȥ@�	" K������5����"���	T�J1�80ǯ얷�}���b��3d|]G�`� �[7�mܬQ��%Ŏ>O��-I�I>�뺧�ے� ���7իi&��%��؅lFOݯ^W���S��L��I�hv�L�S{��Xץ�� �\CU�U޲��5��ֵ��������	[�H��K@��Їq�s}0'��'��֙2�Δ�.O����o|r_/f}��m��>�B��и�P,��-r_�'n��>P
�(�*E��FG�3"���X������SR��A3T��é�q/S�S�sJ�G��3L�	��NecF${�.|q����@jϬ�5c������6�Ւ6TY3�,�{�8L$��춟5c�%0��1_�Uw�x	���w^n��$�VP��Y�Y���=��s�4�]4T�z|�q���b�$1�eJ�,�D�b�tym���_�o�٥��Gk�"Q�эt�ǹ�s�D6DVs�}��\�=��9�s�˨�S~��2�ﾡG�Q/��9n��]�;+^��d��kL*�T		1��MڔfB'H�]���#��*�G����H�m�Q��b��>9Qko�����,l[Ν��Vai�D������S�Lu+������@��B���g6@�+�$� �hkD��<:U�s5�Q��&�6�.�:�S��Y"�b����+S-®Q�'��`�"�p�C����k�p�f:C˾«E��s� �S���N;� y�˲�1��B�׈HRX���oߗCT8���#sO���!�݀����`��_@�Y���ξ;�,���Ke��5w2�!���~Kh�`�k�ǚى�ʍU�S�[�2�{����Ѡ ���)[\Ź�Z�vp	s��w1Lk��g�;�iN�b���G��T�a�n	�aM3��P!��F���}����3������R�]��r����7��-�[�rB���ɟ�+�Pѓ����x�";�l!W�"",�R�UptF�t�@)w(I��e| ���4�gxi���XA��n�Dz�'Iu_���>�b���?�%�����>���FZ�
�]3 7ˠ�У�q�c���t�G�Iy��������XZ���Ckf����h�R�xׅ⌑����		�X����\3�k��Q��VS�@�`�O�ɞ�7Zsk��R��0vZ����E�ܭ��unm�	C7��&z������"F{�M4R����Oh 5���J��y�%�����0Y�7�
��A.<Ŧ3���L�@E�-墈ܨI�^DvY-�R�)���x'8x.Wv���E2>)(�����^�3EY��hJn�*�`�h]5\��ARݽp��={�$��gdIR2*�o�U���c:��4�[�W��y����j���P�����i���?���D�m*���ȫp�w1���Jc&��:��)�׈y�h�\K���qa���VK=�E. G�	��$$�๦_�s����!���5j��'�9�������*��=a��4��N`7��d�k ���t�x1�4�w���i|�;J���tX�%n����ms��p̄1b�����U�/��70����]�ꈚ]��>r�B��B%�M�1K��wPo���dߊ�`)����e�R�9�Rz4&}���V}��t��cE[�v�a6����k��3M��7l�A�y���p�YE���C�o�tؿe;F�*5_y���{D={��ƾ3nR /G����E�����FE<t�����Ƙ]���>ي�Hq�쒗V=���;N�1s�7�5HU�Uo�D�d�`�!��;]���:��{nd3<����� ��A�%�Q*�����9�	�!�v�3EI���&v綉ʕ俕2�W�Rq$�뼻tWyZ^��RX�s����-v�0ic�� �ԾLK�	����&U�R��K��/���}B����Ϥ��8kB��v��y�%`�����k��%?0�zZ������pW��)Pk����� �T��)���K�ɠB�4n�?4�*�&���R�$˄hfj"@�R�߽�_��'�w( CRtN��� 2�L�QK�'�8aVj/7���) ~�{2U���N��*m	����@s�x4$������D����g7�� 8+�cB	�8��J���0��U&�Y��e����(֌�� ��ϫ�t����,y%��2EM��x��KA|���r��?[5y#r�x���Ѣ�\��-৥=��1�	�*Y3e����Pz�Rb[I��������T�s�V �F˜������"�" iQ5�L����Xo �7�=���ps��|)-�&a7��t�9���}�+����������X��< @[�]^���4���O� ��\֑L'��[�r_��`��~�Zv�� v��V�}B�N��M�`BXm���I�A�wDRu��~G�f7���#��(�k��I��x���s�C�2�B c��L����>���}r��F�sz��2�+��GB.�Wy����E8�c�P8Ux�g��70��j{�[�rgٴn���`<R�6��}yĘ�l(�/IŌ���_���@��(�V
�Yť�rg��rO�=!�<�ϙ���@d�G$���ImHb�O���Q堞J������2�fu��O},fI��⹏��(��R���x�{N�9qd�!&x��FhI�rs����'�ݒ�hV��(�����PQ���>T
i��)�[)xm-��P1H���W��\���I�U_r~O?��7g�~z���l���i�،���u8A�r��Mǀ��B]1ey./|!�xd����y�fw#79Q+��"_�^�{�p3v|�6��[T��`RN,yS�dO�wz�F��jR�G�?_��`��B�47����;"/Ջd`�U��. :(�swB�2c'�86�+�a��S�_fd0u���^��ϫ�V;�(|b�Q�^�P5V��fO~�,�D���y�6δD�i	1�M(I+ag^��Bi��Dr�z�
�����R\��I���+V�8���,��t�gNV<�������C��yw�&e�� �������'�?k���)j�*d�[ JV)�c�"����SA�jK�N�v�wah��"�AP6L����"���ӗ���ђ�B!j�?��}�yϰM�H5/`t��e/h�x����dFf��QW|ξ�y�[W�Ss�K9�c�"�aB�U
-�<��<66[rC���R�@���+1�m�V�vܨ��� �R�9;���e"^n5�\s��`��_�_1�7���}(�u�
x�֗���z�+^#t��E����.�	�m��&hy��Z�j*�gP;��Ylĩ����$Q�l�=v����;�|߇J
!_�`Oe���G)��t\gP�[=E`�fO�������Y����[�%��%4�U� m�X��Md �$N�+|TˢS�JI�t��}3���q��%��.�k��������=T�����VE;$���Ia��F�&��n���	+X�P�ݶyZ�W�vf[ i�s7�}����z �0X3���Eq�9���㲲��D��-QMV���'�t��_B�/>Y��P5Bw��U����:��|ܼ8�18�VYMm�D
�-R4=�Z�;>�\�Z�t�'�G/�d��r�	*��X}Θ[�Q��)�㎪�8_R�gI��}�3+�&�1�׳�u]ϝ��鸚�j< 2K�)�{�62BZ�(����!X���{r]|n#�C���m��z�g@OYښ�\��?���V+�4�d�� E"z����,���� �BM�p��m2e�AxQ�d�(x�g�}:rl�ҍ�>�q�q���p��y���[���9�2���~����e�1�ٍ��Ǣ㌎I	�ƽ2�L��3R��2���0/�J�|O.��]��f����*_�6��4�v�����Ә3��dMùE����E�j�K-D6 vy�=D˓ϟ	yٴ,w g`�y-| ������g�t?J�W����BO��m|%e;��-���чOf��	�j�żۼ��|�rz� 4x��L�k!��t�� #��a%Sv��H�Fg&��Fr�K��n�P	���KDL2n����{��k�ze�6S����g�a�(�cB�À�}�l�*'��|<��t��5�e*݆14T)Nw����9�2�1V��aY3�Ԏ��~�5�����/f���Z,:�y���p�e�\3��0J�tn��d^E��К�_�\��ף���"=X����^t����u K��(Q`&��� ����&�B��5ZqZ�Ҫ�̶�<��m�_)��ۍ���CI=d�R�2Q|n���Nq�ry)0�`(��Y��=`� �Y��A�.���"'�C���L�j��X�s���/��G����o� �t^���J?ڔ�V��gIf��(��.64��Q����-�����F}}5��3]�=q)lo!wn���i`�����Nz��4�I��ƴ�ٛ%�2Q�qn�B�	�	�G�#z�g#��������a#J%�*yD}Y5�W:���%��;����:�O�*8�s!Y�hIs��sջW�M���xp(�lD �|d��h2���a��B����N�O�T��R}o�Y�SY�?�b���j;?d�{�-q�d�79�,D��9�D/G���M����OiF�퇬@���.w�ϭt��!�Hݐ��ړ���}�7������8��s4s�[�!����s��|t�	X쎢ɴn��98��3��B�p�D�rRz���(ԕ����3����d]����1������7	�t�}��__q�9�cRt�M!�����_̊����W��^,c}�DԪ�,�S�i�N�� 7Q�?�u��O�� �N���J%�n�,>������!6n^|�S$�T���8D[�Y��V�5�2�CZ���Z�v"�H�<6��F��+S��f�x��]���4{�^&��<�oQ:-�������:��l�F+����찄�ĥ���2����A��#��[+��V��;�
7�Fѓ1�Cn�w6��2�Ero�mj�<��c��)�z5�Y:7^��mjg�d�>�5&̵�M�Rp./R��j�g�oJ\U*6��p���tQ1cV�2���E��7G���������e0Ί��r�c�2>�sg�z>�+�V�m�Z�����Yk���-��/d+���F�(���k��8���LMd�@��.����_�͈lteo�jо��������%!��n?D�	�&���CKG�c�8�JX��ط�o��s�p�ٖ���:p1�qy6��>!Զ�%Oo��3Z2$�tӫ�E���F�޽KWv�k�p�Sz!�� �^�(H�>�f�N��DKq@ŀr��Q��U��o:�W�\3+m4�}���x��y��S�,�䇈a�p�PJ`��8b�1���t�qQز��,itldu�G�I�dic�s!`�Ø�L.a#ޗ��Br4�@��Q�F֥~��~G>�"��Q�y�&F�s�BhZ\GE��ĨHj�}a������?��bvABef0u\^0:@�S��E߉80J]��{'��Vg�,#�-:S#>��Eʲ�(���]�B����n��wAm��8ui�y����>t#�o�4]�Ԕ�:��<�C�1���5�%�8׍6g��x��4���AsmMF��aJ�"yɴaڷ
:u/�;���B�&	��i��zI�>4��pu��H?T�2��Ybԧ[��#�XR

�Kg�@�G�s͚o��l۴05*��/*�)���Ud/��T��D����j>/�hr0�ģ17�k�H跐����K_#I��r;��!m�q��/-R9��z��kܳ"�,H�����M�#z�߬".���O�!��	�4��P�J<S���w��3�$��C�w�0~�2��'`���>?�_����j���yĝ� Φ#��>�����rw���v�b-hE=�s��K�L٢s��_b��+k'n���G'�J�JN0��NܫY�kOsX͝A�#+�%�7�W�K)5���	O?
S��Ҫa�����{MO��`j�+GO�$�;�b��nUf�,����_�������D�t>�*I���Z��-�4�	�aƕ�j��Ӥ*�>����'�m�f�㬊-�b L۰cT ��'~���Ԗ���j�Ba��EÞ���1���Κ��P�q�� �+�b	c0�^P]ۅ)��z֘6�勉Ǻ�O6��5�{z>��bOj��t�����ku��do�����>�K)�+_UW!QM��@��
���ȱ�?J�U��7{nSB�}�7�D\���8T�x��Oc�����{QA��8p-)5���`U&A+ M�϶����l��c(Pkf�)�έ�����یǑJ��Z�$����^��˭���u�f%�ͷ�!�G:'=�#��k��l?�H�[�s$�f���r%��Mq�6��$(�U������N^���8����|d j�ԗX�_�/�Q�d��aT��:L앇�gɐ��c�:�S�dL6/0��˺�2�jLl�9^)n�J�o��h������dz����@c*�y��T�39�yp����pk�����d�<�Y��Y��h��O�N>J��)�&Hӂ(Lf[��=m��� ;.�?Y"�y�m��C�j?�P�M�G<n��6�Y�C�J�{������~>�(�� ~�D��9AN�p�Ͼ3V ��v�(�U���뚠DK��JQ�t.־������;i�&�m��.5�����bW��(�~���J��g�� ��_V\#OH?�#�3�}7��
��Ge�HX�1C�5{���*�aq��О����dM@�-�!��9ͪ��93Z�{
�m����v���ʁ5:�ҽF�����>P�~�R��< w	jp�e�{$�-+sp���^=�����R����A�<�eR �5q����� �^����6�,�,F;5���5���e�=���K������I,�9򴙾g�Fe*[�R����Xҕ�yu���V �|tw=���.H큽��qZ�?�(Hbί���/�K��)����E�5�C��v��ԞW�&	cSlΪ�Y�.�N�n�@���gN���Q�_�:sC�7��:�@�ſkN��:��Y��U�4���C�S�%��վ���+�G�<�k�9w��V���?~N��do1:��D��5�5.�O&���L�	{����̯������