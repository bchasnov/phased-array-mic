��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>,M�Kߤ��S��#f�0q ��aUO�ѷ������\�i� 9����ۼ�KuUΨ�r?��Um+��4�g�a�	��TC��"�
��@)�$�Ϩ�)R��Qۺ���F�z��kf�?���CL-˧`y���~w�b:�m����(;=�n�����������R��칤Lx��A�^��	�]���0i�&V��7�����w��9nήHu��f$���q蒈Fa�E�jsKꀻl��	�-���T�o��${#�6�V���KY�An������$a}����7C�K�:>v��"� �bWwx<2�#²m������7a�D{�`� ���v���:��.�����B��[E�n 햧���E�'���(�lB1yEj�C�"�P�k�=����[�GT��a�P�����n����U=�����؉G��@�+�%F����ct�i��N�~U�)�)��<�$BJ�у��UA�1����4;ݪ���:93��s�E��qV��8����9���qȝJ��T%��T�<�
Qr�5�q�&խ�Ͼ�ʽ6��g͋u�UA(mZ�oڮ���U��MU��2���4�8�xd��E��a�7��REDT�?�h�}�آ�S|ؐ�Z{m*�$��Ƕ�e��|�p��,E��S����?[)6ߝ�3){�o����2�x����0oڙ��;��4�����2�ի'��.s���9��K����<65�[�����{�й?8v>��T$0h���ܦ���T������v:����N�%���'��NuR�+ۨ6&N~�u*b,�An|�8�.\1xHXUc���K�����r\��c�Ǥ�h�j�a��VYU->��fLP���^o�;Z��eWF�U���R��4����<|�Ձ�-��$��iMC8*g?������nþw �S�M�A�� �"�wen��	\��F#=������%S���+�>�8
�YJ������j�A�0�(�����~�T-wc��zJ�R�|K�4%,%��d����GX'?m�#�]����<��.+ǉC�y�ǈ�P1ِ�#�u����iRʶ�f�?� (d�)"�&��kx5g���S
@�B���+0�8aϘф�9ö��
��c3�O�4�������A�{�6ط�����8�v����W���5𾦐x ��0Z;���[�yR�e[���#6����8iX����%��c�2��󐃉W����Ő `��8լ ����#�z�4�x3��xsP��.���(n�\!�<S��[�J�5Yc�O*"+(�Z����g��ik;4����X�P�~K�U=���$X�¯+������!�"�{���}���"�>گT��T_��	���\�3��㏖(2tJ.�b�/N�(R�2��L8��6W�Ǝ�]).��VL�/x��@��[�=�}|�����P�b�ڼ�s���9�#(�����t�v��x��ڙ��I`�z1^@;�&��9�ǡ֫9�d���\����G������#����"�i��hK�G)��lj��{�$�Dׂ�t�[f��D���>�)�Ռ�>Q_�4���r5ꗻ��^�F�e�8 Ke�?�FX����ݦ�goZA8�w��C�MZz���5-��[�J���S�H��v�>ih�>ma6�������d�CTe�$0p_�z+1�ϝ��#�I�,(�c>A�Z���;��`�]�>�P@��n����8la�K ���Ȳ�vW��#��y����p��1�Am���=8q�Q���m���(6�3aF��l��a���ʺ��9��[�a��^[�V&6��k9Hr���`�}6/�
b���f@]x�r�T�2z���{:�F�/�
Vm.ׂK�cl��N��������hv>!�{� �&�US�|J���1/���L�D+	�ZPw��;AD��Q��AR�)^��	�P��[ϓ���5�jSe}�����W���;4t�`����46✧���6���	QS�+;i���E���K�F�����o���tG����ګ���"�7�'�]D��4��r\�O�D��'�Q�Mm���Xl�8�/E%�"ܚ/�K{���q���{�:�A��SVy�����R#��,�����������6�;K*�"�N;"�"#j��؂&YL����d��oz!���E�@;�λ>�(��ꈺ�Ϩ�F�j_�'f�š1��$r�ZN�k0r�ǋ/6ќ�H�����*�Zs��>�*�vk2ue+�x�!(����ފ�b�i�q�~/��dB�uQ�S�g��:t�@�gw�޼���o|��\Ô\J{ ��[zخn�Yy�u�ج:.A�� ̇WK3|�c%��<$��f�Oq����6���b�KS�Á[���T�����m�rs�>�_F���~���*;'��`��x�����lOR��u�^�5��n��jqXݔI9�\���"�����u��H��*k��e��Ze�X\�b�@����,^�%�I�p�T�N��6�J�\��n��.	���M#v�B_xe��zz��a�t�X<sT���jz��&%
�q���|��?������� ��>"���̀WT򦺳�%�OL�����/]Sr��)��R�N}?�/qc�%=q�ic�f�{�GQ��焞�CRÿ��ﻩ�d�E�[^��c�FRk���]���G8<��	F��l(is�ł�;�(B�P��h��5���,Ӧ�L.��|��;*�|<�[i��jR���E��L[�@ߺ�ʭW��ǛOMBέ�?u�#`�4;����M��}�R1Q�g��o��_Z		:�����,J��Ovq�f:�_��)��䷀��9���30�}ͺ�h;��e�o�<�}Aޘ�I��f\H��Sa�����zL̵�z���8ٿ��� �uāZ~�Gq��TY�˳W	7/!���K�?��X?�C�����Wk%��5�;���Ĉ	�:���sKiH��(����/=��!7�
=ر ��gO�׬B�O'��$F�7��|�h=���>��]E2:���|cS�{k�j�Pfn�t�
�(+���h��d�J^͇c;��.fڝ��5Y)�Y�Mj$��Ǚ	%�TҲ7*��8�"�X���j�K-������rɞ*�����9zP웵���
�˳�U�\Of��]�/� �8ۿMe�R#W8r������f�n
{/S('�A�V���n�i��w��:�S��
�R��S�<��#`ct�6M�\�·��v��Naķ�
�JQE��U��Y�a�l�é󮞵P:H�%�<kۧc�}�����~��)96��"�a�N�/Vj*�`�h�Mz�2�!9z�#�Ȓ�=���5�G�� �&�֙���}��J�5��9�9�;�O1�t�`2>"q�l8�t�~p����֭�w]�����k�1l��^����qf��y���#���5!�FK\1q��ו7�O��_�-��R1[50ʣ����dZ����hO̠ó�~'W�G�i���:������Rj=���ƷW�r-vMP���73��^�sn3�m|��u�:��}��
�fگZ�q>��dɦ�/7��
�R	��>Zz�S㼕��U�7°{$�2�xQB�J��%
�ν�9C f3���8�v������HM��e��#�teT�M�V�DΎ�r�?H�\l�m/��7�3ٮLWJ{�W�:��|�����`x#1Dj�7�T/�Y�����e�!����f�YO�Kf��ț��}#�}�v;�@O��&��ar ;�x膞����oj�2��s����K�~\�t~Ff7�5m����LM)5� ��ʟK�N��<�S�-|2!��sn'�v�F����cbz�n�ik��1�vԺ�B�:�af<��2�L)�<Bsm<i�f1��u}X�Zx����G����j0
�oylȤ�C�2�li�l5+�&�1�R�Mܠ�$3�ڧ����m��p��;͚�W��=��|��`���YB�k���9sńJ�J~~� F��{�д�b:A�c��|�Խ��A6�Hw�LG��3����7����6���k��T�5[�TK�\U"�B�7{��.Z�� �B�{�?�+E���(Hx䀰1 �i�3���
�:��}:>����wg�*�(;d$.����$�R#i�+hT��������Ҩ/�hd��f9@��W��:������O�W�@v-Q�<^g.���v�a�G��&[�P�<T�m9����������9���t��a���}^z�u��[�8ܿ]r7SmZ��5QT�<��3r�?6�E���v��U+�z�w��qJ1+�e��|�{	����۩��#��|����ι�wuBs�DH�z�dwx����TJ��K��|{�r�ٽ�'�gZF�b�7w�R_��v�a-G�dW-��'�ʹϊ?V�U�5<౦68y*^"=�
�=+���T�N����l���3k>�N����9]n�^�e�Mr6e���H&��1��E{s��s�N�c��FZ	��� )<��V�Hǜ�sEX�y|��� A�Iϕ��節}��&-p�r^BQz���%$��:o�a���.]�+�E����q݄����:��n�C}����dw�Q+�<;g�d��umk�����phM<�N�B.4T�8��,��:���L�VX��X]�b�v����:��s_gnF}m<�k7��=`=�56�BC-DV��bW����"P�0gb�86?%�������*������;Tr�x"WC��O�em5 q\�(bXa" �D�n�LMO6s��{�i����N���o��r]��jD�JK�Y�س��y��b��Rګ�,dߨ}��U�O��LF��7"n3��.��H�Na-"�ho*���M���#��H��c��U~�� ҎB�׮�+Y��
zvsƨ�a?�k	:ױ��kw��x��@gMO���͵���"/��ƿ%��(��#C�9r�w��{���-�K����a}FL�lI��j4��tP��XY�<06�L��ʎ������mk��������HD�DB
D�;���D���E��kl�2��F8�i'.Ph�<a��X~I/���D���ᷠpq���k�V����$���G�����4�*}�[��G�����)SƤc⵱�ͨ�#�r���b�eMߟw��t�'�-k[e.��Ɉ�qR�9�%�PS��E��~&�I��ތ�i�P�hP�S= ���� ?� �W��;?��|�����m�|*�g�����})j�<<NA��nO��`
���v_������1yb[�ӈ���ܾ+]E�*� B9���O��t��|u;h/�yk��Mr��f�CP�w�D��G�V����-_�/�?w�/���	lݾX:c�يK�@�'�[���]��O_��l�/�|����aA�B�?T4�#�㾍��&�t�Hzэ�1�R6
����;�v"���2$��p����n`�-��������:j�OZ��"����yA���t ~���(O2���_%f]���yg�cd�뜑=l�LnL�6��a��/�y-{��Q�� �Qjq����E�'L�}��6�ET�\���a�v:6�����k�kŠ�*_�����.��6ۅ���y�dD��fI�q����74k7��̟���M�`Au���|�=V�㮒�A�`���P܎L�s~�s�����Ƙ���z�Eo%��d$±|�8�\0��-�0�J$I�'����rn�d��ݴW^E�q��l�5���_��~��ڡ?��\��3�����˪t\�%��Z�������h#ߟ���1>����D��F���6�<����]�7��sR�W'U��& \����V,?%+��'N�c�CX?-�Z02>�┭�ߧ�`Q����X�_˨�@�H#�m4��C�����R%���REhwlJ��|�M����)<��qMPںHX��N�!�)M�O���T@��F�s0P/N�cǊ̩�B���o��D�ۖ1<�۫�an�m�S�rt�P��Rf�H����k���>�N�5%�à�W�$��67�Bc�H�s���F�h����a�HX�}&n<@�ʃy�������
Ҟ��y{(�v4l�3#�2%�5���#M[�i��W�er���4b#R�G?�ڑ�k�_�@�ޘ������a��F㑛]�`┘J�/a��_��q��H~ߌ�4_���C��U�$fw�P~dc��WGEDD�Q8}9����t��qg�L�ſ��%�&���0%��{z�m�bD� .����7cF�,q<>����R�q��0�T��ڄЃ�awTP�`��Ǒ��A�3`0��M�69%\��wa������@��Jȼgl� ���a���d�.+�YC��~������B��^M���WR8��9sGA�T���^�.�|��Dz{G���gcy�d���ͽf���g�^��@iyu`�; ��s���/x��NL��~����5(���`J�}Խ�Q�� z�_4��7����� �u��mr�����d�[1�8|z!
ˀ�~�G09�P?�ULF�邇�����N8��9f�c�P���j��u�4�
�Fu:��)�x�"���&�a�PZ��gb�|�gH�ޣ�e#a�Y,��&�������Q<�-$��`
��G��iG]s@n�A#rr�;���_e]�S/���F�%��Er�l��c�F��Mن��݅�Ű]�����ڶ��#�@u�΀�������_�]�Ŷ*I=�F4� ��6�Hz������i�>�0�QCd���.�y�H���h&�}��&�jk	��p��=bհVJ4y2[TZ��@�rL�U��j���8~����vb�pC�H�UCඅ�i<�c�5
�4Q�������kxב�����=9*���za̐��1��߃��6�	ʾS��[s�&-V��ʝ�RM����������l����y�Ӿ��w��{c~�5�6����n�,�@Q���J!�ܘ�3Yu�`�lS3V�Z�����A[�'\y��i$eh��X]����x1'�g��A�+��&6d�g�,�/�s��rk��u:�=3\~v.j��6�ζ��#�z�����TK�7�4�N�=��k��R$v�_@����j��71�K+���	Z�qz�0E���_�Q�$�^��K��W����cp�fA3�,��0�x�R`�����_�c��a��!�Yj��������F��Ϡ�~	?��/U��0D��2�ݿY�$3P�Ɉ�V��Z�P*�x��Uur�:aǊ����'����J�4A���������
�aB ����j�F��9�0�' "ɀS%ل; �� }X��td�Pĕxn�ٹ��Sg���i��9"�X����Ǫ
N������ ���V6����dF;L�F��Y=�]�T"�	E���{E�֣�"�Q]�j,�|&�f�I�h��xu�A��~�jnP�z	����o�͢IL����G�Դ� ��z�
ݦ�����s�*�R����%�	� �-<�1���-�ò�[��q¢݀+� �C���������N	��[�*�77A>���	��%C9��I[����jW�p\!�K��R�c0��mlLJ�����-��,�GҰLu,�)� a��CW��wc���E]�f(kِ :02������}B
���E��K\��F�]&��;)���2w���@���D�c�Ѥ.�FM&8�[��3���l��N�cL�e$1U�e��L ���+L�2�,�2��Wq]���N6��es�\`�c�����m����k�`��ҕt,�*���h�çZ���ǫ��_���:@���;��+92����ƒau�5S����VL�0%J�{�@ ��T�k+�?PT���ޣ�Ԟ5l�?�v�n�m���VqD���H�d ���QC5k�y�b3�i��LjF�Pň�O��,��`��{(3��s���Vl_۫q����j�������ĀI�2�����E%yX�������)W�d��nNJ=vVO�����BMo`x�)��� 4���
�^s^����$�HX���������9��)�kԱR�3Ҹ�Š���;���s�/W�Z�|��_�o���E�A��:��qwJ�@�a����%l�&T�o��S�c�\��U$ꍱA����T������V��lO(C���j���e*��ư���U�����I��iU��Y�����gp��Y
� 䦫͑�w߯��$3g�C�wͮV����[�f/a����9����8�������7�(�I��{z �!�Z��b��z~i�y�)J=H�r�W�� {�c9�O�.��e�ݹ��8��^��tM"@�za7Cd��l������H��)D�3a��kd֔^��=���u���;�Zށ$<A(e3����P��w�1`O��c=ź��f|كE'��a)�ze7�FީK:�l�^jbK����K�}�����7����7��1C��
�4�eEEޙ�_p��Z����`6�C�I0��s��Wfed@(��S�����g!���,\uQ�)��]2H��-��
c_	��Bd�>����z�s��ch�$�V ����3|�Ά��Z6b�\SyG\��`��oę4�<=?k���Xn\�g)?���z�u���ϒ�
�SrxM%�g|�&ü�b�� @�UuہQ�	֣)��" ԥ%f7�>90��LJ�<^
1<�k� j�i~R^��!9e܉�XI��p��Gm}G�=x�X�\T,���99/�#Ս��겢��xY��2�(�U�=;���I�mGzo>iY�d3�w�EC�������~��B�L�
�8̾3��zCoX��՛�%iY����A�6��|ܙ;v̒���JAI��Z�~�W8����)ӈؙ\�o8���zj��s��w�E��������I�?��XR��5y�����Y�r���-����>�a��6�#�����Y��;��6h�.���G�X�Z�5�b��n���ϟ��CbQ�v�	�i�yd�	׆R�Y�aD_�B"��y/�N��1X��
����X�E�r���tF��}�U�ӫ~��_�V�5�|R���u�X�E"�7)�7+�I�7�W���z���ΥM���h�r��^��5(����q�Ջ,� �MV�	�,m��6�-��$�X��b�����Q���<yCj<�%�Pzі[��[9�]/���U�ɫɭ�F�t�,���O��W��`�^��\��jC&G��ŉy6^��9	�� d*8�)�6��gj���ߍ�:�ȏQ&�θ�N���'���u,�v�s�3+�0PRu��G�fE+Y� �cVo��10�'ǛǘL9\V�J�U��!�Ӏ�5@�T��htp�3�:X߁�gG��Ù�x277��|���[�*��ed7����-V YM�x+3�m8�c����D|g�ZƳ��B�K'���.%M�@��{�k����V��/;z�/X��qgv�PZش��,v8�4��j��Ư���Ynto�>�I�����_;n�ӯ�$�T6�Md��Ժ:K�f�Ԋ�H�c��qYd��*��fT1��!1O"��	rCQA�T�~��� q;����H�-㦖�E�n�aj*4��N�o ��	H���F�y�}��%�hwz����D�7���ih�9�T��/�-�$��R$1�-�
���L������%����ŕ"6N�S�"p��*�֝�m��p��q�t^6$:% �[�� HE $���'q9�B��{K
N�n%Ĕ�̙��D�|�KS���*��,SaM��>Mmh3�ߒ��}���������F�dx�:��$�`���=��9�՘�l��<�w
<�q���#��)#jրd�[4ev��R��1�ZP�A2�0�"����)2������;^�pb�9��I'8�-�����!a	�F�N�L�E�f��'�oM���N9Z���h��_E���к��-d6C` ���9��"���2����b\UE�/D�X�|��Z��jr�N?�:�Z��8��,�Y�ts9XgҢs�C�<`���^���?�r����RP"��x������f	?�����_|0��NG�����~�"}�R��IN.	�WA@���{�R�R%r����N9��f]�����)Q�
'����=�r��Y��,�&�kw��l�#S��%�D0����p�2G����\hg\&�v�#�t���ߡ�y�>�/Zf���;o�iTI� ��ͯ��I���~(xK�"o�47FA�e�"֎��#���e�&�S�-^�u���ɞ��wƥ�j�b����mrB���F��^
��"wQf6R4E~�\@ �9�_���kA6�ݏ^4�F�!��³�\s�PH�|ky��&���X���?Q�H����S��>��X8{�7���7�_L���������d����Lk�:�:a"���i�	��闹'�,S�u�j8J�<���z�����F�D�n**Ln��l���A�N��Q���!S<h3ҩq<(�4�r��O��'��í!WQ*��)x���Li�,��n�MX/*�!D�_��g%K���z��Y{ӓ�����5l�R��6Hۢt,y�������\۪�wh�M��pc�k� �U��@�T�4P�6��0a��|9m0�y��*�J,��d��L����\Iħuѩ�5�j��рE�,��i$)�5��,�3����>����m���
2���ȏ��Y�'��Chs?n����Q��p����!�ri���!�|֛ �
>f�n��πOr�]9��K���|��!���E��/O��}W1 5��i�y�"nc�)NI�;��r����l��?�q�X��[l�6/lfV������Tr����!�A��@���w�M�CK�jѫ×3q,5'4X[�c
`fn���'7Ƚ�^�d�\��db;�q�+��^-��Ҩ�f>7Z��D��ȗ6K��\�����*�*��=q���=�/��O��K��|	EY�Ev'��~���%�TdUX8�bO���O6���۲_^�F�G�H/qU�M�D�GT�{X�޼����0�q	���:�[*k�0<R�k�e����ɠ�����B