��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>�m��`K���`"^	6:�����-',�{�>� <�pQ�Zw̓�e+���E��W�6��Q���c��p|C�Pֶ���rA��B�Hk�>yA�
f�AL����cP�nM�׆�*�ˡ��?N ����ሾ���5����5D����;����7�7?��	T��MNL���/����aw1���O�L�Ȭ�7��5�b�G�U�G��zOw���?uGnۑ�^!J�\{�l�������Դx��e@ϞQ�
�������T��ܳ
�XP۽mԊk������N�J�zO��P�\��LLG��4���>�Lf9��Y�&��V�/���65ӫ����N����˵$�Tδ�3V~èn|�u�86��3��y�x�.ܚG�=�����X�B!VW�8č����Ȳ3Z>�	W��6�oG �l�84+�+�EߒF4��#�;n3ưT1���)-4��%�--Q�������aif�	���4��h�G1�9�}$*�����j#�B����	�4��@4R��'��)khlsDh�.��9Kk�Fk`r
�����bD�bJY���{O���47Ϩn�&��/N|N# ��r袴��&6�L��O������Iā]��P���A�)1.�[�1^����Ŕeɨ�ڂ]I[�˼_�o�$hCFx��̪+p*�2����P�(u��NY]B���>%�7dLEg��2�劻�����m��O�5P�ڒtIXX2�㑿d�\%�5����g�4�\5Ϛcq! �2�N�Hly[ԕ�BNw�3���m4U���u=�J��7]aW�0�3��\ �?�b��6|�w�)�&�94�єQ�T�������]��V⚜�*"��pjO,�{� "�}e_R��5���]��<47ќ���a_�'Q1�;8��>M����v�J[�+�l)&�aF��z��4�i�0��W��p���#���ڝ����ӛ]�������|~_gQ���H�]$K�d�KYZ�թkvm��nvD8� %���*�^�F�o����(��-�Z�]3��y�F�bV>�QpŞV=e>�N�!�9
s�7Н�ReIɩ�Z��r׏cG�� <�5�cF{���΂�(R,�n=t㠱4(�Ck�ƶ��v&�rT���P�f��F9�6x�{�iv9l����_@��}�9pW��gP��_EeKCM��PFl�8� �\w��h�jwT�&�bڍi�䄏|\$&φ���O��Xݑ�U�Z�����c�O�9��鼔g�"���7�}���[��;�-n���B'����֬�c���2ң�/(�Х�/d�Y~���Ѿ^���EAaM:�2(Ș��GZ�ً1"^��1�mIG�����Y�<�\_� �o�&�YLK�hf߽e���}�,�N�R*U�m���o)k�a7��}�4��bQ՛s"Zj1�(nIn����ĚF���3��ۆ�T]њ�Xt۠��(�<?��uh�p.���1?�-��t^��\b.nN���nڠ�Y��A��7�-�|h��僨N�C7>cC�'Fe����~���_�g�G^\�'w"���B���3}� �c�k`l�~��J�mBԣ.������6�/77����>��7�(�}�f�3��ܴ<��
�� �[x�X?h8��I/���Ƚ>�inX�_c]�T: �뾫��d�XZ������,�n����Zp�"�5�e�f�m��@�q �����rw��ّl?����A hIG��u�=[��=̹�Fq������V�x��B~��"�:��������I��8}���`��3'(�4��!��x���h�>��5�-�ت�������_\?|���AX�=ˊ4n����p�:uWW(:q#4׵��=�o�K��L⅘l�������X,m	t�ѹ��a�r+Un���G�� +�"�](�^�i��d9�4�`!�M���1W&f{qu�u�������MJjrP\���c[S]Z�`�����[�x^�,",���J�r>bˈJ��zΠ�73INJ��.���S���<�l��N���nE4b���D��}
�YS�e���++E^��n�I�u0ǘ�!�1Rj�o\
��겻A�Ȗ�r.�_�, �h�o�(��ț���/�_�&ٳL���"y����=HK����c�c�=;��<xE[=ViO3����m��R�|��7O@�Iu��.���s�v�$t�3J����{�I�BU���P�X��ܷi`�ܬ��ڋ�p~h8 TQ���wޢ�����Q�6b�O��c���\�u�?iGz��4��o�@��c-�t��,�kM�JꛑU��k��r�1Z3�Z�\F혏����� �t�3��@����k#Ӯ�N��T�\G�a.��R�ǰ�<5)P�U<0��]��0��hV@eQ��>�
ݝ�n߄r:�Lh��3� �S4�q�����e�9����m� Զ��Z����7!��/ʍ���M�}�z�/�:elVևS٭g�nt��j#T�P;[rI�0:���y\*��f2�s.��"�'E��5�[�k�-�R���5�W��2�I�;|�X8fG�5��Kw�x��}���L;I�fR��,M]���'�����e!@����7�h_Z7	��6z��`H��4VZ4>�Ȓ��$�:�nb��[ K����t�@�$�}�{������&9ނ����J�e�*���"P�PҚ����V�]��I|n§�W��4r?�H��N���.���Q*Na�R1�-9z����T����(��d�ߣi=��&�v�bp�e���d߲O�P�>a��>�0�����&*�V��7J�3ZY��5L��������3��+w�Vi?��Xt5U����zDc����@	�k�Γ�p"t�l�>O�L@�ܝ�\ FB[��:
z�X5��-�3x����D��z��������ի7���_٭�Q�SzA,_�:! �&g�}�:����&��[0�ĕN�^PR��F �ؒ�8^�5� U��Q� &8���_+�	���?K��$�$���$S��	���� Ch:�A��^�@)��~����p����Z��K&q�g�^��^M,e%n�S�ђ��'O"χ�q�u_�+�WR�i�O����3+J����޵�1��p��3������K��׵��jŮ!񄴺&Lq֎p�삟�"�U����.9CoK�)F#e��۲qx}�Pr��(��x���/�^$�SKa��o��A�c ����� ��,���@�]�ݯw����� �D�
����A�H�lX��D�5�qP񪔠O��XP�o!�
�b"�N9�+���N�3�9!0����m��W�<�W�b;Q��