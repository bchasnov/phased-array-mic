��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�]��Xȭ��p�oȡ�;u0ީ�^�)�>vys���2{�L�~|c_Iy�K����-��9!��\�Bi�D��{�Ԣ��r'T��NjH��ဣ]��9��|p���4d��oc���_LG����*k����۾�T>x�/>:��e�=�C5!)f���86�$����ԤE���oZ�&�x���� ]1����V'���Hci������I���-�;����{�gr�HR�l�q����~�n�2�����̴S�c�6�'o����f�?L�2���r�����uq/�Z��a['R�)9"+",��:�l/
����#���U\3�$π��`3��J�,�;K��=.�ʄ1���c��ą�&Y+[&��z{��/j��?|��~:�%��?�!M1�3?ߤ�	d���j"VlVg8��j&84)�|K�\�Y��m���TU-�^V <h�Τ�4XU�/6�����X�_A����W!��i��o��>��B��.��9C��iżׇ�2�%>+o��q�(t�
�%�\����·�*,U��y�oxmX S�`���;�F�S7�
�(���!�e�5�I��Ey·���e�`
&NTv��n�������Րae�m�d�9�<]����kw/��׼3`����ǧ=��ό����d%;�4�����"?E����R�m%���<�:F�Z�䕼jp�j7���P�U����AX�����:;��}1I>�[Z�洽��J�(T��(A���ik�sO����al�	�y�7�Ady�3� Ck�ѐ�9���#O�XM��@ŏ��X@���6�-i�� �*D�ӆZ-sa)K�7�
�3�`8�"\��u������Axw|*�>�y�Z��eDJ��rs�?���P�ι��Q \�f�Q)hQ�&��c�'��n.l�.'I�X	�D)!���s_��@U[%�Q�A���"��L��֢��۾����KJϽ�U ��T�/�f�MYA�����������=��D����e��|E��T��_%�����̸;�[�T�J������i���~��9׾$T�r�j?źR�o��*��C.�������uׇ<V�6�ĳ��Č�z<\�^?�����h�%X7�mp�Y^}Oa�V���_�L��������|fMX���M�T�B>�W�~l���2�<#�dd�9�Lѭ��19d��gTlCz<Lm4n�LV�.�m��7�I��|rO�Ӌ����ȓe��I�'�%�S�wO���b#�՚/�H����Q	��c��.6x�'���OP��G�;�	���)IDd#�1l#<0���I��y�Inw�"[�r]S�<�<��d2z7��RM� !+�Z���E��Y��V2z�f����v����LT��� �Qd`T��{�H��l��1wV��\Fd%R�zjw��[�	�y!/)���Cc��pI��C�����'5�����R?S<�����+�Ѹ1���s�����ؑl�8ڙ���c�!�����J���g�I���� ̏�]���%�xb��.;�a<��o*���a�f���V������X�p	qB��҅I����Qd��9U�񄅬����o|��+����'�#\OPB"��&w0�L�ڷI�U�?=�PUv,]Y)E�f�R�g8��`�ߪ�Y�M2+�̸W�a�V*k^^�^sm�=U��k��`o`��@���늲����B�7e7���x�S�/�(�$@j�o�(o^%)�j�j3Y���`����[�'�/���'4��Pe #Y�*V����(���N�s�C��XE��QI��rZ��L�1��]Bl�j%���q�����������A��<����@�x���-ɴ�f�`��}۾����&I]��D�IU�����}�s	�c1��+�f��"`�Hj���eg��f� .��3{Q����?3\ːT�'����sd1u��pt ��'�I�/;+(��-�&���у�m��;����������]��7D+�LG���Ϣ�߸�.�O��2�tT)_q=�<'k>�]�:M�+��A������UY�|����Z.h�<��O�.�_���%Y� L�����MS������L��)�b|z{�L0��T�l��s������VF�2N��.�7@1�
�R/7�-�s2൨�P�鐢���Ub�z"$EYb^�~��+�K�ԁv��Ǒm��5���6`(�l�$k�{Wj����v�?��_��8%%���K��&����,��{.$�/���t�#�t�9V.��p+3�għI'�|�6���0�\{����iԅ�T�ە������-gm�n���}|l�%��B^{�r�u�&��h�D]gD\���-w���/�e��$F� ���W"ГZ�N��Aw�+�=��%~�Wp����b ��a��e�����*�r�6�i��k=��ǤP]�<���g�e�L�>|����b��!����� >��Dl�.���� P�]����b�B��㰨k2��޻m��r���D�*�f��G��8|�Ì��~�Xݥ)��07K{�9+��ޛ��WkE�3h�\b�ԥ���U�����"�2<w���1�֯B;����=�͂�$������n>� R����\�_h�2�fN:n��ϨeܲjP����S���UId*yO�ɠ�G�~X��
<=]�e���*���a������k
�Zmәt��z>1vH�	��0��H���ݠ)���T��R�!W��0e�jX|�"�^������)� w̑~ᚑ�Y*��/�d@8�q��E� ʗ����??���ģ�a� ,�����⎩;I�����PS��@0�09��E��!E�a��h�Bț�u�4
�X��l�u4`?ryd���nܖ{�'
n}�	��&���v�'o>�1�;���t�����E����m#7t�G6Z���b<�<��=�Iޒs#w ����P��ӜMR�Ú��֩�m\7�������$r�6�;�|��AB�Ü8�pr�����f"ak3�ph��M�3!�����~סş�;b��¦�x���J��?:L�@E����z�jƨ�c46��xn���PţxCQ��כ�V�� q��Y�^�q�/�O�JC�f����+��Hk�A2{D����ڸ4��:+`�pp1�Z���N!���n/}P^��b��q3�'2�E���R1�Bԍ]�R��9L��sf��.� HC��Gq�)��4��^TN�p���؝���O/�׮݄n{��=��s�t�>���o4�7{�h��ᛞR�� �'L0��B��d��r� �d�ᐷ_���!25�X�Z����j�(ۊ�
��e!0��"��
`_L����6��\TeX�!�a`��"$���B�,t��NX*X��<G��緂�
i�$����m̟Aq��4#[AJ�ܥ�PB��2���I��c��=�LV����p�$ ����i�X	[/X���I4s���Ha'R��࢝2�GЋ�>�-���D�6$�Į�����m9S)�u���v�DK*��X� ��f/���U����qF�_�ҨB�E�~MQvn�z�}P�t��m��*І�ɣ���ME��HD��r?l�)ǟ;�AH���u��i�ё��}F�Oɠ!,yg�P����Ɂ��������%�=��F}��/���9��%�ӆ�Ծz��%2n�7@KUi�!,�$O�A)�����UjGw�Db�ө���у����3�8C�C�}�N��j{�Z��3L���=�5�l�bw��s_��/~05�� ��T����UE5v��WH_3yUk��i�,e��G��6���N���������nb���\��|Bi�{�v�M��<������l�JsYE��A���2���qI���m0�ҏ��{$,��u��o�j��lE-�|��.���E�2nb[V�D��u2����t;������A}NG��Y[�q��Ia�ח$�oM�t�~�=r��1O���cu5~��:�%��x���+3�����.����h������'-�=:d����A�f��E3t�H5mx�
!�A���Nn�'�UF���(��S6N�~����׬s=��scn_2��l�Q�"6�xِ�Lāh��s2/��a�c�|��f�(��	�b��4� �ڣ�s�U��vm�R�y�r�D]��	�V��	�v8iteO��%n�%to�69ܻ�s�6x��������$��8ݻɞ�ͭF�>��W��ۀb��v5Bk���:/�m��G7ʆr�W���Լ���e���ܩ���6mA��˩��U���h��A3������oj����'��ē���c5� \W�^D����������%t�
b�E^*��_ۍM:BK�_H��K���jY����>D��{Yp��"w�l�fղ>g�}Yq+�Pw/����)=3@3�m��6�A(��OB�^�����6���R��� =6?g���iy�-��$K��ƑS�_o�*}����1��I���r�ߥg�>�H��`�i�N�#1C%R(d��2�7u%�3G"�8��d��V" i4��Qųb�-#��1�8�b������D[�Yź�t��%�;Nm
g Q��(A[��7��e?�����'�4�����}��|;�:�VOD ��b`DOeu�]0��}z�`��/i)t�#��Y�;���	:��E'GX$|)�^�W�����\�vC�&D�o���嵘�����C����G��q�P�Lu���6�%5���4J��qʞ������`Ԃ�D�g�~�b�q�>������.-sB�� ٠�	����flO@WL�C�`��.W�JX������l�����{������─0���O ��H;p֫Rv���1^j�o�n��$d%�wSz=T+�p��?x��J)or�<��N\�N�n�o��� /�������:�^�w�45��D���˷���;v�7up�(���O4ųSU�ͿG8]�,[L���}�`O:�M��:)0�3?��5�<_��ݬ'3O_O�`��)����Ay�Uְ��K���8Bك�>����<�v�49>Ц#aГ\&Tb����c�����;�cV/o�M�[8�ƒ*GP�/��ީ�zG��A�◼�	��W�|�h%ݩ��ĖP�,
H!��E~�6�=$�|����x7CV��Y���P�y��I(T�9s��O`8�K�Y)XɉR���ϱ^[�+/��m7�R@�ViLMHա��ގ�4�ߑ�"�f�g���&x�x��J�_%={.��%x�%�����\G}:Z�@����r�v�N�� ��Ld2�t����-TZ����d�#�.Dȯ�M��ݽ�w8��f�
��s�,W۠��s����.������Q�~��o)�$��v��	�g<8��z1��!�T�7Sw��{z$(�J�.�4ϟJ��ׄ��S���:��$3ZO��v�>O�x���遯oC�R\���,���"U�2�SL� �F���L��i��B�y�8��}?Hy��D#�����"���x�Z�hQ[�q�{����ސ��bȴb�g�|���и�[P�a	�g(�\�8[%�B�_0�����R��J(X�i�N�>j�!�ﶚ�F���T��U��}�ڋ���"��>��Cٟ�"�	�c��+u�p�w� @0�^wN�t]�����v�.��K+M�.�x��֛��D��@�o�5ǻ�/(��0f�Κ1�swB�O���
�V��}5Ԣu\{hi�V�"�}0�Ȏ�M�h7罞r�.v3yϩP`���A�ۂ�x�~���W톂p�>w��%�w��w·QU;6�_7g�8������GO[���h�tO����y���'e��Pe��D>�ή�H~�@��nbWs��$�(�p�˽�L���or����-����N�Ŗ��xW�����0��Zh����