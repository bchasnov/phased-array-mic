��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\����q�?��e�I8�b�Ǽ$��"����ׯ1�V0����)�.��ϖ4���b+��P��Ʉ�FR%j�qڛ\�<0��7�t�T�h����w�ޙD*Z��L�j	@�4��,8��1�E��b	��7�h�+9|d߬z�z�^� ��t��`�f�Sv�aځ1c�)�;�AX�3eW_�0� *+�{�j�?�] q�i�P3���h=TSO��WX3���C=_��C�ۜ�K�+Jt�7a�I>O<�]O:�>��U�C�xi�@�EGE. DI\��q2Y�,�gNt�)�i�cM�������_�"�0W�������b���Vǧ�X��m�M���7����W���)=l�)/t���d�+#��|�Q�#��L�� Z��l�B��=��������vT��!��x?�������/�!L?�pI�cD�����)UC�9�qaũU�#l.tAo ��1�w���of���%.���ud-���0B�)ׂF�N��1���0q���nB�G9�g��[`F����9lc?�ZZ�G�0�r�~�葉G�C)�3,}���z}���}����gpɫ���8�v_��j��~y��zh�p�|9N'�lF4#�R���n�b_b!�ĝ���t��	���6�C�D^x��ZMP�x�lE*��3�w�h9�N���>s��T���d�53�F�5���@�����D�:
�S�~~q�����ܱ(����:^Ƞm��t�l�v!��gӄ�?���= ?@��)�Ӄ@��TL�����/�E���!��\dhj$��v�!��@h ;Y�+ ���-Zy��<m EDt�0Sݾq_��C�*>�g�� �X�6V�5<(L�l�QH���-=�k�Z��؍}�~�U�	�P���˚� o�������M��(E([�[;DA�|u�z�������^`H���a;�`�d��"�#��BW!�{@r-`SE{�,���,��R=Qˠ�%�X�rD��JxUA�p�� Ӎ�uz���C�p�E�HY�E'Zb:p�9X��X�~̆�Ƽ�RɅ�x���s<��@��"<�'zƺ
9[��.s�s�����ө���u�Im���2�NXD�a�V�٧'w;��nJ"��4�H� �S�w:R@��^\f[@�y�K�uY6�X�	Vu{$���؆���C��I���f=F�/�9.����*�ku|��� ���Q��Z�y�����G^�H�vh��Ϸq4>G��?zw	�xWi��Cd�ǁ�i�}"��7!` ���2�A�=4M!���6��Ξl���'Z��g��Vק��z����*dND���\G�I̶�O��������=�kF�Y/	?>��߶��?8ﺹ���g������z�-�E�����@��]��Y��K��,d9�`�l��3��9����۟$l�	��[��}���#��9�g-=T�v�H�؁-WM��!!���z��|
���o�m��6
Tى�������ڑN�2RlϜ�$P��
��1y���Vw�@��`Fډ �~M�B|��z�4�����8��?���Z=QJ�r�zj7T(�r���,��O�Dp��+�#�=��r.)�L*?�ݻD��_X�q[Gn��4{\p%�hEe�Ɵ��R���ʟ�����H�|��z��ˠt�7���v��Ꮕ]�Ͻĭ��aq����|Ԍ�(</�+�02�R�4�	ڦL�;	���TVBY���,�&��#�k׽zt�sK�'y�0�ؒ����cj}�2��|���ѩ/�����%	o�Ʌ���G����d�+7(>�B�b�y��Q���/��=ǧ�T���,pǯS�Y�>��Q�KZ�$2#���ڳxh.�H�d�T��CuDix�չջNF�'��ei�:Kr7��f��k����_'�Y�<�@���
��KJ�H{�^���bC�P��\�,��/���Xg��5�U�6#q�ڳ^P&T�����r�� �@�#X����M:�qα)�1�<����Ƴ�ml�V�q|��[qs�77!R'�	|����.��4���ɻR���@�)�FI{��Ҭjm�T���T5W7�Z8�*��-��Ha�B:h��)�?�`t*��Ŵ.�}��t�{{p��H�G)lyD���3�A�����x�|�R3�gD��(�{�
5;<A�����^`�
�Zcs���z�#�OХ�����k�K�$�v��B���z����hs�(��Hń?ůnȤ������ղBb�#����К�#"#-^Z�꧖��۠�g�V��ִ+#G���`���`�r�ps4���X�z˷f7����a��`SJ�ز�,ލX!�B&B<��`�}��X�h�@�g� q�)�Qԣj�U����M�υ�r�g"��M����Z�y�	iS����_#D��
iFZ�w��':	[��hR�۶�?-����������(	O0U�q�
�T`��Y��rvxag�:a�����B� �+AOҸ��6q��N�گ����lR�qH�ƛ��V����KR>k���	�z	B���/�Q�(����`�Oo\��Z�-q�JOc�T��i�")11\��)}*o�}z}@ݨ,]�z�9�r����c%�����03#E�v V��P���XD*X���?@�d�0��K'�	��y�w"\ݎ�	�fZ%���b'5�8�iHD9mxg"���ӭ� ���n�P��f}��yZ�o�W>q-i���m�p�K*,�@�RC��j��	��@���v��ؕ0�5)�Nt�A.��I��&��ǜF[�8� <�'� V��;�	I�vn���q�9A���'"��`ˡ���
�r��8�c�����j��51]Q;͢�~֖%�X��I�m����E+T^��[Q�:b��0DW>'�!�_��,�����Y�)w��:��4�rc��:,��6뺍���l�ߎ��t9��ר��{Ge��x�j�x�!��X�Z{���w��r]�BF%6V�X�Dzp:ߴ����awy:��|,E��b����V͈*�3��f���bD�5�BN�܂���z��&�+�2�oj�V�o���jHP׳�񸊡����������D_�D���Ӣ�J�M���.�eV��f�96��5����Rr''(S��	Y���ʷ���q�]�	�1iH�k�ťdap��|��ھa�|��l�|�/�3dS�5�ӺJ��s��PN3��rY�J�#-m�7�d�^�u�u3��ɩmK3��m=�[���aCb�zsXR�̟@UÓ���{���s��yE�cN,��X)`%|�g����vx�k�h�'�_c����x�����)�-�?8���H�i��N�wQ���^-D��w)��2+�K�]��q��Z9�b���ͱ�9S��̓���ٶj���{�ܵ���t	�?L7��<�%6�]�FL������OX$D0h��&`�M�c"�~�:�'��o�^*�/6�]��2��g�J`^|�c�tb:y��'�w�eT޳��f�4�#C�8�(z ��|v�C��V�j$X�@Fc�x���'���45���)��㝫�tӌ��ҝ�_G�l-L٨_יF(���˱%�,��O��ݼ�<�;i6��|�@�\��ͯ�)����~���Ӽ��
J}`�eY�4{>m��jbx؜�셔e��l��}.��m�<�a��dH�Z�Lc�g������zY�_�8�r`L<�L0�� I�z(p����=�JΫ���UP�8	NjS�zY+����T���4C���p��n߆_�6u�?�����JֽO�y]WRS���嬍�#̡%_��Nr�U'�CY��I�R	��:��5<��eKor�J�%�9N��.��~g��r�InY�d���T��1#����<����o/��s�k�9Q�	����z�b�f2��-��\~�`m}̋D�{'���ߊjdpͽ��M�qm�U��Ub�z�a�U�XWS�ˮ��T�l��1a~�׼<DRk3ݬKbv?X�R8,�0O9�T�^֡E(��^¦�x�8��Ӓ�z��ȍ�]֘��Db��p.�n�
cH�-���Re�ǋ���.⏩��8��{^�Xw�^J��#~GV"�N[��_�~�Όp+��[���nU��Թ;�#s�� �D��E������^�i�1ĵ��oW�=*䀎�f��*�^��4��VEL��
�Q���Qr����R�C�6��-J6nU�{~)^Q�I�Ey
@����y��E��45	m��;9��Qڟ	�I�7%�Ć��,��Ǜ=)g}��ɖ�ڜ�, 7o��\1���K���j10
�sE8'�(*\c~����������cx�S8�@)�OC���t�7Ğ5:H
��l�j�����9���唈�J}
1\�mqa/���r�rŤb�x��O�I��Y|��׌qY��e�r���2��in�"��MX��	A%e�ْ:��������2�~��Xr;@,��IDQɘz*5�u_|�d�$�C��̢�F=���gL߬����#�D��|�kUÝ[e��?=�
�G6_��ī��h�1�5��HI���x٢:���p�<����w��P��bXCLO����-T��=��K~T�� �s����q4$��o{"�=h�z��yo>Q��ߨRuyC,x �q��̎D��61���'"#��;�K6�!t_�CYu 5Ir#n�͉�T+�PcM������S��f�k)��vP���QluE�����+)�6�ͻu�l�a2x�?���Z� ���ZN����[�ZT?s�J4��xڔ��+㖤���2DG�x>bA^Z�q_�M�X�Oҏ\��o���<�HíS�>�؆�)���zPf�І��o�Wo
��)��v��P��aw!� ��)G5m���y^.�J�k�pZDrĵ4e�-l6ّ8m�۱牉 ^~%�`�����b!���l�S�i��r��QrSo*Qq� vFs��¿�����=�=-���'_����y֎��	�R���
�P�-�a�[���P(���4���&�N4/����x(��ǜsnX(���wL��������K�R�����S6���l
���\v�z B�9�/��	��Yj8능�Ҫ/�>��`{B�\ԓ���ʐ4d���]Fpf!��Ǟ��Oɝ"}���`c�5kБ��Wj�;a���Π�-�@w�nl�/�h�HH1\L"�ϰ9H#��9uz��wE���e�Y�������?��`��.;���O9�u�m��Yze�Fn$"&���D/�SF��`B���Kq�����j�px�]��`?�4�3^_���ѷ���Zhq'0�x'K�f�1���!�	m��]  S=�C@y��J�Yֳ g���y�I�, rn�X�eMc���۪ERy���������.���$'-��vT���l�x����+��Kf@g��,1hك2�h�\z�k�)��J�TӀ<,r��>ӬIC4}ڞ~�%�E7��+�9�c�I����_f����H �4!P���o}��r������7M���"�B8�:�=�F�p,��%��x���0@�ad��x8 aB&<�<�~�l(nc���:>g����������J����̇R��(IK_q��^ IZ��~���%�ݾ��0���$irr�-���*���t�=y_7D��12��$GW��O!mk�� Zq�Z�M�5Z�����|�1�k8#�~�>+�TX�V�q�w4�jU�$��˭W�~����6���{���i|f+��o�5�|�#�y�\���rCe�:�$��,$�:9]k*�.��X�>��pt%�C�i�S(p�Bے]��^��k^M!��o�� Z�7#�S=��Lt��ί[��lZ��r��;Gnb�H���A��R�*�d���O�����"+����8�Gf��:�"�[�@)Շ��E}�бq�j�T�2!�n�o� ���m7�$R;�"!I�D&Th�JE+�V�n��Kz4���_�̒ĵϮ�%�4�'5�X��"��7�7�}0�mu�onr�@�]J�] ]�ܧĦ�t�OCV^;Zo���O����Gs�V��i�)���g�*ARu�!�o���zD�:���~F�������*��o8T�X\��cY&>��sc��޴�����OO�߉ mS�w��=�8? ��rmc���٢�}#�� ��8�"|�B�X=V"�kC�Kxx��[��.~V�v=�
�����jC���@���j�c�f5Qn��~Je�-Ɉh�~�f75�޽�~x��*��	 5�=TՂ�^�V�˞�N�}$\��8Op/Bv �qotJ�Z���r6�[6�U��5B
�0�@�nom���t�d0��jV��i�[N���0�Aw�7/�7>>�-��{F]�,g/��i�-*��1��h �ÓH�PT��M�H��h=��Z�&S�P�Ƞ6���+���-;L��E��G4C��)2i��N<�[�jg��q�8���7�׍l�rO�H/�.2/8��Ɠ9�K���?-�+:CR�ZՓ�Wꈜz�\���z;�%�)�n�ҝ�K��b# KB�&�e���a������M�eIy`��X�3Ҫ!e^�0�%����]��#l-��� �_�R��§υ�z=�'R����n�) �HrCg��C��!���Ͽ�� �L���D7��ڃ��=��c\�!e��3ef�v�=�W����S� �d$"u<'c?5rt/(�35Ꮤ�.�%Hl�g�r[n/��
��P�2޺s9*��Y>�r���-��Ӛ�<N�*����px 8��J��k"׷n�;Nv�o�Y��O�E�oT�($�&ci4�d*�=�x�1�Ǿ�I������^�;�(��>�3��c�LI�Af��jb�۴���?O-�����e]�4G�ҷx35�⏆�������'Ny�4K5�3��E��sSs].����X|�n�5ͬ}L.�Ѥ%��Y湰�ש5c�ks�FO*�rwr� '.R����j߹Xq�|9�[�w
#Y������%W0�!I
�w���Q�I����UuL��g�n嵻\
�����&~4z�<����q�8�'���� �#A[i6��f-0iuk�`�ۤ"@L�S ����n#�Gx��B݊�xKg,ٍ԰�k��!���4�:�&�Q+#�(���f�äQ��A��t'�,Kv�3�d��兌�F��Vk��Q\�'H��o{ _%a�ǡ_�
��s�t��6Z!8W��jO�����I�H5Nb�:�HU����Gd����uK�+\���Ǹ'�[ч1T�/�:ݰ��Ղ����P�$[�� 8Փc/Ef�e�k8����,c�P�X���'-���>�c���d�Z�=3�L�qn��\'W�#��oӮ&��QV<���b����(�4�ʌOyV!����ڟ`�Y��1�y��Z\�����0ֆ��/�kQ�=e�ݗ6T��4�E����z��jagn�7��v��s�w�/�lY{�M��-�^C�․� �EqMn7�����z@��o��@u`���B�ڗ,��	J�𕿖�M�B�=j�O�lИC�/�d�Kz�c䶧���li[�sm��#~.����էV.	&��d� 3d\����y����No��L=H�X�z�-Z�?�@T�z�E�s�+��3a\�JP{��k� ��p���EIj�ʽE��B���,[�}��x����ң�ӕ�&<� ��r��j��O�pU�EI�f�A�"<IʱzxT��H�9t�ˁSB��'�_]F�L�y�|�sX��E�W67A�*M�;��\�B��_�׆0�/3n���H�eK�GȲ�� ]���!ol�N�T{Y���r+-#�*���:v$YU���~p����r�[%�	�	SRph�����Y�~a�K��袠���Y�ݞuF;DOos^�-��a�R��H��\�l#DDs~	�_��A��i����F��nA���ŏ!@	���c�sx,+;9+����uk�������Y`ǌ��~���!����v�zZjgi��Yq4T0M�¯{�c4?̻tG6��M?F��v�:�1�a/�����ص�7��-5�*�m�D�N�k�a�p{�̥����㋫3X�/��6�~���lԴv�Q�:�lob��,,˖Q��`�����h�� ��N��]��C'����_�^��^NpK�Գ�Z?��0~u_�/�A@�r�Z�.}!h�&�VW:8��|L7�6B�F��\���k�|�ƺyqk ���$3�/ʷ�O���C%��g d%2?;����H�����]M�3�J��b`R���C����5s[�r�D>0 `�C�e�V�壂	���&@�����|���Ѱw�̧��KQ���RQ��i��j�e+z�,X�99d��X�.�(ef|�|&*�(�R=Wb�����1 FNK�jҊ@B�I>MT�aW������ԅ�����R#V:��m5D��T�Z���o�wg_��{J��0�b<�c{��Z�*h�D�h��c�/ +����
O�V�	�1��7>?!:-���C=*�-uĽ�3�.]�^g5���
#e�?�^+�o}O�M
d�ow�88 ��^��*�&N�����wW`%��&�(�r��?���f�Zw��r�7zS$J��6S0\k�in ǿ^�N>��������J7^�S��"r��{O!�YuL_��@��:��D 6{kzg�d�X���W{n�Z�[��@�Y��8%�O������G��*]	�_�����U���u��a�J#Kb�4��)�������B��t���[�uG�|g���C~K���F3�o�^��(�����lw�~���H�!<)�Ճg�g��� �h.��=Yd�z��
�s�~����'�Îxff�0��+$�%8�
�2�����ƻUd��v��Dr����Y�[�I?�f|�5bN�4MG/*�n�B%L:F����S�Hm��3쳒(:�L$4����Ox`r:��%�s�~\B��*�5��W�#2(��b�)��챈M5��6�	c(q���@�� ��P��_��=�r����W��i ڂ��Zd"���E(u7�"��F�4�x�w�0�;�6�����ˍ53Lн�����8���MHOS�NQ���c�"���;�����dz��o�x�{m�KDU_�RyQyG5[	ѥ��ç�M% �|���%ʫ �8�9i�J����B>|F3�W�&�eF���x���&�jޏR�xT����Q���l�i�AW���\c���g���Q��Ǭ�$:�ΘH����m��<e���n��];�Ȧ{��.�o�Aq����"�Ћ~ksm��w`&K)����l���'�tS�c�`K��٭8G�?=��łG���	��0���T�DW/�C��UPOp7���t��e|��/��w�6�����D��Vc?&����:��)G^'T!Y�������a�1�}^k{�$�?̜�ӿ�t��.�4?���=?��2_�]f�:@�Ŗ�kW1�3�p$f�v+��9ܪ��	0̜�0	*[T��7#@1:���"�+��V7�5z{���_]_��x4�ֶ���(�����%lG����q�(��MXE�4F!47��=z9���G䕸��I�QI|c�>�Rr:����R-$D��b՘�іy�Lb%]���X�>y0^���fo�7�1�ll�[G�ľ���tF��c(�o;~�*�Y��M.V�I|^�#:�s}��H�q��N�8)"_���t{��UQ��mJf�<8l��)�.2��OJ?�����\x<g�$9,�m���ٱ)��a�����Fp1�j� $�i�a��ʖUC����?ktX��m@jI��Vb��Y}���"�fMi����_D��
���)A�=��.��Q$�̒��M%{�n}��;2}BM�����c#H`e�Os�h�F�&EpM������pg6J�<W/V�`ӹܕ��w-W���l�qx.�>�I!-o|8���]����&έ��bq'v����3-x;�sS�v(��W��ރ�3x�l2z��ShPp��<�q�K��q�L�����fi:l47[��@�d_���.;(�H��z��_��b���;�^&35"��Wp\��6�>�P��]P@{@W؍`��!�쏞��e�$e\��R�O���D��9�����]rW��/���B\[_�&�}�W�����F�)��)����#�%��>�c���!�veK�����'v��@���羰
}�ĄD�x/"6�*��:<�1soǁ^��U���|ß,'�N�/^��#b���$�S�J,�2���[K�٧���+^Y���+r�e�L%�%R�ԓ�y�kG���M���4'k<aS��x�9���3�����Iţ��W:������ ��ѡ=m���ޡ ��S+jjCW_�>{����f�h����|vČX*ʤxrR���I���	])�A_�ja�bw+8���;p��Er^�\��:#2�5e��kXA�y��kd��d����x*���K��g�e�s�L��}ዅ�o�r�o�k���	%��.���������;�%x���tʩBW6	��78�G �X� �~��02q��"���x wr�(li����x�6�) ��rm ��wx+}:oߗ5�Om�a/�=���(�-�[Y &�(ݭ�c$&*#Ԯ����噮͗�K�[�{7Z`�v�5��CC��CX�}]H9S��on"M���|9��FE����P�j��R�y��(���Rw�P��8Z`����[�X״��Ą69�FY���V��Uaį���}t�2�E�P#e�K�ζ�t"�`1B�*.�|2��h*�o����T��5�r�Ly�\�1�&	A�"�M��0�$����9߇����vR����W��^o��?�hP�O��ʯИ]I�h��j��3Z���[�YLD�V�K����ӎ ��k�#r*Z6o�����1$zy\���F�ĝ�W�܄7|ܷ�ZN����[����4�|s��:����������c����W�i7Ww�����D�(����k`N��L����#iY:��s6���L�ma�Y�s��-z\RwTՁzT��Qnx���kZdk(��V�ۉG�����̪;>xQ �R�����t�Fe,�Y�J3��J>횗��o��+L5��P)b[�05�J�&��X,��y^��闑�=Ǩ��{L���"�S?��t��(�4�ֱ��*[;�8�4��e��Ke���f:�8����g}�W��CX���/�(�\5tGV�o������[/��b�����/��KD� F��.���MI���mU}�25����G��d�"�^�����2e,tG,��ZnX��6�UAn~BX��z�Bm)4����Ų ��.(�M����u�6����&8k�������eR����`�X7�Wl�A �j��|�d��2$'��@/������r�.D�O�g�t�T��@�ꌩ��<��|�*j�l�8�4>���o2�;^қ��|t�
�ݙ<,x�`�D�m����t���ǫ�Q�~���%U�Ae��%I���<H�|�%�8��T�_÷��+v��ج���r%�D@xԯ��d}ѡ�ȯ&�2�-��O~���m��u[Pr^�ϕ�ù�B��w��w�Y4��*��֩*'��G5N��V�~��eA�w��l�G�ƧD���h�4��l���HB����>��H	Z���;Ú�o�zwPPhX��[ /�h����"'���b��C7�KThS����z�9{��A<r,~������ēlr݋6�tQ�<�����i(<�Zn�]���Ru���Vې+�Z��8�H}!LFX����W�B)ݡ�Q_��7k3�0�8��[���H��ڜb8�6i��g]���s�X�|�ڴ�2t��\�P{�Z�N�Qz�|w�@����5�H���v��-�|&��:�-���a�%�����_-.��S+��|���\��� I�6*�b�m���a��:.���O�=fv�T��uޡ,��n�4g�"6��jgEe�?� Ӣg�g�j]q�M�.���(dz�?�)#3�$��t�N*�f�l�;���ON�ے:�m=sv�Jy�љ��!���k�l�~+'"%��"��l.�j\&��{^f��K?]_��J��Б����κᛠ�~����7����aܕ�D#���}�I6]�3����z6�݈�8+=�PB�i9 _��(N�}���/�ƌ�vuU�P�����#�K�RQ��Sp�$0�u�Q�X����,����q0D�@���0�{#�\5��=��o���̈�e��[��/3��j3���}��1�,��Neb�P���UG������<��K���x;  ���)rb�-.楚�%}�to\,�CX����a
֊wj�Y�D��&8Wx�1N��NC�V�2|F�nO�^�reT6П�o���.6�NM��Yp�U��5����_Oρ������l�Ǥ�I�l��2�T|Ȁ�!�ެ�o*�٘&	����r~Vo��͚g�͘�O�G�C�9�*�F�H�E��Q68K�j��q!�u��/:aE�hNҰg��^^И�G�:1�i6���u�V�?.��{n:v��qfw@��9@Ҟ֬�@ߴ�E��d��?IP	Um����^�=����u`��y{$a������дM@@���"�h����ኰ����-��\�x���O���N�XMk�d����4� Kcl�A����Js��a���?�L��P���w����I��m熤җ��Sg*4�q�|�dWK��&N�ȋ3G�}{��C~�}�9v
fw���W��!��)?2*��z��*�\O~��]�0�՟7�	��	qu�ˀmX:���[]�9i��퉣}��O{'g�I���G��Y4mV���'�Cn��{I���9� ޺�%"�zR=�A���>h�0���Y�%�cO.��z?��֝!���/��<"ȏ@5����g�ӡ�_���t�m��!~��6�֌���G�4��A���{Z6k�6]�$����-,�0_���t�~g��)����l���ë����ԍz�Y�q�r�7�E9c,�ʹ�H(�`�9\�]X8��s.idP���=�pq?$�^O����?1ł[%F�8)Z�5�y����cKI��3�#�\�G���U�:�O�Q"�4.���*�k������R���U�
)��T~45�(�°���L���� ����:���R�I����>FP��C�
~�n��K���cDp��l���Z2���ǰ��C���K�6txG�"�%�>�\�M2*W�r�
�>�Lo��5k�.I�K:��Á\��M����^e3���Νx���L�0l�|ؤ��0C�}�zg��W�bqo��T�ɸ|�'R�L�ʢ�J$Դp&%+����nXf�˘&�/�Kc����d��ߟ10,���H�5U{O{�B�^�����*!@�i�Ko�����&6��oώd!7ŉviY+8�ѯR	�B�~9��d戜��z����d��B#�j���/|�o:٣��\��������An����\(��`��w�)��jOo�"C��[`c��k��!�@z}�PX���e�����a��!���^��UZ�ސ�ꟕ�%�F��Φ\���Q)+�s�q�Ե���� �qF���n��nPO@)O�R�y�q2�H1�M�ڐ��������g�sh���Gs��"���*��j�r�e^�9�6Y�#դ�2��.���� �*�
�q�qT^Y���p"I�>�C���c�2E�w�F#d�?3@����)��}t���oѦ���Ht3�z�_��U��sg�f����?;��ul�?ġ70���}��ͩ�dW�'���4ѝ��CQ�͍o���Γ�t����xE�o�_96��8K��s}*�ׇ-�`�#��-,%[�h)��J��I1��;[��n�uEs�~��ɉ���]��>"�o��J����  Q�F[SizuN�f%�fl묱%#��<�2jI	�l�_�۸�:�X�H����Q�"']����p���Kty�H���ֲ��@ᗱݱ�uR�l���ةv�F�  ��Hq��v���$����+�T;��܉�^��ɪ,�}�����@�`
`�p�B�� cy�Jp��L��|���r[YX�@l<����g���5"���E���Wnx
�P�R|���Fj'����\5/���O܉����4<Od�Z��޺�+1�(�}5��Aj{�
�j�B�`c��PZC��#׃Ռ��/RlWπ��c��h��e]�+�R�7�d�g-i�5�u��+��Me���X�q�$�u��	�acnd-���k��',N�O<�MP��}����0o�) #���Ey�{>~��GJR0<�PR�|/��}�\Ccb1o�k���y���4�N�Dы�oZ	x�MEP�r�ח�� �E�H�d��E���?���ܸ��e�0%�.9;KԹp4~���tos�>�A�OV� �+�ˌ��gv�Vk8��:�s�W�R�mV&~��+ ƥ���(�=E�J�|�d���7�8�ۖA��V�I�H�P��1])v�Ԓ{(	fq;I�֦B�]�P`��������P���BE�5g����d��ta���Ѧ_�#@��P�����]U�Q���Xx1t	p���H��Pt�gU-I
��ȼ�I���C�Y������C�� -y���I�0Lo�G�ߩ�幚Q �0+�M~t�"�\��eM��M���_�<�1���g�>��Z)�gZ�O� f�i�G0�m @w���Ҁ��(qn��v���ƅ��m���|G�k.!q��W%4 � �i�&1.���Ԇ�rc�mf��_-�H7�L��;�%���>������j-��������Y��A��$���уK0�{F�%�~U�`H�S���l�b%E�G�9{��i��>X3E7���F�`Ө
\K�Ӏ`"N,�G*�j�,F4����FkG�	����If{e��;j�������W�|��?���˽Ŕ/Ñ�#}�S$�ԫ#��"��x�H����3/ �G͂�&Og�a�3鱂���e�x�P.�]�W���4ef���^��.��
~D���@2��&�X�&�`���9��D�D��;?�}�]E��V)�������E�32��_��YC{��G޶���v�R�0o!��\�.wD��������M�yZ3Ĺ>�2����s�Y�1s �w�3em_9ߓ9<$?J����w8zbDe���5�X)���1���f�����;ya8-Ǖ���u�9]���p!�1d�{�>^���6�����.?���Q%�T�X���͌�<�Fˮ*���rb%}x���-���x����=����^��Wg3~ʾc�j^�_�$��� ڒP�?�i��=�8�N��3ni(�x�h�kR�i���	���\b|�<L4l"J��*�vq%�%Vx��L��`d�n�`m=z��c�}�Փi���)F�m�v!:�R�k>���\�����[��}o���k�����D��� �(�]��J�v�gC>Y��tTpg�bIm�'����G��'��p!�҃�8¥Bʠ�L-[q[�w�����;o��(uȩr��Q8���k*oϖ�3�֧����<ɓDA߳��㸂�&��y�8�� �&D���e�c((h��#��kP\ܑ'�w�C�R��!㭺�t����^�XY��g���@��s��@qv,�'�����9:��f]�D�9��~M��I<�q�p4��}r�^~���ܡl�,
�8iE�!wp�R��1�TsL��:�c+�\\�a6��E������ց�޳��gٽoX�I����S�������
�z�q�)-F���&�k��o.�Pi`I�,�ۼ����.Y@4"�~�c�V):�;��=�*[�������h���uƕ�̪��3M�
��x;�[ӿ2���s��'����/Z~��2u�K<|v9b�ɘ(�Tp����?D���l7��|T�_���Z`��UxQ�3#���W>���W�,S��8�g{�_i�K�}�V��嬽�$�W��֑E�d�i�01�a�yO�� �����9|�����h��0�f5��h�@J
�׶�`�`���T3�A�5��lY}���d�X�K�N��X��G�l�=xx4J���8w�Ѫ�I�_�;\�L��A7�C��R"3�'s�׷5�W�f;3ԯ>����="��4�^��9�����`5���Z���K[�
P���)��?�~���"	}ʒ��K�u��i �>fU>`�pZ�6�gv
�D��Yyv��[��QI�M;�P�L�C����v�T�{9;�=X�Kc��"RX��_xNQ|p��j"�z��_�����1�����HE{
���I�Ln����K9��P>��=��>���>���7��u�-�9C;d	38(��7 �G/)��q1+)��Rt[�8(�58+�T�%0�z.�_��T��`����~��B����z�:�!��/�E�S��8;�G�	 �ݎ`�w	:�Յh8IõXm�ވ;ę���B�!�LP"��xٶG�V�!���:�FY��+����+�"G��vʙqi��yP��^l.��W��DT�<ԉF��y�9����!n�("�V׋���f�5��X�v�K0�2/,�
��<[�9��]V�Av�xq�Ƽ9(�{L���˄�m8��y�5Y�n�����#�Te��>$ñ5�/G����j�	��D�LXq�`��ʺ��&�>!�x�؃����{ekg{9����j���������v��:��O-:&���4
Z���S5T�1b����[*�J��'��Cɝ�g��@'&���UX��4
��[�������1�tM��C�ˡ����ز������
o@��i�_��UՑ�}��L���>��Z����fT�.�b�@��C���sRc�m���B6��jzX�xfݑ��Ϣe?i7t�H�F���y�)7��"o6N��Y��w%�i�����l�i��;l��ގ%�G&�	c�c�)�����gh�v��|%77N���]�bh��!5�2l�"����Y;:QI�l������^���Ä���FNSV�0�x�`�2�Ҥw�_��Jݙ�8a��oUu�<�[Ё���VS�snp����R�Wt>+-�;����l<�-��͵�NK`�lg�-�ޖ\�UK�%�{�D=I��-ץA`�O��A!p�����Xw��\��E���*಍]���l[DQ!�m{"���(n�
�N�]��O,�U;������7R�?���Y�h�ya�#�����anFCI}�X'm7���!ڸ�4�R�D�1�\��0����]-CBwb V���r������Q�da��ˤr�i��RG)dW{%E_<�U��Q�M�b�P��F{�N�+T��1�3�������#��(?o���w����":"v[p��v(�%j���vB�F�d>K����"���wc���
�:V��4��T�͎�@�_�ʕo�Z}��1�4)�[�2e�Q��� �����d�sR����EUƲ�++��W0oVv]�\�����QOa<����y����A?Ff��e��$�v�E��ǉo ��	�W�㣯Y�`K��I�=�ؑ�MKIg����O�[��)��yr�(��G�]X�/׍�|�����(�s]�^i�M�~�w��ps��Brv]�u�c#١5z�CQS��ǿS��� �Ea�kk���h_���������CҖK1��-���|2c�SV����x�/�,��Hy�{���%Q�t↸�"��	��Y���7�D[�*�:ɍP9�b��(�L�.U'�4<���~[������:�h:��aR�+޻`�Sm �b�^�'up|���\h׀.X���X_�����w���7]��2D"nY��7�q{5��o��g<���W�h�K������;�p�*��UA5 ���J>�y�i��m��T2f��V{��m�c��w�h6�����}�9<�Z`�W��«҅�1�#���i|�A0�sSl���!�D��}�Xtֵ���<�x��L���.�Te������@���Y�~r���jq:N����5��������S��$�7��ϫhv�$��7�B�t��f��&p�y�����c��,��;�~���PCŚ�T�����fE8�B�3��s5ʑ�	�$]�,0�Qf��v S\��3t���(�NS�M~�ѻ{��S�Fʻg2�_���>B�á��S>�&�<�Y�"ioPƏh��e���y���#�l��2N["9I�]�.rg^�������M�W�I�����e~�y��%�����~٧x�@�H�P��i�]���@�B��b�z��u ouX���q�<M)��$��Ί��JA�"��8�'J������l�Z? ,�bl'����+�O����b��yVV!Dk�cЂs�f� qc�E$L��勾�8�)���O��uOI�k�h�/�~Lvw�_Z��9���u�9�a��E�i��ꆚo�<>��:etӸ;���
��&��<&��WCZ��=��ǒ���;-�~�}&�.)@�2<����L�_���h�{�{co��!��BW�i����Q��lU^����w&�lzR��	*�����*0��sE��&���=��W'��~tRL\��'K�%��ʯ��:���b��c꒪����xׂ�DL��Pڶ��m�+�h��P~��V61�lj8��P������G$�vP)�L?�7��m�Z�~Hd���8�k�J��-վ��qXn3s��^�x�S}v�����w��Af���jo���Y�Ȯ��e�S���,l���}��zD&�T����N�����H/ߣ��['�0��"�t�˳2��o�%���&�y x�o�
��!":gtkj9����-C2~VbaJ��0�j�����~Y3u�\\�#�&3�<�Ň��;�#B* �K�,� {Br�\��T�%)�5e��ﭬ&_��x�������e5���$���4��/�b��)��@g{~���C����!�O�}�*BJ+�ы̂A���XQeF[V�g�ݡ�b;S�7D���MW��6QO���S�^���ٔ�G^�UN=�\�[��׵���.E6�hq�9V��K.4\?�ѶJ�B˳���C�\���-N���:��8P���W��K4�MV�5����Y��ex2s8ͪ�S���t�L����n ��.^��?�c7[;�6cpتW);��`lUv�z\�U�kp�+��jC��#�"�x�2*���"9j���g���)wB�8�q�8HV%Vq��jć�\����,�!�U������2��QF�^D�<��(�Ad�C�A�49���ަ#��.��e��ޡ��ݜ�w��iQA�<�+��O�x�^;�A��ĵQ�Va���R�%��A�;���P���ܥ�vS�A�/� �!�w�\^��"'	���a��f6��m{h�$ss,7HRi1�]��^��.����(�k��,�@�*��F}�g������I�h�F l�Hȩ-]��d����d-։.���ߞ�]ϗuz���y�))䝄���t:J����v�賘���X���)O[������w���A�j�+��tG\h��
��F�%�(��]�
\K֕��g�W��&i�@��q�⁢���~BO*�Ѳ��u��s�0�!�x��)WĘF��2�R��f(E_���!��)J���-L�8�Q&A�9f_��sC�4xP0K���K�����8R8��u�P3�ϫ��}�U�ɲq����?��HT���Q}<����wuKA���)����o2���Չ�t�SU�����*R�����H޳��<�Ƿ�vjC�\��`�1��̭�;��Pr2��λ 2 �ʙ�S����Z?@:�kK~�K�`6����g�����`"F�,:���w#�S{��<ư�V�`N�n$��{%2�������Z\��Po��ɮ[&�*���j��c�zw�x����9;��b��E�&_
X�:_9�\k	<�2��˵�:ZQW0U��;��SjY@�#~{�h�x/�.�S>C���g��`:X�ٯ�	�-H��Aۜղ�MԘD�^R?!�[�jY�3�B��#��05�>�H&�D�"$Q�#4뢤�I���c��>ܒ���-���X���MǕY��w3M=�Z:�1Ղ�"s� Jj1-C�3������>��5� nbbaK�˗��ӥpH��+�p߂E5Q:7�
�Tηm]���}�ڇ�+t�/l����WzkI��aDY=6$���s����+��iTex�� ޷���9�P�~��J�;5���Ա�����(��Jh��2t��J�|��9���Z�ֱ����3�$��#�O�~q:`&[�8*��R<�p���,ګ@�-BGgYE�se���8�Ȧ�P$��Wψ�Ns����Ik�/)�q]�V�(y�>�9�P\���kZ=g����°Z�l`�{/���MZu�*����c��G]����N\cdq7T��-���	�֖����0�3*�m�i���S���ޡ�{K:���Fk�aA ��"=C�����<~���Մ���"����r/M�<1%˨>����0�U!2A4z�E�.~{���	
�m`|����Z�.ŧ����|�E~&U�;�j-�k����L�d*�M���4{�B7�| !��{H���?�5��$ ����w�+\�b�ًU��+����hAL��!v�Z��2t�_9��S\H�nşյ�� ��9=�8$�������Y]SՍ0ł3�r�o�/�O&����6�f@8Y@� �
�U�l{X�;$QH~�y!9�i~>G�C��6�33e �l
0p�x܄a��E�'��.1Ɇ픿L~2���z���J�]��4��1��ґ׿�/o��x5Yi�}h^�zM�٣T��EҶ'�L��uD����Q|��D�Ƥ?��\uH�O�����Q���ĻT�+�����������{f3ax��녉P7>ٻ訆�j,�-�*��a2��������#p�
�M��	��*���Y�\�ٌ�d��s,ħW�[�P���»M�"=V��3�Ϸ��8��bn_�e��7߾Cn��x����Y����kAMMC_��|1�瞗�'s�!%����Z��qh�B����,������S9ڨ",��借ɼ|~����q86RtM@W; ��b=��0��o�E�7���b�.mM�QW�뛆ۅ���ˊ�9O��ƂQ�qEBi�N�*bQSb ����F8-)o!�;�o��ů}�r�p�9�P��敳%=��&��A�C����q���7�,���d��!F铧-�R�#ɸ��u�w�'��L׀���O���ɮ4j=	+Ԍm���F��||�'*ڒ���_�T�F#R_�ēs.�ʷ"����3��y��O���5o�.]XXq�'��&�`!���XG�0�q��NX#\�;�T]�Ng�5 ��p�E>[RX���]�V�5dm&2��O+���	��$"el�R��6DB�<�@�tޥi�ڍ���:"���
Z�%�< �kQ>s��T�����(;3���N-�pӵC�R��M�Bk�:�`i��.ß`�IA�F%U�N��Iv|�3��� �D���Ҽ�~�	C��v{��:�̘Ĭ��l#�(!�g��}	�i����y��t���y���-�����F !��Z`S$���+��*'���/`�v�����Rj���n��S���G��pU2�� =A%N���6m���.��*:��2Z��gN�����-wk)���8�����F	4pF=��r~!�ś��U�˅R�4�x����r ���﴾۫�/����(��r����r� �.�� ���u]O3ų��+{|t��
�_��Dǧ�mD��ݴa�,�P��0�y�4}������д�׸�jV�p^%�<�4���՜��}��:��|e����xd�):$�<�ƖQW���?&�]c-��&*���olP*��f�f�|4Y��R�m)�0�������#�p���Bދ)z�@Na��3ϛt&(��b���*<����C!JH�"���܇���+T��Ny3t��Zz�=,�dfN(�!�b_��Hkr�_1���<R�kۀ�c��V�\�t�QM�!\���~dĤ��?��۠F����űV�K�WGJ��f:���mBL�
�ƥ#��>GV)Mo᰹��L֎"4���C������A)_�S�\JY�nJ*Ω(��^���/��-��<�+y��G�#K�Bq��l��	����|���U쬉��{��u<")Sq�0�}
'�o�ި��ЪD�#{�:��W��(�� Iux��#��1�f|+�y���}����ᶶ'cdm�N������琜^͆�z��F_Q��\O���t��J��X�lpuH5x2ăO�1-�G��pL���Фi�"�Y/�*�%U\����3V�T��a�������s&:>�@������n��
��Cc5��W��	Œ��� ����[�K
���Ic��� +���(:?0������N�u��q@ '�q���'�|�	0=�g��pd����!�/>��Fhl�O��ι>��!���zxX$603	4�r�q���;d1,9��Mw��:��
���A_���	�ˑ���� ��$ڕ�b�eK굗�,b�C��:��H�-]#�i����+�5&����F�'b_!�;�)��ڡ@H9�%t��Ãe�Krw^|���R���B6���$բ&����|�)
�+I��E�,z��3�Ո�g>vGнN$Ҁ����4 ���ާ��[�m�r���:���5��'\�X��z%��{����jd��/Y9W��v
<�~���N w�P�&�rZ��(nh�0Bir�� "=�?;��j��[����%_ۿ$����6�nS S���{�d;����z�-(��?��R|�;_�{��&Ne�����8��^�{;�"��RHa��i-N�ed̺v��N�EΝ������	�})���5�K���r|�Gi��7F�߼��hS�I4C��Ya���2�@ĸ�������
��:��tY�u����P��Z����� ��-��#��7�A�9��K�e�/^�����`S��5`&%���	��z��)���8�b�8�	?De-<�\o8Љ[�#�(�sä���ecuO�^OܥY��":)U��Ȗl^a�/�)��Er�jj�V�����S�Y��?J�pY��3�7�WS7�4�?7������jՒ!J&�q�A��
�g�V

Qn��W�����ŏ���h ����֏�u;f�������@��8�'P�����gǃ�r�C!�p��N7��Ce��c	N%�_r�{�.�ҙ�_�b�����*l�����R�d�Tf�8כz�i=�u���FM��{ ?�4|�N˿����P�ݏ��6H�pu���4RC��59q�y}=z$1qh	xrtEHB_O�9��<)"߫+~�} �-�j	z��@��6�Y|�B��8!+U[�����&�g��w�0g�2)�Pv�'6��_]���Z�T�Mr�j����V��8�[�Ɩz��%��B����;��������#�8u%�~���V��HW�Kժ���t���,��~����� ��㼤 8�F��Y��^;���gj�l��
��ԏTݰf��Dܧv�ʼ>
dS V��HL=/���ڻ:��̀V�z,���7�����>l�z*�o�Fe�B�a�@��i���I�撗�<Fi0�H�pK�d���A�	U~�1*v��1t��7<�[Ӭ(�؊��j���j�mnI�`�y��<���*�JB��b:�E���:�n�f�&U��8�U�=���+c7�~D�!��'G�/p?S�Q��x:���L���{']΋
�DD��So����\���N���7���.׵+��0�ӌf31��'=���y��:��,�A�Z>k<�b-'Nq�Z0��L�W���@�xQ�L�L@�A�gM����q�J��eBP[G,�F�%狡��t�ZQ��z+M���W
���]b��Q��?K`3��{��m��{�b��b^�W�P����+@���":yy�q�xu��¥V�q8_Z���\#B���By8�ڬ-:i	S@�4�.���(��uM����	�1������<�8�5, )l�f��r�[@yw�+�f�'��	8*VI�1���5U�����8��tk�/�bzU��ko�EG�ܡ�c���Y�XF��� "X��	���������W�*ri�1u��A @HLD��N��D��I�G����m�.��f��LK�E3���Z:�'�I����s5V�ox���K�Ȇ�Z�%-�_2�q�؟M��,�[7՜%7=7��A��U�z��AA	��{�]c��V��$�=��e�V*��ڐ*����N�Ɩ�����\�M���|.�.��=g�l�E�\�ڜ<؅��3HZ�S�$h{�mE@El+��ס)*S/��8{I�	�zRc���c�sq�Q�y�����uFQf2�$Q���-���I��=q:�'���a1�.M�9`��j~��'�τn*K����M.���<A q`�~�w}^����°�kY2��aQ.#�OND�0� �0���A�?�Hre��Q�th�ѰT�=b�r�����
�'J����RQO�|�Z7��	�Tm�#<��,��_�"B�bn���ɴ�@�H�\Kɝ, ?�z\���"�]lk���㍬ș7W��6�M]ꕪ �bn���$&��˗�Ԏ���K���o�?��	]7w��2�u�Y`��#wR���Ms�?�.0dY�2vY/���xf���ҠI�k�H���luK��O���EՔxY3�JH�f�p���!hT�h��>p0L��M�t�6(� ��e�w�Ȧ=0��4�I���{���W�/VN=_���Q�km/�w�_I�qŜ��4(�>�杚(�\��'����V�6l[���a%�u�ЈTYc`�D�e��i��H�r��7g���ފ}cvf93�8�>7R�ԣ�$�����|�m6qL9}� 4@��} ������;�rZ����C4��FM�kiҷ��w�.T9�Y[Ɵ�j��{+�:x\�M�	>_��	EmRgp�g��r(��ߠs1��G��(`8�0�ḰJ�wHM�6?y����|-̌��ƌ;PO����J�l~q-&�U��v�7-���L������|�(M�`�h�
w���O-0�դF&�2ȭ�n��t�&��u!��Jt�p	h�g`o���rE��Ĥt�_��K�f��^�'m���	Xe�,4eKi����2p9..t�9��a���]��o�J����W��J匔t���G\s3���?��;	Q�Y�H�@Iy8�)#�5�v�VH>���	�K��ޔ<��_@��%cDG	��]��KG�z3)�`�;��v���ϰ_-���~V��L��:�	��iԏ��づ�Z���m(�}�"��k�'��W�?��f������松�n#�7;��<-9)��y4@�?��m1/��>�v�8��V���0Bñs]��9��M��}Z�T/a�Hq�@kc�+�	��JZб7�~����n³~�R�V���	 @#��h�~1Z��B -��3& �5����"���M�����V.�x="��`�"�qX���Ѐ�(\�-+�W�4�p�l���B��9HO�n�c�;EW��t,�`�:O��.ׂ��0�kC�ԥ_q3��g ���P�Ae������:B�z�ࣜƦ�S3�nލhq`E4��Brq�l���-�:Ϛ�k�O�8`�b����aUZ��2��
TU���ܝF�0�����#S�f�T�N��|��Vx��φ=e�@��çi����_?��)�������%�~�V�N�,�q�%��-���u+̂���!o��b�g4�2p?��S��Ϥ�Gix[�Br��X*-q��h�X�s$�;-��X�Y;��7j%�L�ߜ��0�\R�>�s������p�M��V���cH��1�<������Нt*<�����=�ׇ?���w���l����>}ſ��r��F�|0����=/�i�(`ↁ�Kך�&д�0�aE�i��
"��'����|�>�8�+Td�>U���Q�˴��pZ�Z�FPb�F����;iJ�%��h�Q�#H�s��­S-�dW�����;	|�s��C����6̵�Ff�&�� �~���Kǫg�U��7xv&�kN"���A��l-&�D�+�W�l�zY2�d���"_ �>�����g�d�=���������������1,�:Z
qʕ�݀#�pv*���Ew��=\t�Цi94r*��r��DPޮ��Ad�S;��FcH�Y�)�Q
���9����.�B���{���B�d�h��I
vB��<� �LKz�����p՘7N�yӛ5����램@�l����"�A[g��k���nr�<�C÷f�d4ˈ�+�4i�a�M��l��ЃZ�+��s�ܞC|���1�'�x����
�����U�겭ei~�o�i�|)����2�h�h��>v�ȍ��lzi{����5d��9~�-�M��
kW�o&��^�6���+��`PC��?��:�P��+��d|��љw��~��?�洹�CB�nE熝�ֶ����Ͳ��_6;�f������{�<�u/�ioR��f1"�L*TZ�$&�*��C��u楺W���^r8aZ5�-��~�HQ�x����Vί^ /2�����=�;�B��� ~��4���$�8X41�> ��멻���B>����TEHQcIҾ(�$:�xӥ1x��s�n"�TܚH;�Q<6b��Z�e�>��?�z�O]AbKf�GK���E�rB�<ٮ#!9��J�*<a�yi�-���pB���[*D�����EPd�ۢ>3��5�-��*��4�]�a���7�H�*l���������L9��x"4��W8���,��5��A���Y�A�K:J�h]R��c��.8M��jQ��%��#hK���+��G�]�����
�E<�	�K��f�M���^:�9K�u;O� �*]��c�)�TS�x5VM����J�ݮ�jnV0N�s��A~���^ʈ����w�ڀ>�~ V���T�s�����屗�-�.����ڶ�������j��6uO��F�1:��7{�sۚ�T�\���D/�<o�g��L��Y�ʂY�3O�	V�'����*�`� ��&T�����`�-͏}x�y̧� �����6�2��EA���n>9]t�/��O���zW��;S���p��j}��3�@^�q,�C����dGĂ�����Py���^�������y�_g̬a?T'ɳ�!,�w�ٻ�o^��&k���򗯩�s�&�5*G)�����C㴀����s�J���0Pg�Xw4���~W�c�v.����h��x�l�.�~'�	wb������u���	sx@g�V�
O)� �5\���/�S��pv�����w�Bҳm0��a�{$�v�!i����5��'5D7� YF ?�\�y�N���!�$4�`&� ��*���(Z�Y�YC;<�E�O�s 2u� 5T�~�.yL����*�N�i
J�tU����ѼM4j�l��D�O�.�K Tg�0&|�'�pT��7�i(a����9�9Q���p�����[�^�/�J���/ev��+�!0~�:�5i��(q'���4�|�.�5��+�Dxؠ����Eg��/)��d�!W�n�aV�T-t�A#-ة���ء����E�J��P�q���S��.��`��k�$��*�D �Zk�mo!��OQ�Z�?s�Qi��O�*�`�k�C3��r���t�zmj�C8}> ��ܶ,�팣)�Ȕ�!������Y�	]q������� �h���M66�MkM'{.���& ��e�U�{q�i�g�x}�ol���q�#s:�?��������&5�4�_J�I�e+��;�lw(��r������ s4P�m��%��ݡ�{��"�E��)�.|{IEzB2"uF���b�i�f���K�����o��ޯWpU~UT��m�) j����kzx��R����,g�&f���cZ5n�_�48Pي*�������XX�92�7��cbo҄
��Q��H�l	��Ȱ,���x�P��n<�}ѩ7P�t�X�0ÎI?���s��,p���^�3&�?L�~��_㷍ʁ�Ko��e8nN��+A�P��OON�a)#e �����!J\M���><�_��%���QY��g� ��R,? ���J+T9��]� �5��mXsN�
��pl�`0kE��X��bV��s���]�>bS��|�{_U:l�ߦU�vA��kN�'B���ST\V�
����H���F/�U��
@ _L�	�S�òy֘
�S�����^��d��6]ά=��H�ǭ�ʐj01��^|Lk���=Mgt�X�H�Sޏ�w"�b�q}S��}@�@�T,�lR��]'_(�m�X�^]����F3܇��p pV�4כF,@B�m4,^�D���^N��b+%P\M#w�F�@\�g����݅�`?݊Y�1t�����U[&�(����+ɬH�[���jg�� �����x)��*m��c��e`k���x�������=(�.yp4��?6�agey��68w~�5$z�uU�@E�7jH%�Z�ӹ����!��q��H�]��XT�ڲf{��?	���	Ȗ��nx[
$-Z�1v��ޔ�@���P�ڣ >7A$��뛲]H����:���7�x�>ȓ�X�uO�Iι/o��Z�C�2U����ED�%�e5��6�E���GZDi�ְQ���<��4��p5�)P�V�ob��˶U m��~v t4�O2u.�k��YoBsJ����T	�\4�4�Pޟ�¼t̍YWFA�HoY'͚��6���8�^(�u��5�axa��=^X[�m�/WF]Fӕ(:"w���3��Աl�%MF�X�����;���o�J��	�H��s`p��L�tL�e�\g�q��r�� )Y���+��{5gUp��;o�}a݌p��Yƍ�e���M�G,�j#�HW��v��+�.?"���0����R���x�X�s����X,0��\���S*Ǡ.��vo�!V]��"�[=�ФQt�6�V��Iń�o7�+�t��3|��-�B�]H��S�v�jD��v�8���Q��1K��� 3����Ϟ���oz!��H�D��H�L�ѭ��h���2�`2�IPQqe����ogjw�^�4�6 � )�WF� ���ᓀ�� �=I�ԼŇ�!uڭ��Z$4MD^�2{��܄o��$f��1m��c��͉z1H��\��_m������x�=�0N��ט2L���V�`�����}����h	y �}��K��J؉u��6�s��\�Q{�m⻂f�ȵ�qFG(¡)��1�Q�t49�KHc&���!�R��j�F��U$�����$��͹���d�$��0>]�&��/����攝C�;���@Y<�^�W݂"����f�� !.�g`���߻'�
tT���������D.v{)�yt�>�M��Ɗ���Rc���4̸k���f�:'��"D�1x��9&r��%E�ޔC�%�}B8��6����U��uŴ5�����
z:��r�Q�gOAZ�	?��1��W��3�(�q�Q��cx�'>�y�� )-�h��
a���UX5�!�\��h��7MC�F����{��i�2�D]�"����	��VWb���-�Z.��9���|��:,�QJ����S�q��8۬��(^t:n�r�n=���n�h���z�� 4�'F�A�Vb�R�!){�v�!H���0l7� ��T��wb������R���7���K&�ϴ�y��m�3_b��zF�y������l��{xl0�B���+w2�q����A[R
��J10c��Gt�f�?V�r����g��]��W��
O;��� ��kꁅ/|#M�>�̉�i�bl��f���{@�	|��:tg�80�(台?�׃�F~X{�"2�qj��q�7��af\� �\�U5#^ѺW!�K[�lݝ��������L�Ƶ��lWm(wM�d�"/�?���{��pZ�e�t��񫻵o���QAy�t&��G7'L�)E�g��Vb�U2/Wˁ���Uҩ�����9�`����!� �(t��ݗ��Cf]��,��k�����K�Ӈ�����%x�ԙ��6��|���.6�0T.J���S��+�-z�<AX� ���N����+t�{h�Y�&����pA�Z�U�/
"ːx��e��H��bW�'-u~N�@����8��#�0;2w�� 9ݷ������~��iR'�j� Åhf1�&g��joiw��L�5�����Ǆ�%R��ءPj<z&�弊�,N�-cfD�a���P���:3���,�K�;��� 3�0�DR�D' ��V�Ol�Ե�m���{\����d�X�]�_���桶?�>ƨ�šL�R*��5��@��טpU�?�wn�*�h�i2b-��FXѲ lD3��e^b��s�oZkz!�hk�Ֆˏbʳ��9c���3M4/�����|�����f�7lU�k�d���>����$)q�����Z;���?���~O������������c��^V��Ӻ����:~	�%����ēض�O�V����r.0�!h�_���7.��w�S�����&.K9a�X�j�x�//��rQL�U�@:'�ǹ^�P�/�E����oI\i�۝�wa��dv��Z2 �f��A{h�"���n��8��� �9r"�2?P�M[P�
M,�7?S-$G����Y��}��	?�ȥ��Cso�,��a������8HB�e)�H���x�A��k�#Y���I�\�b�T��o�qS�q�@�k�4�B�)6+�
��$1�Ѳ@!G&�05�q����e`�Ǿ�{�m�J:��	�GdW�:f��i�d�Sߟp������!��XNWZ; ��ӕ˳57�kX��t���8D���Q0;aL�q�T�������P��u�꒎@kJ�7$���X4�����a6J���/ѡ+a�U��=ηv�)��־&1&Wx$r�Jٕ��r���q�o��[�X�WQ��*�g=B�5Cv7���>�#��:�0`(ª�`(̍��v>��n�Q��f&8���3ኔ��P�R��\��,�g�����a� ���&�����Q!x�t�:��O'���a)�����$	JZ�Zш�}t�� G�$�z�ܬ,Y��3?~`��1vu�Ա��V]�\�5�D{KD�5�s1�Rv����d��Ϛ��d�0�(<���B,h^:g./�ha��Ľ�Uuh�ݚ@�h���.����x��/d/���m_hj���Q�(�����X~�eW?/5YN׊�T�"=��vS��;�-��_�f��*9�ڲ�2ti�u�2Q1�r;p��3}O�eX1�q̊�s��74�?�Ӹ|���P��;�&���ߝ<OJo鴝*�6��%����@����c�=�[�=3B6�(�K�dk��[�i�ޤnHb�6�&af�I���e��?,lj���r��fdV����.���&���)�Y���E,�k'��H@Յ�2u����G���M�LR��Y����N6}Yl��c&n�Z����K��b}U�G�E��"T�m��6҃�wnr!j�ocI��K�g�
�l�Z}����B~�j��ѓ���ק��
gW�k�:7�<5���e�b�Ypz��t#�P�ͨ�K�;�w���k��/�a�Ө�WHS�E�=U�J���Y�|͜�d�"ڑU��H����$�n3G��@�sI	)_�#Ƭ@Lz��B��Ok1\���@�F�S�j���5)7nj\��Ai�Ņn<�&P;Ů?��,�d�v���8IX������C���h�(�/�p�JNbϨJ�t�.b�v�8u�e�Q���@@z漈�c�qk�
*\�`�p���:�\|ϙ6D��+0)6҉�@ O��Y*r�\dfJC�;��C����?H�V��6�9)%M�M�Ƹ1��=v-|E�L��1��t�>�w�7��?A��~����W�� cmkC�鱭j�s��wQ!��c��炟d���b�ݕ��7��s���Գ��ۑ�T��E[8��@fg���[�J�a��=�O��q@��7�����cHv��z�}Ū��u��G���j�.�A#x����!�����r/!�@y��0��Lo��W;���<.�|�Kի�x�h y�e���+�؝�*�R�"V�#�p��Pf�>��q	�=��yL�2�@%�A�ݞ��=���D!�%�(��7�(�J��5)/7m���Xg#�U���pc7����#�t���$$jנ9Cױ��i]G���6x�KM�����j:��:��9	�ĺ�sQVW�Щ��@JY_o�������Y10�{�;<�v�W~��;U�0�؃�N���cv2�Bh��,��f����"���5�a_�d@�\i� �i�}�7�܄�<�������8� ��\�W�Տ�(�Ƭ�:��S�p
~���.�2w��N�Q3�V�����cܳ�a��G8�\=���'X�T����O�a���M�pGn`�)��i&��ݻd����X�i�K�I�l(6bI:�?b���R̟���!��\�4���%�6Vj�T����Ʋ!"�:: ���>�	:j%�=�Cm�J�3�����Nô�7ځ��DǬT���7�u\��T�⌊���o�K3MqB��U��cp����{��1�O���Z���iY��6uٌho��LԘ���Ly�J�$����T��w�;\��XD'�����xn%l`,��X�ٯ"�]=}�z8&���]��/U�|x�v�1M=�A�<51<j��mA!��������G�` S�1Fl�Lc��4�����~�h3fʢ{%�HD/��v(YuHZ��F�����KI��<o"]�q�2����qu=T��Z7Ϻ�P�xW�{�ni^����S^+j#@\����!f��#U+�R*=��Nl�u�/���:2V�x�##��@}�U��1�	��n���w���}̌����5,o:J
�����M�-��3�aj?(]H�#��h*"��`ː���@Z`�U�,�[yO��<�d��6�'=�Hpؔ'|�E��V7�0;L�do!�2 2��n�sC^�����L�D� �"�������A�5$ +*3C^���s������Y�)Y�`�����iO����;:O	���՝^"����L�.Prո�H�6��*S�	�Cp�L��ʖ�z
�s�}[!��TyEp��,�zXB��a�I��l�LZ�1r#���L��9���^�ፏc��8�%i�d&����՜�
��3鲼��w�XDVpsY���v�W���c*@ݛ?��;�XU8���bl� ��ӧC$T�"B�f�b��%p���|�P�Go��[�!}�
��R/1���l���1E��ּ7�ז���4���p�I\.�h�{"V9
k����|~��
����(�:�i���T���}|pR=B�b�O���9��yT�p �}��A
#�A^��C(R�#ߛ �I	�2j�A�s8��o��U����'��O8p#��TM��d�]񑛫b��H�a?�ç�1*c����Z���U��{�	CW���(��v1�f9^�[����p"���R1*��P���m׏*O�C�]Y��}#r3�CY/�w �?�_K��HI�ts��g���i] ��Of��a�&�JG���8e�Ƴ�!����$ ����͎��&h������ù�� ���bfoL"]ΐ 7��U��(聡���fW��/�'�m�ʻ)C��	�?����Q��	�i1z��^N�J��䛁����y��!�u�*�P2L!CC��Y*6�c~,���]Y~{��v����b�=��?yi��y�&�Jd숙o|I�שa��:��������E%/l���BB*�#��p�H0 Y=���]�\�tWD�9�"���Z��"*JHu��)a�!���=D����?i�p�q	c�>9Bg��������Tg'Z܏<ED�
���!_�E�xٸ�L�2D�2�xz�Sг̥jM㫮] �c�߼�X��䟃_d;^ց�P2{��u´��qp��OwN���������Ϲ,x�p��q��?�0��1���a�����F�A/ɱ=����5�$��nB[��'O �b+�y�D�os�w�ݴL��?�p��3�Ns��P3S���e�P�e���2�iD�ӭ�8�-T��<��y�Y������0>g�0�pT����J/��ڴ0�'��f�ɭ�s˾��2Xb������G�G�#�Itr�?���x�&Y��%x|��)��XF�f��z]ikG>���K;�-�� �����Y���-�ط�oL���R<ݝ/�e���)2��رJ�
y2�Z�d�@7ATwx[�h'��R2��@�����p����8�v��̤ؕp_d<-R�|�|�õj�2, �Y������b�%�!��!"+hӽ�|�'nۦ[���e�ɫ�i����6\�������zPѷ�1ێ88����Cڇ	m�{�V�N�t�b�} *��j�}�A��=������;�?ɇ��;7P%��s2������3Z���J�ר��	�F�'�Y����)��&��&�V�N�� ��W[̖�L�B�^��q���R��N������e½�՝+�*襶A�p��ҵ��up=i���g,���F}ޠ�����)_�4{�)A�?���T�B^�L�*D��xE)��KE����Q�65M9{^�la\;�]��YW,4��A�
U0�L�w�T��f��z�U�'c�*���x�h���,{g���}�N�΋>��)X�Z�|;���9װܤ�^�(�\{
��߼d.��.�^4{��)S}LY7���u(�������d���T��K{B�����k�l�D�X�����8ue�m���ڋ�¡p���Ш����f?�Ɯ�$9�� ���6�^�(ip!��g/���춂��j��i�:!��XV*����j�4L�εP?�qm(ItG�E�t�By����8���U�I�w
B�������u/2 c7]6� ���`����ӷ�g�5�zVx<6n}jW�>�R���|����f����Yh�x�_�T$yJa���5b�k�i�<����ޡ�[Kο9�@��T"&���$]z�/�y�~�r�^��ה��ڋ�r76������[��f,��5�m ��߻�U?�}.GZ��"�a �L��?��U�>)��/�C��X��nZ�]�r(�G��j�G(�\;��j-_=n�sE$���1&�� l�].�*�S��Z����2� {<�ͪ��a�+h{����܂�yZ:�d��b�˿�$"�i_�h�:�DYml������JŻ/���%����O������u�dOh%�/��t{x�ē����3�������ΰV�Ps`:�7�}�v-�p�Ԩ���$��$*i5�Q�)�U���S.)Ge�R���q� Rd�:���dC �=k��u{�/jU(��=F�g�\�ۉ��޸���V�2 >C�~;
�$J��������jz����޽.�i+�i,�/�������Z�B{�#4�Xc��v9:O�������t�c�:P�aum(�ިa����7���%�E�Uu�]P����*�/�`t���׻�����:|ё�Ϗ��tFL��X��/y%J��U�$��֬U 0��WҀ��{��?
Ȳ��U��w�mDED��@A��os��/����I�A�O�!���nv�}�m���2+�ו �p=,��&CsG�?U<��o�����)�Gǰmo0*�(�C�I��	�����#�b�X"w�w~��"F�J����l�h��5{�'|�}����/��v�$>(�n��l*�^M���35�n�x��=�3j�4c�_R���&�h���	[`d�`��!��Z�$��_��}�W?�T�D����zCz���9{Ԙ�W�du�GvՅEyR��	�//�J y`�K׉�*����3��`iV�����k��&�ol|F ��ry��ޚ��g���5k��L%Xgs�ye��q�Z_�)�b��:�la���d	Q�;լ#	wA�z@� ~+�N?�P)�uKf�z:��dM �N��`n�sf;?�㻎��	�[�	ji�($lf�E����K}�D�ޒ�h+ɷ��+�w��[���u��Cu���d) �T7@������O01�ˈ)��oG�2��b�{5�Q@V��B��sX�z��/��(hO��fo�l��P��s�%��94�ܐڕ��ho�:���(!�A˟�+&�'���9��O[o�'V6Tj�x�kUs�Z�����*:�<7t�ć�D9�����]]w��L��u�"vJ�/A�Vޏ�;�M��Y	��<��9�	7�V.���^?e��� 9��>��z�E�un����n�'�7	a)�����1T>��%��`��zH��� �t��$��7�L)	9�c�Bd���ј����k�Y��������&h	
���� �փ3n��kQ-<g'w�)�BVie�6N|4Q�A�HB��ip �|�Q��D&�{y�3�gt��w{��9�@�����������9���4��I�g�e ��C�����x��� �`�q���Ǹr!\ �6�ɰ;��W=H��[Ug�y�O�lWav��^|�-G�f_��} ��^eEr~ČfA�ր�8����:�g���	ڨn�w�:��O�n�_}�0�KY�1�P�k�����ib9��jtf��=���)���ٌ��2�, v8T�����Sb#�aT��!���٦@}�m�~�����!�IA�c��-e�xN&�:�q���%�I!T(
]�t�
27K�b/��X�32d��q�I;��Z�ǟ�Y��3E�����K��[������H]P�`̌#&�c*01�����o�rX��-?�����o�����S�1�)Ӣt��P�헊7C3��i�����rD��=F����h[?3��7�T�)Jt��'s��7�M��[�K�zl��� ��36>��Sً��E��\���oO��9=��q�7H�kȿ�sD�}F�I!*Ul]9���E}�Ǖ �-"���`]��X�i*��S>�N�6�����I}����^�ㄲW6�@"�T��ȹ������ݸ��}��iKL֡��� �G2 @�̬�❔��E#M���I�4�U&�o�X����F��Xf#����Z��/�c�|�]������2�u��q�T�T�[��k#��8;-�{C���������<����D�Xb��I�,@G�|�I\थ.?s���K��SY�z�);-������o�At��ҮDM�;�J�gK-Fh��66ޖ�S-_�6�}@*+i["�Ey�Z���F�]�ۺcki�d�/y�.����;���j�'.���<�OP�b�_�:p�B+���퇧o��*�/&��\�C�����@�Õ��QT��{VGFG�|��C��L��ҳp�V���ގ~����ȾN}5QA����D׉@\|�r��F��}��Q�5̞+�Α&庯V���K�"Z ���0S�Чy!��"\�CF������V'��۔��k_�u3�(�SmUk¼��,���4h	 s��=�^��p�;���T�/�S>l���n��F�	eY� Q.^^���������b��4�����<G;�z�X��c�UM��ObUk �+�E��un���Rgl�&�V[<�u_V}���`�<Q�^4	s(�D�W�V:����J-�eB:~�8�*;����{ͱ�jLs�QLM1r�n"y$���L��h��������߰�x���Q�s�V�Lq�.�TL�	B�㪟���~���(c�p��O$s�����s"}�"d���<��#�^P�6k�3t�"��B��	�S)eAW^>��D�F`�m�Jp	��A�()�$���D�ݳ���bHC]��M�Q
F�޶�S�����!p<�_,ٺYfɕ�{���RYR�9���ӹW`A�uO�ꟽ����`�7�7T���J!��Inv�mw�k?�zo�&0��'?���ٔ��~r���>��X�b������1Р��I�9�O�Y77��(doyQ`������0��h��43�����s��G�R�(���I�b;��H�Q�l*�N���k�&��ՒkA�{�,�OM{Ѻ.�k�W8_���b�~�uP��A"0 �I���HA4(�ҭ��x�i�b"\yԁ������������c��o��M�~9P��_�L�n�<X��s�앋D�"g�S���$B����dv�?�j^$�&D>�0�%�w�����?���f�ڗ�Z�T[7��>W�r|���2	Z;:�?m��
�!�1�k���C�����J�ʀ���۲�}C��	���9�؅mVl���F7��� =n��{��������AE��P�������R]�s�5v�ib�3D�KH<XG�)RiS�:����PA�H8f���gt�5�S���x&"�#�B��ng���5�:#f�|��^7�_�+������:���k���4ҋi��(���t-���kfK�� ���d�2�o{�b�9�����ȋ�[kͮ9�
ibN�m���/��Qy�˾��%m��]�~Ј�.G�q���ds>p����Aj��n�i���"���R��(����i����T�s��
�3N�$��G�˻r�����Y�9�q����Z�Y-�)��ՉA��b��뫇z\nM�~+�r���>��Q��Qdߵ;�'���/�վ`�1TDjt:�p[q��pq�g�����ǈ_��xC!���>/#b" ����G���/��T��z�P�s��SO�`�O�n��ة�T��b�ڭv:�[�`��d�C0��YN��,�1�^ST��ECc����ǒ��e9G���2�/y�M��F��=Zy�gU�X[\�����cGX����&o���S+�.��,\PRaS2CT@$R��<��dzC4��S��PfJTo$I�
�V��u�2�:�Ў� �N� ��2B��"q�  \�\p@�B��78u+ͩ{�R�2�|�%��;��᛻�xM������̯�ȒbA�O�h���6!��
z�_)�_�!P�;- Uq�i�'y-���Нp�ღ� �`�9�h7��t����9�5ef9��)�0��!�F���Xd�;�����j�3{�����n:���^�Ce!+����U&��i�����L���	f�u= �(2g��GFa@U��R��G��C[�ad8/�֮�Ԡe�ƐsNS͞����`�6zhӑp���ɭ�F.�N &t"H��ðh���ߥQ���f<�Q��)���2јo�,[�-wf�K(�	�*0$G<|�tk�jf�5S�[W}�#&hcF�mb�Эݙ�U�7���Y��#�:�M$#��-�S��0!��韞1Q�����.���0ϗ(G��1��aș�U�s�L�݂6�/5�4�.l�锜��b��������j-c9ڪ�x�~hS�_�C�oί�"�[�r&�Re��p6y�J})QUM}"�����|^m)��K���C3�!��4i2�*[��?%T$�e*f�%^�x�eP��uW��U3F����:w����R��O�:�TΫFn%���)5�_�3�����2��O�i�Vδ�l�%�����8�ܷo�j>�T{SJྰP��|�c�� y���:�F�\1.Sԟ�W��m\��cf�vF�6�Z8_���z�:
?]]Ӏh�*�Ǚ�r��['�5<o�ZV��TM���7�����`��v��.�EޥP�TLHOoz����dL[L�dFՎ?��
z+��;|cz��["S﬛��Y����r���"�{�u��T��������	hC�&���P�5�)�����#m�N����ɋ#�'��ʲ0h����D�jS�	I�4-[6���w� 
gb�Xg#e�x���m�������NgX>�P�%9�w"�/�I���?��j��]���*C�Uk�6z��.c��N���K�̖������n��������s�ڍ��A�;ك�����|J�U��U�g��F0�&�&-X� �x	�V\ŗ�V,:X�.�����̓����yzBK���B�o�{�6o�5K1ߎ�߅)&�I ��x%�:fs��%��g��Ԭ2B��Zz�j�j���<r��c���>{ �Y�����t�����x�w:� ����kt7m�a��uH�g�T|���T����v,��Q��U�Z�3xȾ���0m�_�`8���s沚�G)�yԈ&#�G��N㾗�p�c��\�H�\bm��2z�y�S	,����b:��+������_���×k���lҔQ;,���%��q�n�ƞk��5�P�D��d�B�Fc�$M��V+�R3Po�vN ���w�ù����Ys`�iC㊖0Ck�O���,Q3�D#xP q�.���TK��"4*F�=����	\�Aa�"�z�Z�ĀLsOU�h������g�cW��2/n��w������h6�F(�MK/��洤��E�b6a���{���0WnDY��"U�%k������<�m�_J]b9�&�k�k�ăiT�Dg�M�Ap�/���#ұ�����@�7?�`�ix��耻-gAQ�n��#��`��ҋ/��D;��9�91B[9�A�Ac���뱏���6�]��	Aki`�)�����o�Î������Iˏ앁�5A  D��	���@$[/>I�'#�4���`T��6	*��j֦x_<�?o|��u��4��i\%��$���H1�%c��S�5>b����)��s���å�[�+%�2�&/ɨHn�5�ϸy)�Qs�=p��c�.�����6�?�<�JݽX���w�_T��&��ۍ�`�[:��DD������ԥ�� y��V�g:��iW?E`.��������R���av�p�-ҫ��u�Hf��";}�e!8��Z:�䱭��#Y���z��2tWڧ�߅��r�t��k�,i���)6�B�惲�w��\��8P{)�� �+J[a�c��i�oҔ�ǒy.��%�Ӊ*hv���-9@[�O�շ���i�c2��(�B�$f���_9]L�-JÃK�X�*M����[�&�C��R�|UZ���[�-[ˈ S��A����p�>]�+'���r����+�a��8�nmU
|I�T����K��aJiVKĈ�|�aN=-�����G�2A���W���0~�-���������+ڝCI5��r���8vKa*A�}��w�>u��ġ��xPJؖ�s�*�O^�xq�	�*���OAx<����ظ"6�/6�,H2$�<Ƭ�Nv yOj�����?{���po��lcd`)��O�w�}����>��E8^_�_���-�Z��T郤��	���������)��'/��:a�z�n-�qv۴��ؠ���G�`%��1-긤 PO�;�>���[�a���ti��ڋ!3�	h�-���\A��[:�O�i�,�i���]�6T�D��][iw�6�2�U�����1ˇZ܃
(�HV�,�?����,;�H��k?*���6�?W�cGS��	/l(u�\0�W}�3Td�;��q�C���z���&��E!i����#��뜪]����fOo����l��s7|��+ZUyf�q8�$����@]�*�No�ueЀ�᡺K��{��	���b=^�2�%Ĉ���ᅿՁ��GtWSR��ao� _LwL멶�MȬ������q1�ݹ��p��7�e(G��@�P��b�V�e��统�2��!�����nr�YnV�*]R��������1Px+yȯ�<➬ �=2>$�c�S,Ӛ���T�pJy��R�j5z�(��%��su��n2:d����d���,}A�U�I�)�6��C�f�n��?�3>�<�9�-Yp��\5�:��܌���ǝy��c�NB���f9}8����x���58�����!��O.PB��H�otb�4@��ǝ�U`�9̲FcQ�UW�a�"���ܶ���@�5��:���R
Ȟ�n�2 o�kc�$t�R��V��Ћ�&.�q4ij���/q:U��Y֥���T�xg�Ѳ��"�ͽ�M���;[��4M�*E:��,��Ҥ���%�@���̇3ltq"  ��<9�8Y���k���;��I��Q~�͡�G����잀�s�Ō�H"?x�
gs�e�����V�/�}��dv`^���݅Ē���a�r1䙣�!	ZP�ݶ9ۺ��Vp�ʴd%�-�d ��#\2�m�dX+���+,��{�ԄPݡ쁹��q��xo��@����CT��g������S������`�dB�~!��#c����q�=JJ'-����xg�.fJ�4��J�0�|i*���g5L��w�ק kI�ŜX�T���1�|��5�B�u�˂�rB�iЀ�pg�dJ��^�8P�B�N_���I��L{�g�@�Fo#ad�/D���p�y�Cũ�s�Ps������YB�
��;ؗ�5,Y?F��v��̦�]�F���������Z'�?C�$r2�ĒIbg9@������<�o��[ohX�F��vV��aG��K����6��,������6M�~|]G��c�>������ 7,���o7Qfr `��Jb���+�+_��,�>R�h��>~�u��? ����к~����H��ǒ�?Dس��3��D�2A��n��"���T�s9�~�ޙ��o�t3C\��"!�rTn��ޚI�8?:Ki�xw���涖�I4�/��6hOC���H��x� ����7;R��bd����]�<�#t��G����].=~A�vh�J�TX,���H�G9��!y�p4��BȜL�(��� ��#N��&���3�Q�w7�Ku\��O��:�ιA(/��C%x4!����� ���b�((���v>�SXyR'	���ɲϱ���>���ӌ>��[#��MF�.�y`ޮ?o���uuШ�%�h�s�9%���6�����ѭ�Vy����J1-��k����"xD�;ĥ~ ��/����#F!N_?�|2�TC� �D�B&��M�4T���3���tWs	Ѹ�K�9.�b{5�֩�+鶛h�_(�Hh���;�p�,��,H�F���ݨ�������i��<��q�ذ#D�
!X�>�]�Yq�
d�5���J~��?-�g2ϫ,�LJ"\�+��T���G�|N���vm'�䧫����!��E��%��j!���
A�C�����\JR�R����S\^{P\�%.�7�-��@�t��uĹ ���
�OG�^5��1�s�]s?�de�,i{����$�3�TT�W&EV�ꬖ�̖�Z�+r��� G�{� S�P3l��i����ψ9������I�_�%�7���#�(��&��<�[w�2;����g�����b��p� �P��e{)�J��A-I���r�����CSS n*s�)���&e��Kƞ(Qѻ����YL��R�Ȗ?a�:��2Z��!|�4W��	Um�y��y��B"�1Ji^5ג7p��r�޿�<��ߩ�����)��(n���f��ݭ����Rz!��������ֳ1�'�츲��zYQOR	�o>�z�Z]ʅb}Qq� �&p��i�=�W�?�&N����%��5�)���B_��_9�xw�u�A�c��D�������k��g=$�n��(��M�����^�=XC�z�L?���x��������N�� �� �6 A��訬����f�VS�d[F��pT|1����*���?��Iw�w-�@�zÜ�� �e��P�;u���#_"���}-T��k�v��sa;����UpF�2�J�X+�D#^X4���6�&Y�m���]�v��^��=N�rR�j��1�I�f
��~���&�PQ�.�����g����)03��35_�<�N���Y	݆l��>1���_H�J���¢֠����u�N"�t��[���l�	J��>ƴg�C�w��d:�]�X�����f� ���%'X�����**L��v��Ø1��Nn�qyE/�n�^�����D���;q�"K�#׾z��CXh�{\��`��%��X��e�z���g������bI�}�ķ>	5+F���c��3�y�qt]�zi-}B�q�~�3|��zx�NU�pU3�P��/���
:ŢV0 KZ��Nh�~���,��i���e��N�W���nऺ\�(@U�<T=�Z���~H;��>2�n�62�:Y��Z�5��)ׅ#�6��>�3��P�B ��ƫI��AUK�k,Õ��1����/q)tO���'���t�VT��1Sg��
� �{�X�Agؙ�<9��4fU�H ������X�T4u�QRh a',������q"� ��[aŞ�b�H 7�$D�����7�.��}˧���4:�*��I��Z�L�	����_���5���Lg��%�;ń�D Y+�}l&.b�j@3��v_|9>:��������u��D���(�93�J��|�&J6���tÕ��<gC�ƨ��)�>�ۨw��J{]�<�����ߎmj1.Ta��R�PW�M��������5�`����8���e*j����.ш�3��(N����	6=�=O ŵ�?x��mA�A��ï��B0�3�e��b���b�a��c1�0,Zv��[�U����k$^7tq�9,�@�\K0u�D�G�5�3x�E�-d.X^�����}���X�#�se�_bqJ�Xp7T�j�����$zI�H]*�Q��W���wF�y�y.�z�w�=|T^����f��m�%U�pk|#x]�Tmӹ�s-�ដ�������G�z��$�k�w�t�����^d�"-eKR��bzp��
����R�X�9�E��{6�ژ0pBls�y�"e��)�vH���Sk��o����#��ے��>}��څ��J����+�xNǘK�z��b�{, ��O���/A=�$~eoѕ��!ؙ��g�{�r�#��j�`�P6@S�]5��L�y6�&}�I���Z�7�a��L�f�Y���W1ao���v$����l�E" ���O�8Ν%`֢��]��t���,��s�cr��vL�3�������.n�~Ke��ɒ�&���FW~���c=��y��t�B��D������n����%+T��o0ſ�j��F��&x�#�,f��w��^T���{�O�s�ސ���A�۫}������:je`���ܻH;��n�k�U�#��M��R�����O-vV_&��.����x��(��Ԁ95�	��)W��sa]r�A�
n��qH�?��J��H��z�X��2�;.�c'&K1!�(��~���U#��TLQ�e)*d.}O?Α���Oe
�Z.G'Gm��\!ք���J6�S�"(�E���v��-�u��A�/�Y�M-)�6��dmf��[�>���6���aNeWz�,���o��>$��^O�%j���>5�!�r>��Yeȩ�}g)�/����܂0�Y��Z�2�O)f�Ќ6�Be�^4�C�K�y�Q& ;P�d� #����U��/��/ ���E_%�4Ǚf�i��i�]��.���>�U��]���7\�w{j��i�T"��b����y
3����<��?�o�[�胑U���"
��)�="=D7U�ѵM"8$��Ug�$e㬠ٮ:���:K��p�Oo�ɞWzl;���H�-����������n��oD���I �r
�����j��FZ��?<LP\�/fa��w�`�\�eF�<H��Z��-(j��U�һu׳+9�W�SiGݍS�-�>R�?����`��� �����oᨙ�5�i���d�� v��P8�TM$*��6MӇL���V�~�߮��'t$�	�JN�����k�/��&¢����ۤ/!L�4=?>J��I�ڈY%$�i�ʹw萀Ǎ�kՊn/B�3���j�bs�2w��ds�=3i��)zo��|�� ׸���w����F}6ݡ_:��%ᎊ��.$T�hCeq�1�.K^eC�?�I{�ǔ��w��0��ݒiaGr)���ߵ�`Y�&ᮃ6b�+x�,�s5��<dE�N�e��ti��t�Ǥ?��_�r��0_%N3�񊝑�u��m�yH!������m@������;fnC�Q_�Q�߼��k����y|�NöOf_ v������hF���u���f*Z���ǌ�ꗀ�ޠ�Lu2!���6�;��f��L�
1�M$� -q��e�M�E�B���Ҡsù��/��T���� y�;�P���� ��W���ABǦS�*ܵRe�`�����o����_��n~O�CS�o��T�e��3���M~����{J����Q#^r��wYx)S#mVvpr�=) 
�x�{��m��"��EҐ�9r2��;)\����D�
�4r�  ��Q��V1"���<�FH��;t׬��q�b�o�=hh���	�I֪3Z�[��2%`��뤪��(rS��hP��"�3*Wn3��l�<	Ԑ\����r��Ş�(⬸����H��Dmw�����	$����Hw� r��KF������$�@T���:����\^�M�hS#3hrG��,��n�|�.l^�M�.��Ye�R����XLND��V�i���=񾂢��`ɱ�䯃��[�!�}�a�$N��B7�Ig����\ݚ�霕�uŠj/����[zr���R�2X�]v^D@x���K�]îG�&��{�Jq�]<*�T>[9��
ڪ�灯�{�)�ƣ����%��!F���*p�6h�`}S�*8��P���y�	G�$�1����ݢ�0�qL{^��Z��h4��Lk8Lak��dw*�&/�S'��~lUi��]�����O���*��S5p�����Κ��N�Ɖ�f@��q�a��;����FW(���ax��NwW'�w��AOH��^� ����z��87p��Y��0�؍I�BA��*y�\lN�x���ᰅ4o�Ն�{Ƒߠ�\�/�"�/�x��p܊UXT|����{���9��y��ZצX�����x#���EҕD���Q7[��x	�������F�3g�|N�LgCơx{YioD� �uϻ���$l�,g��d��@g�|���>��e��\^�?X]��C�j���.�P�Pc��\�뚩Pd�5��r����_ �5�
*��e�i�ɠ�&rV3GN¹��+_A��36���~�&UtY�2	}�p�f���J�Dt�­ȞS���uL�T��^6\n�I��߬�K�#�{�u��N<�窾�r�5g.�K!7�D�Ujָx��Z�2*�����O�_"�I#e~��2>YY)f�����
z�m�bV�'E��M�:�q{��¨����
Al�"�#3h���V,��xJؗ�l�������5�g�"7�,*!�@�����'��QX�f�=��HZ?fP��c�_�7�&��A������1�y�Gk�L#�24b������g�ƺ."�������~bXd4A@��	Ґw05r��M��B�l�r��]iL��-�p#��v�ɞ{��,qQ8��=9�|���龫Z��-���_+�$�����.��x��<V��c�˺�(B_�y����̘�}�����z�)įr� ��&��$���,E���YQm��cɗQB�+��'�3z<j��\}W8(�3у_R�Ӽ8����5 -���WJ��BJ�x~��sl'v�z�)��p�N33��u�L�׫�@����x��ZÁv��/>]Q�m�Hc|����%�D�S��[^�0��~�i4��P�S���1�tX���|,�E�U0���i(#bع�0���`:o����2�O`X��״��D��W��y+g8��ycq���.�8��qf�+��Pܭ~�gg3�>��� @}��'�GJ�|g��T�z�z4�|�b^���5Kv�i��ڪ��|�҉K�Uw�f�����}֮c�=��n��?��Q^�9_�E�6��������C6��Ɨ�)��q���L��5�)j �As��ߞE���4ko�� 9��hx�H�W���5<נ�|���E�����6.�DgK`��G`�7��n���Rl��hG��IEWn&c@�$x�j��U7�<R{���h�O0R<ې��!�;e�Lg0W�v��A:�'�3k�����Y����k��C@��\��4��0��s�s` �p�u.�`���}u�q^��c�,��/zT6V�s�qQ�sĵ���.����,��z���$��^H��-��I�\��<�O�TC"W��r�闋r�ys�ṳ	5��7/���c�;�Q;RGZ�I��	(���kC��,z	��؆��*zB2U�RE}�-C��\��V9����A�3Y)�?�(tq<�tM��4�N}ӷW��	o�k��_G� � 5��ߎ�]6�lЄ��P��>P}j��E�<�_��$�;�*F���y]̸"R-��&�~��%�PΈ��dY ;F~� ��n�o4�������	E�7T���T��-z���-o�U4������*t{M���b"�YC��a}:1ª�j�Nq^ӟ�:���w�v\���n������r�?ś�x$�r�E��f"���~���4>v�"����~�(v�n�v��6���s7�v�{���_$���)�+]����k6TB&�DT��d?.�Å3'�{�)��o�Qc�Ŕ#�%��A�hf�0�j>e'��O��
c�HӠ�"���tE;誈����W����4|s=o�;��0'��W�n�8��?��E�^�ߦi`�0v>��^	��/���[[�K�R��4A�5ʺd{��
%�����鰋��.~YC���d'�Ϧ�Sslg�üJ��Wp2�rMs���EHIf[��������y���k&9#�>i��0�X�=[˞3F��耦Me��`U��IT�A�{ԨM�1�=K��0= ͵�uQ�n�)�)1<��z6�)���ÁbS^i�.c�H�c@S��e��s����rdݦN��X���O�dzH-�a5C���>�Q���{�� �z��G��gh���gf��9�GNʈ��S�w`zo,�D�>�w�}ψt�Y��ά�-(`����ّ��ˑ`27����1�T��uC�=Lȟ��������F��6�ӣ
�r0���da�+��N��K�lc8�̈́_%���w����x(�U�a��t�f�p9p�G�i��i'm����SD�Kg�d׳��F��K���Ǩ�
F�TA���Zh��8��ua��gZ�\"ʓ`JoޣH��[|7ߛ�遀ǹw�2'[�CJ���{W���$Kg���I��ΰ�������q�z�d���h��4�-�Eo+\��B�ѕ"؁`�Ua�+'�k�������*����8�~�QG�ɖ(��9�n΅�^�{*��U��0i>mZ�*��p�5����*��.��`����1��M���Sc��ɍ��N��^ܐ�1U��A�O��楹���\4hɫխ]RB��ѵL�0Qޤ�(L�m"��ao7�Q>
H�T�d���3P����T�e���VZ�P��Na�6��������G$�r�)|��ے��᧱lz��І��%�W{�_y�y�X��~�+�i��kB����S��^Q"�t�ciLuP�������'���%�q��{��H`��r�M�NA��aY�H��t�y�=t�)Ƿ�1X*>�m8&$=j��&�{�@@���&�Y�@Wc�=X��b��c�D��Woϟ���V�*�n3�%�x[ݮ7�
?���`��-���oV4G��Z�yK��J�#a������f��`�m����,�/d9�2E;u:�xm˙G&o5�x�:�zB������6|Ι>R�M���ԸkB�Q�DR�֋~��ۜ�P��n��%U4��&�BMY[\Һ-'� ��� ��F,�"��;F��q��c'�����A�g�~�g�N�Ǽ�=1�&��e+&��:�~!��V�������QS"��=c�����V[\��î2}աq��;ÁЄ��nHQ��S0a��e�z@�A�����l>dY�ų��*kBt��q2Sd��V�J��L3��=A���&����q,o��6���_�Ls`�H��p��z����钘���k͂�G��p�
�����I���Z�p�-˪( d!n7Ң���>b�8*�M}�H$��A��\�/L4QvBR��eZ�������oߗ�zU�<5q��@HP�x��*|4�X5���R�0�	(�
,~70�s"w�6F�q���+a}oo�;O1�mw<����^n��;{.Op꬞�p^��2 8(l����5��l�V���k�t^�ɠ��Nd;4��#|	+�w#�ʧzwY0�a|y�{]�l���d�O���]�7c*��Jas�Uڪ����D�s5'94�=MJ��:�O��9�g�v�T]_�/:ʖD��=�N�хc�=��4��UW|�.C�և@�a�52�;q�=�w�P8�W�&�,�{��̵)1�Pl�ke�5�DV 3��~;��֚�ջ�V�i�m��{��e�}$@�P/�D���)$���t��T)��H��P9���\��}��,1�' �����$~�ZU����kcM~������I)�����jXIЭ�+���n� ��Lǡ����	{ƿ���:��+z�<g)��P��1��c� �i�2����}KA�Bf���w::廸2�/dG6n��O��"c���AA�@���{�:��F�B�ԣ?NW��6�Ļݺ[���K�l�4R��	�v��"oT��_ՈbH�
��c��*
'��9��8H]!Qk������2�c�q��T�=.��*�n�z��_�y���[��)|���L+��I�_���X�z@�?b��od�-Z�a���2V��g�����5αg�����!aѳM��Zi��ʃ��m}:|���θ�K� #Z�����P��ꓕ�jf���Я`��I)3��zA����Mza{px���vZ�qX5�Fd�R��Ca��xr<�S���l���6�;X6��/o����5��J��-��R�����j�÷�gV	���������O;:"�MQ��U�8�{I1(Eà� *QR?�S�X'��c��T��������	f��:�W�>�Hϗh�{B�;�K�Rf�$��M谫�Qo؂߱ ��P��߫>�<�ו��@+kl�P����EU��>�G�Z��}g(����GH�ٹ9<1[$��X h��*�IY��C$��k��S�&c��o�]q^MF�k`)~a�K��Rj�����E�+�0��4zԳr��b�w�����@�_��F���~l�'Wڵ�*��R�N�J=��Bn��Q�q�ȑ�q��=]W��ka���1����Ph��4�BD�`����?���+2u�0�E�X�������$]:?�@bn�����)�Y��:�ᩂm8�h�H�8F�4p�
���� 2��$_��H�|���'%�2���3�5�vR����]��¾�1*�>��!�-v��a�2����\qX�i�=d�����8H��(�g��:w����2 �VK<�ɕ���{�!�����zjݱ�)�vV���@��;�`~GJ��@�PĠ_{��G���	�{s���%��xՌ��ö���rm�vrY��>z�ψ8�)������<
;�}�q�#�qʍ!���G����D^L�R'�ܠ\z�R̡�+�"�8��H�,f˚WC2ŀ����_�]V.EP^>$��l6ځ��X��}��C�r���$���	E�tq��C�W�_���Fm��^�x�tSg�wUWbĕDV�S\D��}���ͅ:��"E�,�y�;���;�AԬڇ鬝�O)�ތv���w/ˉST!1�jѺB�K{Bȓ�5�X)��K��RǬ�@dcdkk��>Y�K���#1 /���~��tsr�d�9${ �F�o���:6
���䢝F�H%z�5L�� ���WÇ���ϙ0�i���p�~rK�Kr�ܱ�5�W�E{�2x�lā����8-T6�5x/%FU`������o���h �������M{-�����c�ԑE���"�VM�(Ȯ�Z���I@�3�^�w���~4W��f��J>�C�EQ��@&+93�4�r����G���$����z)L:�:�%O�����f�dY��H�v�:�xH�~y?�s-�F�&ȍ��E��-��-� �����g��ԓ���m9F�e�dS�`�V3���XH�����;�Q)�[���#pg)a��6��p�2�v�C����
��	x�j5�q�S�3��|ZLI�e��o+p��7޶�@�_?��sh��.��!�.���ɑmO�y�~��c�@R7I(b���.�N#�B&#���@�AR� p��-]�8�Ze~��E:�1,�Qݎ�gT5��lQn��A.TG�,Z:6��Jr5���<����{q��θ�
��4�D�1B�!��~��c�����q�DiL�[��s[cQ �uz�\|������Y.�=��df#$m:�7��!M���FJV7�^��}f�k�b*O\ysW�]���~t3�����]K\���y�/�R���+���[}�u^�_�HΫ���C wm P�^�Ti^{&j�0
��D�J��<_/�.�KQ,,�aG���B|i�ĺ\$N�!�^�6Ҍ�I��0����/y�j��1�+r&�@/�K(�b�J�U����{d���q�rD��e�:$�9ʴ%c*fc��"O�%-� �,*�-8��By��	C'F���#cC]���Kf�ɼ$��I2#��P����A)'�1#�G�u�)�w��^0$�d�� �_�>��԰t*¸c�mQ�/rMǊ��CA5�c���Mi�.�N�:�(����!��)R8��W+�*no����V<_�)t��B����d-�@^�����)�~3���8~�:��� �8gHn
��&�,��/�{�)ݱ<T`����K��6��H/0*�ahȥ�&=�8�P��Bj]�7c�� K���2��dOt=�S�T_A���sjK�Odv��"j�ejz��ҝG���Es����,��v�dn���%��CEO��9V�J�v9[bJ9G���n�����v8J�٘��~��{��t&x�`{nJ��c�>;�/py��S�8�Qa���s��3 �����
���o#��1�]N7<ʞ�/�#G\@���+��?��+%
�l~L�pAe��;\�J���3��(����@o[Ӧk+Iz�������CZgvqme='������򂞣;�ۣ�����6u�l��t	W"�YY�_iQ'��8�������=o�^@u(s޺L^�%9oQgb�of��p���q�r�Ի�.�.m�%���aa��Z�S/S:�Zݠ�� ������(��]�GBʮ���*��V��s�[�Ɗ 	�E7��F�ʗ���#bCS$�D,�<��E��KG���I|e���� ~��Z�z���$����EA�(.����4�r��Hu��ɉ�h�s�ȕ?�U��Q Tf�Z[[�fzA9���H4,�E��a��(�C�Ⱥ�-{)��.���&Ȥ�/wW<߶�V�|��vF�Mku�n��|Jr�q�U�D�����㣼�ﲹ�����U\c)|dXj��`��iV*
�h�'��n�D��h����Ǥ��.ɜ B���K��9��i��L~x��-�:}�I#&��&ji��Z��	�<�Ǳ�@���<8������}Ke���<�k0<�hCtS�a�w.�MM]���T;�[��n`זGz���k�$���(Íڑ�[(q���fք�C��װ~4}C��ޥ7i�v�֠N�'xc7�V��rE#����H�v+D��.�sm�2,2�����z�
�*��~A ��i�>�;,�Z�0�J�r���r����:&]�wՖ���N% ?�B�L�D�B�%��VYΜ�~���ˇ1*	c#E~a=r?h�dW`�F����j�K�R]$K6ӕ,0����
F�AɄ��
�ӞV	�l�j�n|����1��}����[i�ʡ�m��s#Z�'��`4&""�Cɺ�,�S�\$�;�I,���cG��UsO�K/��i~��,�/r��.zѩsy���/ 2Y&��7��Rr"�r?�W���{=��4���l4�ff��I�lhG��F^�a=%���X�� #��~$3lM2禷+��	x���I�2b7��nSz҂�u,w t�ML�|�6nj��Pj��L��PݽQ(���Yj��g��~��a2������<:�5�E�`�~�I�3}�.��N�ڐYr�[+��j����<�j���5V{A���VO5���f����#�S��a#��ު��dyת��ա1G"�(���G�3R���`C�3eK5[��I����������=)��҂ޙ7��
�h�X&��Q�E��;Vh�lF	A7<�s��ۺ�qJ�mX�7�X��n߄o�� J��p+�`��^eaMG�a��`B��t�Y��%�7V\�n���R5QeG�	��̼w�ʳ5a��=BC"�0iNբ�woH�N�a�������ku"�ҭ(�ë�MPƐ�V¿��?Z)�n�:���\m7�iÅ���|�}��C��`c�@�Z����:,�T�R;�\�[4��N�Bo7���ӿ�V
�j�[���q;�*��p3����Z���|2��s�6�#r�����s�{��B(�'�4�$�>䷋����a����z�G;�KW���yY�;o|Mߪ95�a���=a
T
������"���(�4CV���z��t�G�q�N��a�	ӳI�7�B����?��]]3�Jy�R	�B)B�ߡ,i��6b~�y�|)�6�k4�����E���������p�wr��-s�T�:�>g���]q��"wQ1
FK����|��w�,������G�����ȲF!��4��n>�2�zǲ�e���
���_
kW`P
��P �U�>+»J���S�����t?۪_�L!^F������Q7q҉|�j��܄�:_��ہ�F豚l�sHM!Dl1nN-�?KB������XȐˡt5�V���:�$����U4f;�ޙNjEO���!��e?[��)�tr͟���Sa`�X}O�L�����{*���Z�t1Q�]b/�$�i�fZ䱱,���V��C\��&� ⭰b��u��}�Yn�d \������^�ň2�:��F�B4�1��1nV۱�b!�z��>�oқ�9}_��x���rWRo��-uf�;�dP{��2��H=�K��;�T��gQ��1���^'�i�B���Ķ=�z�����	,��Ďk������m/��� ]+e�$�}�L�	�*�p-*oQ$�U���;"m��vқ5Q*�q��Qs/�Ug�5���p�*{�As�.7AM� /�n.v�h/�DH�X#>��C��B��o)���<�C#Gx2;����2��E��q��C�	t������v6acj@�cX�r�bVcSk7'��ɯ��>��v�\�#-�S�7����#�
ůw�d���QQ�O=-�3���]��P5�-�u�2R��e����<v������d�*�n�\��M��Lo����y���%"�S�fS���TC	Q�:}��{s���N{�
�u�t�"�S����H���J"8�d<���E�U��l�X�!x��51�ȅ�ms!��9@�4���-����
��\�3�K>?=��f@@N���K���V�WX.�	>�0��0y+픮�+�(���.���`�U.��,��w"`�\�nTX�-[�.�6�%$a|..���S�/�=#�%��|���o�F�8c㙒L���W��N���?�0A�`�G;u5�D�vm��$}�;��*��ng%��E�xi�֊х1��6
��m�4��� �nUK����m��+�A�f8�J����:N�f�w�B�9w�Q˾�$O�;�S���w7&�����t����Q��uQ`�py�(7Y��C#<b�-��P�D<���eKv�x�A�#{H�+'�N("U���>�AlV	�F�*�N��|B�v��#ꞙ���S�BsH^BXNY	k�b�F�;��=��/j��T@ye���.��]bQ���z��5�������/��R% �uG=�ϟNU�2c3�WP����3�
�T�)����BĈA<�U��MUʂ�E���fy1�~�citt�kz�l�V����U2�����Pz n�~�6B�2!$DE0�6�% =1���*O�֓�sމ,�`�?�^�U��9���t6@�u����/��C\"�t�{�}�4���	!S�~?��X� v	�/�����Y��2��--ht+=��b���؋�&��?D<ũ�o@CIb��WSJ�nN��ޤ�'{��9�3�[���חXb��cU�!{�`.4�]��`��<T*��U}�~��8vg���ֹ.����N	1���tH��P�|�\؉��oz���TW���5�2[�\�������LA�%|Yc�����9�����Q��ꂴ�ʶ����UQ���d5C�gr(w�R��Z�l�e,����i~7���"U7� ��#W���"0z]������-���9��a���H-2�I���A��^�\ 
����4�/MXްݚR��T0��^GF�/JL��>�LzO�nؾT��b"k�my�A�D�ZnW�5��*Q������x���WQ+}�#�o������ �����Ȓi-3�y�d�?1(g�e����[%V�>���@6M��=?��0�3�X�>݋ ��u���b=#B�T�.�]�?z��XϢ�}��t
� P���cH�d��%i%�_��D��?�s�%�+,#�����D�rg����s&�+�SU�v�Om�y�Ƨ�|X�N���(���?�luc*�V�!�{��
�$��p(�Z׍����Z��rv;���j�|WJ��Z��M�F�i�*1̭A��]���n�������^0z�F; r�A�O ғj� n��:��8���+��?��s��P>Ad�Cu�:�i�q���N�7����z.��W��4M]�nq��;�Ԕy�i�i7L��jrlv�Ņ�����:S�#�#޶�E�eWd�AS� ƃ�:H%&=S� �&�v����l���C�����4~��Ixh���ю�_x�עG�B=jܬ�9�I�2zÀ�rEn�[�� -H	\���r�R�׊+î˒O�-����/umb����?���a;�����=�pn�u�z��fd�����,��hr���dҹ�qD��?�0-�ȑ�`��/P�G��gNbn���0�"|Cd����3�jk����R�?�֚N�|���K�->cd���)[R�י ��X��}�3����򢌏8�<�M>@�Ac'���&����4��\���P5�Чg:{&}Q�o�I�H�T�4M�
4�B3��O�hf1��l�᪭a�k�y�[�+����Ғ�͕�_Ym퍒�� �t�g�u��>�Y��8��yh'�B�V}�]�./��t����w�V05�ԅ�N-$��s4,�`�ޮ�l���
m0����2I5��KoOc��c�:b;��������Y���J��˵U���p&ce����j}�Nx:�q0�_��9	SJ���R6�Yb&���I��'{'��B����b��^��PO�E1�C}���U�\?Fu1䓭���fb���ȥ�f�T�������	� �9�i�Պ��8?[!��h.���
���3o���rj�/�v��e��+1��8(CXwPa�����-+G_��;p'^�HԘ�A�&kgov_�H2V�CnCʙD�N�����_�-���z�?LY4IJ�������n��l�� ��ΔjЕ�o�1\��ɓ��x�2� �M��9>Z�$�iP Tw�H)��:KP�
�xڔ{�_Nz����� j��m���:�@GO�B6�B����K�ї�o�;�DC��_�$�ց�����Ly��Ϸ�W�=
�0�;
�F�T�,�Y�@��f�D�uZ,��X��B����pqHl̝�#�t�3:�_=GVrY�9g6�#YI^�0x�tT�y��
j�.`6���|��cOî1�Zz�)e�ܦ���� o�4_�����&�M�Ĩ���_y 	���T����0h�M���0AV�ZY,�b��Ԩ�H���O��5��,$`�6U���܊�I�hӡ��-mm�9��]:ϊ�ׇ"	h�+n\E��
���'X��`��N�]/���f[<� ȑ�<���u�*E�N�������o^�܀�U�j9/b]cO�nQ'eB�:�?Tvo��'���� T�Hu��Q ���c��OI�k��Y-��\4MT��QX�ɢ����.���p�ٔ�
��ǠQ=� ��O�{; m� )Ynm�0u���х�������������Ͱďm����a��h�8����'�I|�Z�Xz�7f�e+������h���(�T��bW���ɚ�r9�7��J!~�l�B�
/�?s�y��S0�0��o<O�Rٻ�B���f��g��=���g���wOl���Ǒ���(r�!e��	��H�#��]�{�C� �	���Y�,�8��
)�ѩ	P"U��T�wE"�$2}�{
J��2�G�y�1<i��ωw`&�Z�3!���Y¼��sщ=��^��\�*Z]b�!N�6��u��jc�8&U�qW��Q��b��W2L\.�Q"�����}'6z�D=p,�oDԅH���d�Ĝ���E@/�$.��?pt�:���=w��j|�`r饤Ik� ���|y��,^5D�l����1�����@ґ��<P�0D�%�����Ѐ�#}�$G�;��� M�r�zt���~>����4-+�b��j�����6R��]C���L����ۑ�5�0����y{l�e������Ǧ)�J0�#��~���P�2����5�̍D�j8�Q���%t��c�8��.��[�,��7��Hk2�aLJ�o�U����-)z��5���3L�� �$7f����C����$��T�v1�v�[���lr}`{�5�_a�o��w?223U)&ZcG�{���`������Ou�1v3|�a\��uU�h�B6�2:)����K �˕R��'��1-� ����Bq�|.��Ką�J��4���I!So�4��;��SN�l��;�c���U���0��C�0h3BI�3V�^�I'��y�����eCÀ�"��f��x��U*\Q � ���\;���6s��yJ����1Ս�g+U	[����h\�a�wǣ�|�Þ��OG��'d{���*�n�.�t�,��Rߔ�a\P�>�!$2�̑������x�!��� �ehi�4�H�ߛ���V�Y�;��&��?�jLE�U�����g���P�M��Q@�D�R�Sd��<`Se�	�Yr�)���(@�u-�A���m�����ל؜�R�E}�Ӑb�U�2�N��i=�斯'G�miFy!ƣ�h�W=L�7��AL�QAwpiܦ��fܘu��0�D���eK�-�'�Hf�˰ �)k�y��tH�j0t�H��h��u�k�AQ1l��t�=q>�9s{ԫ4���$��g�uASM�g�(/D񭉈0��,�}��-a���Е1C"+��u�b��:�ԣ���:�ڥVz�d���dh8>xq[(8R��w#�K5hI�Irê��V�0�c.=T��א�?A���M)��<%�U���]H�3���]�6?�8p��Ƨ=lg4^��iw�3��Q�G!8�eQדP֤�
������C���X��K7xgf֎���]��7cl#�3��)p�6�ޒz���b�X��V�L��$���LJ�X'����$rB`���W+�`�<k��\`�ti��Q�W�+jb�Ԋ
��]ݢ��*`��_P�N����������r낤�5����\�m� �k��O-8�a�s���!	2����<\AQ(K��xI��EE9�1��0o݀/�Ő�Q��Č�A����)�+t�:d�'9=!��w��vn��bISv"�Ȫ�"�"Ϳ(/̨��[#��OfVMr8Ǖ�N��Z_��Զ�{�Gv��#�W�r�G���"��4�no��.9�YߥY�Z�)`g5 cV?ij��`���s��
���R�m�8I�7�bx����Ec֏6]�WTGE����w�d��R����U�X�ku��>Al;3,���veBO���[���whj������MQʅ��m��a�*J:'RP���6FL[���p���#�3�t��45
�eF���fGd2��C[;i�� T�c��(�qrة��C��N,k"vDF�,�-9#��}Y��/�-��`��"�,l�L���VW�Z��O��G�vF���!�>��F�ݖ&�>(XB�0S$��ކߋ+ 	�[�Q&(lN�iT�;��q�����J��u�������˕H�"?p��e��&}S��gvbJ|���a�u�c�Ga4�������Y��m�M��¡E9<� �<t��,�7c����@�م�-j$�&Q�遲�����ہt������ռ����.����d~l��a��ɑ��MZѧ�a3����(A��`�A �����u^v�G���&=h>��3�H)�!�s˰#�z��SJ��"�yn�(�)���:B|��l�b.�m:�}M��f�v~r��T�A!jP���V��'8�-�ۑf��և<%Ot���e�H�>7ۖ{R�����hY��A���1k��V�~�J;���t�3��Y �2�S�SVq�;���Ge-�z�໽�B�;/6g춋ԏJ�Z7���e/o�i>nK��.�+�����|㟕��5��U�a���InNG>xie�S)�7�?�ÊLO��ٟ���lY�Yr���fN���H!��R2`0j7���,+Oo	�r}7S�é�zL�����;	����y�fk�m���r�VC�/��ǅ�(�)�mRu�'�ť�0
{f�2�g	i<!��d�uX(�9���>�,�ۢ�MI��4��n��e,ﵢ��AM	��^��92y.%,�.��A�}�\�$���T}���g�S.2ӏ��i7��2���u�N�aȄ�ŗZ`�|��(h���݇W�&���h*����ʋ����a�:��W'Mi�-y����؉�-s'N�I��ȎhI~mf^��@J:�A��	R��pL�J��GWxq�?�}P}��'A�"s����%��'I�h+��lg�C+��I:6�e�*TH���<UuY�h�T%%}�Ւ����N$'������NH�ul��a��D2�b��}���FW<c��4�	��V��D�X��	�*�׷6�nD�v�P��/K���<L��b�]x�Ό�� }�z�&k��\^vs��s7��;�QQ�w·� �y��^��)�T��ghٕ�����4��F)�8�nÎM�w�ZC�է&�t�o�H��=>���+gť`�1��?�}��q/5���"�����9�$��{A)�QQ�C��й��R��B�a3�x�B��'N��O*Өb�p��$5U���H����&��j�ˀ��L��ݕ\	+T_4�9��H���������5*�;d��`{9E��y�2�Օ�?|l�2�V��#|2�4�@M	ƍ����\S�e1ᑍJ57��N�d<�4Y�M����z'ⱠP�U��]3����dM���;!�V�����<ƕ��m�q��͌��%�j�N0U��\"u��}2m8{禓'�q��8�̋�h-ya(����}��n��#���Q�^�d���T��e9e�:� C�!�V�*{�=��\��W�� �?u��!�!$�+�d-p�΀'��J�<$��B�w!ʖ�,��̊�ϯ��@p��C��k$�ZQ�s�8�L��D�A�a�_�҈�7�#�U�����a��pДM�]of|���U��XXg�p��߭�P��))�OLq��.�XJ�-덴R��n��4�5��͸�j�i��F���Si�QGE�~;�n��^O�3ȁJN�£k��( Õ$v��1"(t9�e��%�Q@$��^�aF褷�L!���>sQ?�?X���{�A(�O.�S�"�����ha��v�����yK�Wt� �@��~�@��S,�w�9x|ɼ#��=�� |���#�e�O��7y�� �ϯ�8��2}tᜰ��95E�i�;rh]�� J���@���0Hp=F�������(v�KReV&dٕ��fr]/��e�VFxX���f��`G�Q�E����G2Mԏ���E�'X����5v>�K��n���1�`<��Z �}�jR���<m�
���_�=}��g7�b�a�K��korv�'�`.x�"7��_pe/��f��զL�~�o�ʍ�	��R�����{���~O�����(k�D�g�q $�N�����ԣ)n��	��.�	"6��O�2#0ɫeYU�_�+�	ԁ8�1.D1��w�.۵#���a��OyH�uY�(#�֘^
͇������8��TBJb�����U���*��M��c�}m,��� ��+.���\��`�{z�n/Y��LZ܍�}���"�FK�|��QDԨ'%K��^�g:ː&Yf,�u@gTL�c���(C���a�����pr�GE���ԑP��vȴ~�e���{�8�vFD���S��_QL"��y��)��v�^���n�mH�ڙ�=��B ��3�է-tNO�D� )�*���8AܜC<�������G��
�N�$��}@�I��6�C�Ȥ�17�YJ�^/�:�-O�J�(ٺW" )Ϟ�5��?���Z昌,u(d�qx�ȯ���!hQu��7l������kjm]���:� �d��W�^��-��o9�C��ɱ���[�1�ѧow��S)2�B����O���!���'<�F�̩
}XHl�B���6(�E�I�5př�.�J}�͘?!a��w�F+��i��yv%� �[a�+U�գ��$J�ZW�0�9K���!N&�Lّ��?����Yn�(�)aJ��P.b�AKR�;�9H���.ay%�e��`��U����>��=q2\.���p��'�d�ȿ��������<.G	�e��A���d� �z���m���:��ac���A1��E���������am���7��Q�Qg�UsUc�y���J�
)�(q�/rh�U39C#�KБLe2���.Ġ�t��7L����5�j*�aP!�6`d��%���>�Z�R8R��f!h��L_kf��,fOnC���G+2Ur�v��ʄZ`߲�˰,ϡa.����/��{w�왹o�uP�r9�<y��S�T��H��l[7s�J&�τ�`2��Et��w�����t�|I��l/�ʑd�R�pD�l��$� d/�0�_�f���:��-^����Z�־o����y:��j+7�5�R��mEa��#���I��o�A�����;�^0�\.7B�ө�{桧R9�GB�?�ބ7h!���H����E���E���9���
��L���ġH�ǩ�\��0`M��]q�K���[��,&@��t쩛L��NW!W��-~�ow���o���)��y�h�i%a��SsjY��uN?���c�IGK)��z�l˄���1N�@s����8ԑ��,	��y�M1��3��'�ju��"��A�\w,�~���J���}*i��Q4�:�A��qQ+qtQ`Gb^*lx�Y���5�2�����oc��&��L��Q��[�����*Z��w���6y��>��Wd.����<�˪w��&uN���_���f@'�XJ$[#��}̀���5�˷`�k#�WAy�Gq)��6B�=Ct~���ʤF�wY7`�8�g*,��E��G'���M���Y�@Q��[,��!p��Syq/�6��kY���6��-�-�6d��8�K:����o�(e����ړ�Q�g�U��_ٽoP��s�EV]������E�_N��)L�j�T?�
?n��~������-��ރ���������
t��}�9�%r'�i���!?u��zTk��Q�����S�_�8`�L�N�l�J8�ڟs9�5�EJ��t�RZ��`��H�'��x@k�e�<\�FۙY���������+U�ï#���a���C�D></�c�D�`�aώK=~���)C�BW�$�Z?��؈dʆ[{�䡇��0��`Oϩ.�fs���VU��:���W��@���:��u�
�%���W��\7YU(P3�P�����p���~QHP)�	�;�s���[���)~q'�+�LB8�����~4�=m~S�κ*a���Y. ^��dN#�����{&��f���-�+�y�ط����J�.ny������(��'�:�.�����"Zg�V\�eF��,\��ny���Ü0�I�ϐN�'����^�kI�/|5�D�گ�
����)yL��)QP#bU��w���q��]��61����Ԋy_�)�ς�ϺD�֞��_�-�0�ީI�pOM!�&���}��^F�l!�<�`�5�ޮ�!�5vY߶ؠ�Y�ϗ�ǘ�u9����k��bWOϩCZ�H�D��;^�H�(�v�����.Z�%hJ#׉�ӫ](��{�8��J�:aӗ]W��Qh3��CՌʘ�	9�q��i��D-`�P�A�^��=�Ԇ�:��?�'*���reH�ޤ��L�Fq�?��d�,�=t�1���)����v`��/�ֵ̎	߫]�S4��8��E}�)E����A�g`��$/F�}�uW8��W���e���x�ƹ J�#�wY��u��EI�'�!�hP���E��=H�/�W�0��:���=g#�mO|c�
�tȟ����e�o7^-.�ցn%�K^!���"ܲס�7� ��R}�Ջ�����%?2e�XxH�|�*��d�Ǔ,N�w"'�/�o)��I��1yb^��yZ��>�Y���.�k��C�9�c�z-���9�oAu{�$���Mu�������y���$(���y��ͧ��D��&��:�$� K�Ի;v����y�_d,ޛ�#��r`�9zm�4���$����f���ޙ⵸��{�K��M�bm��q��#Xμ�:����3�"W($���H;�P�4�p.*@�?�@8���H�ϐ]���F	�qJ,]��en3X�]��B��J��-��{���ު�����*0l`waN
��t U�s��3��L&��P��o)x��!i����X��Ro����?��p9�7|�<�]�n}�{�wd�mE�Ӂ+З"�����S��2H|j�@���5��fwĥ��͞�K{�����.8�,{�CBıR �aXx_���r���#q(^T���}��A͹����iZ �	(ٰ�tXZ�w��$��}����	�tS�>�����4�g������&ci�n_�3����p_(�Ѫ��>��G}	����}O���q�1��>d8&����L����xl<�����ZA⯗Ñ�+��Egk�e�7 ��;[{DY��rg�b��NۖJ��I�����k��[;"x%pk�h�&9eq@~=��
�ߢ^g��1����n����a�hUQ�?n����3��E�>垊?�*�\�U�U\�z�3�P���X̉*�t���O��ç��dQ�,{�Zk���˞1χ�]ok5
����.2~6E=k�Бd��a���hy�A�:�xᎋe���0�b��
�SA�~Cq���{��m��%��Q�51"}p��Q���	��2�~��ְ���^K�'��G7��i��>qbb��s��9�H����ڬ�1�Z��0��-	_��f��g3���RT�Pw���$c5��F��,��L#�n�(
����*��F��7���j��&�Wߥ��0K|��ڮ���C�t{�/����%cR��}H�)Nq&�1���i�\����C|�ߟ��\[m!���	O'�"UH&��rkw x�/@��E�G�(����LAG�������:q�w�:pW�!.-RS�x"2�̸�Ej<�ܸ�B0*�V�n\i�ٟ�Ia�
c�X�L4;9�"m7�r�י�'���	?�cA6 ��>SO���X��=�Qx}xz�yi���k��?�V���G�g���������AU�{1�?��{Ym����M��1�k��uH�$��d	)6��>9�E����朑��x�),G֍A�\m����2C��K�fR��,\7~���k!vQMf�Бf�>�h/�����03U2����L��V�8�A)B�d��[����d-l�/�=9^�۸C'.n��]��%�Y���iˎ��5ω���~#����f���q%`�V�|�m�^ܒ�y9J�{aZvA���K�Kn���B)죗�As[����!5�H��v��,EJ�Ь1(S2�윆���*b��?@�Y�?8{�{ ����,�J��E%^��i΍����j��9�s$�+����S�.ǜ�y|2��QQ<���(q���=`��^)�:E�.�T�#l�W�a\}Ũ&�>����([{�YN^���sQ���~
�>N��s��9.~��e^uە��%��N(�i�G�ѹ�����)��w�*뛞]�Zk%��"F���!	�L�W�=�Vt��0[��P�E�Ʌh&r���VhA��2�)��Ԥ�����;x��M	?�4��f7x�dM��Z�V�-���B��N��-ºI��aJ�d�@�h�盳�L,]q�IhM���_���m�V9t{ٰ@��#�hs���#��ֿH��	`^�Z}��wP~�![a�'��.�3�ԇ����/���B��Ϝ"Ԏt�<og��|g�V1�>��()=�QLδT��@(@�� y,]��8:���?��ŋ�S�u�����S	��6�B�vW�B��q��15_O�QC(�Ki����.4d;���`l�a��h#Z"�#r���!U�PLQGf�zSKrT�/�L.�7�s̐0f$��W5�^�݂���?G��hn������&���~��M}J��%�����JM1�jk�\X!�[�<CZ�1�(���qco���W ."fwRV��++��j�̀5��p��m��Y<l�$6�ˏ:ی=c�EĂ�5�S��������G�u�j)�G�*k�P��X0��02ge�Б��S:Y��Nbu�(UG�B"3Z�6�UÌ<��2'	��)��IW�u7���ЏK�2qrdB!9��g)�����L�#����.Eֺ���f͘X�V���`��7��G��e��-ԩ����wWD��3X�J�8�1��ƒ�-�^�&����1� ��X������w����L;[>�=H5�U��M��A ���x���#أ���e�g	8F��<E��ŀ�"���|��4v����4�4�97,���^���X�%��_���DM�?��ߏ� �/����i�㓛�B���F����_׭�X�����Xʴ\\͒�ý��+4�מl��1��*��P����L5	]Vh'�Ҵ����7�P�(7[�̦�[�h�>6�^8'�Q��ǋ|P伽��͉q�VYM`D�m8��i߂��6B�8�ϫ.$�x���o�7��/��0�
������|�s��r*��
1��H:�wK�h{����6��M��r�'��ޥ���[P�>H��Y crB���<Bo�.�>���@�j����$-]�������մwb�a�� ��	�������N���3pO�,fW�RB���i���z
��I���*�ut����~�?�����6R��AZ�Y���2�a�!�d_�/x��H'P#D I�A�JV=l�8� '�uV����ʪA���i�#4���-�m����`Ӈ��kyJW
�����T�=@��Pm���@�˵D��#;H�Ib�v��x� �t��ZAMI�X�a�^=�p��@-�V_zF��`#*j|{�������