��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�x�W��$�oC�Lw�S
�,h�eԀ)�CQ�_���o�E�'+��l�����qz%�[LըMū��ş��Yz�g�#Vz���E���_�����/��'�w|g>ѐ�=dC6����	NwJ!�
�PΙq����F�<hŚx��#��aT��R��`v����*>wEb�3�4��	ηto��b���RQX_�?+��M���C�ӛ��/�7X�FՃ���W�"�Wa�'_ ���0��a�ߛ߈"�|J�0�g�w���r�~����"0-̦_DoU �0�,���-f��!3�!
\/��M�;�P�[ni�s� R F|�h�[��UtNi�qDۏ����F�N��Q+�9����f&D�����Ш�q�v�.x�a󖷮�]g$�3��|�jWu�m�lB8nB)
�
:�$�y]��Uhֿa�dfp ��:��b��Y�ٻo���i1߾x�B�i��F�"�<0A7l$&������y�Vk����1 F���C�l(*�]}Ԓ�*H��*PPm�>�Z;8~[���Z��{H���^��-���؅��ʫ9di�����K�vk�E�:�3^t3Q1F"�K����>@�H#����]է��檹J���7
W���Z��c��<?��_�[d{�ч��Ϩ�lB�����A�捳�pf4{T\K�:j��.~�����l)��r�^��y�u���s�:$Hh>���	��'xN9��yEySSKҐ*���L+C�4�]j���*�ŒqK�KYeU ��	���X�Y�C�v����]!'XK��q4"�cE>��q9�����2įP����?(�"�{�����,l�{�?l�7�`�@k3L'�����2u[�*R�����V�YN� g��}&U��KG5��[![�@��bH�<	�� "����ޡ)8��0>u�$�U ��F�Zd6��E<b� &S�|�� ��c���i�ڑ�A�h�'��vS��y��+,a�OG7M�ܪ��̮2��x��y:]�/���>5t(m绶Q��
NqC�M����a3�@IHb�).[T�|���L�ʻ@��rk�6��˨�S.xU��x�	��uo��Bf^�-�;��J;���@^��I� L_N���̀v,�Дm����+#��@�<��0�!�d�-��e3����5w��k����T�q�HAX��6��c+T:L;���7ɀ�O��O	٥f"��"�1ش��\���~ˢ?,������Z� P����*"�����L�}��v�0�#�9�)��C���w�.�e�&c֙6�I����Bތ
�h�b $�z)�d-zJ����m�H�-E�s��ٚV1��ܙuy+l�7[�/��Y/���L�h�Z�7��<�<�h��Q�%gB���6����,�W'�J�_�4��Zru��F�[�V�I �z��j�7�JC�ֶ�r�I0gӒ���55����e��z�NI��F���{Z��,OV��Op����!�| ȗ�fY�>�z�h��1х徂�	�Bw�ެܾڪI���r��j9����ԋ�d�&"�:�1��'A�@6BS5I9�z��w7���)������إ�|[Q/���.�||a���F!� ��`bY
H}�����^C�������*�|����?�Иa��2�(Bg# H�d�71��}�dP����N�I0�`��ݺ]ƽG�D��P��7�'|=�!�\ĽZ�}�65l�� )t8Q�d�̬��%D�綤��M+��t X�c�]���⬟���Z#J�O�Z�����r�_�iz@��T{��,��脡Y��8`_*��Kv'���ٯӐF� ($M�C������݀�Jt?�\�Γ���U�5�M�bWi�⟢$�YLg��P�YX��5m-˾�l��D;H��'3X*�W9�G���?��ɩ�1xV�o�ٍK$�[n�UY�d��^Pe��;^�՝��b,qZ3��9�K{�&������yHp߈�1�+JR�{_�R�p�T���wUs�Uj��n6��p�6�i�����]A�C�tv~jwy��뎙�������Z��a4k��҄�k��'����D)LR�)M��� "��Xʳ(�X�%o1 I/P���8b�$���f+4��A�r
lW�T�J��.q~�I3UkM�����5䬻TA�����g�GsjኤZS�Yt<�����h�Y��k(<B�Ы�/�ѷ˅�8{>�*�uf���|�jI���{<"���
�)�2��]�x}�~8��"�щ�x���O ��|��Ea��_Ig>̗C�=�l;c&7e�����{d�)�Q_�v'��$N)��-ǘ
��<݋i{9\��a	�t�Ro[uz���C��@��?��4E���}����1�Ə�U����|��h��!#~r��r�34��0P�JL�UZ�B
Q2�J�(ŕ"�]k~����ø�����[�0���7���[��Ig��K�����&� Q���/��b�;ņƲA�We��$���KMpD4UӾ���O\�=��/3,<��x����n���^�,R�Q>�u���߻K�S�D�U��s�&g[�/7E;^)?�:0K����;����G�~:�5�m#�О�T�(��n�li:a���s�U���]s=m �(GΗ�{�/3wp5sg�;4�����~��EZ0���lމqlF�+�`��դ��&+~D�H��V�PA��)����qMP���o=Q���:-h�B�oBv��)̎Qq�!�#=�i '�������*Srojt���'9MUD���Ez����־I�&���+(���� &8��s����yxa ��r���0��C�p]ʛ����r�d:,�:�_����Q��X��/�g,����]s�y�	�؀JJ���7� ?�ωe��*�2L!�<�ɴmg�r_0�.�O9Ϩ~�@�2�A���a,��k.i��<l ��uY��	�����R�K�~��[������
]S2nqD��$��oL�#UH4/t�,Iv�"�Kr5�&Q���ESyS�h����%<�E֓$�C��D�$�K��Xq��2ηKk���00��Bs%k`��y�����p���^\��$aa{ ~�?t��z�^n��zI^z�؟~7QZ����8G�[Q�j_���#$a�~�~�(�d=q��XU�I�,pK����x�\=�H|���k!��l��\�J��5[�U@Մv�����Ib�KL����fZ��{��Q��1(�H1 �b�J^^�6�	~�>/FA?�v�ed��Θ̵x��>���GA%x3RJ�5�pCa�]�t�������V����dxn1l�����Xnw6�B�x?d̿+"L�VN�wl.�C�m��eI�,�<�YL���)N�N��Q���ހSՉ�	��h��g��Dd�dF�e-M�W����ӵ��b��&�{�i[�GN]k�����Zmt���W �k��e��|H���>X]o��`�~"t�3Q�qh�}�C���i��k�إ�^�8j?�B/L}�� B��B�W�o~�"�ƥHv8N��s�g���8Vrg���%���f���k�/-���G��Ұ��D���<�C^Z[B*͡�0�5������b������� ̮�mR�z�o��_�u���r��i׆�:-������aIS�ԛҨT����=�#��m�m0	�(�,�������0�Jə�}E�d�G�;mCՕ5Rbn�e�x��>̻����/
?���##���Q�(�_�D����f]5��T�p�@-�_:Ĵsh��'TqE�I^��,]��#��C�SX}c�zKS�=VLnC��e�C����_P��M3#��_4�r�ؙ'7��隫o�t������r��z���e��n5�1�I�;�#q��9Ò��3�	���	�Kz����#�s��d0i ���Ys���x�D�3� ��X�a7C��HW� M2�}lR
�l�K��*x.�F�(�����t��;\�.��1��h�?iyK���z
�����a�D�9�w�� \����Ⱥ�|�|�%YJ���e;�������v�r�T�M����%G{{��<#O�R�#��Y��Y�Ĳ��?(�?jQ�4Ę8�.��2I��;�0wȚc�D7Y��;�1r����e^Sb�KQ�����A_��"��+;�F�!���I��Aګ%`P��.J⢃�K �Q(�%"���tq�4�b�K;9�%�=�A�&@��5._�!����vK��S�����1�S�l�`3���2�ȞVz�
I?��C�/݃�2���y�����~�Ɗ�������l���q��ݫ>�ӗ�T
�ғ�Sp����M���R�!wﱭ?Tk�~��(J�xΎl�tF����z�n�d�0��v�]�Z�ZLݬ�D^sy�L�`���"�1	46�H���̛ɋ��;�

�@�@��?�8j y���a���,:A���A�zm%us<�+Fi�I{p�#bBz-o�KU��?��;Љ$�h���33/7T��O𿶨xx�����@��!9���ɲ�{��g!��d^@NZB�O�oP43�N�K�4�{�>R9����t��\޽v���
+�B��M��jE�{&�.G�?`v�8�:�A�i�a ^���z�$C�+mR��	��S1�!���Q�~�K�&���փ|�-f����M�������R��>u��?�w9����Hi�]�����*L}���ز����)���$yc�����w�1���/�K1�#>&�w��In<hkm����Ξ�b8|�D,���e�"kC_bJ`���<C����z�9�ayv���ܚ��C�	�>e��XR���Ρ#*X�v��'�F�f�h��	&@�ƚ���C�o=5e���^��
З����Qq�~�E��.,>[_����ģ�%9��Q/�{Q��q�a�h@��4�2�{�'��� �86&��U�l�Z��6����������e$gY��;��BJT�C@��<�l%��Q