��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����)n �n�NP/x,�Fu��D,�C�)��j�vR�������|�]K�U;���A@A�qY@@բ���e�̍�gF<E�0�z� n��Yaex�1��p�+ [�B��;$ţ!
�_�c�>�Ή4�k-�e�M�}Y.tצ"[^`㻬Kg(5�f��#��D-s�q:�0eP�%����+���ݐ��j\�8��n�p������xo��|�v ��o���o�4,٫'.Kq��$�q��\�6R
4�q0����R�R� :P~�آ@�����Sx,[��0�$���E7ٷP�g����w��Ϗ?\x��%�2Ç�n�Z������eʔ�/�w(¦.o��z�2y�m��#��S�F:�..!U1��#U"�SF��A~S#��?;�
�~&�Ҝ*��N*D��bg�K�JsL�ql���dD���p�1�79F�ryσ��zp�+���W(`$� ���Mk�S�<6����%ү!LxGp�̓\�J7M��d��$ �)�.$JxK��\)�ZU�<!�R������#_�r-q�HJrEѢ�*�C:�&�D~�/���F�������^����S�C[;�Z�5����RŤ�Q�a��ߺ�b����+t��h�]�*Ԑ�;��C#��]�r����2���?]�g��Ϛh�D�;�<��l��W��4hJ>NeH.ř�!?=x,����p��dAdp��}�X�=���y �w�S����0C3U����&;5E�� �����>�ݢo��Vr�����m�4��q�=��Ҧ+$�HIgKp�PB�F}6��GXz���x��b��)~#�_�U#�=4����q�ȣ�&P@ ^\����(L��V�:�������e��`�R�Q*���=W1&�ݳ��C��b�k�,F3��2	]�]^�-��ʯ;fg��GG�7f�.��~i��������Fچ����I$�Y�@�Ӈs�d7h�)~.���0���t�h�:�����8m�Z�"��Oޏ_8��n�B"kk�|�TƢWv�S3y?��ߨ㳦D���2e|
���Z��"ĭt҄�X�����Z�W�Z^~wx]b�[�+i-ja�T/�"(���Ѕ�K<e㹌��N9���Q���G���e<�ˉbbN�ۀp@��1�s�b�����'�F|��>5~��e�PU����Rmr�퉺�UC����l�39's9ܓSi,�&(��9�'A?s���͠�"z\X������I�ű{�����V��� �t���ߟ#��,��`@� �a���}ju$o���D�s*o��ݨ;��8�?u��R*�0?�O�8|�C��$`��C���b��_�5�YᔧH�}ӳ�ͅTˤ4�����'4���G��{nն#�鐴�mV�Q��b�&�kɒ��=��z� i�����4Qtі��X&�0��/�O�o�i0vX��þ|�jr�#j6�ǧ�5q�m����4A�
-6�n'�l2y�p��LF7�Gl��	��]'��9����ଙ���r�+^�ƽ�<��}�f�b�փ�󿌨�f�ݭT*1@�j�Ma�"�N��<�	)mBܰ_C� �mU���uk�%��ez|]_3I�B�Q(��UeҦ�"�Yhv ���2t挎���2�ˤ�m�l��PFR������'�ڳ��'�#��/e�,�G^�L>��呿�!�R\�'�'�׸`?�!9�QG����sM$ߧ�.u^m"�&i3��(t���T!�O�9a� �O?"�V��T�+w�J��/
�\���nB����̺B��fL,Wt�}�Og6���3�_7L2|c�8I�)cEg+%a�v�yݧ>�;�&y����	�B�O{$�\�P��^G�lU6PQ|�|*e�b�߇����ă��A��uE ����B�) �d�9`K��d)�Fﷆ|�i�е���߿w��c��2z��\����7h�FAI�����DN��CEikD����R�|�k�H	_���0x��Pz���~�vrm�� H	�{�Q��K䕨����<2k�U��L�G�y���\_�F�]�������(��
vuG�y[�g����Z�`���F��A�Xi�^2�R�����u���̳v�&vԧ�_�G�=+��X+����\z�\�;\�-e (�~�Α�d�^�q�1���;6Av�r�y'B~Z��v�P�'���v�I��Ւ_��N���c�����1��p����ON+��2�RZ���*r�=�n�vpY�p&�"%+������_�E�S	�ܯ���-���!�M=8��P.M�@ّ����,�Ѱ�II/�V2TW��l���W $��q��l(yU��b5h��s���/��������6��'��~s�k}�-(_�>��[�����]E�w�$�*���sunw�"_(�7A���i�I4}��i��?���I~�y-.b#>Rf�P�u��2EW*����J���/K"p�6�:��o�?�����l-&�� �����ra�VI��(��S;_\J(��d����r��%]����^��05�����k]Ds9~u�A��s�x��3w�����볪=Dy�(��b���&��T���xnuF��K�����}�Q��N�,)g<ʷ�j���@��D����c�[5�Nx�[^�� t�`0��;���{��aBU2#ε��=5��g��ʖ�N(hD9�0�x�*�i^G��[��[�����r�V&�ӳoF��u8[u�� �H�8�m�hb�*�%�b縋��ݫ����	��i���y)�����Z�.�x��%��u�s������h���/����Q.}�6NU+\�����P}2�	��%˞�7�Y0����Wud�Ul<��z�U��v�*y�������cc��_��kU�y�m�a6��J��*c��wP&rJ��[ʉ0�"��XyՓ+�s�Ԏ{>b�o@�pT�3�8h�sWZq�F�.>����o�b�1���'9������M����Ң[�K�46e �x{]�JV�Ǿ��j}$�w��94�n��+>���eg!�=��:%�0
 ��#�/����(�H��L����
��6O��N�1{(\��3�G"��)���m�qL���ݫ��O|5<�,���.e>�Z���^)KG����$�b|��)���p?�R��
��9;mi9�s'l��7v5��p�G��Do����Ւ�.k�gb�"����S^�a-e������'���El��7��k�
Ի�����E�7�s�-�@z��}��zR��n�*�\m����HS�~J�0��><F����?�Z��؆.�ح�(0�_��%Y�)As�oj�i�&D�ks����93Sn�N(j�4h��	)ͼ��<*�Q���F����Pi��JN
%�T{��Ɍ@��[��Msj�C�q��Xn�Ӊl�"5�`N�Շ¸�(��M�����C�a=�Y���������0�RL��n��`�5Ry�}���-���c[zG\T��>��3�Х$��^FИ��g1P�\�<����I���h�f�	�<��W�+o�ZL**�*Bj��(9hZ�!���j�{��}O�l��u���Ye�������ݻ�)�A�k�t��������vE�s�J'��4`�Ψz�K��E'�����!���m���`mQ��,�?��v��aJCo��ŔU<��LQ7�f=��Fo��9仛u�\�@F����u�W>fo�o�`X�m�I
�U㉔tfF�.{	���'~Y]D4�O\'(�*��M+y(�
� �U�@���tU�����Q��P��t2�_�8R�#�V��Qt�sS���Ҿ��ϪtB���*l@� � I�����!P�����ԓ8���F�1�D8x�?M6Gz�V�:�oW�ꪝĻg�w��'���D���G�y&T$�|��ݸ��J�l|�K�l�ޑp���\�C�P��нA�ѯ&�~/��VI�b,y�n���葂��&��I��И�E(�}M�\{Ed,�K�[�j��%"Vd+9�� 63!��&H�5j��B9r�|p�9S���%�炏��U����7�,��f�ic�#��agkB��r�����F���b�K)�]�TȼB<�~ ���ef����5��y����rLN�$'}��,�z�1}w�0kcH|P�T�g\��fy�.2�yg���_ä���q1�����</��2J�&)�ر��%���N����?>cU9}��O	����C��6�K,���WN��W�jSS�$����^m�z�8p~q%I����yU�%������:�����DP`�:���=ZJ�Y����'2 @��[E�
