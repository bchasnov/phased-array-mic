��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ;l�Fv1�Lژ�O���3��������F����Q?���b�V����Ţ� K��Q�G�D��i�o�Yʫ�|�F�V{:�� �{��LBB���Z��^sӽy/��[����I����k���'_hx\�Ƥ�?���ƫC8�r��j���?�[�b��Gk����s��$E�C���Iv{��Ϗ.��R+!9u@Gf6�e+~�7k>�_3�T�@�@����58fW�o$�T�h,|���z.yhb+�[��>���W��Oѹ/t7y����8�A?X�Xw��J~���k.W�$�'��(��ꉑ'[J��TF�S���o�z󷬓�I�UW���{�|�M�a���@�F�J�Q�tx�tEV��Z��i��lzt����#��I ������T0�=C��'1#"V,���)�r����4p1����Ɠ��LS�d�,BbD�י��)�@/
X����0�9�C�'�8�5��I��*���ŀ�К�;R�g2�9B}������Qj����F�5#,VF5~z�wY@�g�ږ���jbY'��&W���Q��p�>��@牣@N�#���Up��]���ߏ����\c0�4i���jK�tƩ�H-c�����d�@+�FRxY�,��~F��(��y���^�)P݈�k4<�w���Z���?4���E�}��_�á��š�0ޜz/B��Ѽ��#f�݌$��3��z#G �W�fĨ��H+hnؐ�&�,�Ɍ��9�ċ1�(ֱ�{��v�RF�T5r�����F6�}6��2l����Ɯ-pw@���
�O1���3��~1��І6	��v�A���@�e!����� S-����193��n���2aD��T�=��>� �롹[��x�eo�@ev;��ޕ9L
�#�M�q���$|�1ᾑ���Ż?�#�1Uq�w��I�_�xS�+�Dj���<��!AZ6R?�-��E�Z�"����YM��5��O���R�")HG��^>�����d�s�НƓ��jO��1�l��5-̡㚁�po�W �kB���"\��T���y���Dˏ|6����������ʚ��s`����FЄl��q<+������^�� 
�| ���h�"_9���P6q�)'@���QO����T3��!hƉo�����2p{���}�c�5�׍����m�0.^��M��J�iC�a��ܖҚB��I�k�J
��Q@eW\K��/�����ڻ[��RK�e6ڡ4�~�4}{��	�$U��Ҭ8^�
K��j=yx��s��LP��R*B�.�a��v���z²�T3y�<�`S�*�+ +�6�������Lp4*ĵ��l��)Q���v�Ĵڼ� ��q-"���*��aё�i�*�����E�%���$I%���M��4��J_^ԇ/{*Y��Ǯ~�=p';��o�t�������b���xs@]L��J��[�~��ro|�a1��f#^��"�Ս��֗]�EPHf]��`�y߮�{�_3&̛Z�9�;�(X�p���a94ٖg�F��ֶ��%EZ�7�%�/EzY>������)[����8����O5�S�R�6>=�������z2N�C�㚢mE]q���]���q�C|}��wL&���h^ї�H�s����Q�E��{��t��e��b���T�
�[l])Q�_�N�L!�-����a蚳�$����������!�$�����1�g�o"B���g���h�\�t�o��ޡ,��Z�.�:����Ձ��S��ѭ5��)N;{~]7��k�:��+�������d�F��Yi8���P�O�)�Z�� Wr�Ԉp ����Нc���&�x�޸X�k�3I������	����@o�����ھsH�i���G�B�7�Ƚ�5����m��'A �H�|�M�Sj��Ix|���K�*Bx���?R�`6�_I=�˂��Ҡ!P{� RGY�p�jT�$��d�������-܆;)q$ٹ~j���|>Q�"�jg��ՔG��>)���i�
�m��e�˸�4������_�g�)f���� ܾx��x�{���>K�m�"3>T��z��6Ip���`�a�4��2�	�Ч� Yq��<=�m;a