��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>hs�*�U��Q�����vXH�m��h̟���}%��Wo�$�����(1����)RP�Do)�c:=�lM����%%9M���}ۖ�xj"�NU2��f�(Ϳߓ���8�`�B&��<���^H����T5�ʵ��VcѿM����%3>6Jcɞ
Q�s�",�4���tI�p�����w̬f�J L�m��Jo�z�K)RDq|�q�8��҉�w _�����#n�+_&)y���G��P���_>��Tx񠒡����KȰ����qq�%�˨�V�@�.qG��UO6.��^�t(�1,�u+q�ǦO��;�]�]z�RvB�tVͱ�y��(���^�4�-��Ն�Vd���>Sy��������BF��:/241� 藸(�5*n^G�>������Фby*�<����9�~��)ԁ��_Ov�nHk�;@j��
�{��o�1������s����E����iԥȋѪQ�rg^����]}�|UONJ�֙�g�F�j���H�5b_n������yn�	*qs`����*���Z��)ޒS�� SPa��O��]<���tr���4�iN�����R� �N�K"4;�B3������b�T+���$�`NQk*��y��/�ו�(�]�>������Fi����HK���_��C��`h�AC\*����x�b�T�۾�0�B^1�7´S������ԃ��-{!V��2�}!����Y�^����[^���Y1��(ym^/������!VX�ZnA?Z�:��.}�R�"��^P��|��N���>��
��BT�X3�m���^�ΰ�(����i�w�] ܷU��H
���ߑwc��h�s�N��dNp��BD�U���ʂ��2-Q���`[�h����yc�YG��.Gy��[�q�-��l�� ������/��*P�\�ԯم�_��W��`2�>;���m��6�iN �	4K�*��>���֋�l|�������.��s&s�c��h한e��D��F�,h������3���y�M�]�u~���ma�����VŶ�dn��e��	_gO��lG��,!.�x�E�W.ޝ��*���G�?"���S��K5�J��:��D]4;�c��{���Ɇ����#M��5s�:�r�ǳ�\�Y���a��F�1y�[t<���ܝ����cD�c��D�)�)�Y����o[��h"�lfѺU�
K�JqfDtg>���<�*j>�q_���xZd14j��X�|a���6�C�5SL�Ʋ�5r���(�َ���d�Dz�KG$*��U�o�Oy� ���h����ѽ�냭l#�7�f�H3�j��p��)��H��{�9GI{�q��Dk��+5�1n+�ߏN7TI�[�r stw�U��o�Ak��D�`|������B$��i���9Ŝ���l_!�D�e�@�覀���a�9�K�Z��q�^U-�(����	�	KD���r
�@�:�.�N����"�/������مΉ��2�z��U8���������F�
��<����2	5��ӯ����) _����CkEs+.�_ l8^V¸9-(3�;t�B�F8���A�?I4�ap�DxI�EH�#�đ���
�.F�1q	̅R�4T�b�����U�'�/g{��1�^��SI�7��p%x�X��p�p��<�b3Iˢa_�� ~�'�Eq�2c��o�"Q�r�n4��\����SB��A>��P�'�?�Y�K�/*�F�����䩇�a��K��?�t�v�zk��!��3���~����s={���=w�ط�� �h�]�f�j��E�*	ʜ�>�;�ѐ(1���Uw�Б���U���e�N�S����hA�sO��yJ����>�R����%3ձ8G;�'~�}W0��)���V.�>QG����K��`��R�R&� ��� ��^ז510޹�eӼoTF���<d�E����Z�W�m�V\�Y1�m���k�GM��U�B|���)�i%��-*A��`�J~��kLFΈ��|��F������S�Ps�tW#u0�q�U_O���5�uV����F���Wzdߋ�^��f}�mR�d�Ow?��L|"�Y{a��G�$���P�@V�?��j'=_�Nt�f02�j��h��!ƋL,���\X����r�H��1F�w�}e��Ĺj�d�{���wq*y�ϯ��R,�ݪ �r��=^�e�mW/������Du:a������>NP�6j�����63������8@�M����T��;���*�]�|�1r�P#�����[or�υ4��nI|����W�'��&+T� (5
�@�_M�2� �+z� �e(?����R�����=�H5fɨ�v��zNe(8��5��<��zN�8$�\��#�=�3bqv�X$�����Zl�^�v����F�dMӋ=B��Ŝ�tE-*�w�nۢ� �%T�2u���sH���pf:V�ӏs�?�C�"o���
6�Cf��E�o:q2��ܝ^�NMT����!3%j]�'� �ȫ�⍠�) ��mi3h��l���
<h��˸�\t=�\�}�u�����p-�[�2����o���UˁwC��:�_�~�],.oA��/�����<D�	��W���ɖ�X�<Fz���|��!,���H|�B�4��g'ʴ��Y�b��pqZ� �d+y�3��G�Jf�h����A�s�l�}܆����?7��C�S��&Y�@�4U�Uei�я�g�3���/RM9%�ܯJ�RL�o.� ^Wj��k���`�x0�aeTo����W�o�|ˀ����c�Xh4�!v$��|�&�:�S�n�ݻ��a�9 �JV�M��!C^뤾�9�_7�u�M�� M�<�FoA�e�S5K����݊9�3!-�O.^��#[��V���+ �Wr��]�! D����=Q0@R)l�{n���
rU�]VO�����7�x��aF��e�Lx�����T��Ã؅H��3�_7)��7L@�־�G��qz%:﯋�0
�)�_�91s���|ڣH�RH�6��X�ELW�����2��,:x��[�ANs�¥�J���ؖ���k~�(J�����t����9�Ձ���%ٵ�\/^R��ل*�i�,��Ɛ߃�G��k�����_�/�"���
Y�֡�M���zS�3�.G�=껔<	���y3)��,��3K�Al��c��xE}!�-m2|It�ɻh�pO�T(咵��p6��]�,���|���8�|�hxv1W��g_V���+��Ϗ�ԡ����{���|�WНQ�8�W^�Y���:�=�~]��L|��2l�_˰}�.>����B�O�s}L(��C����v��(ķ%,u���扦/<1��r�@ �?��~��g�J����xC�f=�)�ꇩI&1�a�vqp!�����bxQ�r.�3�%� ��N�k�KZ'�V�	����t��1λ��͎��C�o�Rz���H��G�ڱ�������x���AG��N��"���Y����>��("q8�
ޒ�"IK��١+����o�W]��R؞*�c�RYʉ�z%���5��*Fq���[�'ڼ_���"�E.5;��j����h�0UWV[��}�5��N<��a%�?�en���Ow��u|>3k�p.�ci�u�v����N̎����c%�5�C��WL�:	��2����J��P��.k����!�dŸO�):,��w�X�<�2���<�c�S l���;o	����{(P���X����DR;j�}Ĳ \�3�X[X����!	�M` �u��wAij�M7|O�| vA�R6�~ш�����U��n���'�I�gwY�wf��h�d֐^2�@�U3$��,6�qp����i<X�\����!Vj�jc�za�hF���<��H���M��y������x^D)�4�-{;��@<_��E��^z��s}h�_�y?v ��FѸ!���>Pz�LI�JĴ�]��5����薟�j�H�3@��%4��-�A4�� ����5��T��j	h^�%�	��P�I���/�k0V ���c�H�Rb|��@�|a�|�f�$��&Q�����M61���#B>hB�����[`�^�R�`Y����* aE:@��,Y�	~�BW��'J��m�����iɺ[Lz�G�����+�9�f%��z�u�5!�]l,7p{�v�~�Ø�C:�uHѵ���c����8�KE.*G9�/�J��Ǎ�.E�6��s�b+�E����-����Wޑ<tv��Oң��N�w�K��Ֆ��s�x����S��:�mB;��wW�;��N&�N�r)r��o~�X���.�m�1�#�u{d�W
�z��6<C�s�G�𺏢�;7y�)�v�1>뎁����Z�R�FxE��}����q��ݨo#�,�e���d�T�Sis_�7�G��b��o����W� DJ9k��Lʱ�a|����8�/r_�B�{�p
�7�B���l�x6'!��В�����-�����i��?}j��`A����m�C�>�TNn�+���am$TPQ1�PGc9!�Â�R-�VtQ�"�l�X4hKpӤ��,�c�#d��ϗ�v�u=�S����.����<vdJ2CO���E��B�\�(M\�.��E��\
B��7��6�6�-'����|��2u�G��f�u�,���	�:��v&'Ȱ��c������� ���d�Z�l���oJ�M��Kwd@v��@�y���U���^��0��h�yQ�eK�L���y���� w��ՅϵP��'l�3�Dqn	��ו�IO�/`�U����_� u?��P_�j�7��o$0�[�|�8�6P�T�#��k��櫩7���ko��X�J'%�Ǐ���
#�puoű �44*o�=$s�˼��,ޭ�C��M��D
��Z�!5�r#I��,�a�U��Pz��牽��[���������tA{�<>�����^WƣMh�\�	O
5$� �K}���t�osëA�Q��Ly�l%<�f[ʽ�%�5-��770}*E���>�T��<^��@$�U����}�1���?�.$�ߋcR���K�><�'�S�X�A��\��@��3j>6�Vu�	mI_7p�_<��9�Nݲ|�\��o�]�X���0�{�0�zµ�+�(��K�pB�JQז�b�#�yc��|n;�?���OO��κ��jv�"+�Y�4�Q*Ӏ�`Lp�Y�ݒQ��ž����T�#�su��˨��5�D���
 U*X�#=]))w{;� +̪D8�����߲�ܴ_�F��no�;��9uJR�{�7xad�ev�ݪ^�H�~x�����n�/��"Xv�
�5��Q�s��p+�R�*�S��O�c�Lj���Ƕo&�\�`6�T����^	��E��%M�	�Lä$��M�ݖ���[Y�4�x4+��n#p��K����L+k{Qd|Mچ��1� c{��Gc;PRMI���� ���g��/j���I��a�c>& ��`�8�,0r@5�Y��#3��g3n�רk��0[q�<G3���JD����g>�݊��ަu�)�צ��)o�Z�_��������+��ЛT�+��Jc���W���%�����꘼{�2Rk�棲"�����Gc���G��{i/��"�w�ͺY�!R�������.	bb7�0�*#�����hK�� a@�1��1�2���)�6��|�4����7wJ}��:��P�X!W۠�G�w7t��m��@톉
{�̢p Qk�Nj5�����b�	�P��\_{`���w;+�6���9���R'Lֽ��6g3(�/���îm|cg�������{�<�#�ྭLۉ���?�=b�#7k��PFK�]Sr��©cF����m�=�n���R���<w���q
�)̢mN�X� ��"Eb�@��-'��d�=hjgMAk�1mN��r����W��\0'���m���ᚬy�ۡ���ڧ�L��¯n�dR�l�O����@ �p�sf�y	��/(��� �
��Z��ɺ��A��֛��CM����Ҿ�F��pDx���R��~a�k|��A�M�"pEL0=�s?���������g;���')}�:���o��<�Kp����ګ�5�����p<��l���Ʃ<RVe�(���/c��a�ȉ)h/}{3y�Ki��}���:�L��ri��Gp�Z۷a5����8���m��D��{�w���w�T�6*��e|Abe<�� ��)��>_�HB?�Zoa�8����'�К�D��co,d,S��T�9o�W�!R��<�ջFߌTO�c�Hb.)g1ʏ�Nc�5`�r�k�����-�HGb��$����B�5u��yEt�x��;N��W<U�;�b����P����J:�C�W%�����v)��A��h>��Tf̕�ɶ����<)4��b�Ŭ1�����H�E]��.���Dor��V���r��J?&�v�L�m�E�A��	� Os9:�>��G0�z��J2*o@v��4Qy��3 >о��@����Bho�>4��/�S��ePUoT�m�_�_�> ���W����B6s�_2s8� O�p�io�6�F'�6"��`�Q:�*=6 `B�P��4�y�*/E�'���
�UI'������S�D���LI���gGgL�j�|�Q�ةU@;�؊e
\�4��4���f��X��G��,s�D訠�&��w�@���q��H,�5E��a�/��h�X3�����n��E&^#nR&d%��a�o��g6榛�rAG���`9�@�V{(��^�n���Qj��Ҋ��ͯ�~I��_Ԛ����Y;<�����np�������ܨ(�Q��N�q�h;:Xr��#��FX�{�,��ꀃ�C�sq�@��������3�y�-S�i���:�F��ƨJ������(�P`m=�����S`���`�'B�O��x�j�@�ڋ����#@���5���"�K��%���toޅ���(���}��$,i���v^�`��JƔM�s_�2�@=�q�m�R��=�����˂��~y03�)��@T��m���Kٿ�'��oC]a�uml���2�L��~�!�#���Y����R,*9Y_*v8��z�cu�u�KD$F�\
P>��bj��t,	\�����r�]I� ���0��(s�h�J�(3�O��$(��Y0`&��R�5!={ŉ�$U[�	Tn�zlT�o�6�ӓ"b�R|�}`?��Ж�����g�.apNz98�ظCn8$P�=΍$��8��z���)��zM�����}�I�V\mE�r���P�c��]Cq���/��`�a�9X������k�T�2�,إ����c����y�<v-�z�i�/���_��Qr��Q�Ho�ʝ,9Q &FfS0bC*�p���s��D'�FyHJ�$U���ˌ����<xr���/(�S�B���-U|?����ܴ5����%`}����~������KY �1��S�"Б�adfE��X�+�$
!�T��ヲr��nI;�q쉖:{�4	��j�J;G{w����<*�.I�(� ��iſ~9��<:5sL��[��.�&��4��}C��j�~殰�