��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>>�Htd�η��$Y�_�R�K��z��Ui]XM�%�T�O��I�.����N����Q-�!�W�� U�z�����y<��W�<j��s/f�W[��_pr%yp�ԑ�iI�����q��7�2�f��!0 Ù)����#/�}�����$�o�ܴ^w��r���C���$A�E����i�W��(��*����(!dq�a�gd��$��� (�Fj}+Ω)�6��y���s��\
��� Y�ϯk-��l�ğ뇎�"8*���u	�ే��'�F���y��;8��5��""l��)�Ȃ�6�E$ hGA��}���"@LF�\�K����RY�@XV��/��7B�oF�8���r1�(<5>u���n~��Y	<LB�#�ԇ���km0Q,�Ͽ<���1%����ĵ�.�ϰn��ߏF2����H� Z��j���m��m�O������Sֵ{U����P~3��YYW��/X�eG`�^��u9p��2�0k�?��]9��ca��J����Ic�w�w�0l�뒪���?�:��:p��TR���N�2� ��ssw[{�>1F�vy:��],�.�4�0� ��@�q+��ٸع*$��ýJ�V�2��u�@�m{�js�%?-�
����H�^џ�|4u<���i�����(�Gc���)�@J�
���T9e�j�A|�a!�ŉ��K9z�������Chl������ӆ/���%�	g|,����炼�-���< ^�ޓ~�OV�'2���ǊB���L'i|'ǩ��܉�u��"L�Buu M%���x���i�M�t	�f�<�(L��B�n������B8��'�ù� 9�m�ߏ�T��c���n�|J�`�q�I��J&T	��Ӫ"X�Z����TbuZ��drv
sɤh9t�ܒe�K1���xZu3mG�X�(F�� X%E���d�0EA�rT����the3?�_��Mx�[�Ժ��N�4���`W���>��S��������p��mJ���	��z �e)�p}���C\�#�b�H��+��sz�=Z��>1��48���
��ɳI.$�g�����_�q�vs<[��@C�ZSIA`8-o��,bhR�����l���ƅu�T�xNH%K�k���~���?4���s�x;���;���G1�%?��)������2��se;<,[	�\�V�����k
����VZxő��#�-�2>��ūܺ(��2{`iT�F1�ր��)���4�F���H F���"�8/f�C�v���T�lRXr���|�h�ML�+�ߪb����:a���ѿ#OP\)�C��`����7+��ZvY�<ݷ���Uy����e�,=迴�w<r��0�L"�%u�,�y
/a��mV0rH�5!�9F ɠ�٘����r�/�^�rܰ7�fn/Gi '���#��r���Vh�qםd��05�����8��^�"��	�.!_p��e�Y���M�
P��g
�^f7��8B�ٞ)j��8E�BNM����ئ��el���@��MS	�$�����J�+<����G�- B�˓�s�i:<. �t��ԇ!���c�<uL� �0�k�8��O]NW(
J'HͰ�j��v�G�&+V�$��O�I��*�E�*Bb�Ho��I�`A@�H�C'�$�5�$9r�U���~m�бAD�?4�G{��f1���~��z�B?IKR�M��2�C7��K7_�W�䰕ӥ=x�JJ�J� ҝ=&0s�J����7^����@|�r�����7��R�W�7y9��a'�V��i�F�P�J���o�v�C���}PÓBU=>�?�WJ-��Ԁ��\��;] (MA�15a��c�M��WcG�BA�P�E�{9���W�@L=������?����V���&�p�4�RNH^\���3�ag9.�����)�֟c
c[ҋc����W���x�=��Bd�Ч��
td����Q�ϗ���K��\�p7-���U����8�D�Kx�=t����Ӣ��/��M�c�%�z��D���:�8�=SD��f�YGO�O��TZ�i0��)�ƭ���Eg�8:0j��m�K1Qo���J"��8��U�,&�7X��	$�j�	�[����U�}�o^�3�2�<�KG�W�ҁT��\@�\����B�Q�X����@��Sj��D�58B��ѱ+HΜ��A�7+�� �1��#�C�|,����v)��3ҭ+�;��ĩ�n�}��%E I�QnyO��H�����!��2\5+���]�=�F��8<p���{�q�]�_�~\Β9(1V��3�Rt��	�Y+i��!|^�Ӹd����ug���a�����2(�.z�e�f�j� �)��t�=�JNT��j�[�u���n������X�[W�[�,Ic�f2xĴL'8�E&�֬Q��]�pA����\���_a���e$��׆�����_��V��6~4P��?�3��;�aL1+���d��.�����*��'ׅ)L�O� ]����\�� �ƿ��rf�M�Ȧ��Z)[ŀT7��0tP&�8f�W���d\��_�É�5����z�-���*ʹ�#�`��z��≑���zݔ��k*'wx�-�_$��$o-R�����>q�)�Ԁ�!/�!�tG�;�8�fg��T1�5��Ur�*��Aa�	�������[mzAw� ^�*���ţ�fg��8�����\�b�]�Ê2���	���&3REg�d �k�!��y1��m�s�� !��.�3�\@?c�lN|��TLp�_�t����h��������|aҶ[Li+R�Q�a
缍	�@����:���N�>�U֟et��c�X���x������A����l��א[A�n030#cQEW���Q�4d�G&:8HJ�wD��k��q#�.��v}�%"Ɇ�	����Vow�������X���H��xQ.l��c�X�V>')�Q���5Dtq����3��tǾ�3>(���Pl}�x@Tz(?�K,*A_��yV���!�ۑ���s�T�\�ƹSGݘ%Џ��]��-��
�^Og�/b���z3�:�8~$�T��2ff;T`o@�Z�A ~k���;n�T3/�� �Fb����ʅ��]j���}�N�y�d5�"ܺ{]Sx��?��rԟU?��K�����ם$�3��ӂj�*��@*���n�۔`ͮG��We[<�:+��{����R1�6�\y�R7�'�ώ��m�)�2��6�����'�#t�O�!XpKdy� }���8Ⱥ\�N����-4U��
�ݙ�x�昇(V�.y)���e,��:Ҝ˭�m:I���ʫ��Cɶ�[U�������������Qߛ{��C