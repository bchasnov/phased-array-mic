��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\����q�?��e�I8�b�Ǽ$��"����ׯ1�V0����������w�Iߵn�>��Ã��g�y�t�U_���1���V�#l���{E(s!Z�hx9~��Xe�X=�]t'����IH��}�ݘe���(qt7ص
�9ݸ����P]՜,�Pk?��m�aLi��}�%�������B"�t�n�&^l$h� #͐�:Ʀ#ԁB7Z\�����+��þ+!d=�Ɋk�����bx�9P��x�hH�u�r�I̗d�c��OKc���%"�_#g���t)�*h�Bw�4�������q�aFc �L	�1���*?M�f��۫ e��S� �M�y-�çť?#�=&Y&!����t������8��~p⧆��5�}Q0��Ě�����e�5xo�u$�����v�F,u4�[7/�;M��K��~B�<Tb��y�4�+Ք�w y+� ���Q��{��2@�ô���Ƭ�v���S<1�r%�N]"�Zig�w)̣�T�S������*��@�Z�[�[Ǎ��f����x?����10�w�
�B�@��O�b)���rq����uYL�N��G�	r<i��Gx��WW 3��)�]�"鱫Uq��O!��mC"]�Q*�=,|��p�cm:S�#��5tB��T�� 	�=�	��;�Qz�Y�N"�A�xi�𸫗F����I�o�k����XB|<�ο�'����+���h�k6ͅ�"Kat�ч���hI����J��m���X����W�%ԗsN����W%F�oҸ��uQ��4|�$�6��ϕ����S�������|7�&y���gބk�@�],�o�V�.��A1�;M{�oޔ�pU�u=RF��f�� �����v������dAJ�j>꙯~���}Y�8�Z_^T�����pj�"�Z���iׁS�c��{����@B]���Coc��K֔��m�m�R�#�rY"vګ7`=��VP4�O f&���Q	Ng�=�y�5��p�9I��s�z�`� U�/|�
�����q����_ċ>gpi#��_B~yG����(��î����p�V6�<$4c�L�;	���J�������LU��� 0b�ĵ���SL��{?'6�q�X���8�Q�&�d�/��z�n|�韒����j3�����]D�P���6�ˇx��Ў!p�k6A�@�v(g>��K����HUPa
n�}S����^��WI��\a`U��us��Թ��W)t��}�b�͚%nbz�usA�.��_�˃-�>�&������ޠ��<LK''cZ:g��g��	60-X������e���I��Ya�&�@Aې���A@MQ�}�)E:�ֵ5l3s��tR��]LʅF���Uu�ޞ_����E��"v� �B�S�v�W���b�Z���ɂ��!H}G�@Q�J�m��uQ�a�����\'�t�4&�#u�_W����Ŏ0�}���籒��j��}�"��&���ʉ�E3�1��P1S�4�l��N��<r͏�{���{Nf�7��-f4���>#�1t�J�S��H�w�Jä��y/)}}�ٗ�Z��D���� ��5P���? �'�^�@��b( �*���-2�"Ђ���[h9YEDeY���l�Ȧ���ZY<]e�_�K�^��>^�H�@a�^)^YKc|�=�����ߐT��m� ��+�qB\�/rDb�2�����C|.S6^�D���o?����N�]z������Ǭ� �r���gO���.��S7���k����*�aPp�TQ�^��5g4f,�R��,�Ī�I��f8���ृ���l�4�]��坐)ހhNuz�(8��Dea�_1�&E�/����p�.:�?�Yx�����IJ�}���Ǆ��t�ʱu��{y�z�E{���z���x9�*we��3:4D�gǘ�nj����+C���\#���C�L�ח�e�~k��ry�?���vt�!!1�x`v�&�YE��^t��G��$pQ%�l��<�.1�N��ʩ�0G�FY��e�|�����;�M��G,�Ş�fj �Y�7�:���?��9��|���)�g�^�?Y�Sob����~8�hȰ�5�֒\=c�oK��(�+d7�Ն��@��;���������B���\��y$.�gU*Ѵ��� X����Y˾1 ��Z��Ƞ�*3ra��f�H���?�r���]�}�ԌJ�DN�qx�b�A*�'>��a����ZX��17y3<�����[��kO0��
�N�S�)K|�􊸮ۅЩ]�ܼV ��#��钳Ҍ�Y��:��������`.�$I8S;n���;��[�+�X�h�R� M��
[��7�0�y�N��(�;�(�J�{��9��ƫKkE��L6�zW%�L���ie������v��V4��d���t����d���HM�1е�I���V�&�����EuaD�S�Dx)?ƺ0 (�xTl��W�5�������L�����&�Qs��ъ4��G��h-����A�F�֜띭,�G��+p������<h��m�R�0�Y.aޥ��E�M�$T�D�
"��E���4AH@v�xl*�B�#�SO�g��M�&�[CCon*�����F���r�>7,A3�[s����f��H?���˿���. %Z�ԕ��w�Lz�;�ť�J�~�Zo1�7�m�n�O�����Qi �
��m�3�I�`+���CTke�%9�*�1�����LaD���
�����r|�{��-|.5uoZ�����E�-�7��0o5��^����|�x�A_�&a�a�P�a�+=mπ���d��+�3��[:��0YG��0����l=���j�(�JƲk~���ls������BL78\�CU�g�%��+��%������o�{�~��l��;{�)�7��0���$&�������kW�E;�o֒$��[����_����ђ�^���$��d'[���Y|�8B�����Ì�/r�s���k>;��ޛ%�6Ux��^u��ln��J�Q��Nէ�ݸ~��n�HnPK��W���pEGC���N��R�����R�>�.%ZPn��Q��P�e=� �/�4���GJ|��%�"�ξ�=�n��J�w�����F$�U�s3���