��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\����q�?��e�I8�b�Ǽ$��"����ׯ1�V0���wR<�ozr�����G�LדL#��9��8Y�S����R�XO��/L/IU(�xe@Ϡ
}���k���1TNs�],c�o�EFd@5����u�O.-/��}C���;^���d�x����y����N�Y��/��x�)�%b[D�߼䭩Y�|!&�;P�C�U^z'[8''�
I���y�C�-X@�1X8�s>FZ��!�+�z$&,�ot����ȭ��lRI�层���B6����7TF�$S�C�Y4ފ݂���py�L�p��������O��_��mӐ��?����!�Cẩ��\�J�+k@ͣ��e�p<�gײBX޶�I�3����t�k�)u�_	�9y䝖*53Ɍ��	%d�����Yܛu4�Q����L��Q��~Ӫ-��B�S/)J���ҷR�`�!�)���I ű*,`�:��j/�4��ݞ��ιLޠ�Z��M|������Ũ`}���oO#|c8Y�|�[�Ѧ�B8�r_�-���$yN��AS��ˡ~�!? ��8�(YY�K�FH�m5�ݭ��|&��mK�{<p�F.����l��W�c�uRe�Ӆo)X�������a����_�N�HZv�
m�Ulv�ɐF��ËM2����<
���� �,y�x�c��)��h�������wI�`�97��2���d����ب��Q�X����:#A"-�m~�(7�o�ʳi��:�O�XN\��(��xl����*�����P����aC�X/�$1�#g>�_��K�)OV�]\"�s8ȴ_�l!�g���6А<�Iy�ç��vhe24�;�=j�Ǩ߉��g�1K�b�Q�6B��*�"U4�f���F���u���Ѝ_۴4��TL�����Q٘0��	fm���^Z���*��k�ˌ�0{�����%K���z��C`r���ް��Δ�yM�	�T�f�����x�ap��q�?8ܿE��Y�m߄R���V������#s$sؒ���k%vU��w:�BBo(A}�?\�R��T=���q�sO1�_�A ˌ78ʅ4���͋A�Q#�؇jmt;�^G��6J�b���?hj�y�Ǟlg���iyڴ�7�])��@9�@��0�h��G����싔Ǿ��=���J���V���$�*ʹg����)��s��$�T��or.�[�#ƿYDN#�ء.8�#����B��j��l$I|��t/���J�&����������@e��5������ʌ�lƢ-���_��\	;8(sW�e)'�q	�K\��l��=��8�7s�Z��~N�p�����w^�u�1$\�ŏ�\��+�iW�A.�ܠ��t�}�$o��ЇcP��VzC�*�Ι 4b�<)@�3�4�X�` {��<[YG�n��L�Nu�|�5"�����ݾi���;��F����à?��!�!1ƌ5�yV�`�y|[���d�7W��tq�]?J�%ys��Ԝ�ch&
-f5N���� /,�L�WyW)VTf���V�@>�d��Y|w>V�6����#�a �bɐ/�Tb[����Io����s�ڗ��4=�����}��� �=���C8��B�=��g��Y(hq��o���=��n=�	��2D'A8���h�k9^E��Q h-�i�0���U�ɫ��SxoH\�fW�\��p-)nU�����G��?ʍ���7�G}�T#�̼�8P�я��FU��u�~^ÿ�D�=wL+�m��� �z��b���]:a��+�(��&��!h��^�^8bK�v��G����7���s��w��&d�	�i���StPg�'���^����=p�.T����|g=�3IY�<N�S�,����嚑�nh�r��%�r�i���?bw|���E�������	���T�T8P/K��^����A�̋�t0��f]-m��m�2��Gg׏e�&�^y���.e��	;���ck��&P�x%�fͫ唠
�U.�r�w^�^��	A��7n����a%:���
/�ըl�m-o�PR%�T��d������=ܚr�����$a%�'GI�o���u�N@	������w2���]\��@z9}t>����v�8� ����n��!�wO^c=�S�E�cBc�%��x�����m��R� N���)'��
��P'os�H�*D����?�rJ��Yg��"���G��L�|�	uW2,T��������=�W4t؆�T����e��K
��sL9U�%7>N �~p|TN��&���	2�<����<�۷-~�Ej]��`}~(��(�����xF%��F���i �&���]F󛣢
b�m�I��N���f�N�rs7b���,�Vͻ��eA���C��N��f�3�D5܄x*b���6��[��|L@��9:�o3\��~.$hH�"X���/��������̰����UD��<,`;�*5]��{�u��i��u{�9;�u������TM�reׁ`k>����f[z?��kS|��}�긇I���Uw��Ki]�0=��2�JA��+�ǧtV<h���ԧa����]�\�q)��\�Wu֕s�{��ǿp�q�������@2�.wL���8�.@N��i����[,u'7f�����؜Ei(�-:w}��������wJ���p��r���K<s�-6�`�ҵ�ݹ���&�O�<A��H��?0��,�`��rE6ܤ�fk0P��y2�ɢM�b&V�^��ȵ�<�8� ��~�F�ʳK� K�e�<�-_��^��وE���+�"�T�)LF_CI���$#T[�^�`�-d�|��xf���d���c^4��3"|J�pr~��eQ��H��nՀ(�������}{���v��{�7Ay� �+lc��������
���uB ���3V���i����U���Y��@�=Bi�v7�yFե�\
i	�2�C�3b�o�c��b��h�����T,�Ƕ�O��2Y"f���xPf��E�].�M��G_|����~�n��o�cg;��D�>o9#��f"H�|�޳�@�}��]�J���Ţh]p[��Qr��ԋ�*�3�420E����p�Y��� �����3�+E'#M��#;rNQ��GJOC{)Di&b�/`t�C�ee7��`y-�SA�ᕿA�����Q�b���?��6;I?�O�1b�|V�����!��6̺{��g��)�,�U2xsL���<s�5���H��V��BX���$���Hb;�>3��Buߐ�>��]p�^�&�y�֚61Z�D�7�"�a[x�j�� ۙ���+��M�lР��>]^�oǾ��3���* �7�|5��w��ً�DÖ]OUD3 �	O�^��dRr��U҉�U���3�[9lJ`7�ނ�Bߪ9k{�ev�>Ũ�!�~+��}?
���R��^���Q�&��߇4� ����
n4���O|�c���\�p�#=�	���q��(bm���3�P]�br
�hq�t��Fz*��#.��߫
��.`a��c�9�%��;H��K�S.�w�]���b�w\-�c��Dzļǥn�����,{�ac�r"�*�b����E��r1���zZX��x�q�J.�D�`v��b'ԳȢYʕ�#U�&��b�nQG;�o��(/�1�n��/�Kى��x� &���F�C�vɈ�0��eaϔ1ئ���,A�}�	(s"Kz��L�O��%B(��2w��k���T~�syB�� kӖc���W���L�}ҝ3OV��������E��Fc2��n`��u�%�Ye��uI��aU��٣@!�_i4'�>w�BՃ�����RYs7�+�R����P�?�b��fK�����G�7Yս��HFju��ǟփ.��^�zX��d�!3��l�\}{T�������LQ�)��sM�;�9m�����;���i���M��_kR�]��[����ɃW>�@iJ��>7Ҙ����*l���s���fo������DÐj��'~PK�q�?F4zy�Hm=��}Z�7Z��)7��"I�4";P�Ȉ�;N�R��+�X�Y�'$ᵍRht8�HCe���	K��֘����ւ)+y0r�c�v,��˞��y�H)��&��[��W��)I�Uؿ롤K �c���宀�mh��k��a i��5	�b���}�\X��ڼ�E"�aIqn�ཀg�Z9�5���u��@�/���7�ܝ��-s� G��9���ɏ�Ic�F@ϻ�wF����~��+{\�܌u���������}/����$�{ρ���,�F1=�o�4�W�Ƒ�s��_�o�@�.\R>X;6�8�>5Q��Y��q�%�G�O@Z����Q�6r��.:0�6����:弄ʐ�3�M�Ao�'[�X�;j��u�]�8�L�s?^�D��w����������ԛ8����k�KM�*G*��	�p,�#�� �w)�0C�4em�����|u+���S��pp���yQ�e�J���F�ǘ[���-���"�]q��HtH�kv��a�'xX��<���}�+���s��~.*���� �PӀ/q��7� Vg!9_)�n�ee	8���M������S�3"1��ۘ����؆�%�v�?�������˄d����ɮ�t����d��s?�}��3�Y�c�pB��M�3��oO� ?����\��+^B�RD��K�W�r=8"���Z$;}A6C�	+��\јI�<���I�6ݧ�Ga��F�Ϡ��K���w<��q	S2C/WWU=�A�hS��8���̎rUR���/�T��6�?^�B�v=����M��}�Le:��C��*PN ��zByx|
�l�"W��|������2��WT�L��E��u;
q�b7�>܁���{���!�%��,0�ʸ�za�{�6p�󠸕T�p�x�t�Ӿ�P��I�@K�4��8Ҍ�"�Jc6$�;8��]��m�ӊ+�D"p��0;��c�g
#~�o����EM��1uߖ)��V*�TT=�Y:����Gr �y�Շ�)�m�#��/Va�\��q̤�W���������Mg?N(F.���ȷ�c�0vYe	]���|P�G�4m�N��ָ�������]�k���4/L0��$Cv�dIP��i��+u�wF
L�!�~�k��|���^�9��C}�DuQ8�}I��B^R���҄_��L��Zx��ԞFC�!�]�W�=�p�zv+5�P�U���n����!��� =e�����N8a�+������Bj���/H�9WTa��a%��� �3�l;'�y3\Ss�m�h�x�oV��o���n�(�5�4˃���_P������{���e��t�'��`T��Aj@���f�*�T���p��n0�i�J��I������ҏ�9=`h�~j��{Q��,��+�T�ÍE�[�E�կK��/bf����I�c܍;^<���Ky�/Y�{=��$'}�>M+�	ڠ��&�������5�hz�9���C�$�}��ڑ'��	ѽ�PE�ڪ80Q�'���Xet��[������M���ki�����x�����oS����i���EɅ�������@�C5�l���*�i4��i#����QA�I��+k^O���c���u+~,Ks����}��bYU��(�O��=�>�9�WW�
�rX�����@q��վ� )_���S�]/�z��7N���Cxܽ�77��i��4�)Ocf%;�_�U��~ޔ�[kqw9_:�aЁ��-��M�%�T�)M=���I��*��/Vi���p2@��h��7N��P�|�f����J�9]�¥0D��)W�!�qH�
�����^���K�l�H�\_Q������,��o���m?6Y~��3���pu�>�17#F�DN"���1�1������'��"Q��^ךx��]�C���V[d��x"ӫ$�E�m��V�Nz�m$'���7"���':?��Ќ�����lw�dc�Kh��0/��}�sǘ	z��}�N�nz�ݥ<O7����F��t