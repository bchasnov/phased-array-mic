��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1���e}ʲ��cg�t�ϙ�a�:�KR�%���ݧw���ȼky��q~��9�W�k�����{e��bֈ�*���Y�3EA�n�[��_���6��qd�JD���u�B��9oX���q�a���a�D���z��닺#H}c-��>�o��#�oi�b�KXf��#�39G�ܰi&��,R�[�i�5�Pĉ�0�Q��2��O]�|��<[!]+4�WekgI�_�&(�,����p6з撍v�z�G4\��	Oq� �i�oEѤGC�٘-�rZ<�O��M���I0j�u��*	��P���j�H�{�-�E�i,]��U���^J�K��oY��yH�`b�q@>��K��}
c?�L̒L((�լ1S���'��=O톴�Ү��c��5&�=I��@Wk�A.��)B��#z^�J��.;R�ܸ��&L��ӗ�'1��/V�)�i�֘��B�cMop�����K��>*��Oװ^��/d������W�\85z��'�F�k�Boy��d�U���q`3�q& 5�q׷���v��ebQ�c����~���.x�*��_��?Ȋx�}$��T�������ʡ�	v��BS"Aڄ\b}s�:���%��&�B�q�V�5T�D���ł��y��� �Xj���Hm�mj�T�5�ګa:h�p~��/������o�k�ڎ+�*|�4�ߧ4/g��TxW�&~�������;\���U��Â��io��X�_�L#��8L�ھh`�TB[�T�R�,(f!X���+��i���X7�Y���?�j/��F����uYsq���E��@W�#Q��
���Y����#�P+'�|f�hW���l�	��4���$z9�>�R�C���A&.�=�ԅ���3;��Ew�48d�EOO��i<��ۈ}�ЧX���W�1.�����84�����`0y�5}1u����3l��7�����ǌQ�v�?�`	5��x��[�%j?��ta\Q��R@H(Gq�eנP�����cz��y��j;c�����~5ǰp͠A�$�@F�#4;*�6�r(`���I�/q�#T��@�F����b�T�[��!�*X��fݖGU�����<����_��:�_�ԭ��	�� u���&P�z;������<1�mC�K+���n���*�ʩ�:�7b���t%l���͡�.�V�� �����X��(+���`��@^ghw�Oy�A8#S��¨T�l�FH"{r�MI�=�l�1�������\��
��LPF�n��l -p<��`V��� �
�Q��qs����ikT$���J`Ǳ<�|rBv�B�aR�1x�=)�U�}"�皢J�C����	���<��=�5���Q��7'�8ǈyZ!I�)���Y�Z����μ}x�8���W�#����J ���Ǌ�w?���y��If
�u',��k�x��O<�W��F�| �����.���G5��������{�'���p�?--���Q;H�q�#4�y ����}+�&�������X�,�F.��]���L�zD������E"�h�tl~
#�.�.<�Di}�_cx%P䳢)��<`�q���	Tl2�M�[α�p3�c���ɼrav��n�ilT`���X����Ĥ�$�2O`a�I�8(&q�V&��"DہG7����Li5K���c��J��8L�2f���~��,Z�t���@����_f"%.�O,+6.bR�A��Q���=��h�� �z8g�
�h��"#��TA	YoZ���C?Δ7yzj�W~M`�ڪ��|�cAq7�TO�*i:��5�������qw����jD�xn�0ĥ{��Y�~r�"O�f뛱qd�����T ��4*i7���<9��`��Қ8l%Ƣkû,]�oFa"�����=�'{��e�W�y߲"�a�>�Ҩ��M�!�1 Q���������(�6N�K��~4@NF��
rț�i�3#���>�u�p��6�&��r��z�~���1�Z��<^hq`�@f�mEY�qu��ml/�b���_��W ��h���|0oc!�G0�@��:�����c^X�D4����Ԉ\RGc���B+���{Y��@M���o	 ��k����1Қ����Y���jZi1+�d.���%1!NwY��AU,&�P�c\�2á��V���-s�͋���B�=�R�)�B�3^%���pA>\�nʲl,��^8ܡ�d~"�N�K��Y:�Xm�;?b����dv.t��R@�O����!Ex�����Gǜ� ,�6����@R�Jm���-�Y��#z5e-jS5�����yH���Ɠ>�ˡ��p~�Ug�MUs�'�� �7dۿ�z�����4�`�u�e���w���)�S����Oo� O�|YM�#	u��r��G�߮(�.�Hwg�o�5��'e�u*3�EK�jAq.9]�s�]���^O��/�g�-9L%�ks�n��<�V3�&R�隍Dnز;R��������ߐ|��Je��Z=}��'S6��B��t	��`�|��|/���F���F�hjK�FG�Zct�5t��q���b�&A����3���(f��[p������H]򽟻���@�q`γ��eL�_	���b�sA�K3n�5�y�-Ӿ�6m\@��l N�fp�L����g�����{ε�a��{��{�D)a��3mJ�=��H->�He746������8,�qmXo��E������5�R���58~�VhA.l�>�NC+%x�\�\N:�+-ք�&�m-H�ȇĔ���	bJ��м8qت�\~?c�'�}g>�
k��n~uo��q�U�iőT}4^,$.S��q�Ͽ\��+NY��;���h��J��@v�vm�����������U�N���~���R�c"�ϳe8���kU>�E./f�W���B�h�hkO�p�sc\����W�3_>�0�x**�G�������M�s)�=T��c��!n6خ���	��uʾ����5���V�o y�W�L�Eu�m����O��hٙS=��w�y�n�R(�jL$R�{��C-�
?��!Q�⛃�+^7��d��`_%�}�PRVk����G�{������$g{8�D����A�w,[ĬT�sZ{s�'T뱗G��08×�d������ɣ�
��!���b���3�J�Sj3�b <;��: oQ�̯�q�-�{��X���O޼	o��l�%����%ު�p\��-G�۹�	�l$`/�K�� �e�|^L��_V[��(���L�6}2�	�j�6�zX��?g��s���_z��\���J�+����h#����c�i�H����G�|��I{�·����ʉ�%�BA�yV��eT�]�v��ӛ��yl�� �&������!�b��E`=��n�? EZ��ǮaVm̩������	O��!�D���D���� ��4���7���xt����r�=JU���P��END�HF���������93��>����eI�n�D8�JS��_
������6-PY�F��ݶϬ��f����	��/u��H��C�Y:4�5-��Z3W1��4�΀�9���7��B
!֔[_�>[�&}��D�ڨ��x1�n��ު�L�2�+p�hD���@�}U6�#�8�N�����Mp�{�qF=���QN��&`}�A��#�y��MJcyv��L�����B���C.��Q���iP^#un�_�3�(k�Cx��u�R�̣m�T�R+3�*�x-�U�+�ȯ�h ����������
8��]�Z�9h?��Ƿl�r[p҄�R��}@��(�kHV�'�85����&��E "��=�!��h�mR:�vDvC�f���KOR�.�^Ru�� ϝ,>FG�w&0i��(��'�2�0b�ɼ���iʓttl?���
��G��Q�:��lۯ�Ra]��x����)����@CVS^�9�(� �A���r����Z���&Q�D�Y�˥ہy!}}*���na�l�	�B�I6����.��I�({�qС`�"q���$�%X�M������S��U�����y�a�Ӳ�ΑÆ��r�;�C��覐L�'y�*V��ƫ��;!xe�0{�<��~렐��:6��R=�u�V&�N��K}�<�9u-�j�_.�5����ل�F��2ӶMÙ;�Y �~�^�3��JL�(I&m��-w��/�2iLl
��E���7�����Z[B��V���i�ѧX.D�����F���Jc�ĵ�\\�t���h@�1V,�M��*� �E;9�cŒ0]�ؚF����~t*`�ࣧ�C"�PK�e��q��q��3��i���`�rfͷ[��$���f�59����[�O�%}��Iڄ"��t��}K��J?�MF冟TT��LHhH�d���k�ڱsk�WmSKn�x{�Cg]�`�RG͐�L]�Ty���1<��N�h�H��8��)��j��t�Sŭ�Q�^4n�'"GbB�-V�U
����9|����z�D��aD��@��bK��Ĝv����M�:^�Yw|��x%��8ֈL��-��_���>c��vd�Я�@n���3����\��I`�ϔ
����,���Q�2�������e��
��j�!_2�����6#?P$w�L����.� X��Ř����|	X�7���4�kl��T��1âK�h��Q6�<��7ױ3�<Df��Zg�DA"8#���y��.l���П�m޵��
3z�U����H�V��Vo�q@k�aY<K�o�%y�`��<���E�$*��<�m��o#�v���l����cL*�9E�����`;���[ߣd�D7b���?�1�{��4��4� ���"����*/�h������� �ݥ�
�$*?]��L��IR@��ʺ-��t7�9���a��]!Ҙ�/y�-�A�<qcƑ������߁�naw������Y;{���OB��Z��
���	��k��~ޱ�Ƃ��l���#�#}���V]#f��J�����Sa ���홑�f������i�0,�@9� �e~	���;9�"І^ޠl�n)�X�܋�^W������"�6����y�Qm"6�\�i�8B`S��KQ㭢3��})K|=��%
o���=͇3w�˚����g@�F�-�Jqۤ�m�lB�����o��S����3+"�޸���^u��U����k$�#�����.(r��\���^=���[$�7�Ad\c3�ہ/��.'^|��F����5f\5�}ij���܄�.��1qk��)�;}��ML�|X�8���R�H����v�b�qO<�এ?<.M�ʺXLք���\g�3e�]���C:�.0J�����(��u�gҚ���E�(���KSE�d�*�¾�ͩ�� ����
���g���t�к۟@�u�������_
d럩%�`�q�E��Y:ǰL��c�mA���u�F$����[�J|H��B������G��R*nܽ/�d�n)��ܡ�0��N �
miU�&���$cT]����'�[o�
��XfW�쭉^���I��C�J+��'ک�qm�C���Z�l��1�*�� �>P�E�)y4J�T��v�c�w�}{̾�� �Tկ+�n�#~4�C�=������R {�e�\��,�T���w>�r���V;B�4��*b��o�����Y�#X�_�-�ݤ�ֈ	+[�X"_/��a:<L �s
��������|ځV^0���]N_�������=StƼ����9�9�)c���B��Y��2쑑Ym��C`�!3���̔���������[��瘉����!�lm����SB�l.L4�a��
��Ou��w�����6{��o��x{��� �
�h_��>d3��s�2	i����e����r��/��`�E��(?��Z�ݱ��&���<O�e�F����g��Gȉ��4ٶ�'�D�h=��	V����Y�5O&$�L 8��!��'�� W��v�`��č��r"�PA�H�˞�����zd#y{O�
��[qo��.��o��~�
��b��Ɍ/CZ��*�d8�����1�����bգ�u	���`-l��T�T�]ᦉ�X&�Ju��H6N��1�,��]ӕ����f��B�[<�u�h%����z�c��0����X}�_���/��\�P��]�/���{�F<;��g���c�dd�n�l�Z��1���a��s�!��&�	̻ɞ�d,�ۭ�1�$�XwAm��#8�| ���㰆���.���+ ��`�7��X��a�^�3{疋�Yp��7��g���`4��c���ϥ��&&v����)^���~�mtPѵu�w��Q�"a��Ry.�B�2B��7C`�u߫E���qdA� g�����"����G�w�X���$��#��_vf��w����� ,)a�O�9�j<�I��}����J_�(�`�.���-�"����J�T?|/�`�όJ��|�mi.I���n
@��Oȅ����`�BJi]�;/k�(j��X���J��v�[O��j:�x�WFb���̀�K���h�ni́3��;G��.��e�^]��Ou͠�%���(���V@A���>O�˅�!�S}�'����@3�Z��+�r+�jDNB��q541P�3P�˞^A����VBΰ��ڒ�zv
]&P�R��P�P��>\Зy,����N��:=��D�X��nMd�e�82�"���Q�����-v�4�e�j>�a�	M�����s>C���A\,��������G�$h����_��wq�}�i�j V�.�2�kX�^C�k'�;Y���u���d����DM�"��_�L�@K'M<��1����x9�����lF�:z��-�b=?����N�-5Άq��x� �+Վ��2�|:�E4����$+5x �#�=���aE��2v7��S��n�,zG��&���k��6,�M���	���:�w�����;^�r�_�F�X��c��W 
�!�%aG�r8]��2Sŵ�� ��q�������� ]�}�=�"#qf�-�L;����Y��D/j$�H�������c"u�Hsln��������Xh*���$�&3	Ô�(������&g}(m'3�M���MΎ�V���0fc��9��(��q��h�$E0oT�!1X����G\1��}��3"�q��M'E�l�� 6|*=m�M�O-f�'��� ����Ʋ���ґ�v���I �#��9M��(�h��>�� 
��#��o�̝�� [u̝5j�� �,�;M.�k`��s��:\H����W�]���!���IB�oE���ȧ��|d�=���I.fk�_��!c�6@r����l������ר�L��U��>3��Q����T�A�����#ɲ,M��>���C^�gM�w�N!��)�犩�x��,�R5�QJ

2/Pۆ�C��h�p|��F.K&He�N���,e��u��S+��P`����n'�� �T�p��1��m���Dh`�󰻢�����L	�����'n'���k�/��eB�-����\��Z��2Y��҃{Q�vĝj�:�!*�o�p�n���}�]\��t������ZHQ�%7�&�{���B9�f�L8��\4�o��+_3
h��w4t[�$4�Fͧ���6"�c��<t�z���88�&���bG���%ۇ�Ĭ�=��u�e^�� �Z�O����Xx��A$��F2�ijFf3"#�IX+�Y��5��M���D�f�m�����n������,�k�>7�%����3+�.�٩;1ްbS��6"�<s�A�W~��M{N���]aS�ST�	y�9%jQ�W[(�������6L�`��XW��P�dV�5
5�7p�u�����q"VT���#��e�G(L�e�)�<�vu�]�6����fk�Y�_s\�x7ǈ��
�h�tw ����p��a0�s�~�q�Y����ۿ��WA�"��w��i���G㤾y��"�<F=%���fÖy�[���D��
n��ڟ��XT)�¥y<vk�9��p����(��$�Z�J���}�GR�@W����v�{-�4�I�Ye/ޢ	�H���"�/Z�C��t�z|Zoow�66��Nh��V������~`t�!yswBi�mمny�CN���'n�x{W�Ze�-��y#�c�{��γ�鉶��ѷH�j�p���z�8X�O3�)|i����fuSX�ј�Jk]��RZ��!����a=�=2߽�R�fD#�;b��o��T�|���v��
��0R��A�ʋd*��us-�U�nC���"�����+z� �]��xt�/=�v�*������o۱u���2ň�#q�Vi�Ll��F
lߊB�9e�P��]#꼑��Z͎��]���b�\M��/ϕ��겱E]!4>�ƫ�2�m��-6��0�w�ы)2ɳ�v�  �>>�ײ[�ݮY���9�$�J��1����A�sL�j^���G؟ ��5�
�PW�H�U p�l���4�[b�[�l%���S�RMg)�G�{�,.+t�@�Y�>*�OR T�;����lh��;���Ǉ�զv8oRM�*�v9B���3�
hܐ�S1n�ɏK��XIK�V����1m���b|N��S-�,���<07ԟ�e/�Vt�Dlp�G{��au��5j0&]'�:V�Da��7O�:K�8z�W!<�c���+hU�{��(������A�K�r�fV�t���X���Eüs��v��::}��l��b��O�=�XHz�gW�/(㮤H�EB�����ȳ����w/LcU�tO��<�t�^,i��ӡz�r�w�L5)B�--i�[˨0�m�]��*n�@H>����j��wk]����ߗu�T���8��:�s�˫sG�@���˛�&�;��
@�¤�{�v��pNa�&�2j��D0'*d��� �~D܏�3n �|@EI�0���!��l�^�`�L�gdР>��#c�}�k���#dĩ�������j��A(:�㋭��Ne��dPMg"_2���%��0R�����SU��C/ث0%a�`I>����u?�ib�{8�[�w��0�,H����/�4N�.�Qj2�ax�z�����j�����%s�1ڋ��2�i6�1���ђ��p/!���Rp^��ۅ�����K~��+�r���L�\t���R1d�Զ:sD��4�����\�79z�d��6�Kk��SZ�@ܡީ{�l���4B�vs(%������A�]����o����e�o�R���s�O��A`�e�ļ Nb0�o�X��-�0C2uN¨̯�{��H$7Đ�����
,��S���=�����t�3���b�-F������M��
�;�Rn.���Q>�����)r�!`ڹ�݆��<�~���2Ta3Iw��J�Z�V�ϥ +~c����|؈�# Ur�p�� �F���64�d��@�뉬H�Hn�S��F�Tkz�i���.�V6�9d�RD�B��09C���~ $�n��y��Uڬ`x�=UŦBd��q�󐺉hCѫ��d�&K�0�;���I������@��ǵ5H���������cٛW�lD%�'5�a��ʷ#��b�.�,IgTv�P���-|�b��6�)Im�<Xîʽ������5�`K�r(F<���a��_bqb��x5mPu�мE�:�Gm!�c�n���2���-�in��j�U�D�p���,�~�]�i�9L�a[u���
^��麶��A�-��5~&Uh0��y��F�Ϸ���::�nO^���!x�qg���ڥ�fP���P�n���.���eG�OB@�ǖOז`>]� :x��N�gN>b�C��M��]p�c�<Q|�����(�imgI��U��>g��S�����F�o�I�?��]dt�x��v��sج���mҼ5����֢u�>��H._�5p����4�y���7o1�;� �ri�D)���U��w}�2J;�,z�,��3�$�on}Of�L����I[{&f��u��Ww�";��3N�Ȅ��z��>*w�3/���َ�'�=n��9?l�L0�k�Oj_VÒ]����E4��݀�IC<=��A�/�
=SȢ��C�zr�/�����wG�c��#+�0!&?���aא��.L�}��җj0M��-ͷl�)�L��«�%������[)-"��X_+�ʨ�A��n/�J��x*^�Mܗ5+��cN��Y�?�1'g��_~�{�����Fq$�4��z�G�U������\�-?��.��PQ��^29T�+f� w�U�QZ�a_���EK�]]��� @.����HdX���8����b�7��w^���6��!q���D1�_��n8<�<��5yb�����4�~ fDMܦes�H�!}�ܺ�.@;"N���N���,��LRʿ=)���h�:Py��?e����Q�T�D�,NO�?�2F:{�ڧ�+6����&S6W�1���?���5�ov�L��^j�x�Tl3O�w�й�7Q�x�x�}w���
�b�a�dC�^�)���� V�mV�F:܁�ծ�d�WF����΋d�q)F`ь�u�D�h]��.�@��v�E3Qg�i���-�ѰZҟ�5~ѐS�(��7�A�2�*��Cm\$ͦ��׈��ڛ�}��t:<ks��' ������� �N=�W ��4Nq@� ������[��O�o*���2!���רS�9h���(���7����Z�S��c�@� ���@I�:&z#�B��f��O�\G?L�N���XO�`�n-!"���]�?�p��y�D�{���8� ���:g�c�tH7tnt5��΍��q���!��##��6\W��
��'\5��#�>�L#��Q�1q_�]1��ukz]�P��Y<�����vqd���ݒL5���4��%t��̱5�)y����%y������ 4*W���T|&%l����jG�Z>az$�.��6�딤��P���[���$g#45�B-T����i�N2🦻���v��B��#�~��Z����D�2�S�v��l�%ɪΏU/tQǑ�V����&�iĸ $�Mg�9��v�{P�����L�{W��"�-�w��s�B�H�A�9>�$&�y�0�z�je �<�/E�Jl���&���ꔋW$�/[��(i�ec?��x�f�y���Ɠ��?�ZL���=�%����^�V�D[n�A��L�;����-F�2�	���1��
{�
c��Uw-�n�9�E D�4��;��/��Y�l|s� \P�X�$$w�>�����\B�a41=0��5��ث����<��d7�N��)��(���e��3Q����z_ꅌ;K�Hx9}t�E��u���L�c��x�<|��hی���SVaZ�(��E  �2�@���u����wbRN'w��!
�c��� ����N2䄥7�B<Ӕ�Q&��T���ܤI���_z%V���RWr��/:QpgML��Z�pL��-��U��8?JYhb
�|(Ąc���sH�z� ��Y��H���X�s��-S�G"�ɍ�l*s�����P��k�t�W�̢��A:���<�='>��E�L�uz����Y5,����<t�^e��}��������c���)"F�o��>�K\�w���q",�S���kE�|����QZ孁�L���=����+_i4��T��Bh�Gf�k����%�Nz�Ѷ�D80P�9�^� 8�d��@�bq����0\�x\f|�]���]�#T��]��S|^W��%A�zLb��7I6g{�P�0X=s��1����&�ԡ �h�I��TE[Ʋ����\��[Na�1"h���"�%��n�iR t;(+�1�$d��F�N���ڭo	�T�g�����B��f| o�����,�ρ����e�:[�.���j�><>�t����2�}7h�16k����|joUS��5͍麩v*B�E��_0�
*�iŧÖZpm��K�p����w!���n>�u�.Q�f�x�^��>sT���p��n����O�`�#�1�B���6S=皬̸L��6ڢ`�`��Ly��[	� Ա%�&<����g~�iJ����xF�I�߆7� t>�];.���`��J��7�b׫���lV�M����~�
^�i���ьb=�{�Wǰ���C��,��'}����m�5T����9��7������V'�6ε�tV.)�C(��ԗ��dtb��uk3��M @b8$� �|�\;10��fk���D�?�䕍x|+Y�3�jP{�o�q�R���q�yTuB}�~~!�D7�z�:�͖�j���yU�?�
�k(����mS��߱\�TC~3�!��3_��	��{i���v���ZN�D�Y᧽Jd�m���>���|mt_�p�D7Qu�D�K��� ���6�����Nk7���hpnU�9#��T<ٵY�0�S�s�.�xvNq�n? r��مg'�A�B��;��n��G����r��^u�"V���Ĳ���G��ɅR�i{n�D�T�o�t���z�b�x���n�$����$��y���%�5g[�h�$.f`)Pz�n\5ׇo��VW�W�֓�T�{MK&��z}�C"�V�(��6a���cX1�(�
� a��Z1M/�GĴ��U.��.�]i����/Ǌy�!,G F�n�~f���1>dJ8M]�H���� :���g�q3�:�O������p���,r��{�9gQ+u �����[KEc�t����O��rȱz��FT�a�S�J��pf���\hDJ��Zx)J|SBh�J;^�NFZ�j�0E��+�F��_�o����j���[yO���ױ 9,ݧ�1�=LQ^U�J�Ft����q� ������3�X����ݔ=���'>��i���p"'����B���C�Đ����r�q	ံ���T��*Y�z�~b~K������?�CAv��ɭ-^�&�ɒ�K��~�Yx#�����A�;�)r-�&�qhٻ�B}Ю��bK*_�Ӽ�� ��G��� ���V�;T�Ō�ݰ�-R3�*�>�Ӭ/)������X"9�.��HZ���؇�9�����X>n������W�;��`�ֳ�ъ�ؠD*(,lve��"���'��ã��Q���m���L*�&�p�҄����peA���G�D�����4�Wuu�z��j�~��l*�r�Z�|�!ނ��q*Y]{��pʎ.O}D���~j!������y�)A������M�*x������\��v�J���SٹIYW޹�}�'THd��D��r��{V'|m�1[��t(��e�T�qŸ�{�a�]Ď�P�^�VS���!.�ÂR3|3:����,U�L\\w�i����"mQ��qWRख़���[�򎮲t�٦�3�FD� /3E��x�$a[M^.AZ����,�ۇ���t�v�����������z����OB�HW\Ne�C 6�a9�T��	g�_bE.�~{m�e�U4�l<�ؓ�tYؽ�T	/�!՟�,�"?��=S�@�$��`S�켭M����j}��d��j�;��D0����M�l{�֕�����B��=|�.��F���>q<)=��"L��C�C�j�P��+��/�\���b��Y3�5֜���[1�^(v������AD��]��"�%�B�|�--�@0��h(۪tfH�۱��+P�����QK�:S�uwf�"t`/熩u,%�+��~wQ�[:���0�]�;y/��_�Qgd�#1&�z���.#�U�&Js�@`����N�h��h�|F�,h��fo�aH��Vm@�uA�y�uܺ��
��\��A��x�w�����|��m���G&iK1�m���-w#w�U8	F�:E�!�#�Z�EӞ�d��yw����ϡ�Zw- U$v騑���	e�S�_q�N�fUr����h3�$GQn��`��*���li:�%?�q�(}?Q^93X}nioW	��$�N؃��
`�Ã�c��h��!���C!6����c@q�I�e]m���T��f��'[=��Kn$�9)	�{s��ƫ�l
ʣ�ٰ3����2��ܑ�>.ƛ�ǋ�3�|#��Ȁ$J�r�K�}��HK]ci3|��`�`�=����/����{�cB_����d#Q�z�\c��>�KU���8��FLo��84�ܨ��B_�)n�����c���-H�D1M����&l�$����Z���g|�qF#����(�򞜡�v��o6��*�c�Lҕ
�����%e(]�D ^��=)�6����� w� �r�K�8%_�i�b�P��t��>�ަ\�$'��.�,X�߹4��1�v�L(�������2�.\r(�%�{�{8�[�M})��Hᐺ5̞��I��x�l�ع�=ǈ�UR�;8�j0���ݟ8}ɪQ�s9�jÖ�VX��p%���K�Գ�k+�_�>8��&��>�m��� �E�ʕ�Gu@VĜ�M�T�_O��>�z?�����Nn�h�K�ٿsj��t���Mk}պ(�t��PYk�s/�r��#�]by#��C�� ���1��l':�k�ea�y��/�F�N���	 p����k��U8��ܶine.$�Y�h��R�2���ҟ��?�9�i;�(=�-�R,m諓,O���k����sZ8�3r^�||�	N�O@ņQjQQ ���Z!?cb|�`yX��\�7�֓�;صTdJx����:!P:�2]Z�]��
���/F��Ζd�x3CȆ�����x�@���s&tZ���;�X�HX����,|-;"�~���f(i��%�*���+��V�C0H��zM<���d���$�(j4����,ܽX6%�(�y�ޔ8��=
���\
M�"b�
l%U�D5+��z��� a�ؿ�A�����_�3S#3�"Lw�#-
w}����ֈ��	�<5�ˁ���'��-~��4x<K$K�3}0Y�����t\��j�����3�|����{��P72��)�"����^���
�=3�n�}NS&"�\.� ��Vʾ%s�;����yE�s�3�[Wc�ԯ�����A�����̛L�&��q��tїD���Vّlx�Ž:�6o��5����v���k��IN��1�K"�4v���!��A��(�L$
\��L^��nJ�*�%��;�bt��<O"�(F�΁-�7.���tC��+6wQ�l �̻�L\�Bᒭ<~\��S�󜚌\�l܉�V�q��¹s��o+�>�)
@?�=��/��c@�gp����7|�_�d!Ct+�q���"���p,�NKjB/4�)�QFB�t�k
X�~�*p��/.T�yGn0��I��B �08�=�SZ�j��ԸU�x�^�s��y��Ĉ��rg��9ZG+�� �U�zc�_<ٛ�`�K�w�e�ұ�Ʒg��=�e~S�ӓS�yx�j9���6���['�4۾
G˦�S�?9΀Gc�������:Z��%n�gVYE�Ҥ����l$�bv�Ԙ��ܟ����4�cy���@�@OZӲ_)�A����/5>ư�F_p�j9�`��*��$���Y����<�E�g~C��z�����>(j,�T�Pjr� z��QBL���w�<Ç�s�;P�4ܥM����� �q�\����ↀ��m�J���㦼c��!��֋9N�W�m��B����A����G�������� �����޴k�ċ#њ��v⟨�8�� u��6A���4H^��N,a%���υ���`�Zr3tC�u'>'�bO�t!*�N��Êw?�� �B��.q~ظ~3�B"Yd�E=ָ�&X�m<N���W����򿣁�a�i������zb���d�T�S���@HW)��	��K�
����Z�(�!sr@0����Ey'/ �Z�Q�q����#�,||h�=�� ��ı��2��������a���3�((����;qR~��?�t�?*����V,ZR��J���3ЫҪ��-N^g��}�cO��+K��*$q� .G�.�W f��r�b-PD���9 ��Zxvmܾ�Gl�g�h��}�X��{\Ȓ�o�;�b����>\�rQ�,��b$�{����8� ;)
��{d�@h�GM�(�V:�����:Ŏ���AV�X�W�_�]x�yq^��8�zC���uÿ��E�]��Hk�n��c�Y��5܋W��u�d��_��Pm��U�өJ� �/�J��g�6�mL����蔈��Ѳ�45�{k���s�:�Wb�e<�aޔ_��WX6�����\���X $�6wI�zr��Q�6�D@������3:Xx�ÿI����C� �ĸځ��IL���d�4 ���B^ '����g�Ö�+����q��}
�Tτ@�(ðt��%{�
�T*�}���j7�A�3��J^3�8Z�2`�U̳���F�o�_�k��y�S��$���sB�8\Ӑŏ�8��W�,�����K�'�3��ѧ6�+n����N)ܸ�X��2ie	�� Y'���h�S��'�X ��øo�qW�Dt`DO$���8�kE�|Ye���!�&���b���5"�}��K�����؏V���,$��V�cP�a��l�����9��/��3�5��݈�&�<�D6���-.���AC�E!f�H���g��/��4~�4����ysq����5\ܤ�s���upu-H����;я���ο�>I�.���q� t!�K&���o���e6�i�ު��d���㨇N��w�n-��JQ��ٜ�	�OAe�x�=������}N�OU��#7�ga��G��	�� �U���I��[���*��xҞJ���
}l
���� �HX�$��k����Y�2��ɣ��&�Qrh�f�l�g�TV�7��01-�7�W��K'NB`��Od��~���P?���}����C�,4�������K�2����U�8�W�D0�<Z;V��"�+�C�;8#�t��@�Bw/����t�f&�U��0���s+���{7s������oe����������,�� ���^#�cq�p0���!��la7a�m�>�c�Vߵ�{�F˙@����!R����p�$���=���R��iv��
���M�ǚ�cЛ)���S�Bq��NǇ"�v��`�3�dg(�^�������������@��ϲ�n4.h�Ǌя"�	��S�Ѝ�!\���l�F�^n�b��]8)�aL"��˃��o��-�d04NѦ꘤IOJ>#�S�B}pw�d��Q�K��R)q=�U��!�g#��e�>6pu�M5m��2����
٭�S�ј81�S�5�H�|��fC{��|�(Xmt%��N�WИ���a�����х�����Uo2�� A�d>b�:���}~�Qw�x��("����3q���YYYo�8�b���=�>]�x7�P��RRFwF�?f��R��Vp2N2�o�q_�v��隉c�!O�@h�Pr?Տ�QR�R;�;*45j�@JV>��Y7�޷��ԹX�{�nQ���6vK�ӄ��VEN�j$���=82�~�K%��a�s�-{�4�J�>3��.f���˒�o	*�u���3�g�u%%
�9/F4�� |z\6��f>����I.sa$���u� FA�f��"��[�C d��+�"�&�(�~��K��f�oxX����/.r[S�C[�W�i8�.��\�↨��Vk+dU�
��µ8+;��8/���Ū��ҷn1d67b���.�,���Bӽ�x��W	U�e�)z%�6�3�Q��K��<�f�RDi��Ƹ��Bi��->ł��a� �j ="z$ tx�`U�C"r&��D��w' Gz��ӽ�2<��\�.�R_�����ݭ8��>P*�4KDQ#dx��d�	I���5*=Dio)5�`*&i�V��]��j��Q�v����݄:9�
��Ƌ������ ��Z����EU=(tf�̞G�z
�%����Y���}�z	��G����rãҕ�{��Y�͸/I�J �*_.R� q���L��h|������j`;�)֥������SIyF-��H�Y��&�4BI�(��խox�������3,�q	�Ě�LL�GׯK����UH�E��[�Ǣ�<�q�ă�ΰ��Dޢ\#;e��|�Ǡx��S�ȃ�"��{.�˽��kxeCd.'��3"8�R� ���#*R?a	Jo��ٹ)I�٤u�=������S"}eu}�>E��7n�2�݄Nv�-#��~rˇN���8k�rR˻n^��_��
���35����Êv ��m}�����=A��0�{���~7�j'��D$; �7-!���^(G�����=7���)�F��3l�Rx��b�^�3" ۋ����8.���v/y��8�W��+м�Z!�#:b%Q�,����؝���#�d}**�LH5�F�y8^8�/2��V ������閱�EX��V�������f}LYOW ����O��.��p
��"���Ю��}ї�DuA��U���Ir��������i�Z'�������{q~��ɠ%�'
"�)���2���i9Զ�,���]I�3\Twx���gu�M=����%�܁�g8��֟��)EзAh�p�u�����Y�	":D����Q�/����u5�M���;G�wx�wɦ�'E;�m9�M���v�?�ag��G�i�2Ŗ�����¿�C�Jk�¬&�8W��V����U�	L�,�����eg q�I!;���Q�w (��9�'��3xbU-��HI6�ca��^��gLT�*?�m���Mi�b��㜖��ʖn`bu��ȯl�-�3��v��p�	�;���ENRt�Â�ٵ��k���;��ʲ�ӶA���$C/3��莽�*���KzV���i�JJ�`��qJ�ʌOi��+��7M�������F������8�U�-����7ѳB�O�9�J���,ȍh1��#s*�o�����x��T�Aqz<턻����!��-.|5�?�s!����e�j���mA"f?L#E�S�IFN��N�;N�	�Bg��ЙIJam�"����*���@l�O!����dPI~^�J �ʞ�-;<��l�"o{d1��c_�rp�p�)����tو}.�]��YK��Qz3��]bw:�Vl�A~����F	VU��C;��)p�g�zh��e���6���6��D��f�me���(P���zU��#��(|��_7L'��p��E�~B��'l�3l��cؘ�c�!ڵ�Uy�kO��+�qy��k�lC��zI���A���� E���Y��1kJ�\(f¼z�۴�G�L�`�~7����崝A���ي�����6��@��=�{��I
�Zs�e�>��'Ldm��	TN�DO�=�M�i�CŐ�>��1�qU�rL�R��6�m��Y5�~�4p�Q�v}ď��Ҫ���U/aƻQ3]��I�2��߮{���20ޤ?%�!ܯ;��A����NoY��C`�/T�qk:���M�lQ��D����$��]�����Sg+�[b`g(V�J�y�g��5�	aTcY�ᶀ:m�i]kQ辛4F�YN�S"}7��!py�|f��r]��X��C^e9;(��Ѽ�W�>@˃Ͳ�QZ�K=l�t/��5g��n+��W��6�TO���a�*VaSc���Aťb�(zN��~DYŒ�ǔ��j��>`0����Un�Q8W���`s�v�o��+���	�������L�5D�C��;��)8�Q�1;�,h��q�0d';u�=����F���j!�
�z]�@h���T�z�\K��c�G��0�_�zb��\eg��f�d���Tߣ�eB�Kժ���quW�g�^i'�߯�6�ϫ@�h��Evi� z�En�xzF��;��ag�onߴȕx:��$~1�2�V^Z,���<��yaK�A���A�w�*W?�矶˸)�n.Ir���,J�;uQY?vK+�o�"��r��3�W�����g`%Ç�dS�Ph���	�C�&�-��	��,����2N�I쇩@�Vp����\���Ӎ��-��`a�q�*�TZ�X��o�@r|�hĦC�a��ORrdT<�s{+��-�-�I	`y�G�Ti�a1��G�<�5��o�+�Q��
��-����s$���M��y?��?\q��`�"Yܓ���T��z�O"��oơi[���bz"V#��$���/i�>ʸZ��)�����վM]�ȷ��ُO���J���=�Y�B���D���%��"��%��#�7�}����i���x��A�%q{��A�}f�*�_K~,��1*��<�$����:���.?i���=�6���=Y��`?Èq�����Q�vW�r�ˉ��C�g�ک�>�\[�EN����B����'�����|�=c����,�L�Q����zq�E�j$`NHb�to~�e���sIDI�a������1=�@B@�����2�-Y�Z�dN5�*���b$wU\T�+S��,��G�0���Oʁ�5��9�b/M�&����G��<���t�3i	��:�}�'Yxϕ:�:�����\[�:�(NC�����X~봝��� �q���(]>�y�~�"�eZ�o�JY�7���<�7Y�q��D��5#/>GVF�(�����Z�D��l�S@���Tu�p=3��(�ȗх�|�[�ۄ��όO���}C3 ��v�$f�e݁�f�Wp��.M�������[�E��>�%�-�8(�-tJ��~���qZL�$��L�By�mB���\�A<��N��hߏ�~�uP]W<���5R:+��+	B;��<NITJ��/�B��H^�#������v��Fr^�\�8ܖ�"��ǖY[�5��4cB������|�8���>x梥3%W�;Djc�j��Л��ί���M3�P~�Z�����Gh�e����/�l�s\4J�."�����4W3\le��~:�� �����4XW�]Oa� �2���	"���0��E`֑�����P�QMU���-���i�j��k'��%D|І�g��Ι?�*x��g��B��'uz���;��.�lPuIy��y�偎����1q�1
۶p
�eѭ�d�nE�WA3�ۿ��@��OǶ�~�/����M���ɳci���j.����=�3��ߣ'\���|P��&W����a���oXU���_�L�k0ź�6�Bm{Ĕ��i!�AXD�3��;QH��� �
tW���:1n�e*�E�[Ddc���3��M^ _l0>1���a���v���E��כ4�u��},gݾH���T����
�9���H��KƵ��t��x[�b!�Q��au�c��>S�"�=��0����E�>0��f���c33�lez+`�9��wmLh������c�����9Ë$9w��g�~�k�V��r(�M�Z�K����ha�K�O���DZ��@x=a�� �3�k��Ļ��G��C� �S.0�"�Q��9�����C�?0�^�:gD�e�EVRJP>�|H�L�=��sD%��"�bC�b4w��{Hί�j*g��$+r$��R�|�*��x�J��b�b%6hj��y�����f�<l)��}�\�@��W���ZˉV!ku�i,��:��T̨��y���ӟq��"]��V�~�eM��]t����ןl0ǀ�\��v9lc[3揣���N��!��M^R��,L�PY'��d��Md�L
��:6U���w��BVC����`�E��4a�ͅ� D'EJ�nZJ5*a���.lr�ݓ��Φ\U�hp̅�\����dr@{_�0����!��kh�^�6v��V�z�k%�ŝ=�'Y�qem���n7&UV�?�.�T��,OO�L	�x�4Hlb�/�W�6������˙G�.]oáe�I�s��آL�b��勛(LZ��s�k&�F,��]*��(eҰT�'�ߗ�W�}s�3�K���&�ZI�`�	Wgφ-`���[��#���+����`s"�q�w��;�z\Du�!YAf���EB+�#��(��3{l�2������^J��|��J�^���Y�,�2�eZ'p��P/W9�©��J��=������H;�+#	��0v��X�yb{-|<�;[��#�&����ʆ������j>�����]�`UM:m��e��p-�Y��R�,re�\��{���9��pp�ļ���Ǒ�hR�K8g���pڋҎ���yY���1�0�TI���Ftv+gojt�����h�Uj�c����t'�iHx���!v:���eA���^��[-4J�I5�6�M}<�߭dV"!i�Wp>i�QeDu6i��z̏#�};���9��z�>\����+a� �>Q�X�Gb��qR��d>Ϗ9�����N����T�o�����e����i&6�Z
c<�ݏv&�-q�m�^��6r�C�QDr�P)�(Nq�]��/�Z.�"�3��(]�jA���q����x�\j.]Fob��#A�í���r��t���̫��|6�9n��_R�n�X�,Gf��rhe*Yj��s��ɿhtIϣZ�WP�Z�j6�O��mU����i�e��a@�6ȟ�[mQ�ղ�v[�-�U�J�'��(�	B y���v��1'�����|X�wd ��͙���\��nP~��VE��A%�bc4)�Δ���ߋ��˥�5"�_e>�>����Z8���5q?G}>ly#{�M{"�	FyJT��7��D��n�t&�J6
�^�k���Oŧ�x���Ԣ�~8+>��5|����ح��]d�(���.u��d-��������4�Yy_D�9�=ݺ�b�{Y��29���=�+��l`���-|��E�ےN}�Y� �����Ĉ�\�!p�Q}9����� Jn��+;]ń,e��L��a��@?�'�h  ���9�A��KAmP�z�".�W$@��]]"����3�'3���}02������9���=l�e�����f��47��JQ%h���7pH��E�ɯM�-��Û�� �\9[!��3@~��
J��E[L__Ϯa�?h��<���Ca^�_'���s^W2�	`�Gt����u�K�q ����Sy�o��|v4A�Hr!0Ƈ(�Ja�����v<��6�(��$K6L�p��j�-r��R�+����h�R �R���Z�	ejh�O��G{{H�3�����bV�ga������S�[Iqo��� 9����>�C��f!�����"��5!�ۢ��@� �>F�ؔ�D,;J}���`�*(/ݶX�J_�������lҾƃ�#�'��?$xH�'4�a��}�i��Z�t����Ö���5F��>�I���&.nt~��3Y��N����;��� R@���)��p0rQ:f}�C��y���k��]K���U�q?#�
�_fz{�N�D���|4� ��g7 ֧�'�}�5���W^b����q&� ]4O���'g"l5QF!��	eU�9*s�~e�N�/���
�whsUHw_���KA��cU�To:�l�[�c���@��j���B1O(�}��;uc`x���Վήz�YU���T��Sw?���fIi��0�+��� y�4�+cۯ#���������]���wF��s
�C��E<�rs��F���,��D �|.�M��6y��]}�Z̓���TK�`���uT�.[�)f�!V��e��䝂�8ϔ�)��B���xߊ�����$1��s�:2�ַ�K<���hd?��JĤ���w��8Yy���H��w'���6'+��{Gn���\6��dkd��eBu}�H��&��L0UW�u�5��vmy?���@���ѣ:��E��@A���U�WV�%o��C��DRӧ�P��Z�t��� ����]���0�Br}C`���RYYv�R����Jw]�4�_;ͩ1�*��C��u���ïR�T�v�u�/�sˏ��G#]Y����� F��I��Z�=z�5����&��W�{�RF枲n�ԓ>�}�G���j��R�]P�0�ط�)jG)5՗\-�A���|P�9b4Xm��L��TN�n��Y�>�(+:f�A��S��?���9��l��(�pH@%~�[�����"�e�[��i��t�Wv��	��,;#� Ҁ�),9,ߢ�n_kW/q񧽝\-����'T�-D^A@o����!�,��&���T�x�n�3��Q�e�yA��u�|x�E���᧕#]�[|5���c�2V��OW.��aJ�Ly��C�����X�ƻ����f� �V���9Xw�T��ӹ�،	avBTq !D�TK���E��cw��Q��4�݊��b#g�I>�#�C���e1l���n�F����]ÿ�X�!�=��&	`��hj��up?��xDg�`�ލQm�T��/p���p�%�tD��1H�ba�ݢ�u�=&�/MJ�h�':W�z�cD��NQ):>��~M��Ӝ!.��2��YN�73����-���g����2U�;���>��]�vp/d�>d#�3~N����L�j�qu�����!I��N�|��3G�7C��q�/�ʀ2�D�������#"Y��6���k�&��f�+@�(��ߟ|3��/�ɯ��$��X�EC_�"�~F��.��P��1t��YH� �a�u	�o@,<��k�����Ѯ�q��`��op#�^ :�Ԅ�%㰚".RKI\~p������u���phQ� �?�V?�Sqp*��ҦW6]�gG�FØ؅+�m	z_n �;\�Rc*!�l�6ot(	�]HMK�L{�"e�����ЗT?�s�C��ѬH��% cm�*�:8��W�c����:�͘�B��޸��s�U_�
e.MSM���BS����m^Xg@��Pө��<9t��{Lj��r��ѵ�cpc�Qd��;-����<Lc^|G��vR=����8�	��fRS��?�,�R8��	n�T���L����&?���!�8v�3P�J�B1��)_\ p�MQ ����Pg U���2Q<�� ,��3ٮ��6��HB�B��C��#�T�?�|a���W��IP���_���&��5�=R,@`��|(��yR�=�«���������}d��� �0��hr���	o��+�-���T�s5���(���{8���ѕL�6���rh���K	�5�����)��ō�E"O��
bt^��l�W��=��;h����o ���/2U���zK\N��Y�1yq����eg
��6=��ZD;�z+>��������KQ��_`�l�oo.�f�"���F@�[2Ѡu@���Aؑ$�ߝ?R�,G�80'D�&�Y�C��d��`T�G���o�� �y �/��<)jwmJ�[1���֝�J�[�)�^� %�]!,�Wβ���8axC�.��l 0P�Q<A@ɣ�a�{6z�����ާh��G�3@�\:��	K�7ۈ�W��;����ͣ�
B3�A�|����w`��{��쟱T�I9U�'U�;ी�姛z�mG�P/@�=�Z�XWJ��3R�E�~�P>��
�u��4��l��9ǿO1�2�ܫ�%Q��=��"bV(o%{���fM�h�0�|Wk���4}�@�y\��iz��T�|oT��j�k���[�w���U+/��a���2@&òI�0���MF�^�.:mC�;s�E��B8'^��j���|�(Bu�х�z`o�k���B2h�]��ۙ��]��5���^J�男����M(/c �:V���Ğ�l�OI�5�t�0���c����Qndt�%g:ވЙ�2O>�J�Yn�Ϛ�%#J�,��:B��(�.9�j�����]�4��p���`Ϳ0�N�v~=�m��~���S�}�ha�/��ԋv������)��ީ�x�������I�2��ա�枴>��a�X��qk����X�k�-�V�ؗ�\�9����2��U:"<�eﲳ�̂Ip�wC\7��
�NT�2���a�wg��ӗ���<+����x��N�ɱʮ��Y�����N!�	j�Jp�}�ܗ�:;XVYp��a��Ԝ�R�C�Q��O����B�"�E�hx���`q�&e���T�@�������j���/�� 	�Y����d_����6ͽ!��� �#�N��!io�����tS��+v&��
�H8�i�����\�����5ʶ�S��qO�
��LH{4|I��)��҆<���d�t����v�Q�F��E���|z�6j-�H��5�o��%U&,����E͡s��%�E���z�:x^\���2�O���?��CEky_��v�l�@<}5�0�+'s�j�FI��<�CJ+��8�'�^��ƆW�/~����3M�es-�o�\�fMW�*��;N#����$�68K��O;i]8���>Z_��N�º9,#��%� �
zܹY��
���0�	y��	�r�|��βֲ��/�p(x��A�p��Á.Z�o��a���2�aL+`~�j����4�/4���f�Ah��n\�n3�f����==�Lbi���4�Y�C�O'!����:h�<͚���_X�8��Eb�/I�D��GXU�x)��0����NۏX�p���Z���r�[�	io�ߜ�l���#�GЃ�����sŻ������ �ٯAwzӘ&p�
��j�8��Hg�^�|��\B�T!��mb�Zb�P�{6;�Nv���������d	���o��4�!��(&岔��S�OC	p�	ѵ�(7�d8�x}j?�����5�K�����}��.�?��D�7�������gl�R�Be���뮦rӬrN]�L�£��;��F�z�TQ�o�s����i�TY�����t���т�����Zm7�q��)�V?�� )D���R��Z��L
�R��p�!r��வ�ꎼ5.W��B����/!���H��H�8�}mezpO~�����U3����U��� `RX���Ͷ��r>�5��E�!��ߵ.�Q!�8</�+iA7ltݜ2�����N�S��#��PDI���g�A:���[7�tH��y��컞�'��F�Ĥ�5�fdt�b�]���!�w��ct�a�_O�HX�C�$LO��;:��.f.^��&��r�b��%ʲ��U������>�'�@Ŕi���Vlc��%�1P�m\T����a����h|\h�ᑣ�����^�<<HI������#�F����9Xm�����G�s��5� �k��;�������U�@�z)����ù���^����-n.Hv���#���z2����h����X�2v�Ó��{q��k�~�^zh�-�D+��HH�|h���{���\�9`x��c��(W�����-p��r�v�6�|Z���mt/���֞�"�o疽W��fQ$��!�KlP�T�Q~����+�%������%RT&����5K)>��NO�>�ǥ���5���7ua���-dS����
�����j܌"�pl:g��c4���d�,-�w��2 ��}���V��uHD<��%�J����g���Ɲ%�S_�S&/AuϪ��4e�C�����\/.M��B�eX����K�Gn�W��I2��D*���hls�m�;��T�M�n�r�zy�"8ulA���Hv�A��_�4+��A<j�>M��A"��[�`'��Jٰ������BE�ܚ'���u*�4�?U��f`���m�S�~�B��������*��w�u}��v��O��mݩOBaj�B5��駏S�V��uF(�qߠ����L=�R��C�t�u2Q����5�w[�s�X�"�.!�E.��F��9�����G�z��݇�ij7�m�?��{I����o�Q�WRo=$tҁm�]�uo�i�|�pJ����L*��ђω����U�D��J�e��r��2I�g�Hg�j�My ������aUΜ�{7��P��s��\�XY���.�S��M���㖱��yA0�y2�+-�r�oY�J��F���Z���Y��Sv2<Ґ�mx�� Qö� ��5��Q�(�sr�E5
cz�݊p�����M̑���> NR�!V�Q�No�'�z$5��?Uw���#�\G��P�"��S����!^������s�7t�x��A=�2���~�½K^�Si�:2@��3���v��[�5��/?3�V�9� Q"� �&@�������4&�u��d�)�
�tB���5ݮJLx�8>�)�0��S���»Çۆ.��J�D�?��.+H������ղ�����^�(��-`��f³�a`#�n�2�]�;1D3'�$��8S&xf<K�;��cU���N�%�������I����=hVk������ث�}����2U��ju��{�mR��n�X!���Q ;�#Gtٰ�pD4��
�$ۂz�X���m�v��Z����L$z #g�ևf����W�[�����2H2���K�{Rv6��ܾ{��;}�ʈ�_ϥ��.�{��6��U����P��<��n�i��ċ�����7�!�D��R@d�̽뒂G��@"�&|�]�@i���N �\�J�3�v�N�(�3���a#l�zn5I�7`��GBפ.?2(1�6Q�h�G�[�Ҳ�+(�����A�#�u��M���*~s���bE	���B�ev���wZlE^vgzœ�����nH]J��)cM�9m�,+���H�L��W�ت+zF�Rs�$��u%��L���/o&ø��*�`/ Q��P�5iE����B٬�D7�PsPF>������T놁/���ۺl�v��^c?��%�� r!q�~���/�	'ʂ�ܞ����|gu	m6�U��΃��`��Y��}e�_]��"ꅬѝʤ&W`p�1�7�Q�1�,ྴc��o���1;��;S�B6��U,yJw�
A�~_���6���6<y0��ٵ�6��&��C3�88T	�pj7���;&��n��N*P��!��b?7��|�8/(z�9
��1���5j\��w�apn�u��r�P�%S��#�C<����Tit�뱒
f�!�JUi��w\�c�DM�/y�Ŕ:)¤��4ѷ�~��a������|��k@M�W*�5$v*���3�����)֕���鱑H&��&�kR%��`��gS������XT��_n�����ZXR��*�2{@s�_ᨳ�.&�M<ym�n�@��V�"F*�x�P:OPl�n��� �� BU![�閃(^�e�8+�⾓�k�ȥ�U&n��Yy�3�KY��ta��=nɂ�S��D�=�-2M<��3��|#�;���~gB�;W߬,NM���G�&-Ă��~?�,���ʖ
O�g��"��U�K��*��B�k�R+�}�
[/��V^mM�Q����<|�����O)H�\�Z�xuɇ���3��[a�4�\4�U�Ӑ�)s�?׃��C
DH@��?��I,��p������ '�LAT�av}��r�G�l������ql�n�������j���;q��>�G�Aͅ��f~�`��oA����#!��ǧNEN�%��A��/�Q�VB3\�EDZ�(������&ʻ����26��qb�iо�@P0���mPzI�ec䵒oᯠ\���l�J-�@�UIx�ޔ�����l��2�4v��T�ϧ��:�Q4w4����>�*�H#a�r�� �q �ډ%"�a"���BTY��gN9gQ��&p�;A2�/yp�GI؄9�^6v$-� X`�V���.N�M�x�V�s4�8`K���<�J#�__)�'�8�MM��V���1ћe�A����^�v"��k�C 0���a�;i�ec�f+�}�(q��X��`n�>��5A~=�-����o��:�*�	�x0���q���p�%�&�Ϲ�|c6�L��b��)�e � �da��p�j�d�ZG�%�1�cX�*?׻[�c�j٪ ��0r�}H�E��H�'_�V��W��WW�a��gG����k}�Xu*8�:]�ل{.m�*������J���hW�7yEP�ī�
ц��IY�PV�V��a	��P��g�^'*�杉	�樂b{���=���b�C4p`Q���[�2(���f5P��_N���2$u�A�(�d`�wVZ����d��H����^-���Gm�K���r��/~�y��#��c�%��� 8�]�Zq��R7�V2c�)y�B�����=��O� �?3�$�����.1:�g��0���Q�����*W����w����L�:���-O�#�p�"��$i諘>���]��\h����Y7N)�B�����^c�\F6V��μ�U��*�+��QXV1����>���X�:7��A~��p�UjF��w����*�q����45d�Ư���*��e)U�S&��b��k�ݢ!
��*��p�L68����3�]���>���ǒ˓&�,�*`��\��%��F�FmK��8(�G��=c�_�B%���w9�_蔑��5��$2{��N�f[�Y��W5�C���gc����0�Y�,:O%�]&:���H77p���HKo�%#��
4���1:f���^�'��,��_<��$׌�5�hI�jl�h�VX�{���Kz�`ť=<�Ɲ�R��E8�U���­M�Xu%�#N�1�*vszj��h%)`���.S4���3����H����hS�7�NU|*4ݜ�|�:F�EPe�(�H�����m���(�*soz��|��I�%���Ӊ���l!�ً����|]�i�������w�����A���w����[�y��<#�!�q�l;�����'�K޾��S��(RN�~9F��cI��]��2���y�e_n"ݍ-��Bu�6܈؛&��k����}��p�qoVC�3A�o�?��G=�tRɦFwl�W�Г��\x�|� >��ڧ�b�Gv�-`�Ѫq���ή}O�,n�ie�l������j@�ok��ܶ���C!�\������Weɺ��x�tD� ^۶��Ԡ?�0�(h?K�:��-cT�bX+�Y��7�j�3P��#Q���9|&��ׇ�2��C����!Q�D8����d�P���s� ��N�]+~Gnm|�񼍮��C88>Zj�i��y��Õ��p����@gŷT��A�2jO�$���`�j1$E���k7��KV�|D�5�pd6e�Qԟ�iK/�b���+Ño7�N�du��<H7�@��84��	���޽����]�^"W]�F����W�9�O���F�k��W��ŲJ���Y_ؓ��SΡ��M��o���i����*̓�{��/,3�'�f�1F���C�]����]��W��S}�cX�v����C/ ȴOW��#��C�szS~0��p����H_����}5�|_��@[�1��Yx���3�����1I�t�_��r#���ؒ�J\E,��㠱���;+��G�}����M�n~D�aЕ���q��3��0k[���\��1��M���О4�#!�<�b��,�ŕ�^�L#8������+���T`��C�S�ƙ�Bo���1�2n�M���}�I�����j�]�Q0��ë��.������IS�4�Z�wfɮ���������������?�5�R�pZ�̈́��Bܗ= ?��f�_��߈��0'�~)���;��.#�Z�ۦCX+ۯ�2���0�L���u����l���jݲE8~a�B殜�O�3<E� p&S)�s�^Y!%ҫ�u��'q��a�� �=Ɔ]xK�Mgh�/�1���m���޻��EB�`<o{��������q531jE*���2Q�]ן���*�[������M�jp�O��(Z7�^��?Oy<�z�G��Fq�&��e>��_ew�P���'	h��y8���6)�7��������e>�.Z�(�}\'K����~9P�鸬�
�������\P:Y��m�"8T��)�����(W�'ز�y�|#Uא5�7��be:$׭�4���W�C�u�e����M!��"<��8Ɯ^�E��*�k�F��^X��^r�s��|�D����J�elF8��1��D��MpWV�i�55ʶI�Ba_el�y"���vO0�E�uɄSU��O���n���}�P��v˝9�c�.En���<�X��QE�����'{��6)v��J�C'�jֲ�9�D�}N*��9���>K���5� ��!?�v��t����d\D��H2����&�������A1I�L�W�V���[u|qR��ٯ?��?\f��:��b�O*���㞹����l��y�)�)��܇����:C���,�m�
_٬όü	}�h\�~�
�Rf5�`����gr�n�G�L���a&�~�0׺�{���VU[��H�I������Ӡw��1�ݜ��X�=��[|m�Zz_Z'���A�2����:ɬ~G� �[Y�9�^*����i�� 1� �RL+�p��u$#*��D���w|w��8�d�Z`�`?�V?8*;B�M	��+x��'rD*�B�� &�	���b�S%�dONTE�R��s^���A5Os���lQ�#�9�s\J�G��'�M1?�8^�!R>�mW4�O�Β�����w�Բ�o|ӌ]�,d��H4���� �P���E�+��b�4�D���ڐ�P\\�WI���ԣ��)��l��Q���#�w+�Op��V����Lz�wX�3�e�#f0�V�57ɰ�;�:e;&� �M�xԒ���o�ҿ??|(QI8��=S�m[�z��K�gB�!�s&�TZ?np�tO����&s��-b��nҦ��I�#��ڡyG�cԙ�Z.I�e	'y����IŠ$2K 3�#$8��AM_w��/�����\�U�㮟�C�;J���;8(�PH+kX��&���ʩ�ɔ�gTSO���B���]q��]��$2_t�Թ��Z�;���e�y��$�qm��}Ͳ��T
D�z*��G ?�^�lS��;�8Œ�r�[�J�8D��m�O���#vp�u��,�+�MԀ�b�m���Ld^$���1��%4�r~RbA� v��֨��̗OT�3����'�E�*�������l���E��h�Y���� �;��6�Ĺ����,\7F�*kI�|ı+������-c�J��d˼����8y��8�H���/��P�Mi�3{[Y
��5��~K��,e�fc����;��;���V U�ġ��&ȶ��7d�3���������UQ^��}�TH��r�Zb.E�ϕ�1#���ҋ]� �f5�#)���^��8�Y(I"Q��bU�.�&d�J�(~�r��]Bb�%��l���1��c_䁄�'�63����Ǟ��_����1��V��ŕ�M�Q# ���Rɰ�9��Um���O�s��ԕ}]����&E�0�
��� �ن�c��!�x%�$�rVe�\-w2.��)eJDj�;ЀO��p�vT^���s�!��q�俛}{i*Y�P��!�����}�0��i7n���AN��J�+	8PF
}��-��X�?�K�BX�5u_ �L����:_z�߼r�p�3��~y+�h#�J�!{�U�xw�X���8& D�{�����ςYm�q��M �Gl�8�Db�Ǌ����l^��R�C'xTy���$j���#���qTZT�6LD�I֚,7ʠ1zV������Yj���rQP#,w���r��H��eZl�ؑÓ�D�]tn:sP�*Jr �̴���P��&�Ʉ��z�6|��P��n��N�3�!�����'a!�g��ίJ��c���ZoP� �5[��"b��l ^�Uu4_%n�8��J���9�@Rc��%��_䈐j��"�M}g�˽?��7+���G�9���E��fl�2&|:���S*�h��)֏�����kY��/��\dX}���C��k�4�`b��P�o	��(��m&�c����'� 7s���ٻ���z�In�ls���[&�<{�����L޼�2���3�J�"���ָ��	g=�3i+��@����I��*�R1L�&o,����g�W��>pYRM�Ѩ���������rpf�X�V��I8J��i�3��R�ְjI�'o'�$��c`��8#P���9wL�����H�2S�%I��.���%ɰ��ȉ:W�mO�{���Δ�)2p��4Bc��ݐ��Z&UH�*��:���q9�`�+�_�y��Y��?��0�)���а�OԂrG?��v��/?W	���`EȞQd����P@>�OR��rM/���!Y��uI�̣�G���|IP#�Xl������r� ��/^J��:W\+��"�Z�	p�hu	'�lS���k��˷6�:�@��b�ϕ}w��L�!.�P��W����@��6����[�ġ�BBj[��d�A.��qx9���')=C]A��x�Ѐ��7���2/�W�5��:��@�Z'"�T��