��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1���e}ʲ��cg�t�ϙ�a�:�KR�%���ݧw���ȼ�iV�� ���<jՒN���\�MN+{D���TF��;U�RB�K-����N.]�u�^�SɆ��8���ζmC���x�V1��?�F���)�Q	1����i;)�)"!]h���EA����*Ŭݦ��k w`�,?d9#���=���?��^��m���j�!F�> �b���Wn�#C�І> ��ڠ�����&�Y^8;�)��8��^��4:0�wz��w`�K%i��h�uy���I�P����W�`�e�|���)E>�C�m��n�F%��h�&�4�B�xp���~��[�G|v�.���S�����EZ�Sc?>�}\��ꆣ�`���fNg\Z�d��V�xOP	(�&(�5��ehih8a�q�d�_8.��&�eXIN0�&��^�=�<��YH��Q0"�-�v�-(��0��{%��4�T�K5�����&��"��3}Tƽnz�G�s�$���z�q�d�{��{/�У�G��m��.4S�0*,]Q�cᆽ�%,��'��;��kC���5�>��V�-z�^�H�I��U��!��)_��נ�d��*}�X��iM9-�/�rN�ζ��L&�4\k���grzN��n�t�Rd�KA1<yDB������Y�۝�6��$,��U}w9#'��He���KvA"��E� W!2B�-2�3|�4���/�g΍�6RK����_���^�ˈ��}�����.��06��]+���Ca/���֭K|�r�9B,�W&�ў�6&�A�vQ�m�빞ۆ``�8Ɋ�?N�|$zN��G�b}�t���l��1�޷�H�>RGN�6�07J�et5�uFS3�"zh�̰
�5
��;�	6�� tȿ��!?$�/�i�����O��;���k�	�F����3Zz�߹�*mg�SxD�.�;`V��dj�f��l�6�'lI�d?4�`�v8bs����~��AKx����E>����sŐ͟��ޤ�}�[��بO�ƭp	��L���T|�<:�"|C3�u�CZ��S��C�.��"��9zlŊ��/]��idl-�}� ��,�QY��d�����`S�����XC�;�)�C��c�����I����#��2r���R�n`��|�K��R���K}�<�s��	�>ՐYZ_܆�=D��F�YcW��Eyr���S�e�.�H����}0��r�2M�,(v����Rꂞ%��c��>�~�N��'���Xlg�py@�h�f�S����ל�WF!�B#7E~,f����g�<�-:���@ �����(�>C�[�b�C�^c޺��+����ƥp��,V���A-��bw�9��q�E3��И�������ŷ���e�x���Q���E�=���2�D��Ξp�/���[%��m��7'�n�jR��z���MAŨU���&�d�,X��T2�-c0�\��,��X����d#s�-#H�TT%��H��NY����p��L]J� M���Y�g��_�'�����I ��W�!Y�y�k1�w�?�u8J�w�c�kUe���W�!��pr_KD�W��G�mםpIQ�˝9_��q�ph�����Wp�0z9�M��~�pE�k-�Pe��-9A��3�?9��k<wL���my�	�T�
OAȁ��D��f��C�Z"�t��T������Ul�>
G�Q�De��z[�D�>�ܬ�Nh$�`����[����,���g�z	w�]2�6� \�'5���g���&�R�ݬ�B�XA-�s� ,�#e�4��G1������
�]�FJ�'����Kf�����ᙂ�ѽX���$B�=���Jg�F���NU
���$-���6��߯=��a��hG� t�n�*�Eh�IĊUIW01���9_��},���"�����z��1�R�V����]�(F�%T��sY�E=T
��P�S�,�Ǉ�^���A���!t��z���*N�w�Jeg���Z�ɲT����x9bOl�h��	5&��j,1��	�I�N4���/6 t�~��c�2�\M��iNl_��ӼO�Db�,
q�i�~0ǁ2�F�^��I�'#t���!�o�ҳp��w�l�(5�#����3��i�s�[��s:���q��������K�<�@��"P�:DeU�����hBjl�5k�%JpO�ˎ�FXL0.X��O'����[m�GR�V��M:Y[{[PtJ�-�F��:�qK�0{~I2eF��v�i�Q��D�}A#@d�ʈ˗��`D4i_�!|��x�&�a�����@�6+%�p��f\g@h�P&�r0�!��������:�2� rZP�%�$:�v"2�i��Z�e��U)ϵ��aH'�M	��N��L2�ɂ�㟅44��Ehl�zwc%�CgD�ʡx8-�'(������U��b0O��(��;=���3��6�iK0�v��%N}fuI���+f����aM!9q��!��jO��N{�p��;�Oݎk^��9e42qhg�}��ƼeRb?���`�����:v��B�2��QY�>�V�9wXυՁ�Ԕj�����	(�-CKj��0�������Š���B�r��Z*�N_���IU��5��$t�٠��Q�g&Җh�`��ʵ�,jT��8W�
[z��VY(�ׯ�&��'m|����X;d%��2B�_N�f���~�(A�wo�*Wi��wz��O�9: ����ƶ�o�üP.���;#��}���X*�]�l�2I6Q��hh�H�
O���޾�/�51s�M6��&��c�fĝ�E�����D8�C�ͽߖ����)1qe4z�V!��c���~��`�M���J᷋"sj0��BV=�����(����=��Ț?(B�<���K�/��I纺�f�0�j�c�]Wo��5����h�OeD����J4}@�0��Vf�[
L���=*�����g����	���#BA��+4���R��3��vk��4DBG^�1ǽ��ЕDϢ�p����z�J�A��4qH�nަ ������B>��gP��Al�V���ؤf��Jn�ʦR��%�!���U�#�T�&5z��}��=d,߇�� r�
[69/
p��54�3I�����r���0x�0IDI�O*J�h䓷q� �����]�L��'�U���W吕�a�x��-e�[��R��6Tǡ��lK�F �M�gS���4Lf��,�,�䍅����C��⮜_lQ�v�woi��]*�u��4���<KKkϓ�#��n�9S���ނ3�x�A��M#@��3f�a՛Xse뎱L�������� ��e���f1T"��������C�&v0��ٿ���� �.�
;��Z�
k���z:uY�M���ZZ������ׄM_�2jm1��Ō��M	��67R�"M]g ��7�Z#�Kۋ�1��F�I ڃǳ��F��V�{�~J�0�AY���R;�Er%af(�Qh*�S����7w����މ�W�eU�:�2�[׽X��y8f, y���]���c��p��DOR,f���7u�YYq{sHN^h����hj�	���]��[�5�OY'��Ǜ_&����[��?0_<Ԧ�͙�L�6��^�s��q(� ?�y#���2rփ/�5���ش�\J�	V$��6�Q�P��d�{FH�PIb��iXW�A ��u@{bG˚OC�]6�-8��_���Q*v�� �G��,(��� ԐU7%2�ǎ)۳�uH�$�=������9�X�\}v�w�6�z�Ѭ�0��Z\�u�ISLi�k暏h��W�H�
Sk.�K�򺟛�_.uV
���5G������]�g��#+t`���Φ�?����2�w�rh���H2�!6����	�o)��A�AT�k
��o�	��tc7��Om'U�*H|���p��WT$yG���sK��������Xǚ�}2���:�X I���v4��؄_JB��k��S��5vRPV��0S2�֨�����F�y�_�(�p�s��X�b׬;�&f��J�U P�t�6�a�����>�����)gd2&��9�%���D�\�i2�=�ʄ�4�>���%����$�r da6ӆ�4̎ƃ��@���"<f#դq:K��R�I���7*�С��p}<��F�������zy��当b�i��׊"2뉛M}��;i'{����#=5�n���(���_r��x��!;$�'���n��'p>߃,�tW��y :f�䵁����/E��C�4��S�I�QG�Y"WC�՚�}!fn:�]ί��/��ِ�T���c��=%�'T3<�U��fƘ����dJj�cNro�@AY�5�����3ͻ�2��E)v/�"
_�tb|�@�c����4?H��Mf��+e7��	Iw:j&�?����_�E<�&wyH�<����cRb;վ1K��-�41�� ���Ҕ(>�K��և�2\�)9�%�b��=5
)���J�jV&��T#�OǢ&u�DG!,s.���� [H���0E0JT���eB�ĉ[�'�~<o���rw	<�qy6x���J���������,�8yF߈��+ RNV&�2F)N"Ku%�)��6 �0\�$�C2;�H�p��:bP���������'��	��Lu�{�ۻ#��x�kȌ�p_A��#��i�0�KV�ʜC��Ba�S�*�u��3�q�/]^[��C~խʆ[p���q��i:㓼&�Ԩ���,���7�s3W�u�\���K-$�K�D�����-j��gz��Q�:�E����qp���&��>��$K�C�i��q$Y��[\N��0+D��BK'h���;K�6��}c��+p�{e?�
�^��
WTcH�z9�B��g}����(
x��)G�,d����VԪ�����>x4��P�Y	SQ�?���hI��Gs�A����b
R8��V��+�<*���{�3u��(��9�{�L��Mr��[6���NN m���������P]�Z��Q�,�����@:�f6�czl�n�����h��d}����������������<������*�,ч<�E�L�$�l�T
�K�͐2��1�$���L|� �} �_aB��g����u��j�j
x�~C�R��=4�E%�+��ż���i�+���X��;��C&�q����-Ć4w%�׫�����.��Ո���ݧ�0Ul�Kս�*P�Jُ%� o^�B�c3gR�[��U��4�@����}��!�h[;�!~��P9R �^d{v�ΑY��;b>�E?�r6�x��ؔ�o���{j����K�4I�C�x}�k��)��y���6�z�8`B��9Щ,�4�j���!f;�%;����_�w `�����'h?�3-f��B ���H��ϡ��>��Fos2��M���"� ����S�����<O,1 l�N�G���'>��Uc�!G/:Q�ғE���	�uzS����Y���қ�}6p��f{��d��b]�wY�Q�+ps���*b?�p���~�?4��f=g)���V��p��ENP�f���ph~��9q�*����wS(��.���e� �'2���9]���g�N�Q׻y �+���&Sb.ѥ��*����\-��W�$��`����GA;{��W�(g7Ihw�r�Щ'o�6�x��Wf�P?�)��5�dˉ&�=��S����tT![��'��#����G[ڐ�,�? nKa��=!?�GM�P���w~!Aa�O�ێ�1����m�4� M��=��g���=�������+�`}ˏ�9)C*Zf5���TQp��(��3�o1	��k����"��!$��}���Qz�5M�G�(�1��l�BѦ�8"�
E90��g��T	3���V�{$��ԝ�`�&�C<N��B�t=e�	�.$��Ԣ-�:D�>1��`^my�H9��ݦ����C$�§��4���z���fy��P�5�
>���O�*�m��\^�:��.ij�AjD�C��"C>eƟ-̼��i�?���������D�o��O&""�Kj�x��~v��o�mvwkT_z���Ur���vI"��RPޤ��_Do�s+~��UE��R�H+��t�|���]��3