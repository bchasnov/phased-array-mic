��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|����z=+���v�����G�o�����$WD��^Vi%|a�ћ��,���u���#f%�j9$�� ���:O����}�7�$oҠ�W���5�r�:wy�P�ᆹ��i`L=������rnk��{�Ԍm����c�AY�0��>�:c�&��bRDY����Z��mM����)�����%�t����k���3({bz�&�[�kK�rqVP(V�����3���R}
��Ţ1������2����I2�*C�T�}g��<�!C�	��0oH?0X�?��i95�ઘ�Y�e_��֥iyQ���c4�E=�k��]���>�G�m�'�a_+F~���4���:J>ܔa��C��Y��UqC��5u����1��_� �#̳���z�S�����ȳE�-���L�ھ�3�Ʊ�4��#CW��Z�nᾗ�6�
���?[��Q��	ż��,�`�n*��ɶ�=Q��)�6�E�I8��H�K��� ��s��B<r������+�50�m!s�E�h��E���I����c�L���7��;������pץO��\�fzwH�u
��2��QY�C���x�^v�$'�f�؏ĥ���{˭LJ�����n"��-�{��~�W�`;�D�TN�o�c�[�Nb�$�ܸ�y?-�!�?b�3�)Vj+�a�6��C]��﯇��\ x��������|��fL�`���� �^0����7P��h�a�ܢ�ף�Ԯ�������>��Xx�@'0(1���@ ���E�V,�hb�d+ݰ�>����D�*�$��ۜ����ǞQCV��CO�V[w[�,����m��\�U$�\J��mu�I�,
Gjv���*!!�n���xԓ��f� �G��0�\fh��<�RH�g_s������y��r��A��T�[fcY�Y�q�r���As�,�^�b����8]���m%����'W��?'{�5mh�Dfy�2�����5ܫ#��M�\��PF~�	I�%�
o(�[e�P��M{��!o�H B�0��i��5�w�4�7Pk��aΚ	zs2x�zY�ɐ+�z���i{��%w�a�@>�������ʉ
�,PwN���h���^=7�:<M	�݂p<X�{Qc��ܷ*�)p�����&{��M�n��e,ox����8�<�ߖ}iw����T���RUU:`q5��e���R8��%�6@i,��)p#����*TX��u�9Z��1R�N�-N(�%$����u\�����R≕N���toT��5W�6�Tp-��ǘ�
�^�f��.�����ޯ�C��(�n��H�g�?|��}סȎH�n7�7���E!Lra�`�h>J����"�\װ��^C��RV�>��b�>�2ke�g`�Ca%��bh���l��K<��*�F�#kC��­Ƭ��;��Ӟ=BM|'���b���,�S^[��0S�C�^�iF�<u���h7��GO_�����㔇W>�b_�#t��ն�8��<�lr����$�},��)�����
��}@����w��H�>�v?1�[Zeq������5���t"��wD脲�v �btZ $�&�K0��4#��1��!�MѠ��5��v�,�{����Ʈ�pP\ ��T�zI���OeBd��N�') �g�t�,�yN1Z@i�z��%�J`��A�B+�Z���(�����*��������FJ>���m��(!�9�:ߣr!\��E%K{B���1�,�k��Z�}�6(��,���p�Ɛ_���%=Ee����Jwp�"�>�Z��X<˾��C�]c����LӪ"��W"�{2o.S��M}
ٲ5EwiW�hb�4�<swZ"b�y;<������k����7�wϨD�����S|�I5�Eϸs\M?�!�.��0:�f�Ʒ���u����`��0�|m�$������bƭm�N����v�ڢ"��s!tJ�~������3.C�?�`����)\��YC��М�kQ��p81llDT��-IV�)ȉ�#Pu�Xa�RG�s��ik$���:7}�	��B�Q��t�a����T�Uj�w�BZ2��]@1��D���m ��z���̈.��Rs{	:��I}(Q��G:4���1@݆*�\# ��즘d~���/�~��6��`)g���]f��!ߦߩ�gdj���v�x�4fW`�Ţz>��W�$y�3$X֔�Ő"� JosK��>h�0k"��ԏA+^ߩQ��q�KT4��gt%��f�sk��2�"����\�C�hh6�gL��p�8"��O�uH�*�BF��ˡq����b�F5a6J�{N�w��k�Q�*;�L�|qT��5������,�>� ���C��e\'����#vp���,�_�,�S�T&�3����� �IvD��[�?y�����Gxe����0�,e3G7%a��H�~v�f��"h�cvX:���WVf4ԟ�Tj�����;�O�п,�����JK������տR���qEz�����N��Us���.����I�'	��� #k ��b~`1`����l+hw�(��K(�n S��%A$k'�+����:�����m��h,�i��+�ޔ�D��o�����LXƸU��$r���o4�� )&Q�^���m�l��2�������!;!y��DV�yr�H ���[V��R�`xJy����&!0�n���~��!I��%Ľ�vj�ma_��W���+m@�1!j��a>�$�&��L�R��d�Md)41+�)�&̀�b��LF[�/a?�jNF�G`�CZ%���/�Z؜����2�ȋ���=�x�>X��m^��|3��'���5ryg�
��GFsO)޵����X1�Dj�ʔ�\�]�ޖmF��p��i�-!�E��[��}c-OJ�v���eq|{�(M�$��3���	[�rw��x�ތdyw��t�i�4���'�����?븰o�A�@�F4+È2�B�b:�c����j}m�����G��S��`�k�^}=I�����Ϋ���M�"i��0f����yaX��|�x{�Pq�"�.����ı	��]�kȼz���([����H-,�_䳝�,'�[��Z�M G"���k���/�_u�2M>����ic�I�%%��q����J&��YDv��5��D~+��{R���O�Iߋ�Q�/�S�_h��+Ъ�Q��9>[t�6����P��/��{�?�r�l�0<�cXn�saGS����������َ�D��G�l����w���n{O�gt�I�.���C����A�y]��)B^ ���2����yCj�KD|�TW�d��i�����n�A~@��I�ETp�ŐePt7�ؚE���������k'!�͛�����8t�����F�.���V���mQb��D�n41|Y�0�-�$�2�l��FE&�9d�CK�C]��U՞��Lq،�7����]7��ND�u<Pǃ�(5�iC�X��ͿXK+���@�-`���x��n���v�o6��1k+�_<&�;���KwH��=����<��0N��z�>؇a{cr�'�OR�'��"Ul*�ک3�n�	'�jAl�\$c�z߾