��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\����q�?��e�I8�b�Ǽ$��"����ׯ1�V0����3(;g3X�����Mb����9���:���UlN-X��?���GUQ�]�J�P���s����4e{�M��T��3n�8�<�'ywo��S��T�a.t��A5[�=��y���|�j��T�Y2jC�N�KP� ���M��vI�{��5#���JK�pm'v��p������=����f�<����FJ�ki�}�-H
�FS�º;	�v9���HPћ^O��޶�z:r,�QX��߾S&?Q5R_��	_{7���6%}�I����g�<.��.�L�5�e��pM�u8۹������� ?�z\4�c#�ΰ'�e��F[��-��*0R�z�q"
&��dNa��i�]��L#��L+��Ѵ� ����~���(�M���7*L���ZЪ ��;��$��D��=��sxT�Th�V����0�P4<�q�
���+M�1l �f���U�ZJl�tFV����7�8�o*]�BD�u���}��{J�f�ԋY2���o'>�͜��dHQ�p��wuM �������Q�[笠��MyO��$�mTC�l����`���U�>�\J��������~�����#ovy5�vS�O��:�	7wa�f��9�ՆF�=t������r�I���j �sj3F���\s$Fx"�����������V��~6.�-#�Ʃ�>Ƹٴp�[k�7e������3o��H-\őU�b�A+t�+�fCz�&�x��qm*�
L��QY=!8[�_Z��TВ���iK��'�[�N�J_A	�\�4�-ެQ#+�N�P��?��N�Bɺ?�?�~�:!��;�Sv)c��\����})�i�U>o��K4B��CL����i5��_�W�i����x�3S�=�|GS���*$�D���vOf,�p��b-��l3�+�0��BX��Y��ܘ���
��SAP�q��PP�H�:@[?��t�49^7�t''y�33�[!=[R���It'�Jm봧��G_K��ڽr��@���_��=�@r	�9@�L<{�(q�����¥���K�͡��c�j�;���O�i�A��r�K��>R��-�(�I�_��R�N������-ۣ��
��*�'�=�q��d�Wx%Y�&�|+O�'j�Y�DvŇ6״�����xޕ�+��(�J$|'�թ)�T�������᫔��Nԩ@�����^~gp%���D;�W9H�b���mD��%H֓L�;����u��q�۷�����V�+qT%�~p?�Ţ���0���i�ﲩ�+�F��<�Q�I����_D_�m�-����ⴽ��R�.�r%�����+3$M��ŝ,}h����J��)������t�ww`� ]n��Jɂ�V�$�潱�!#@_�C��*k�a�ޜx ��m8���w0�B��Y� ��"H���!ݴf�Pa��ڈ��*�2W�yay��`?�s�d���-�߅�['D(���hG;1 �1^�402�^��l;H�&�deER��<��~
!�5�z��Ѧ{�/S�+�E4���\I�2�؃U�D��R�uW/�$9�:)�cV$�ٯ�&3R�����1"��-������.`e���?�ڋY}J�0�����`���J�U㼍�#�y��<�a��A��	ꡱ7����3�*��&CQ눣����l=���m�����A?��1)}_���8n���ہmZ�Z��fs��#��!�SO�Ѭ�N��<[�/Mu�q�>l�m_�{,�Q���rN��-�q1�e�g3v���/��s�^j8�R>QlR��TJ��Ia�@o�tNM�����8��ܥ[�~N�Ĵa�x�� ��x߃�kϼ��9�g$����%sp=���&3~��4�z�BZW����fbs���#��8����h���2&��e�,�[͸��?-�o�	���u�|ڦ�~W.Wc_)II���~"����-��6��H���v�Ǒ�)Y����K��4Z��'��CUUCQƅ�s;@8��c���U(��9MzU�*j_��E$���j|e}�5ܮRG����d��-og~gt�6� ��4�ʪ��|�7�؄k��;KN:%�z㴹�s�Zy���1���633�c2���X��-�Z��I:���sd����E�������}�s������<&�g�2��W�xlF�N�}�����gMB��+��B�LԕI�,t�a���i-Ʒ�ӆ�
L:m�H2�c�EGh#�w�W�1�U`�����@lĈ_)&���� %��� �;��A����t[�2\/�0h{�qĕ����t��MN7$Z �VL�Nn6k����lQ^�~R?܁4�|	׊�{�ıCw��i���i�2E�q7�5��] �#�CC.��@�F��\��i(e1U_��L<��h�wP0;p
��E��;� �@׈�������1��d��c�+�ƹT�
M���U^�`67�E�"DV��%�Q�?/I����1Q���;��E[F�mO�Q�f1=�̱��8��1[�������z��`"ϻ���I*�&���}<U�&�������4qh�wݐ#@����8����D�[�ƭ"^V��'��
��:�����m�u�$Vv�x�g�M�nEP*�N�*HȀ��3�u����{��ŏ�T�_>��[�䠂'�1�v����uq�7����G]L�O��^'�
���p h���6���9$&�Y�u��Od����@ھ�>�� پ��zT
%Zh[7� ⷫȁ�Sg����� ��j�V*�w�iAQ!��=>��:���`rQ��$��+�4�r����z����y����4~$�}��*�������E@������}����w�����Ji�]��J)�^a���Xl`(�"�w�iƃ.m}.��&f�&y��|/~#�6�/��f?Fo�'�-�XZ�#L�D���Ym�(����!l
L��~���e؛�]�B���+��X�A��4��a��8	���\��3� L�ya)U����m����_P�N��G챾Tn��6���{ĉ�R����^$��ʆ�y�}'Vk��RӐ~��ۃ���2oB���6��=����fV��Shr��a�L�+�Yf��P��pF^y����l�v3yZ�M�S=	ŋDj��UG�w鷬��7QY�G����(	&���#{S�����������g���pK;�<�����[���}��x�0$I�%P��P��e��Y5�F,-N�m|a%ۼ]>��o�C>������Y���#��y� �90�( 0��#a�G^��T�6t����i�O�6.��ۢ�Lg�8��m-��	�V:�tD��{�IU�Mq(����
F\���XSb�Q��$�p$��R	�v�zj�R6��ڴ�p7^�Bp�﷒�d_��������׆Y( Q�urZ�Z(�A�iϰ���^�o�z(8/��U�3LjXZE@J��m�k��`Q���8���"1`�5� �9���Z��:�)��y�������.	wqK���� f,�(�|	j��V~���GS���=pS�t��o�H�M���7G���`L��f1Xu�p�d�dj��mFǪ�2$
�#��(F`(�Ӵw��Q���d����-�����-,Le��n��U�0���;��5��j�� gb �6�Izy'Wm�l�N�<��Od5��I���*hV�w'KV�E2�;���]E��@��A��-իX����A�j/�<#"!���֍�h�G/d����������F-���l␊3a��*M1?�n���Y0�r��8�
L��ѢX&�+��N�u�E^�M��.HK����������j�q���9H�%J���:���W	�^<�n n�OZw;�5L�sJ���p��K������oX��&���i�����ƈ�M��W��ϼ"� +5���2�^�R���x'��,�r#�߿�t���<d����q�l��c9~�cy��ذyN�`/I�p����,����\��]:�	�MQ��E��Z#I ���I�j��`�A"��(y�aGT�!�\�z��+r+�a~�,jh�2�:Y�̓g�U�;W�������i���W4 F]�ݬ%u�]H��Q\�g����n��4���[Y�i�۩y�,��opF敯Q��XQ��J��-��v�]�w�K�9Z��h���	��|ީ3�C�S
�A��fZ��_w�xS�H�i!���V3��