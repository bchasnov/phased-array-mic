��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@���$U[H_#�/8�y��,��F��`G�m6f�f�aiI`������tC����dl���=eZ��^�٭����B�FYĸX�G�����݁�]}~�s�cC�_ �c��2)�}ma�dظ��v}�b"@@�c�
l�bx���,���M�4A<�r���w�$�S߇��`w���~p�lV8���
��%�4�0Q�Hj������8�Wnwx�5|%�B4|y��<���C�bA��T�N���Ζ�:U���J�::��;��B��O����k�q��Q'�O"�h$ZrgtI���IB�Q��s��P=�=�F��Q�4d�mM���v�#��D����)0 G<��^� �_�\�y(����¬.��	�y�* ���Ob$�}h��@y��y���ѫ��A�".R�]�hڳ��2��}Έ:�g�wQ� ��)��E�w��V9w{cJ�d��(�	0b�9k�X�� mKٺf�רZ�[4D��<0p?���T�4)G��L[7[�4�l+-
X�tv{Z����N�8O��B�埑{�	"�=%����Q�FF��bi@7��J�5V��n��fo��; ���Cn��m�s`%s�*�+u+��p�m�|:��d�%Oʴg�6�A� i��8��tK�K@k�W��'��X�@�0���K?n{ץ4Ej����=��l�=
q̤��+'<�-AOU^uO�����h��E�!A�M�]������w�l��C�h�a+�����?���{��}e��_����9�O�н1���8����J����j�H�R��T��f��ڛ�.}��դe��;rJz~ل!���̽v�Q(����O�i:
I>{��d��Q��r�D~;�������wB� �����AP��rB`�\$�Bg�E��Xzy#0-IA~2���A�K6Q,��z������JX��	�����%ӟ�ݙL�?��f"S���s��w0�ۜ!g���S�HK_Ư��lF�%��6�6�,ѓ��ͨ.�,��r�(N�mG�����Z���/�Ci?�˳d�?�[+t܄����D��E���~��s�Y9ߟ�HN���=T�H�b���2=w��x]�� 5y��ț�Xl�F? 3B�N쒱��Pk5�@g6[-��P�`�d{�gY��+������c���5�n���R��}*���{��7���"���ەyOMk����F���8�K Un�O6����!��4K=� ���@̑��[O�6q�H�/�o3N�4`���
׸ Z�+2�5�@P���4�u�ʳ�*�'�ћ)�(��^�+p���Jm�|�h+��9��hx��#���N�dŴ�����ǅ�Cgٕ�<�ڡ|z ���*��k!f}�Gk����X��	�z��-&��D��u��}���n�4a�?����%��r���4X�b�j�J͎%I#xA��b�sl�u<����	�vr���"PJ9n��o�I���5��hFg��~�\��/����	#�	L�?H@V�q�8Ս<�n���r%oK����}�CԠ���A*��(b��9�G�-��4��ѶW.Fz��>�~րrz�o�U�j�`0X��U�:�DG�,SM[:���B�����CV�@��׊_����pg�R"VSx���4/��/#�"��-R�ime� �_��xwf�7+�f��DD������ƚ�N؛�)��u�/�Vʻ�� ]�f�L_��P4#��,vjH�w��e�W=10��$��p�|�F�W��ă|��-b���a�y?"�ܕ�����՜�Œ��϶��A 	�y�K�*�B*Q>z��FJ�4 u��W�?��Pr�P��c"��1"�8iCC����/�J4�S���Vz�����M����8�Ө����ҿp�Ł����`�+}.9��`��9��g�,2�Q�D��[H�۩l:{`	!�K���9� ���=7Dٔ�!�EM�s��9��3�C���u���ܘjxҊ߭�?xoC�U�z�F��>/qXE�I���{����W��v�yo�i��ѥ�7�j��^(8��}B��p��˖%�u�����[��C1*"�U�45�{�m��Jbz�-��Ȝ��ɑ�-�n=��Mq�Rzn��	ߡ�#���[��yV�$?��)@_�o��=�1
2h�S�u��_T`�)`�R't��S��@fƙ^5��Ӕ�������.6�3D�jaz�"��Zm��(k�S�0�d5d��NBq.�dpm)_̂��;*� ���A4Mn$�%�[-ӄ����L땈d�1���#xsE�gQ2W]��9���}�~��H�0���9�:|��\�t�O�Hy��Iix���S22��!ޟ�3��',2���h��xcA�E���q�R"����\2.�`]�{i_Ǵfc���."�Ɋ�nu}[�I�3����l$%��,U�|���曝���q���
!9|��Y��^ T��:�!=��6H��ѹGr}�B ��d�~�>"�+W���fW�����O~p��nM�z��7�5kj��E��_	���]_���/?"cG��w�F�Jȕ����?V�Zs�O�[_���2��+oϑ�ƣc���PI�J�=3N��V�J��	m\����`ѩ!��"��q��K�1O�����}��p����k��&�q�����3�t��{�zW��������k����U��0L)��4
��S�R�ʄr�O�
�@�O����)+�����wO3�h±�b�7B����4#�f%�0��s��:h��p�~g�`���SS���9��hR��\���c
�n@&t�V)�tu�Q�Ӑ!A����Ũ4��[�7A�Yo
1�aFqD�4���5|>��i��3B ����Y�%Y@�{1U�h"H9&�`�(m�����;!yV�U쌰�x%���C���i~��B� �NI�������;n�XW��-m;��zf�k^^�P[�&�q$2��_�%W�?�1�9��{Ue3���Ȏ���}�v��ҿ)����&^NQ��������0_��,�9a�\7�4����i&_��,X��[��SQb:�ܺί)��!<�8�#�����֚[�ә̰�J1i�D]�z]dd�ٓn��M�N�}�[mN�y����]���񻒒���lbc;�X�)��ۉ��&F����}�sc���/8�Ȇ���Ö�qPێ�T�(0ݖiz�
�t��7���@ǉq���=��*�^^^<����8Ga���//w��@x��J�`���qB����SM%ˈ�(ˍ�6�}�^v0\�/aa&5����(�2v{�Et�T��!�p������G�o��-�*u�;�O���^��ᛒhn	A`+/��8�z��T�b���W/�O?:}l�`"W���W��و3tX/��Ne�����<3c��f9����/���#e�`��\ק�&}�ີ
[.�o��M����w�9�E�6�~0��� #a�\��E�c%�F1��9��s�֤'P`6Oj���3V;��؈UH�;��sh,ϕ(9���HD_���K�q��8�����t�eMti6�93�h5o�lg�]G��%;���'�\?49*�q��E�x�V�: x��8���tEA<�{l*��GNQO������̂�4ѤI��cM�F.ç^&��RR��z���"�Z�۩��y!���5�zG��6I]N{"�O��^M��XG��~�g�dA�U�m>&Ta��F,�|��a��}\��Ϋ�@n��\u"�TL{�	C���g��d`��:�6��I��^X��65!%?�~��Ċ̛|X:��G�A䠝��/U�u�͐��1wcc�aj�(0E>+˚-e�XG($֕Qn�9���iyJ�Y����r'��H�#��T�a�\�MP�lm�t���h�;|��<��vRt���52�?��=�Ê�"�:Q
���'��$!�~}������?�H��@�fB{���+ڄ��MH�˃� Φ���$��Aɑ.�E�|J��x��y�V�j4����ݒW�Cࠅ��� �9ެ!��NlI��C+hu�Q!����=��{��'�1���
a��I[3��h=j>�`�zE�L�N��H���/@vyp��[���#yo۫��e����\a	��