��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\����q�?��e�I8�b�Ǽ$��"����ׯ1�V0����r�xQ����ez ��ɥKG���t�T�L�=���Q��W[�吀p���Fy`5�i�ґ�,°0r��P	�S(:�Ĥrhl��{�}:!�����R����>����o�A��~JO�u�L��/{�^e9�#08+=a�ik8����E�R��t��j~�Z�����!%��ˤ��)��݆� �[9�3f ,�m_�d-�#���e��Y�
�Ne����;t|�ğ͎C�̌\5�6��cYq^G��a�TwU��`�X�$T�F���$����R��1�M��Sh��|�s8a��^v����l.�j��
�� HN{ت(�$O^��HN����� ��>�[:<�8Ȅ��^M� `8�h��g��6�jaÓ
���Ԩ�v̉��X5�������,��#�ƾ0N��@rp\T��)�vk��1;}�V8�1��TU�}���e��$�5����|��}���Q\�H�0�d7V��_���n+v� �I
ˮq�Ǆ.���Ӎ\=g_h�G"��[��yb�U�p�""���~�s'�ɩ��uw��(�F;6!�l���D�a�[q�[��i܉YϣiW��O�&y�g?'P�Z���j t&���<�7�ym4����QSO݋�s�a~c<�S+;���uӂ6�o-9z�����Ti��� ��d���:	�y�[�lol߳IyZ����[��S�q$��v
���[#�������AcW�2�UbuEө3��%@��"��g]�z#X��*¬�b��/����)I-#|+������X(ÃU��xm)�m逤�y�X�����' �m��$.��\�E�z�p�m4���-�8����:�m�U�_I�C���v-��qС5�
���Q� �+�	m�i���9r��Ȑ!�{LI�h�Ε�fF3� c� yj�h:dY�!X,Ҳ.B����0���J�R"h�����U�V����e�<j˴����I�O�K�.�xC�� >+��ଡ଼O�1:����V�H�H���.�m��c��P{�\�p(>�o|�������c����B�R[�C%¤>�C�s�ݤ�Q5ю�^@�S�ׂL)O-f}��d��S����h5�ym;�)u�왓������5�����f�M�^}�˗ԡ���eb3�8�د�>���rY"?��� ��zCZ������䑸O�<��J�����P��D�H`�~+E��|N�|��s�l[�ͤ�prj���1�B��{��U��.H�4��ߡ?�*�y���p3_~��>&bm�=��Ԍ��h�����A ��qP��r 	�b�pr����a����EM����\S���y�(�{�s��$��Y��"*��V���b��K}y]ۙ
}�x4oA���4�K��N:O5A��Eeu{f����o(���`�T�od�\7���v�e�SnN�*�%8|��?9�\咾ټ�rN|n�&�����[�ŻUG�U�qŴ��K�`6�$tP+U�a���^���]C?+���%����j�����8j����ʖG1����c����%���/��t��D���G�HPjg�q9&���,���9�۫��� ��$w�˗h��������K�����UУV�s��{E43�ę�񶕸��0���yӭ�IC�EĠ�>&=�LH7�nA�1��C��#/���Oa�v�~j�H�E@��Z2S@a�a��mruש��R>p�;�r�-FK�/�g���E�vi4�F�W�����c����a�tq�tBf�ܸ{�D�|8|0c>���+3�
��䘼D�Ā��с.Z��Da�r�$hf��K;K�+B]3�~��+SV"��U�} ,��(��9�0)P-��&+!�ڏrk8B�z_pBt1Ǐs~��w2�RU��H���wiR�_�O1�NR��=��XV�Ξ*�A� �d�u� �YL�N�)��YO"r�Ω]߅���;;��,k�Z�JI �Q���P�Dm^� @��:!q6��Y#�%J�Y]!�/�h��|ٵa�lF�����9�3�p��L߽A��(<O4sOuJ�W����'2�%��.yH*��!t ���'��3���.�;�|����Ïz�r��[�&R�N��`�u�>@`�Ȳ�P�D�UTǜ��@F�a�a]�O^x��}� �_���Ǒ�q->kVœZ�=���`Y�^j�}jHԔ���,�����6��}*6��8`?G�� �$I����\7R)�ց�o���X\@{�u��if{���dk
�gUEa}e��Ώ\��%�zI��2�X��W����95�pq��SJ�[�fa:^���[L��L�tqa_(X�O�aSz��8)��&dx�7} Cft�#S�*������)�
X�Z޹**�@:5:��x��&�(I�g�_��O���)#�3�	�y��}-IՌ�%��%B�gsnfZɢF�(�x�;�+OF/O/����@G]�׭_i�<������!��x�
$Q�	|>���V\�����*ք5�^����t%_����onYK�*��M`�l���Hv�,t���şE���1���_>=x�|�f�������@\)��P�E�m��L�ov���$��V���<����Q��@��5�� ��}X�z�s>��!�ٿ��� �II�;�@L܁��]W�d��B.�p)ʑ֡v�% 6f���[��\�f#CFG����!(w׻A:����O�����ur�Wlf�%v�Ѥ�KKa��dj�=�~��E�w*0��"�X2>	�1j���b�5S��e���IG^n����x�7_	��٣���f�׺��6{�L$E~i%wtr�!�s�Pt���?;ST��JA�I��xB�,�IEB��5��w�M�~�o�=*2��N�FX�)V�}F>.�ǟH�j��~0�Mڢ���)�6��)r(Ոy�o�6n�E�J�h&��Y� ��?s���eHX����*�Xz,��l��܅�ӗl���${�Ŧ ����4N��=�$�7��\��~ux����O�鐲��5AC�R�Fa)���
�l�!��om��(q�贫�A� ������W�2�ί�\e��q��0��Ǐ�~!Ƶ�0������Ш �ҾF3�`�|ew��ae$ՃUT6I{m�G���X�=3?�z��o.C�/L� a-�y�	������$�ym�MV�y�z��!:D��OD��;ɯ�����$:aV���"���<�7��_E	V��/�q�d�=V0��Ck�S�4� ����l���4h�롼;��5rM��ʒb�����} p��{�� q\�2�F>FQ�n�~$Flő��-�n�Jm�<�ݮ|�ĸ��>��x8ma�B�4|h`���l�26���?�:2���X���vK�o3a�˟�����*��zp�B�Z���5�y�>�<�(,��E�����|X�=����6����sv��;���]�%��Uw�u?g��/"M���쁮'��<K�����e�P
�'���є�;����(�/���cNZs�0,~5������z���w�r�H�7s���y!��}���.���=�� �����Q�Hq	��Ԑ��6���I=���O��|��ѦԼ�P�jO�N�9T�� �i8SoXʓ-�	s�fj���dą?C��Q�`�r+d(���f��3g�bv�3�jMڍڑ������ ����wԕ=Իw���w�������u"�a�N9H��6~)�����s�'�	m�vi���<�N���x0�nqq�CH�Q^/��qC2�����tRfOY�a �5}������m�q�O5à�F�۝�-��iV�R�D�s}��E��ZkO����c�����@�q�P�s��!��4k)(a/�rg�G�ҙ�����|8ܪ�jbȂ�4"PL�>�V��Tmv�[��:F}\Ԇuz��쩭w����y	�jc�(ó|�ow�Ӕ�Q�c��5F��)w|��l.�E��Gs��۵����|��MLǵoWA�(��|���zm&��*��	� ����<�������<e�۰ߵV[
���t?n7����QJFތ-�׾;[_>uy���b^[�!E�Bw�촗4�#�LH�����8hQS��W~�{ѝ_4�i?�Q}��ϰ���p�o��<�vE�hn��W�;�
�;&����;Q�o(�4@Nk��y�m�+C�~�r��⎝ԧO�S�d��ڃ�5{),��{_OJ:c����	�i�� N���`щX�2�� �oΐ�<�_�9��,��	QX��p�p�N6D�OZ�.K9�,(����"��0�:���]�A6�y�ح��q�iG|e�U��	+�E�������#��0���
�D� ��1�H�H<9D�X�F�m�$���9<�1�;���)bf-��;x ���~wu�̨h�%v�!��ڣ��p�Er,�?'�@���p�g^˹�9*(�o���D9A��+��6�>��F�\>ϚM-i3�|ԽsC�K��A��^>��&*�P���c�y�0�� ��nx������R4�E˝�sN�h�&@(Xxu�D��p�v|�	3��5�?D����Ǘnn�nR	�B�
��������-Ҩ��F�ԀY�Nx��<H}y�f����U�� �����ɕ�@98�s�ʀ��|N�8U|��aH�h�H �q�k��-]�S�G� A���M%Y��yrP��JYZ�@�p[��C2A�F>��U��DF(�<�"���7Pd(�"�L��� �
�\�M�?Iʞ6���+
��^�KlU�F�����,�o������=-�����wo:��q������Zn7���wE>rc�g5f��%-��o��i��|�Qc�O����;]g��˪Y	h�@��8'�q\�x�n�����5�e~k�D�����y����#��Z�%�n!7N���2
�;t�>t'QN*�&��-��D�ܣ�������i��K3�]دam���bؓ��t��w���>#