��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�k�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������H�W޵α��wԊ�6�a�3� G��λ�:~7 !�v sh��~��P�'|#��x�C�[�~���{-چ��!�:���)�#aE�C�;� ���&�'��c�w|�:�)��$��Sއ�Y�K��N�4uFLN��6n���)G�Kh\��V�x��w�!}+0��M�j.�"̃�����p��V@��׆�+�ŗ���A��8���e����\� Bx��%F_���*gd�pFߕ_�U#�E�75!}[(la��M���+l�
�J{�����O���/{x��c������x;��%S��!�y����������U�vX�iS	�}�ә�6���6{r�b8��M���A�
�ׄ����y�G�T�����)��(�A"?5���J$m�w��p�{�b�||�� �W���=�$.6A���9��˶g=���`�YI�x�4���`l'��o�z�m�8"pa
�21�*Hn���ivG
��I���_�U���I�)dpd���P�� ���������lG͔3�Շp��Vf�uxSnYB�/ґ2��M����9���X9����%����=)�����}�:��94��d�Ly��Cҧ��}R��տ<��͂I�}B_[m����8ų2�9�T����Z@{�o?�R�ts��c�.
�����-����$	J��� G8e2��ݞ��ܖ.�M��0�)3�E�"m7��K�DK�$�˂�� �>s�^m{UX*�K���1�J_N���@[��3j�!��	-4�/\i�B�P�ڙ"�>=��U�ٴ��}����2A�k��L�,.��t���f�o�R�����x�4{\kύ�T�6��bi͉#�~�Yrd;��!�z��'`��*�SF�q��w�*�|�_�%T���r����aW2��w�3@$�	��ՙLە �:�ln��c3���YOq6!�R�:���d4㢾�0�ҟ���O���X���g�w�u���>��|̃�Ql�[)	9�~��Q��P��M���To"mԜ����q��
 ���;��zЇ^p�V���E��D�#I�<�8�-���O�rR�v���{������q��Ȫ�9�Х@���9��#�u�H�xo�+ͫFn^��ĖI�����z/�zr�1h���t�N*�!;���me�K���Pj�ܦ�s3�'c�_uAnTdQ���?�f���ElB,�|ԯ1G�,��qr�i!a�Kϱ�~	�Sۇ?�i�ͬ�P��:����/2���\*JG�r܂$���gj�K����Dum\8u3���%��2�t9�t���nlM.��Lk��U�X9ܮE�+�y��p0�����_?�\!�g)�=�KȽԏ}	w��r9Ԫ[�u�e���S���oEg�S\@��~�_|���_����������.r0�=R�JSk�k,�n<y�@��I�K�H����
0Qz�3�]8l�a�ꤻW!z�SII�fֽ-]?�����VJ����}���F�
2QH��XZ�SE�I��h88���H��ȜΌg�p�����% w���05��W��V���fՄM/:��=o&҈�3�>k�~��e��A ���������BwHO�e]�R+J U�}sk��iN�.��R���}�A�nvwkc?I7�]�'�W3��*�q%Y~���	Gw��uå�1[6�wf�6��l�#�B����v�2%0��ʩ#����p��e*2�ւ�S�f��,.���#�<����8���}_�3詬X&�1o�P��ZF�&�k���]�h�d���"��{��0r2kB����+�E�ٴ�����D���*�����i�n�L6sc��E�"����8�2Y���׫ѧg(�Zn@=Q��GΉ�sr}�Gr����l-j��b�l5�.Xz������~�2�3J��;׾G+�F��䦂��ZTd�	Zu���Ў��L�8.�
�6���IX��u����`p��I/ϓ쭈_W.6u
?~�d�Z���v����-���.bֶ�]��i)0Lݔ�S?��09�ű� ��	��H���ȴ����}.�融��+:��af_i�o�3Z��\0,��z���/�j6m[�P%��N&Z�����^
�k@�c!4�Z1p�f�Ț=�}�W���9�ə�b0��v?��1~:�UP����p�G�t�S�]�w�n����9;8�פ�v�P�sy��MƤ��,��P*ѩ�n��6E��_�4���j�ʦ�#�!��'���B>�D+�-��+��=y�Q��_2+s�	T��t��W���ì��Jr:F?�״��7��X4-�%)���l��b�擛���o��S�k�Ѝ��k��0\�rCR��>��i`�w�G'��s�ߋ T0��eA��/3{�QE)2q��,(tם� ����&�D��X� H�Z4��-�n�k�k�L�^�\�`�Ӷ��Bߠ�V���O5�]��[�G�r�C�[բ�]_�E���C�t�a���� Xv��>��F/�L���.|F�P$4G��91�{�d�qI���h1��
V�[=�p(�E�h~�嚔0ԫ��!f�ڶ���^����,��iW+�+6�8�`�e�o�%��oM�S�4�Mt[�Z��.v"��U���1KEğ���C�:���S/��ͥD�<E'&-4w9�V�Z�����E�\h7YTu�Gl{`��N����7�y��~����ue+�����{���c�|ɐk�ñx�j�Ոwխ5/.r�jRv�:y�O%�E��������rޕ��^����}I�v����'� >]�ty �n��ý�rQ�^_���چ�M�=�����a�qh<�!�C"S�,� #a܃�!!9[���%g��,��k�Q��9�V �\�P�[-�j�ֈ�08Q�[a���k�n�p��$������h��#��^obD�Oۇ-7T�~�%Fa��7t�*��ʳ��R���Z����\SS�T����T� K�� L�u�e�{�c(���YHG��������ՖD�Ή�ȏd������b�՝�:}S�;z��1 ��QB;h�xnM�f���	ZCe�(ƨ�|^u��D� D��M���q��M𽭿� ���95D �8¯�