��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1���e}ʲ��cg�t�ϙ�a�:�KR�%���ݧw���ȼ�B��~Eвa��S�f�ap���&�[���OմMɪ�,/dY\d �ʚV���]z�:<��&ͼH`���3�5ALz��B��ʖ�Y�j��)�&�T�<U�]����r%.���{����0V�![' �l��#���G�ї�/��+M :P^��4�A��X��Lÿ�|��b���h�p�8�//cc��}&|��w����z4 hTpG���K/Y4V�����F����Y~���m�o�O�0��ԉK"�T(ک_�-�Rr��ӮE�Ō�L�g쵵�Y��]�jT�eňO�O�+���!o�#Y[�Q2�\$��fH�L(�R/�?,�O�c�;ѽ��.F.��p��,vc۝�؋�p�#��M���� 8��'���/b�A�6�D�8�D�Y���"~K�ғ��A��zȒ~�5Ξ�˜r�������>�~���>65'�F$�����(��E�b
"=|�川
B.`�FʆF�_��^J�w��<�hN������A̸�7#(=�`��Pf�}�5�5*�Bn�2��	����aGS�iΎ�U7-tbC�6*���P�����v�~=B9r����~I��gLS�K�Vw�@y�[��z�]L�"s�2�Q���4:ܓ����Uo�vh�tAL�nD�2����"Rnc���Z��j�NĨ��x��d F�&Yz9�5�K�M�b�(^�.����Q=�[73&d��z<�(u�nS��6�ѩ��6��ӑ`h��/�Ļ
��@Er �m;�>��J�H�2�ix�'�a�{��������S봹7�.�xMIFL-��N�1��2�z�}�p�<�<W���ia��Ҷ\G���#�98���B��$�j���[�zj���T��ߘxA�
Q���+��Ƨ1��Z3�}��"��s��؟�B��o}�6�kÛ_�KE�,���q�G_�]W���Chݿ�C��6�>T���M���fXП���Ȁ�������x"��H�d#�߆������P�LL�ځ�L�4����8[��_GˇX��a�� �աP�8��4ݛ	(V�%k3��=w�B���,�ώ��\f���4Γ4��qף��̳I�����d���p*������a>ɷCr�Җ;+q>7:�nކ��"�Q�ٸ�Mwr���E���VX�L/�<����`�?��;��f�V;@t�����ѥ��c�o|N������]-��@[�o���HO�F�*�k�K7sX�I���c)JsM�u'��A8�&9�������Bz��	���pF�D�IL�= t0�@fl��o��"�E�ܙ�l(����2���M���mY��ѝ�TĊ���-x����Ѵ�:�:2ա�Gbߊ����F�7GĈQ�E�ܥ;	�h�4ŉ��z��r�d��� }?����5}AR�#��@�I��O`����neu?��C'���Ĩ1���#�4���:�$��u�<��ɡi�&lM���r�k:a(-#�=�?�ZhC����P�#��L��������@��(��s�7��к+6e��uIu�ɮ��l3�����'�~��7>k���֕����`z�������ϱ���i�3<����{o��מ��}�}��l��֙�+�	i�{7�'��W����V�������̸��f����U&�8X~�/�(����)���߼nT�g���TM�=�7G�d��r�0�Z~�!@��?B��'�\#
O�7� ��B���h@�v$6�&�&�Q�ߦ�	���7Qs�B���N�L/i�n)q	!��q�#��`@�ȅ=�O4C�s�����鏑�ok�eS�NJ�cS�f'��P�[�[��Ab�:��$	�`�'�雂��g\�k-9a���P0P;����a�C�ǖ����N�V,T]M�+���Q�r'�M3#5������!A 2��##��M`'��R��;�{C�l��Xu����y��4M���J�ћ�C�+)(�q��k-TB��N��;����M�ǻ����Y�V>��$bP89,�@����ָ�=��_�r#*����f;lw5&b9dR�� f��?�t��Z�η9�~%a[`�H�J=�xk?�7C�zwr9�T皣�=4�}[hT9 m��w����qvS�@��������8���ln�|�<WL�̰ԯ4�-ʇ�s5�R>���b0C��>�UF�����>�<�����#PQ���]mТ��h��?��������@�HY8�������l� sXȹ����!r@Ĕf�<bH���Åz�j�yLb��3X��ՙ<�~�����eɋ��y.�j;#�ŖPB�g&�h�I����z��-�H���L��%v�j�n1�!�o�g�Mg�\oT�1�h�|�+䨍�Lj�B ��.}.���dh�I�Z�Z?4��鈰_��y�l�&��3�}J��6�͓��6�ώ��Kh� B�W=l��D,FdZA
¤���AY��h�EBC��*�
��I�kq�.������	���ʼM���2�+���y�@��:���� �a�67�\l��"����o�D1N]D������z��1'�'�rNШ
���������x�4��a�L�����tOc��.ǂXimRdc�`_��p9k1�XR���)d�@r�q@Rl@	;Wj��.�i�U�(�.^U&��x8C�B�a#���>�UgN`�U�h`
�գ���)�SN�� ��hf��zl�t�MKO�6+�r!�t���������"�q��ы��lw$������h���z�3�T� �JN�ʂ'�������ߔ�j?J���t� �QPedso\�|��Z3�Qe2��ҢX��w��UsO`;o/����q ie�	�G���\U|'�+y��ңjf�'��֚sU�1�`����!���)�*d���m:��bu��������_�T�R�����>}� �ݯȼ��E�Y��Y�̾[��E�\�1o���@yC�\��$[/`cf�'5�c��D����P͕����Jy�q�^R��S'[����Ar7m���4�ᶑ�M���ur�F��SY��*��Ϊ��2��"�z�MP-,�4�����ƥ�:�85Ò��h�Esc�Z"7j��U<���3.��il�@�l-�F�*zf��D]wV2�i+��G�ЏwX�ᠴ|��*.q����Y��ƶ
1l�~P�gn��y�b�#��hK4�啬�C��L[�����mA�Ԏ
�q�3n?�k�%I� MGmw?���XI%+��Ӝ��=ZbZ��K3=����b\��D�~L��K�����
�v?��y��M���m8�;�����PUS����8K�mŒ��3CAj�?<�,�<&!dcG�#��)�Z%z�S��g��(Bp�@�x��V��j��������]���j��G�h��Hۥ����.j�0�>��+�ͬ��O{�Aet�������6+�/�K�x��G*���'j�����z��J��hEB��
�����~��FΑ�x�*4�\�^���D�_ ��1 ޮ9�7��D&v��)\H �7���C����^�S���7b$n��b�����5F�_���o���O��j=�E'�uY+�����~6
#2���A訜BC*juE���9�I�K��Y��=���ɽ�\�����o8����
�H����c9�J5�rY�R���DW!6����D{[�8lH�;�;��:H�+�j0�ިS��屢ոy�,�-Pp�dR����*:�u�;��H�Y|%�
�:�������ÀB��E���>� ��	c�(���]L���/�R�7�CT���N^��H�d�9�m�1�O��}�ؾ�m���$�5M=La��UXÛ��=��?�E�(zy���g���� ݂�ɴ(�-��]1ͷU��8yH�FoSjJ��8�
����=��ʂ/��$�����a:!�K�C2�Ld-�� &Ǿ.�g޽��	��$�7��Z��Wt���u��R��Gȋ�,��ج�Ū�-(� 
T�(����i7�!�4*��@����0��?�4�#S'���C��y����Yѻ����֭r	���ay�ئ�*��7�~tGyu�n�x2����/5�N3�(������b}����a#�wqk�Qq$tM%�yf�8��	���$����c�D;�ym55���~B��NZ�</7�x{��n(���]=����-|)��X:�ǁ��m����ts��{���`�,�F���#��O�����fQ�|9F2� ��`@��G�DN�Iؔs)٧ƾ\����3���:%����j[�F�=�Y������}�n����Ն3+��;8�:�Jߐ���~���:�@}�U����Jk�jI�Y.�e����o�E��"�xv
��,����T�����ciDJ�C�Jf{��(�	�%��"������"�p����L2w���E<��ZE3��[Q�ͤ���ϻc�=M2�v)QM�H�Lr�ۈ?o�T1ND�UP���Y��s�z��*WR{FR�
�M��F��Gk�E�p�,�.����
�,��޼��d���r���f͘Z:�c��-�{���amղv�/��	��eY�\�en�cX�;7[r��l-a@�aB4W`�Y'=Hj����ӊy�&)"rN#��Pϔ}H���[���Zx(�,8��S���إuT��@8L�@g;���Q�h$-l��xjsv���r�!�8���k�H�w?ܜ�Ky���Ǻ)��Ŭz�K� X����J=���6�2��p�>��3K�_�#��+�<%ʧ��_�+�NoR�A�A�i�T�j�Y���_v��@���1���R�;ӾP2Z��FP�<U���������a�@�Z��Qa:xE���5��:�B`w��tj�[��_�ާaU���@�@��{�f	��Ձ&� ���$��s�W�Y�n�5���&6N�ϖZG�#CU@�N����L��.�����'����]E+q���>��v��G���K"���A/�Y"��f��3v�f���4�Dk�ߑe)�����[����`K�@R�%�jU�H����	K_"R��AY�m��M�6���X�p�eZ�=E�p�@g��b��܁���)�¦�v�K&�,m0��N__�`K�V��4�E�ܽ�g���)W{�l���'���^�p��+���i�{�iEc2�(�
r�����dg��d�|��D�f�f���,+[r���
��Ў˂X��2$O�)��[�5|��V.���[���2m�t��FxO��}��9��X,�o����"�!]�=��c�
P�Ź��&�����_��e[�aGujf����s6W-8z�?��#k�ϰa��]��̏�p1�7������R��l�����&6�V��5mR'�X �J�Qׁ���0����V嘃y�i�������"F����� �@��US�Y@5'�c�xݙnlچ���⺧��fM)�<�d���_h�g�z�bR�d��{]���}O���AѾ(MEL���{� v��[�$��߽zu^�L͏��!"$[��O�����sO'��J~<�Qҹ�[eV��B�Է���U��+d�9\�|̪s�%�OI_4��c�t������^��c�){�ٟ�j)��W�f��B�p'Gj�x�x�������w!I\���eȲidxf5�{��*�/ 3���:���H7�*�$�]��F��ȆԤ�T��IED��<��֫"�H��`�:�J8̀��!���"�XѴ�r�绐?W-cFd�r���7���.�L;�Mn�Qk��Ýɾ[}I��kO��ӖF�C-�Wv�`i!��[0�3�&e �~��{	�L���iF�����������Da���3e��Ш����al.����k��-�Dy��B��ƃWQ<_��:o���~��%⍙�\�����7�Y�-U��8��F�>2�2�f<t��ɤ ʣ�̸ӌ��U�u2����W�b����wuj7���P 	�'2c�TU�n�<��B�5y�����&�(J�&����^����(��_�Ü�C���4fr��I�Ol��]���a��@*U�0o,(_�<��`]�R!�,�^L�Sk�S(����-v3:b(/�#��Z��=�LЙ�D��X |if�m6�B�W���x�KI2���2�x����8<6r���2�D6e��}5M�A�U!���q�`\��m��k�B��8fӖ��d?w�o��d����!�����9^/3(��M�7d�^)�F�z�Ȕ��*Њ7����~��¨f����BWG��kG�q����{m�$@���-_�Y��>ƫ�n�'Ii�Pޭ�,p6�E�0�>S;��>C�s�j��M��NMCr�Xo�M�k<�	J�V�ȓ�L/�7'M��[q*�f�����#"�ƍ�ۇmVd�òy������$ע.���ۇM��3�6����킈�By*t��އ1L���b6>����r�RM�vF�5U�����F�Y�6��A���J����nǊN�?q1�`�o@)�+d�ꥅd�yu��+&�<��k����)��MH����d����picQ��!K7�bN�������BL�#�Z(��zgȣ����ˇm�q���|juv����؏o$�_l��iA��5���/mNՀ����"�nn}�02�a�L�3^���]��f���Zt#/�!�1)#4�Qz3W�rY��@͒Tڑ��]��!ᑂ�Z�p���~��i,�װ>�U�{���ōN�=b�r�6U�c�b�Y�}�-Q�[�깊��9q<~Fl`���9)q�}Y�W:�����*1����yr$(�.��:�����;ĉ��s���9s���c�UJȧ��T^(�k�&�[>>�I���Dj�h�L*�ᘻ�<*f<A6�=P�_ll�vʔ4��+�;�l��	!�(��>�����X4��5��ͧ"�"A^hM������.�ft����{��l���<*����g�<@g)�-���X���������$3�жYi,�_l�h�~'���J��h�<6��u)���%��e/���-�}���Z���d�F�w���*�(i�^��V>��|<����U~�{�"M��d��^F��%,e�u���F�*.m��Ȫ�r��FYN����l�����%�k����_������F;���$�0ݾ��s�b>�!�q�N0c��k3�-�xH�t��y�6�c������{�VA�T��y��BNo˦i����զq.�G�ru��s��j(�H����dK��7\��hs�4�!��l�����H��u�E3�=�L,� 1F�\O���z�o��A�Cۃ�s����Am��<d|5�����D9D��r-&��4~������h��8A�pws����]���_/N]Av�"�IPL�1���l,h�{����z;�FN'�䀙�h3�ʈ��g�3��b�E ud<XB�������$&Ȗ���ux�3�����z��	��:�F(lb�IJ��~Z'D�� ���Y$^�H�/�`[rLf���5�?�3�v��n���bS5��ncq�|����	HG��ܒ����z�SO@�q�R��hWr�,�5���ZR�6��fah���n�[�2�i�5M6�U5�0>�o�==B��wV�S1{C��M;�sj�x� ��)��q��S*�!�ؤ��X�͢���,�ʠk��a�'�Ks���6?ڐ�(�fu:�u���;1h��F$����#���r;�wr�T�8`�j�|&B��TPm���Ɔ.������d�����N�J��c��(�� ��-wD�0���}
v`vU�I�Zk��>n������;%>���DP�yW\?M��o,�I �2s6)�w�^3S�l�q�;��4��La�`��Qj'.q�ln%:�����v�o|?M]�j�V����s�j4fD��0�SU����3��Tod��0Ͱ�W���?f� �t5�hC蜶~��qü��ά�����x�m���,B,vs�#��1%� ߿�9� ���}�v։}�� 'D����Ыv�`$���<~gBx�s�?��S�o~B8N��F����Cxpǲ���5m���л�I��C1C�ѿ������w��ӫ�pf<Pu��9�V+���;�`y�����Ԩ2_�#�m�Χ$p�^�T�.S!��'x��0GU+^�7�όx�+�o���D��NI������>�m����E'����aϦ0�~��N,e��uP�@��9,_����M�X�2;�6f�|N���VLX�LJ|���5k4����(��L}X�'>jL��j�a|!�s#�ٽ��k�h���ܷ���I�Y�!�]�m�h�3�Z�Y���1OH
$�r��$��&/.Kh�9���`���̈́W�D��;����}Qy�îd��(�K
P�oZ�n�M�r2�0@K
���PS�=J��dG���SnC��&ĚC� _�Mx�@A�L"yQ�����NasN��\��P��H(F�0~#MXͫ3�XWc�]{b�vp�!Re ^�c� A��y'up48&���7"��o��R��A��a!�D!��O;k�ི��J4�[P�;T�Hhka\!�;ʡ<^��D�I@)���A�DY�k��������#l�rz����8WD)ǐ%P�_Ǌ1[�:��Z+�'���5;�[���r8`%^��s�����:W�l� @�t��p��q���+�P�^W���*N���hNZ�Ｇ�x�JO�Pq�3�cҥ(����������nϬi8�Jю+N�=�д���K.��'�I���΀��/�n�����
�Y��9�$���NS%qs��h����ѿ�B̥=3\�I&)�^�`���)�ǆ�6@?�8���}��Jز{2��c�X��?ͣ��o퉣O��MEe�-|�<�K6S�C=�)$J�E���YXRHaj��*D�Y�-����80�x���Rj0uVB�����W&M��d�]���T^�=��5+�I�=�h�3��9��մ���Wo�u����p��9R�*�?�h�3�O��q�8�/�}}�n<؜�}
�Z�>~��t��+ˬ�T�jk���L�m�\W<*�*�w.�32�T�" y�U�i���n{-������"<A,UM+���=�2��7�m'^|����F���%ix�6���I_�6��h����wh>:?��rZ�t���B�1ݼh �ꨱ^���;�����$���c��G`�"��v�@ <�>�z�yW� l���Ui�+����sVp.��e���3SE�����cnp�v۵Ĥ����֤W��w�+�����R��uߨ"�np�8���HB
'?3����^�`^�C�:��ƙ	�=ӱ����mM,ׂ�%��Y<L�k�{k����87��s�%Α�7�Q�X��[8�%D� �K��5�aӏ�~�,�y�:?�4�'���du��l��{��Z�8������������|)k���[P��`��f���*Bh�K�XK� Q�����)j#ן�i���OW�?��&�U_�5:�p��֟ȉ��E�|���qr��;9�6�li��q��k�Ƽ=�^�dh����0͂i�98|s�.��V�W!��'��@�����z6�"�ޯk��hh/g�zE�¤�[E�/30�y����I~��o�\(�-��6�:7�3�
o!:��x~0Q�*�f �t����N���*WG�cfWG�1�peЬyH0Y<�����/\`���k��Bi�7�����hn����|� Q��'�Z�D���E��[f½��33�~d��t����}'�4�cU���h�{��X�q�o%���܉�����J�G��#6�O���E�g"k�L���?�J��4ܭP���!�xA�n���f?�ZJ�|�A��~�GՖ�B7�J.�a�ʢ���=�l�L. m�.UOV6]�&�9���F/B����F�	��##z���I:�q���� p�X���3��t�Qޠ�jXgjbz68���N����$#,3�lL!=>^���>�T����H~q~�Z?�H�v���>
�AѬ�/SsѼ �啗?T0�iA�z�/lW*o��p���j.=�~^uh+�>��m�S����p�����a\��7ѓ�*M��o��Vi���U٩�!h�$�&{P�~�	ݧ{��Ǚ'v�V0L��ܵ�.+��_��(⽤	u]�2���)�m�fJ��
@�"���:Y	v�y��8��R���K��vm��2���R]��v������SdO�_!��c�`-���8�����9:h�X�$$�h8��'�93<(J��a���џ���_�7ϑv��x���u$����!XႴqZ����!�����f:9��e����'1�FC�9J;���7�~V�a�]p�0�h�d��Q�v����m��h�j{��J@B�R�F���t�Eqqt�K���-�'�l����o��1��5��7݇��W/]!��d�����E����P����l�Ӱ�+-��k�#��z ]34�`�S�%�uNN�2�	��f���/��<��e[�E�z�v��,��9�Tl�^���b�فߤ�^��|*[84�.F2m���
jX�+�X�g�ũ5
9�@�d�aV�׀��P)dOh[��N���C���r-px������땤8��ۗ��%reF��1�s�	��T���J�s#�dZ���n�1�>$4�M��M:Gl!	"�k�,ԟ���ZBzt�%̺S���l�MS=�մ��-���Գ�4�_A�<��.̘�7piN�5��x՗Y:b�A�����l\�ǵ���s�J����}�W₭�!�b�N�|���1�|���%�%g���4�,��ė	r�zcZ���~��-ɮ�=�e�	j#�E5����~�D���W��(��m
�3 �;B�A*��8��92�R7^G�M�Ҙs����z�G�v�k �$��V�Њ����`��R�MXF�64� 5�L<��l��qLE��iZk�5�]�g���e_
!Ω��L�S�O�'��s��%��I;��Ҩ�7�Q���1U��eϜ�����e9e�z�������+G����^�&W�C�����>	ƭ��-,_��'?̞�e�ގT�,ܢř�W��������ك�K��ے�6��,Po�rּ��$p#�Y����U���QLr7�I��]�B��j�>i��GY�"�g�~k�}��������z�8�pV�hFxG+�y��ˁ��u����t�z;�g�����wt��W��G;�ݔc��u#u��Cڟ�~�x��O0�<��.��r4<�>�<�M淂fJ.|�49J7�!<K���0��u����/?/��g�/��~|#�~n��e*���pu�7K�/K�΃	���w�����_�B�NK}�C��e�Wg{�\��Δ�X�g'|H�zS�؏q�o8�'�Y�'���d�e�r��kk\ 	�gmu�a?G��cYT)��Z�H�J]ɳ����=&	gyR{��~����m��!�MsE�4gEQ���$���� -/�D��V�>0��FM��#R�,q�[^�!��o�����O;�)Ej��Df�C�o�{�/�:�~؄kMڡ ��ឝ��v�匪�L۝�c�Lc��z�&�� F>��UQ���v�-�
XV1\W�����w�:���������=�;���v����5��Q:;.�R�_�lG�����[���T��b9-�3�a�S��1?Y5lEb����bEWyYiSh�='�1KIxj� ���X�Ó�XlLr�i���|���(Y7b&*�-AU��m�8�7�ųC�w��+df����|�&��!���pmKy�7�B�
�v���������'W��f=,k�w�b�47e薕Z�ӯh��&пW�v��f5y6�Z��̛��i[>�=��Z4�Q��)S�TL�1:�*"�-5�b�#��G�'�!��6F)28�£�&�]�˶?q)�|�B$���B�p�b\�Uo��M%d���K��T�1��a���XЪ,������f����Н�}�<j�y�4w�7�-Dy��z�;m���z�c���pk��3b��U��rV�R"d��¥������s&�W�>/�0�.qT���nhdXBQ3$�^�4��·9 XZ�M��v� �y�Ёv}��W���@��A2m����]�?���D�n�'%q4bu���E���E�f�H�놕Զ�jC7b(��[I�����G��_@|E��dA��\�d㆕�+��Վ�f�o�ޜ;wj�{FeA�s�H��C�ZzhU)�p�9��id��|��Y��;ҰQ�LH�P�7SJ�팕�%b$,�ƲW�]�h4��y�-��˸�
�WBl��k���8�vI��eM�~n�W.�Z�'�,��'`�=�@{E�C&�)ؤ=�t�}��^�wW�H�I�b� ���_�m��ItO}�-_O�'v�b,䇅E��s�b�Oe�w�k �Ѱ���)Bw���KЎ,��`��61.���}V��c��z
�5��!g5a�a�WoK YU�}T��Ed������.ȗ�C�T�q�߲;�ء�Ҷ_�L��P�~ޘ���^Bt�h��f9�i`w�<��sM���
��3�7���*� ɱ��u.g���ْ�jܢ��ĕ�)�<�g=&��X�F�L�(�B�TTO1g��y�?���6��=bK|1@a]�J���u<�ǝm��Qd}�Q�-W�&�t8ZH�hɳ
��\����Q��uC��盏���s؃|�U-B�U6ﾈ�������(��K��� �>v�T�n,T/��Xv1��ۂ�&��$�;Y���u�����5���tA������;&��Uʖ������)��ݍ����r��4(���x["}1�B%��'?��T��`�K2�h>{G�F�Ѣ�`�%�%N$^�v�weA�5��٫�Ģ��𑿷ޜ�
tО��5[�4j�7�y�5sN��?L��d��~�W~��`�����4e�6"����)"��1 f�v�O���MPe��Lj��STIB2@�����*r:��4�]_�6�ѡ�`�g���}���f'�UP ���hR���)F̮җ�8��`zsC����N1($
��g>�$6�J�D�~����ʋύ�H�.�&:�~����XO����<H�O2�La�sؙ�k$y�3k
b�Z@3�t���=\> x e��X$u
�l��%EQ����3^g����s"�̘�KⰥ��
K$J���n����2}�:_S�,��L$���6X(��p���?�/���/�F���(ۈ�C�'p���M]���鍬�ƽ��-+�Z�Ao��ӵ���{ �\>�ݾN����<5$*�h�����S�(�����YZe\c�p�(݂����ۛj���M�4@��R�+���[�ԧ�N��W�X�t+ٚ'���y�T��A���%��T(4)� rז���	;����tא��H�W�>��FԵs������T>9d�����c6ꡀ��Y?1���Qj�˯��m�v�I��F����z� �mP�@:���1&����G"�o2���-�M����>�4107_֣��i����];!#,,ZЉ���ج
P�B���"�%6��j���5.�s<n�H~O��nJb���\ꁏkPN4q���C}9��n
¯/�I3^LC튑x���$.ᾘ�6\�)i��Eid�$�����X�}3�B��t��i� �3i,�vv&�`V>�c�\Ogց@ȩ�)!�r1&�.5��ߋrm��ԗS��_�UC��7�9A~��w�[�bB?=����%��ON؎!�IIC�(��[��3��
#�b�ֻ�ņF�΀S`�9���!�l1ݔ��d��~��_f$cX���{aeǠi�;�	5���ȭg̴�;4�����Yf���U߫ ��%3c�̀wp����_�\��O"��8:/���L�x�_�j��y���LI��T�x�[�Z��E^n�g`
����Ǔ��ڟ�������;kq�Ł	3
 M��O���
+�Q���
��Hl7��ju�m��@���QP�W��uUpE�K��F�BU���V��&�O�vP.�h�Z����C D�';{ ��� Cr�|8�/O�_�F�\4B|~��@�TC���B�/�9cv'Ϗ1F�>Ȗ�f����%W5f"��g�vxH_�@�4���j��^�t����
.:��+�Z��Ώ(�!��X`.����ޜ�������g��ͬ�s���λ*A(c>�N�ɷ���;�T�����©�]��]�a�u���� j�Qsg�N��y`9%E�,�'�R."MRo����-��9KBó�i�`я����������%i1uLM���ΰ���^����ᅕ�]G/�~nO���!dD��D�Ko�E�#�Że#�V�o���mL�) �U�7�7��Zɔ	�Z6��~K�������]���+0�nҔ���2�����*�n7/��"/���Ց4~䘬��b��-�)|`�h/���^	����R�����hIj�?���J��q^Z� \�@�W:U_K�q�>ŧ��ߍO�ea��Uy���di��6���q[P�?j�5l�ˋ��i�!����c:���S|m�0��d�^�O��E��� ��l�qXL0ܗ"W#�'����] �Bq��UL%��t�z�ba�"*��>'9au��/';>jA���a�"��(nFÀ��1�Ә삼�����-��mE
�V���{{?JzD����{��*��;���R�����O�x�]ty�GV8荢Q�� ��Z��s��pS��N�+�����#�4�Q�|�K�׿s����Vh��`�#�_�a�����z'�S�����#���,����D~�੹���k�N��Ir�5YnB��
�Uo34��Z�#Y�u�5�wÙ-��u��4�X���5
M�hĲ��1o�����B޷
�2�G������H#���v��U���T)X�j��}iÚ6$jߗ/V��������'f��_���,�sXc��>����=mG���~��#��M�m��n��#��_i3g����:%#�h'�ܱ|j����������D��=$��]�\�PH1�h�	�hPɾ� �ɣ C���v�=Y�#2}�5��k#��j؝��\ԥ��.s��w�VP4��m����*|'�#ݍ�Z���޷�Rs�䓠Ke7����_�_:�&d2��[�z�[��Ҳȱ��Y�}�$���wi'��G�e27��E��`ٳm�O@((3�Q�5N�]7��s���{A�r�](�B_X>�u�g�o��X��q'c�9#d�{�.�-(rt�����d��P�ں���Of�O�O�ێ������eh�\��c.`��ΐP�z)���IJ�P6�x����Ƶ��2S�`�� �	R� �{��$�h�n�4\����Ƅ
qgSW��E<ˇR���`�nХ�I��Ư?�4I�B�ɢ�넦�"����)YU`�@�'e��ƞ�U��𣎺ĩ��SU�)w�K��px�a�F�ނ�]0��T������V)�-�i DaU�A�yz;`���~���o_Y�ԣ�%?��<-���{fS�ͯ�4j���1��,��ot��&AxUm�REV)�~�VZ�&F� M��D�\��r��8�^5q� �'a�U�=����~�T�d

p��0�"�_�9M/��<3� ������*+���5e���CG�=~�e�b��EA�]i�ލ���8 _D�I�ڴMX���-麋�Xۉ��Q��8��˩!O��_V����L��|��ꯠ� ��N��]��A�� حKS�*�1���(EY��G`WJ)�e�O������JI�\sͫ�n���bn��qF�8���i/�l�2jw2�l5�)�:�Y���8��$�ۑ̒A|QƝ1$�;+´Ը�ȃX\K6����%CE)�1����jё��D�q׸���8��P�ĝV��m�+��8��KjN��E܊����x�Z����El�B�,���O@"�p8Yz��Hbb���؀h��21����#�z�a���Z�P*�g�θ�O�+�Q���(��}�s]u�_om�'s�[e����L:<8��wkDPcϠ[>��=ֻMYO����D�6`ޙ^����t���5�dCq�|]�D�Wu�i\G�մb���f�
�c@������ǚ�����7�鏞��Lկ3�,���$p\yg>�
����kV�請hh�r �5��hK�Ե��N�lCB�P!-z��u]��E��RJ��>�p gb�*M�a��>)Ά�un�2�𨳺�K�f��e9UB�(�*]7�f-������[���/Dq>L� �Bu���S�5P���/�yq�ʽ����)��s�o�W�_e��{��~�<��A�=|����rRaݧn�\ۨa.ڙ.r�w���w<��)���$ly��z�<F.iʲUO�|�a�\�M��2��#���&�/Hj��~�a�����[]�Wd�\_��̣��I�Gg<�zWt������C!��>�Y+{�a��h��"<�-��ǃJ����i��3+IN���Ë1'$�z��E���T�P� zp�I6�0[T��~�@K����b���MԌVQ�ai���뢠eDڃ�f�?R�/��lnk1����)���ݲ7>�`/y;ʙs�;y>�	��IS��1t�Y˲z����4*�7+e�E��з�Z+�Λ�~�  �3�O�m%&��=��"!!~DWd�)�>����b���1�ț��
�� �����t�y]'$Pͪ%��z�=�PuN��J��i�p�2��3��&,@�ԗC�~)�u8�ʰr"������0����K��ՕJLjL�5:�TQRu2�<pJ7�O!J�=���&���4�To��~�?�cK�l��$;r��S��/��W�P&~�y
����捧��8�n�z� K�qD���4�v�g�MϿ��� ��Um�ZB�8 �WY|<�Zn�Y�}�|C���)q����M.������pT����۝=E�y��S�%�譹�!�2��Y�}��)I��T�̷�ǐ�!}��o�5�����ic�ɂX�\�{5]u�W&����,ap�B��hX���0���t�&`�O���R���̑�b��`­�p�|��Z�ۯ��ՐȦzĴ[��h�%�ڟ1���Wy*ٕ1Z~`f8Q���!y����WY�s��T�4g�,��US'�<^�এ��(ӟ�s��&����4��=�Z�V��d�FDG��F��k<����z�`�����Ѷs���'�ClY36�,F�����Ҭv�*�Y���T��������/�R΀wD�X
+�P'��Uj���L��sP�&�w��$�w;�+�E�D|�R�Ư��<�A 8����0Y���TX�E7��B"�^�T~T{OWUR���r@���x0�.��dkV<�Meٍ�P�0H���g���׾��X��Ob������Ge݃0�2n�Bc&x�!B�����n�����֠�_;*�&oҍ�Y�㼈!��T�z=	��C �@��E*��= �~�YW���8���l޿��咚o�ry����J��ⰳ���rՒbQ��z�=ծ�YQ��	Mh��
�=�P����o�K��m:&~�L�?~��|�:��=��ؗ�|�d�3ug��yL*��MUu�9_z�4 �Ю��:ujsJ��o��w.\��d�˙H"a����Zy�θ,�a\�V�`��=Lգ�Hn�]/e�c$�o�^�~�`�=���!����Ǧ��HE�W�ʄ���W1"�|�fzѐKͺ�"�͆�*����7?��O�B���F�iz�Uw׈��N�s�<	.��?GW$IA
���,tϰIY���WF�̿lD��6��܀���˼��q��l}�l���~CU��O���N����0���q ��{��Q_'�&L�����z��(}HǇ�/���������A'!p���$�b+'�j�-�������$Z7T�=�Uҍ'�Dq�f�
�$=��6��#^���i�N��^���ӡ`_O�Uڮ��\Fͯ���#�Tc33�2Ϛ��h�`�f��]��h�v�lTAJ��<�8#�bq���Mᤒ�)�vy� "�E��4d�W�j�YPG�<^"����i����y �1���L=EF����@#~u�]�$)"��ٱ�1ńU}Kq�H�z���5Dq����b)�@̲�}�r5	k2zW}���9D<U^� f�wx��y�<l�
�l$=�E�W�d">���'��������:��a�(Q��D��%�4?i�'��L+~p��F�׏������&�m0U����E�kL]��؃�,�ޑ�ȭ2T^��[�K���<������6����ɛ�ra8�BF��+J�}OD7/�tϙq���=gC,U���Y_�H�k\���a+L-�l���˶)ܭ��1�_�G)��5j�v�0C��v����A���촙���N����z�yӂ���!.��(�&F����"u�ź�e����P��sq����/��xw�S���"�]2Y����Z�Û�m�\M"驃��;��x&Z����Jv$��|��<E&4�� �ZcQ�ێ�:�*�k�)��u�A�������T�\�H��X��-�8��߬�����ҩ'�U�&� {:w�������?-���UA�̊v�\�f�!5�ݙKLA�Dڵ���rȉ�v�|�_H�6����\;�~pL�쯱����L���c�^+��e�*�%Y�0]����o����>&C���;r�Vɢ�4��!;OK�tJ�%�k�}|�����/V'[>K�ظr�결 n�ƈ�9�Sz��������'�Kn�t|0�!|�s������1z�>�H�*�?��Vc��<�ʡӴ�*o9Xn9rh	��9ޕ���j2zy��q4�	��_]m��ǜ�����w�Ծ4�i�F�7��u�
'��"&e���V�I�m�8uݒy$2cΌx!�t��>�(Ex�[;ذ|=nf��ovkmp�?{���(���=C���M��� �I�(^�3j�w�[Cc�L?�$�QX*[��!�3��:�|���JDfw(M�$ d"�FFб�i�R&B�1΀��y���p�:�� ���3Ǜ����yaޯ�@Rs3jCd��dr��?m�-�'>���.:�p9��.Ks�F���fc�ҧkn³��~��겏c8y��іL���yar#nEwk;�!�V��s1��]Z�G�>ʖ��sclSvBN����'a�w�B=͎����J�	�Ȏx���א{:�[qj4<���O|3��|Z���� ď����j*Μ�1�;�@�J�<`�ܰS����E����BF(�ίŁ[�Ri����?1�0�� { ��1�[���_~����fi%��*'iR�[���Y�*v��
Rn�R�6'�c�PF�4�:`��E�1@���0!ڗeۆ���"{Fk#LU��|�h�ڴZo���[Z�|1��OCY�$���b��e.,����+:OO�ƌVd@�	�a[�'#��dmrM[f��,�T=/:D0��x�	q�u��{gɟ�3aV�s%��W����0�U(�r�>��wKA��O���.8~K{���SVn���F��:�dգ���n%a?`�cU:��YY�|p�ڔ���Ձ���3���GP�I��7=� t=g���Ō�1���Q(-=�=�D����a��:� 9�J�`���c�Z����ZR�h��]�&�<F�d�r��͡����lQG��:��Y�ů���5=߳��a��T2g*1��)�av=ք���6�@�)�/:�0��7��[R�Y���dNϟ�>�/p0�q5!s�^���l"��[z�~�K-�u5WG��hHa�w�&���<�4k��B�F��uwKH��;$©f�]h~�~����'B�	7��\,����<H��4w���_�m��bc9kÛ�[�NT���STߗ�Iosm!e!�h�f�I％���xAֻ�k����t뉯�O���,1��2Ɯ�(�f�yr�����UK&��U5KO�D�uHjъ,&�3tn~T	?���k7�%���ju�7�{��=����x�d.�Ŧ�]-°�gZ'3�!�[��.�̕Bh����n�j�_HëB����l�kL��ţ%�r�Bڶ�9�GN欝K�z.�0���
I��Nn�0��L=PJ���+���Ep�D���b��,ǰ`��.k�-j�ׄ����^E
*S�p���e=V�6���/�\�#�m/�ӡ[�����	d{�2DX����W��ِ�5}!�%n�wh��=����q�ʸ�J|�K�޵��{���F����8g%Ҭ��6:3ge{�O4�5S��R�;��c���!��O���}�̌��%���ubzdϤ��V��ך� sz�㇭[�t2"?�>��=�I�y��=M.��YD�[|dl�ָi+NK鞲�&�Bϓ"��q��dI��z����!�_��ܰY�y]I&�:�})�D��5lƗ�^����U-���f���";<�@��P?���Q�D)~)���Kt8��kͰq��,�n��\md��[ ���X�7`�+�H���H�9�M|���0�U|��%/C����,��Pz�QN>����ԿthY �y#�~	�=�?�u�HW@9ujz'�qo�#ȰpN�����%�[2/*%��o ����eɖj#���@u�~���l��G{T��:,����~�+}��ㄣjU��5��U�7}N��S��	D���Z�efπ���)������<�=� ��U�T(���e��Qq�6����!Tԝe"
	�P.j/= n`A
�U&��0U3���i��}r�v�_�Bqu��s�P8��}�5?O�*bj�v���c�^�Q~S9���p\�R�hb��Lt�:��H�����+�ȫ�mg��<a���b���GƐ���^���Ȱ����ͩ-[��J$����� �e,�c��ː�0�O[�5RMr-^�L�@_��hP��>4�s|�J6�87�	� ��\f�	�A�/��1�T�tC��xy�0g^��^2�->`s��h8�Kz����z��8���v��Ϯ�,�" �5� ��?h�N�H�������	�5�ۤ�*�{;<��U�ȁK��Jz�s�q�1�8h�0�̂�b}Ǐ"�H%�?���"�v`���0圗�%�9N�a9�4Y'\L�욥m�7d$�m,f�t�#�)�p�z����Ԯ�O��"B���T��� _��Τ�sgR���/\�����ީt��r��qh��u�Q����bzsU�>����pG_m1D����#Q��,�kb��W��ᎪT�J�sf�s�ETi�����["�\~q��b�����P�ER��2�@��R���jy�<��/Qp'3_-ځ��y-�}W��#�?�8�u���Գ��Y��9ׇV�zo/��M��j�0t�#r4b��ru/	��4�Dl�8}�پ��-:%�r���'��^턍�t����������EF�̈́_m��fZ�2��Pj,[������kQ�8F�:�M�G�rzƢo�����
���m<E{��,n叱9�#�WV�f�7���������t{G�\zN�ĳ����o��>+>�SJt0�M�qO=�θ��
q���}��͂�p�*�k$�0V�3)��p����� ���0�<�����A�q�,҃P�3��R���-D�3�r��M0z�a�����f�6T�$|���J��[�ݲ�`��>đ�w��}�dr�H�;�+.��?�	�s�vch�+:j��*Sϖ�Jǹ^�������\����?��(,xJ�f��h�X��E�%qH�78p��Q�\��ϟ�ɣ�������RS��2���FN�Zb���w �g�-
�x9P�����t��FX�`�Y�dӵ��Rh]�`� O����ۼ�c���8%>�6�s�6����cH^�)aU:B��y�4U7ᶳ�uҖ��9��F��J�;�t*o�w�mH�x�X`�����Z��K[ɤ�3�}�]mmx�t~�6ؾ +�&�\Q����M�'���y��]�<�K�B����a����Rj��3l���$LPQ#a��9��/���׷���7�ݥ�|HfM���=�+7�Sd	z9`���!�U��6O�59�i�FU��>��I�2��&���I�C�e���؉��7ū���d�S�߳@\{�$s��
� Dr$mي}%���IN�㪲:����8rr8Z0ُ�x�be����ȏ0��{��'S�^°[�湅��h���G��i��K1�K2�|���6�2��7�q��1��
�\�$���K @K�����W�>X�R&-JK[�P�E��F��D�	S�:d�I����e�!��b�z�7д�h��`��<G�D�C%Y8E�؃@��K`�\k!�$�>��)C.a�����,Th�����9�>�	R�-ãIk�,5@������]�����ɉ�Zs\n�X@�Z*�� د�I'tz�A��HSj\7� U�<��U��R�قѪ:���\V�ѐ�͚�Ek��Hū����Ň��g�E�~[Ȯ��41!�.`?~s?�vt<HFo�%�1#�K��m� av.	F!~8�@�m��`l,!��o��\�ь�|L�2��?���dh��0�_%ѡ�jEx;��1���A���Mʆ�gυCNH�R�7�q��}
�خ���3��l1ڂ�y�w޵�C��x���b��u��5�Q��,���
���K]�G[�Ĉk��0�p�IDv[�2�.Ԝ6+
����&c�7B<'I$+ke�|�C3�s���y<�Fл>�\��d�:��l���=�e�2�$���tp:��J� ��S�.,���	�"qI�n�ʣs�(�4N+x���˕V��[�a�G̅�_�D��gd��"qZ׸U�M�?M�aJټ�8Ҝ���*F�!����8���eRr���5B9Fhs᧘
����X�����el�i�E���CC<0���,��u����0�ӗ��u�
��R���ERXw�s�}OU��u�Qm5z�=[V�i��}�������+����8}�:S��t���/��l��|ٳ(��r�������t��CX�԰�}��
\ޯ��n�,��N����[�"��1��@VN�%[�-�P�d�v�[o�wz���*�H�8�������и����-����j�$������4�n�ȷ�����sF�4\�C���Ψ3�f�h+��>
�-]�����2�F��!���| S
EUcLn+��6�-\&E1M�(��Cy����N}Bd}M	�O���'?V�㽴� ��	+hs�^x`խ����),�uF�9|�X�Iy$��w^�� n�.�L���M�H^�]x��9Bմh?����ͼ�@E��q3�ho��#�N�{}Ȣ�8}�rLA�߱6�7��4�b�Q�d�",�?O0�#ʡv���O�ъ�0<v?⚴�d'7��UBX��[�L�J�,��/V���D�s�eLW���S�֏{y	��M 9�g����U����6�R��+e��<1S����?��Q�!�l�x��Y�g��^C�QF��� �R��cPkL�#��&���]�\��y-�Də,)��i�I��>,��='�ӈ��������w��S0p�B�?N}��+�鉀J!�9�!���.f�NB��h|U���g�S��5��1�%��wMl\`��߾mhUX(�ߑ�ْ��wUi�w���D4ՇD�nQ�B���{.Mx�5��u���X凊��kvB0��q)J�7��g�����1�:�f����+/֧�Q0j�&=����Zs�4`��Ÿ����kYP��@>��H���%�qAWP��9�S'�����nT���<W���hiv��l�,���G�z��ݾӽh��rt]�邆��꙲G�q�8�r����}�Y�� ��_hj.�ݡ�r�K
P����B���ԦT&��6Y,�]�&��ҩۚ����b�VK�lƈ��^6�b��� ^���k��b��H#�f�'h������popp�!׮D	*3@*!+�ѷЖ��eV�%�(t���O|�#�������)�ܾ���܎����ioC港��)8��-�~?'����y�)�|;.+u�ě��t9r��~����Rr%þ��Z���?t�RX��b
����Ph��>j��~�Ĵ���%�f�KǍM�������G��RS�3+ "���	�_� �Z+�-*d^AZ�$51�sdj�7Ѱ�J*_{�zG`ɱ��/Ưu��|F�m'9��$�u.���kπ$ɼ����M��jɀ�4c�mG�7I�W�:~���`#����;�M����1����pw��w���
�x�ksX^��q-�T��4� <��hų���c�pd���|��U4�a=�Nk;{l���������w��G��-ii ��@wV��[�����8I��p+�����88	�@�?��1X�V����6�;��V�I!Tӗ�]���$�K�fhB��+�!��[�W�8�	ϖd�E��5��d��*?��M{�̪����<��,��9��9Ծ�O���]Q5-�(�e��g�:UH��ïeb)�	��Y�Յ Kx�[,��<?!�&��q�!�/`����EVP����M��Puj�^ �`)�0��vr�NJ(��`��2P5�M���P�Wc#.r(�K�8�_�����M	:Y���F^P��Ey#�xuͷ�)Հ�y_�K;�>��fC{e֤�c�{A�j6W~�T�t��(�-2.�g"���5oH$�֠u�L囍�{e0�Z����k�\8�Uj�S�H�[�� e�h�+�T��Ι�T�s�)՞|fɰ֧�o}�����S����x��5w�66�*�/�(��N��v���D�-�}�C˽h���}CDe��F钅�z6W�<�ϣ��R�k<�.8M�Ok�6�aD&��| ��AJ��^W	�������"��S�z߿.R�a��D�1�����
Ȼ����&��a����t���c��ꦛ�d������d�թu��P��H�n��D^@ko����,[�!*V���Ρ�[(RYǿ2�)���țܰ�й'ܥ/@�D��d���2^ir3t%�ɱ���^揿p��K*�#f:=v�aW0��68�?a	s�
�k_ى��8+�f���BY�Q���2t�Hds�tO+Aِ��I�Mf\�qv�9�Ӎ���8D��'u�1�-��*���&+b ����$Ğ��S<YH �$�ޅ���>�jR�B��P�/���p�2}ɯ��]P�B�ִ?���(w2,rnޔ����s�>i����rP&�)� ��u���r���)� ^����	�5��U����q�fXq�n�ABF~l{�=�>r��!j-�愠�:�G�EtF�����/\X�bŌc/@<���9J�a���*W0���ʏ�����eP~���xB8�ɟ���U[�
YE�zL�f�+a҇�/�tS��Q�i�_�g�'�d5(#�X#]w�YF�[����$�q�M:o �ր�c�ND����� ��bZ��`F܃ݿע̻R��=�ep����*�+VFůj�	�O̬,�]i*��e�ja��{�س����u$(7Yc��R�*��pH?���d��F1��5tC�"SR@��U�)��A�o�H�K3]�3��nUaM�6�+DB�қ�E�5UTNړ<
y
`x�����T��TCe0Ό:����@Y�j;�6e%�ﰂ3�<sD��jm�� *�ϖ���)���<��.w8���HY��"�B��@�	����2���0�'X�m�#C���`�}�<�&��)a�L���B����s2�H��f�9K!���s_���`����m�Y!�JT�"ʭВ:���?F�Q�x8��ё�~��T���f��q���?O�ߓN�Rߑ�d�J��m���!-&���<�I�\������N�m��5��(Mfi��n�
�IeC3Q,1����5�� '����!� 	��0c��\E:�e�w�0����A��䗝ȒD�p�tS�h�MOW'�v�y^4^�֮����˟�����,������6�e��1P_�n7nS��Q(��5�>��X�u�Q	��Fh��@w�����S�`���7<᲌����93���$��{I�y6?#�l��\1[���������BM?k�&�����D���9L\Vx�ėE�j8�p���`���1�Wc,����BA'i!�?aǼ<n	BȚ(0�|ݒR@���W֛����Y��l�X����������������k����0�FiQ̆�k���\Uu�~7��^?Ks�7�r]%�f���6<��@���G�N�/\</�䎵rq,؇�lɻ�e��(3+���
hG�5�iq��ܰyn�;_�"���p��<R��&�'�}�x�~z��7���֝�y��T����^7�������z	����h�A(��r����޷a��rQ�.�T�u�҆+:)��۰��Y�3�2h+3�;�o�QZtkc����6ӘީN�B��<�uy���C<q�?�WOi���V��(�V�n�~�1��~K��={���|�q���~��w�'�'�o�((��/�d��m�Ϸ�_���c=�����@��*3H��Xɉ	P�6_�֕�+�aX�u�n#� �д3-FH�G5����X[�O�F��w]lFމ]��;����J��@Ǭ���J��O�e����x�� �4�hoA��/#�-�K�X���EO��m�pj��Q���  �w\�Z�1#�����Oa�k�З�X&1�C�j1x�ϝ�i��T�6�1����N�%�C+�<�U�'�kU����d�:+�5\���ɰ"f{�B���z�N�&:���	u��0�W���L��՟��Or9�<��:��D
�O`.���Y��q��n:�oWd�@�Dl�V�����X�4v���]eb�#ȵ��%�����'�ߖq�r�;���BX������`_Mu��(��!��`�	��eD�2�Oi;�N��6|,��;�3p���~��+j����&뷼Hv\��hu�Vpy���BO/� ��9o�о�9h�F�.����0�qb�3���������R�!j��Gvx���l�F<���"`��40��0lB��S�^��TVA� ��h�ri������o�����Fp��;�._��K s�P�ruw*��]Xo]7u�6���t�tvn��5���c�&o@Y=�C�~���q���A���b.޸\����<5o +Ku[�ih���c*��ˤ�vr/=\�RE�n�P��t� ����61s�! 꽯��Nz�o�'���6�d� ����u�W�y���E��PN�
j �.�o�As5i�~m����#ɞ�Lb�0��NSʆ(�?�mS�#�:����{��$��$�_p�/�iũ�hb����tH��KT²]ҏs��)��:MR��ޑR>�!x�B���0fd�0���%p�]T| �u�����ʬ8`P	ue����K�D�OE��}�Tb9L�g���d�[K��޻�������A������Z�me�����oS�� I�� S0`.9��/�'ynK& O�؛���m�8˺�@jA�PDh��}�)��~��(��Ӷ�;M�����,�ޮ���H���{yF����g�>,�Z8"�A�e�fM�	z�Uv�@����XV#LD�vU�K����璒�[`!~3����@Q�m%}��A��/W�Av��soi;��(�oa��d�P���Hj�T_dsT�b��$�k'X�:� �&Oc�S>
�C�T7�ILD�'I軶���g����]xk�����Xo[M��,#J�o,�M��c�^��F��H��U�~��Q6:P�#�h�w�h�Q�B�R���!n�MmC��j��?M��(;H������0��$8���'���x�=���,J �M�����8��t��~pQ�̫�c^(��V�v����S�D���;8��ӏކ��펏��3C�ѧd8F>�����3���U�5瘭�)����2�%`~d��F(o�"s`\T:20�spT�z�
�8�2�����z����J��«2Xl`���V��@��(T.��C&���<�������
|�ڢî.��
��)A�L6�H��@�3�]���A97)������~�Y���3�����3eF����{`�F��7��eF����9�.*�V<Gn3�l�m��f8*���p�<|���X��I��SUl�$������'�m<~2{�f�GQ�Y�n���a`$O�vm=�_1SBXz��ݯ.��JJ���rуM����S�}����	Q�u �[Nq���V�f)��0FvT�b�q��]c;��r�9��$���"�/�z*�F�P�f#A'X"��J��`�=��~�ȍ�A��a�5��T�7�Mr�}��-�0�9y/�y5����t�t��\L�%o�o�*��"g���5,�n��'P���H�`�]����x�=�F�l;�շH]��^�T@�c�����J���R�*]�08��ߋ���[\�F
�D�C?|��qF픬t��̕%nr���$I%�Xe�f����� #Q�1�]�A@f�u��71U�@8SEV��X��1�����MJe ��Շ�W�����}�e˔+�FfC}��_�}���ΐZ'�`Z�8z%Rcn���h?����nc��bL|!�ٕ�D����l,2v�_�ƃ���p�r̞���J��'��Iq�TX0�=����kU�˶��|(���̵n�y��k��	�+�H2�����c��l�4|�T��LdvGm��X�J�Wtُ�� U:�nh�2�&uvF��[;ֲ�d���+��c;똪#����R���MQ�D�Ǎ�^(�B��>^ٟYNWe�H�a#�������c&��QH�A������OF�+v����EJ����#;iLJl{k\6���Nt>ƞ�c�*��\�౵hg�J4�V�Q�G��4���\$<\~��s��:-HKl�fDY{gm�*I��91/^L+��p��%�Z�~&g@_��\n�w�DH`��TΘ�S��0�@Zf�r�}��(H���4�J�3ϐ��oe��*�脣Su@��6�p�X�{���dȚK欙G� 3�*�j3��M)�ۓ����z�el`�zuC2b�	.�c��1:_��Y���X��X�k�S,�7��|�m�| �<�I�c����p��F��@G�����=�m��i��O�/�_G����Iz�=��Ui�ݎɁQ*:��p�}C�S�x� F�ɞS��)���3��.9GD�]�*�o�k�̂�S� �Tר3�W�]�LȌ$���7m1���n��/�cIF��j{k*W{�Fx��i��b�v_�PXtp��}���G,2�l)xOi@�u7�7h�d�!NfG�G�w�ƣ�	;�"?1���gٛ�@��iB{Qei�y �0|�w\+7u�6N	�ϲp��%�u�̨+�P]�'mT�.�������!��W˥ѥ�r��tq"�.Qdj�э�	ނ�,|j�R�D�dXn��v�I@���H�+���&��_9 ���`f���`4�;=�~���� �<�������ni��
<�༩E<��٦��U\��0��(�n�#��:� :��;�gc�~����}�K�3{� �k9
m���__JJW)�|8y|����)�;a�<������V�����,��-9(��A�6!	7����F�J{3��/57=��8,f��ݍRâ�I��C��9z?_���U���A͂�Ó��-�A+ʛv�.�y��U�/��n�%�w���hP�Oss'�F^%߃gg��8fiFi}T-LBf~��8�SSOcX��i�&��N��omm�^����p,#b^ߐ�}��Q. #����vl�aՔ(�����>S�xQ�4���11*#���[$��]"��L(�0�j����/��p���N�^5h�U�{<h�lך��'P��_'��Il	��+PQ��̥0�2�&�D�����P��h?F�{$.�6r՟�"߱+N���FU!I� )�I_d�E��&L�9�XK����-��{��2������Rw�n��Z�W��lR53�˽%�HP~x�C�kDp�x0x����pȽ�7�x����$��55��N.�(�}��J֫׳�z��$�]�礤�_KWG{��m��6���O/se�K$��l�(�RB�u/Br/M^�F=�����cI*s�z�T^�DeŃ��ϗdTK��d��g�J@X�?C�g9�G�񁊏��䝛���+�i�4�ź�W����,��������� 0��48o�ȼ@�ξrsB�pI[絑���#�[Vs$�M�!5�Uk&�ͫ���:�ߍg�TC�Ɨ���֝�v�b�����ʳh�A������ݒ��ޗ�'�@|�������e祆���w�[�h����N�(�uS�銮�OL� ��bC������(��l���iDPiiUBO�"lvF&sw?E�j�� �2F;�=%��1Corc�{�Veeo�qE1hXF�F���J��z+����
���L��_ٙ����NL�j��\��9�|7n4Vr{VF�x��:3�X�6|xp9���`�墴��$���*�z���/��V�ɛ�e((3٧��8�4K��ҁ��	�?�԰��?ݵ(͘���T�����npe�kJ�?�͑�^�T���9
���%m����U1�=rTW���#1,�.�Ώ�H�*c��Rwq�Dp��X�y��Wa"FS��3N�X$�l��A��B鵬ÀnL��2���;j�NKî"�w�|�Jc��0�g/��X��'~L=��\��4*'; ������S?ő��n�=ouK��T�N�gP-ؽ�\�\	(���Ɠ�]�e�$�(I"ӷ�ib�-Q����gZ� ��zhYQ�M�[�4a��;e7[W��n��J��5�P� ��C~k�3DP�����'U�͞���w=ԡ4ޘY���9�+L��'��!�f�o�J�����1{yn�/+��L�2��]/�\	�zm'�Q����|w o^�:��j\-zg�;i�$�i�h�ʕ.�0��H�W�w�xQ�VR���6�a3�P�����Λ���]e&���bx��N��OՎ��us�6VLW��U��?��Wm���~'C� �Q��g�԰�#	�_ʷxM4�3-M�w��i����k�A����7���nQ��ANR�OQ���e��"���.�����9�vQ�};v�|¿��ђ���*��>(�9œ�-�r���[��+rT�%���b����&�xp�=	i� �i�J��?�Y���@�a�N��Ig��#i�,W!��c݋��V��@��������f�O�a�t<�H߲\U<c��<�[�LH/����C?��Yλ2W�tp*�D���5�~�G�����&����i�p�)�t�5m"��o�G�=5"+�c���ĺUD⭴B�E�g����hȆv���
��.+��o����<}���%Z3!\b�?�qgh�녪P���-��h>�ZB:��R���)����Z����P�S�s�E�+��6>�\&-U9����Nab�lkJ��q-�G�)I\�����Ե~�hN �M�1�����!��q�Eñ���i�4��RK����ݢŤ����0��$����;"^-'dy$ߚ��{�3����8|2,@�Sɿi��h�$'���ǹVy~�<�$��
q*S�̧�^�}y�Z��T#[��m�b̢�&�#�ٗhp����	1q�y#g���h�Fp�?�w�k$���=� �p��5n�N9�I�T� �طm����b�2���Li��ђ���9D�߶���P����Eb�;"BL��x8�أ�׵M�y��݀x�,���7BL������p �Q+7.��멢m.���������)���)�g�aQOy����̈�y��2�'����^�ƐK�"?+�i�vNa@`)����Aϭ+�X͒+��&�K��F�*H�� J�9�x<+�ܦ3���t8���6c�����3'��$MEy�(�[Y����ަ�y)"����3ZA=fʔTD�T
 v���ǭ,�k5at�:_�&t�:%�2�C2�Z9Y���2�O�2f qn�`0��F+'�j���s�9�C��	/���	*6�t�(���4Y	��g���s�%�z�(5g)�nS�`%Jҷ,�L�d�]1�l����8�]l�E��p��I��ƾ0�ڰ[)bL6���G0f�lJ�8�B�"��:HP���x����&Z[� ����d�G8�T#�s;����?��O�T8�!Hx�d,���V�Z���GW���>�6�}����H4��c
?�%65ʜr�e�^�ShЀ�2�X���ˬN E��d�tR���7n�v��9s�p���v��u�ItD9,�����"�
���q�Ws�;|�ͨ�\t2
�<��V�"!���9���!���!<F�֊�I�qr0�+�Vmp���(n�[��D��Bc�3�@���t��{�|* I���a�;Q�1��e��G@�78Q��/!5c|��d
d���1�.��c��=@�f(�����tWUf��hUW�V��;���8���ؚ������m)X럴Xm0����yM_w�%c
�j�TdѲ:&��4�.�,ix�v��H���b��CL=���1:d�B=�\�����_��L!��{+���fN}SEW��	�w�0T�<���{N�
�f!X����e
�y+Yb0{4����6r����[�k���~�p�������u� #�]}���������5�����]N��S����;I�<�����w���|8���'_�!x�L���[����k��a0�$��,O��E�6��� �sɵ�zĺ�|
�U�?�w����P�������X$�YAt��b�+�n5��ew�>��ծ0H-t�`�i���wa������%�k�#�nÌa��$���)1��[��ktN
�#��+���*��Ǧ�t���g��4sl�6�O��$_�V�0$N�P���L�����pc�t�_�LI>�����3��I&4��]G�ə=a@�[h�nR,;x�V�v�١5���ːQ>)�3� Y���)#��f)%쀰������4�"j�-��kKDv�`�Y#�5��w�������	��'n��kB������p{=�@�>�;���_�W\Uw��`U��j9|��ҵ\��zw����oPB*�4�gW�9ztS�3�e޶)�
�e��d�γn�J]u�{a⑥ؗ�>�b&
V����&��$�(w��o&_=M���!���`���_e���T`�f���t5�����s4��Ҋ���{�E�aY��m���_�b����{p�8�VR"��"�h�V��!���\΂i�2��� *
�}@�dL
d�9l�^�Z���á �!��7*K76$7e�׊���x{0ܥ\�<�2BS���P�}m�jXJ#�@nADWދ���>�4�������c}@��L]��Yi7fWڸ|��{v�L81�^c Ӟ��7�^��� ���$o�����V�U W���|��DB�P��Ё���F�e��j�K�v�JR%XdUZcg�P�`DI�VI�kO���L��_[�5���_�q�f��|�k���×� ����[Fϼ���2�(Mݙ��p���m�F��>��>`@"�P��ڧ'�+Ф��SG�D9�ȕE�Vji�\c����({3`���z����..� ȵ�6Ҫ�����R��Fl���q���Jd ���4����I[�y@6@�����N�����'�Bn�l<���<�g�ۚN!(0p`)���\61G q�@��t�������I��ĵr�:�҇�4�N��G#�{��4�r���$k�[��*� ��mk��Bh��)g�����M���Aej6׶�՝�wL(�ʘ7T���+	^C�9g/�f.2m�M�$y�m�)o41T<;��d�-�`����t�%%���٬�#IB�Ԋ*�j/u}OU�����6��:23U$��qf����$��	�|�h �`Q]�K!$V$k�{%�r�����mb��V�������'C�����L��C�/)	J���*��c�))^����	��L��q@���<{,^)YIԬ�>Z�#���nh��1�X	��n��թ�ޢ{��\�A$��Q��(���U��(�w-�j�Rz�̀�f��7Nk�e��
x�r�ґ,'�"#,�V���J����b�-k���i�����V�X�ಜ +��z���J?G����� a��W��X3^Ŕ@xJ���Pl����$;XUG^)�z53{����:����ə@o1���u5#��m?�T��ܚ)h��~��)��h��:�z9�y�0��{��vI!v���0�&j]���J�^�i�ɨ#T���F3��Q�����:[��Z\A��.�2�U��[<���B��wU
�����o�WE���%�칈b�?�������[v5�('O7>޸���+�-EZ��z&X������}=B���a��6��L�i9�t�C���Y�Ħ��^2���pߢ�l�8�1E�L	S���(<w��N㵤F�X�N�И�F S�eX�j�W����E��m�G���.V.�+������/hl��������.��R>�(m)?>�<T���U>\c��� �'��h�&3$ק&4o�Dڄ|�4%��)(��K(CS>ckk�36�Ll�!�]3^-#��
\�1��J�D�mY���
���zO�7x�n�,VSW�� �wS�Z����Щ���mFj�%Υ�Zjo�M�Z��}�S#�;툛=��2�ΚK�Rŧ�h�ɶ��*8ȞL���$#����ݵ������{ۖ�vn���>�ڤ��0�F�z%���I���a��M�>l�hv���j51���Mg�������ﴒAGY#W^��x�Ξ�Ła�����3�{u���a*q7��*7_����hTKpm��S�"q�s�g̳	����W���Y�4Fo����c"��8��T`�mq
rU���U�~(e%�v�5"&�U�	=&߸�wS�88Z1@)��Y=}���s�t�{��ܛ��B��k�ĭ�ՑW5��5��*6/G�T��X��n%D2���g�B�yn���5��};JMv��ue:�#�U�P��J\?\��cҭ�2��[֐�o���E�����7
#+����%~;��\1v�~~-�:f9���?:&���!j���{8�E��Y؟س�o�P+(�	CV#�%Y��{�?�0��;�ɉl�U'��ؽ�r2�`���d�a~:90O�	f�@W��9ʝ����!��e�r�bZzP��z�B���S&t֠u{a˹l롁��u���(�� �	)C�l�2������^�~"�h�i�;�����ͳ��b=��=H����zH]Z|}��q��hkJtXALԔ�$�"2��,��|�*�G��Cr�C��@�ھ�C�}�+�N9W0��y�z�w�8M4�)�0�W!�B�bcK���mk�ɘv/�?�� ��@�{�t&._�IN/���8dMT�x��j<�B �s)�s��d,x�[k�9�v-[D	f`��ųT)=�Ԉ�v|Jp�����Պ�lr�lzӟC������/���#�P����uO�x[�
�#�y$��bp���)��-i��f�+O��ψ;��ہ�4�d���w3*7L�hp�S�tA}�f���: 3����d����haD�Ʃ`'	�G]:��ȣoW���zm_D=��r8��[��y�`��sE�K�Z�+��:�1j~�;x��Nmc9Yb;;�o[9³;�]=4�(t�F���FQ�]V�o��0��33�Xv@�����U<�Ҵx$���Λ�:.��Tr2r'2��U��M��t����9�Q�7|�!�a�+��#����x~�E�������
��U��S��r��F�Rg��>r7<��re�`"x��&��(���`��F) L`)���2�Y��'���2�b�t��JbY��2���sv��H��h��z�����b��J�����l HU��C��	�X<�\"���:;czE�q);y�;~�� /���E�_9OR��*W'SĳQ=�oߙ��Nd ��%��),E�wH�|Z`�g�_Ĭi��|Xe��Hj�.�jh�1�
f�ֲ�m�.�јyFh��S�3ټP�5�q����*�g2��Ǫ�ˇF�!KҐ�-�w�����O��l&�֮��h:;�R�K��^���o�gV�ՊTN>ڪw,���D�㹯M�����8�	H?l6�rҮ�[�,U:|<�����*hէ�����V���[��MD<Kxjp5�(%�9�����t��I'S�2D=�p���_�F��N6>ln�AN(�狲Fu3��d7��	��R�V3�9�p��_x��S��K򙶉{��<������P4�(�W� Bﱧ����/�yW�쑅Nހ͜��ƪR`���ԧ�f[�僁B�!�?�N� �ꗤk�ݟk����|,��{���@���V(���L��V~��%��U�{�t��T�O�3��S6�Fzt��(��S>���h7�;�Hg������]D<���i���8�#��`�o|���=�t���3#������-���moً�G�+��zE.8�%19D[�Z��!�ȱ'�A��fF����9� :�k�rvd�o�:U�`L�$r47ԻFS��0��	��Lw6SP/˽1����9�g �h�/�����GtJ���H���%|�
��LDr�l����49��0�F����9�6�W��d��V�B���ÌB� ^R�4m�6^���E�	�_�n�*@���A���Mӄ����_��	<#�}���(���S2�����^	��]?i ��r���8SE±n\+�m�p�a^Ƥβ\4I�^|�����De�}���%fV������_a��%껉��B(�ig,U�Q4�F+��~>-�ߖ$,]�ѭ����f��d5FtK�wq��]�b~	��8���h;�j(ZOW��]�@c��R���瓩��G�c��9����#v��e����GA���{��U�-Uxl�v� V�� �_�����쵡SS��sd�r��6$��xZ��Ib�I!��Y�zH*|%V]�s�!��#F�Vl������c��*)��{س�`�GA���Iw���a�����Y��i!�����P�\�rF�Rr��_�>��~��U��/g
v��	}�e�A������Bу�CV�
�L�<F������?l��?�t�'���X�{@�(�><���/<j�%��`z{�}���o_��<�xh#~DE�4��g��t����� �Ƽ"O���TyW�Ш���a'��F���v�t��B��JX�mN�@��u�Ĩ@�#x��άJ�M�'���m{�����o�T������k��L+A
�;6^q�W0��G2;�d�z�܆T��Bܨv��o`��7�����P�۲4��c�@��ו�f��WOd^������d0��q�aG|+�9a1��^i��/1�	2�u4�_b���XW3'j���tN��)F�*ݓ@�lh�l�/9i�? �
oE��ޣr�K��?�V����p�#Jm��X
 �'xO�/�C�V���So�a.`��Wf��I�*'r�0��eVg,&�����ꄌ_�Z�����F���qG�$�9�Ό�弊tc��e��T8���^��8��뢔"��ȧ�?�7��%�õ#\R�,�x��x{�?ا�n~�q���c��f�z��ec+gMߡ������{�	M�����4!�6m��UA%.�X �U�{G�X��_����<e�������	����DO�}������&���ql��√��h��J v!Җ'��M�Z�<~쓽-��������Q�u�S�"����VHWzV�_v�1$�����41�Ƿ�8�"@������D�b���)�;Eby���p�r����O�JAK	�4N�s��-�}�_}���Kl�V(�r=����
<E]^׼Й߫�J�m��q��!qV�ᣎ�8�}�˩�:¹�>�5S�K�!�S1��e�mRk�O=Py�� ���-�� ��4����Y��9��d�`�WF�v|aݽ��¤L����aCK 1~��Ǎ��-���,΂ȫ�lY�
N�7�t���P��5b-�+c��X7�I�Ql�"���gm���{��9��{u��j$�_jLTY��Q��qdVSv�x�Vž�!��|�Z�@�B:%�������p��Ƥ<C�u�?yhMf?��e�P����a2�m9���p{��K2�8:�!���w�'����o�A@,��Đ�@���?�v��dkAŅ�_�%x�~
����
0�Qc�;�t���M�����ސ�
�W��^��&�13Fv��^��(j��x��Yc�3T��9�f�}����p�a��JH�i��*�f��RmjD+�h�<R���h�POƚw�`D1O�w �K�>*ph����
<���oD�l����ҟ��\�6��b$Lţv�w\���l\��Sǻ�<߃I܌ N�5;z�D	Q�)BM������И����*����� d�V�8���R:�zzj>i��8�y��;o�H��Qcjj��y�ʑ��]�h��Mˀ�#��y�nkJrN�t&�,itLK�0/g��y�����P½H�d(F6�ԥ5��ԕ��v��,��[�={��� ���z�ޤf�8~Ą2N�!���d�D��m�:'�"T�kp5Gb���շXF�i�^K��W��H"�z	���{B��XZ�cw�4K1���)��ђ��bl֘���J߇4T�[�����5�8k��8I�LJ�:FA߷�w�\¨7݄=W�e S&
�݅qb�BE�o�`����ŷ ��F�|����tԷ?<��U���Ej��u+�1��A�m�~/N
�f���]�8qv���3�B(ǖ�g:1>��,�ss	?YO�n�q��U8}�A�B���B�Y?N�h����
����R\��hF�n��e��Z9~Z�����K�nθ1��L
C.<G�JH�+�%�1� �E��J�v�2%E�L��CSoe�f��%ԑ��OyV��'3C���z�>�a2̥�C�mV��������0d�*�B�}��(�!��{�c:��a��Қ���+=6�n	�W����~GY�\��V���@���������܍��?�H��D�������@βe�L\��eǮ��ɚ���G(7VfD2�b�7�������D�=e�����$`j�D}`(4���4	2��`���+E�_r�M�8I*ҕ��Rc�"�!>�K�C�'���i�'pM���t͂?4�g�ʥ,@�;}�� �J@�t$a�h��@������p�诗���V�*�+0R;*)���x%�U2���G@��#�$1�������MJ>�����% -(A4�o[���mQ��/I����!ϓ��}��8��,�LHt`��p�	f���o{|��O�ġҧ����ݜ(�ס��s�фع�f�"����!r�g��(6��*�ֿ��v����/��
}]��L�C�:L&�ţ��"���|��\�P���n7��P��e�������q�?�嗗����3��Q�d�e�!������+�{З�
�h���n�se��"6���!�7�j6��n��v���9�5O���5r���Y#<	p� m�����+�i�>Q�.w�'�o+�2�]������B�6gv� A��o��t����������gt饌�a=$���K�R��97��tk,��^�Vcj���|��x@�l���Y��ݴ�Q�OP����}�?<rp�7��f88?�!��C�&R���%1���VP���6�S��yh�p��iE^����q�w��{�(>)��an��aqs��W����7Y�ωt�[&Eh�ž�(��kP�a0���5�UR!�x4��d85=��)��HS��j#�~�o��Ns�j[�RU��/�-�`/�O���_�R8�F���ؑ*��^���cƙ|MEZ�fs~+E��ը9Y�דB���@��{��	�9���:�YK���Յ|��֐�`C� 4�?p:��#�_
�}FH�¨%/�9�4��_yW|���ӬR���B{^�za��yUGZ�FƵCF���H�a��5���hd��_וs.�������(y�jHQ?XkV���{��EՇǊ��Iv�7�s4���A��PoȘx�WRIe(��IV��:���m6��2�'����ε��OO�'��5�%2��������z:�����ŕF~��1ӹN���ō�[[�y��X� �9T�b�5�3���&M NKIS�-�pU���˔)g����j�������ԟH�{<"��	�J?BUla�@�2��	��9�^B)��ˮ%�/�b1��1?�����R�>â��,�)�lpR��n�e���p�����wE��9>!�<���H�<tͤ��
�7���KT�M^��G�:��b"��Sk�����?�؆0�����]:�P��z85#����]�IV��EƓ��|qt��eQ{�h�=�6�A�P#?<c�%��>���t�	 �pz6��������x��eNK<��#S�d~">׏z;�E������TjO�l�d>+��b�xu?�HV� CMukIHk%�K����ƙ��+Q���
!�-��""="���pq�m�',m��4��6,���m�[u�������F�Y�Ͱ�<0�:��K����0���9G�"2��\�R���q��E��B`�q=����u���e�N�b)��_�g��Iq�Ş�j��K=��'8	]*�kё������T�JK!�y�C	\�p>����)i���>�6H��y��i�G0��C�9�4����ߠb��	���L�����e��W1S�Q��YarU=�kQ��n[��i0�L�����k��IGe����,�Yh!���Ü�ɁA�a��g.ɿ:V&�3-�Σ��xm3gH�w�=�d��ds�f�?�W�����X��ސ�{}o�h�Ďi�@m�|����#Q�
wRJa����c!�p�sֳ�o�zEu)X���i����ԋ�F�G'S���3|��O��5 :	�U��	��\��U�D|�Ni8%����ښ�c�/��Q ��H{�����S��O?A��6�-��ɰ��.6���L��g�Ӣ�v��|�\�0� ϘC�R�׍�D ߁Z�2N��z���ʾ���������<�a��=�y���3����������mU���_m��fǈ�Hg���<����^S*Jd�Z�2c
����d�t�]���q>���n��]���bS�q!y5Þ�nr�A�ܲ���]�xP�x�*�1�[P���r]��(��JQ��"��������A��J�>�8�v�܏o"C�nER��d��ʢ�|�ߑq�T��+k\��7��w/t�[�L<������h�~�U����8����ֲ��Կ�I+eⰘ]G1y��w���ze;�c���q�g���$��)���s@A�gI�����H��]�x�Q���3���<�N"�y�rt�_*Њcs��S͉���X�c�Ə���S���S`�5�����p�uZ	����?��&�%'�n(A`�������t�5!���:�iĻ�~�-��G����0m�qI�3a>GlL�� ��T����J��3�Ǆ����`�"��pM�P�������݃�1����ض�6��)QAhwr��z��-���l������O��֣ȉ�mYo%�֣�&�e��Ӣf�NPsV�|E䈶S]W��|�HIh�#8��7���́9�M�f�^�Vn�;��`�Ao��d���E���;O��v�_EE���a1 Ǧ������h�L��F��4j���u��6lb�5Г?��~���#/4W�Bθ��}&���x���B�l�r�<Eb� ˣ�Z2��[�q�$�*m(��-${C�_����q�3V���~�,�k�@�+G51��a��B��JO�}��XY4Dխp[})t�;�k��+\�K5�J����j���o���4��~��T�.t%6����i�WHsBٸ_va���j<s=.-T��De��i��7��L�FX0�����+b� �9Zg4B�N$E��Lv��؜��ZZ�;�re<��"����d���6��
��~[����6�+6m�G-=3��2�	3��x��^�
:#(�󒼼�WJM�'�\΅�~Q��ȓ�%�D��	�����_��h�q�5w�[�X+4���G�;��� 챬���N�JX�f$��+AA��rDP���<ܹȄ�tX+�A�6�n<�WhR9F���9n#� )�;wb}��hRm^=� ����S�� ��wgY�s�W���1� L#Yn���� �/R��{�G�z7O�m��_�����`�[����i�˯D��(�*�.Hi�n~+�\�P]�l�~is`*�B;:� =��H{*QenGJ�7&�"�pF���f��C�������B��Ǧ#�fh��K���x���I�U$����Y"�=h=��i���	���*��04E`�'���'F�4�){a�(���'��|��^�AA��Ȧ���p�4�����W�� ��c� *��'�K�g@�VBލ̥H�m�}j�[��lLX�'�{:咽��Xo<�_Ka+�@E�-�ŧ1��[������w3�FV�����Y�	x�Mm3�3��"�{�[Y�I�h�ʜ��{@s�4lL��o���7ԬM�y�V��*e���_�Q$>4�i��~�t��@�we�Lb���If��Za��S�p�ͪ�+��R�p]j+�~�$ʓQg�x�/1� ��.���#�Ό��d(��f*�p�0�� ĺ��
5B>qm�>�_u��Be���X������i��ٜ��dw2�NGq{�f/RCk�*��9�%�&%/Ck;�x`��ߑ�JJA�f��5U-�.�B=o�O"7A7>B�2*��ZU6b��t���0�W<�D��0Ux$��B����[x� $i.��oV����!U��F�e.0*�볠B�sӾ�u�p�����+ʔ0��dX�`�D|� m���;��h1dh\� Do�#���a�jq3��i�4�h<ٽ��jz��dK���o8�-����)�;��K�����X��Ps�=�a��A�`���Q����J�o,}�SR|��󝆫�ޯS���c�u#�����48��?r=UA?R��y�%ó�d�0�M.�M�
U#fP 	�Ht���̢ߨ}��w���'3��������$�w�_��?�)���wJ�P�W���h�ᯞ�~�y���;�҈;�Vɍ���8�͊��G�İ�R��������y��i �unr�/��}eT_H<����������4��=�y9��<��ѿ�dAz�喇кS���g�}��'7%�WN�E���&Rw�)1�m�������$1�m���uJ_'7�G.٫�RQ���Q�pzu�+�A����4r-չ��\m̵H��L@L; 	B���?�6}g��1l�<E��h��/�Ŭ�zA��ӿ��R|��L��k�d���3���b��C�5���r�£
�}�ɟTPJ����_�e�4����q���$���?~j¤ݗ�
�z�
�̃���Ƒ�2���Bƛ�F�~mr�c���s�C��B�}V
{��}z1�!ف��y�)v�qP�����H�?	DD���g�*Y��"�u7��Ӈ��X���QtΕ�6<��7�X��Y�{0���y��WQ�u��;��Z�f�%Z������f��8��k�8��A�ǀ�?s�I�Իo��wf� �� k4	��h���鳤���83B�" ���`<��U[����%GZ�]��;�Y?�!E]:rT���� 픢_�g���*;'2��RP���� *���ؾUg?�2���Pb�关�����(����<l%�nF�UPp����}Q;���%R/�"J�#d�)��;x^v^k��:u�z�]�Q��-��Ů*A���	Ta�(#�� �g�����Ll_[���2�%�:[.S�z�M��6��"�9�SZ�Is0�:���+nG��[ꐢ���8}/B��*����#�����R�H�l�����T�
�V��a�����UM�v^��4o��1P�B��2�µ0�5��j���)Zov@��h�Μ��P8����sx�sg��"Գd\#Y�k{񈑐k|�p%K�X~���B0�$b�����]��H� ��T��f�bq���� H{�3�sBü��J��M���0Ew�K&�P43����m�����wHA\�C�>��L��Gp�����g�(~N�8��yJl�U�Tt��a�C��.�o�ͽ8m�4�@��ܮ���Fųih��h~nzg�_�o�:g�G�!����e��۫��!��
���p��;������-��%����	��Y�n�h��N��bI-r��(�X�Qjqx>	�ȀqE���d����>V��`hS����D�r^�� �F��茗Pp���M������f４y�#���Q�kMKe�z8�q=m��v2B;/�4]ַK����~��^║
,�k��S�Hd@;���p��h{]1��^]X��I������#��܄ٓt7,���`��� �ZGB�T���=I� nBZz�D���dl���M�n6���9�eF\�*k`[��&��o���lF[OE<�W���`}�&����1��
*��A�����LH��E�,o=�^إ��tBc�����^j��ǰt����n�7��*��,���e�.��u�U1�F�7���1d�?Է��`���p�Z�����������qN׽�tF�~��ߡ�����XnɆ���q��'�&j@wz�L{r��t&*Z��;6�ʴ�2�.�>c�W2��u���{,����b;�vL�}��F�����~U���,��:��K�@��gmu��*!!F��/���\�DS�c�K;E��h4��uy�p��y3�������Hz�Xk;�^7���5��~ޣ�<� KZi���4�˵��7xu��<�_����>	9�ٯ%~�0���v
��󳊃��9�k
��y���'��ř��ZM���5��
�)�xSAQ�4�"�,���S���Ĝ	�C6tܰ���ɟ�̯��buWcP	9膴�y8&�	+�,�����>�F�8�R�Ya2H]����y[��EZ��XH��Y�"TVɉ���P��=�ݙW�	�Ee_F߰��K�D[���\Ƭ��qF�v0�����8o-�ʥ�bϋ=d��磛NPް݊�(�4by�!��X�80�4BW�֛c��� �r�$����羅q��
7���#�B�@���ꆡ�� �/B���Z�>����1��癀��ܸj��]����gh�H,Z>V
�&��{B�:�gF���AW��6<ݗ��i��V�4	�*+�?�h�N����l���I%�r~�3�Fs^�>�s.D�H ��A�q۵�[��q���3{��2�
"�:��_Dvz:f>5av���k�<} �`;>�����
�R�4���wh*�sCK���Gw���ɰ����j�]���]�ϊ�%��h(r^Q��4��fĪ�>�xǋ�^� 3h�o�	��D��ݙ�7m�]<�&�O���t�к:*���R�m˃0KU�z�`�JIaB:�!���cM�P�nJ�g����0�,���}0��ɮ���EӉf����[�;�^CÄ*����p߱��z�j�����iW������,t�	I�{���'c�z
�޺0o�fz`�}{�$� ��OB%��B7 ��v����ï8��"G�X��_5��`k��hG�ޛl���O���
=��7a���+OE�<���tv��d�e�8B/g���e�1A>����P>]���0DZ�%���~R!�4A	B���[|���`|��g�S}�J��Uk�E��0���څ#@�'��Qz~�$f����$72-��x*8xBm�r�p_DS�G[[&�VM{�.�Ԗm�bOU��"4|��s�[�������gh�D��fQ9�l��C��ڶ�,��*�&.t&�l��eE͚,��K2���Y�,:@�c�c��9�� �S�W�-'P�K#}J�!�g�/�<A� #(pqgS�a���K���[��ºݪ5-�<vf��7Yc,��[�ql��[H&QL/��j^_��%���$��"G�ow�Z�4��+{7Kw>��H7:�>)E,��*��3OAh	��o��c��L�N�0�A��s�A���F��W�����5�gx���R��|��[�6�,r���IK�\� �C,뜯]j�"�C���`���m7��9���g��!7|뒕���#�w
��r���}�b|�\u?�U/�4����T���'y/��2��wб��}��ԧ�$.#$���agnk��5���h,�År~��g��9t��`e�?ߎ'���c}��-q��������3{p
��:z۳�p=1��1�jƖ�h��������O�r�v �V�#z��gwd�1@d �*:�Ea�</���;@��J� kS�� F"NI>{�	>LMc���e��h�6�Gs�?�����rUt�^b�4,|���u� 4�0p	�L�����9��K��3֚��OB�Z�7,6H�\6`�ىׯ���p����3i���O�rh��#�8���\��	"��r��瑗���9������N��V;ͻ>O�Q��@���\�Ҳ��}� F�?�%�/x��:�shɮ�(����*���Pӧ�E��Gh\��ks�]���,*��a)U5x�o�0�X'H�=5�DdU�?��,����ާ0[Ӯ��3h�����ƍe�B�_C�o�_|���w5UP��ك����j���'G���T�0��t-�K>	{_�����.D�Pg;2joY�=��uC�� 7��h�<�����*�&%��;=�O#�����h=)��%.)�q4,�g�X�C�� o!G0�@h��o!�9+;8 a�h�;=�5dL��r�;��S;-2�ԕ�<�q(�+A��0���n������{��\��k���� ��D3�h9({�(�X�����w2���ˎY��}k%R��~̗r$Lǿ�4��R�2�ί��N_�x ~x�U*mA�2�����̊N�R)$���}��hө�h7���ɋ�����q(�B�G,>A��
�v\�pR3Kc��"<�'䵒�̧�H���t)
���n��N܃�)i4�'��6�'��M7�ܢ������7�A{�,]�[��ww�S�(G�x���Ul�ӅJý�lԙ;�}��� _ꐲ��Z��,6����W̝~cW�R�D��?�a.|d����#-��'�'�q�mi�[�Z��&X�E�f#�	Mw���W��ɗ��1�5X*hZ�j��kM��œ<m�c_���3z�Qb�S�{�|���`�a˃K�mf�"�h.�RqۥD�/�7 a�IݜLJ�9�9D���\ڼVy�5lq	�=��S�̯==H�#@+�t�Yp�tz�Wr�q�)��}4h>�z���w����	 �B����϶$?>z�Ev���#��X	tP'���\+�]�]7,=Հ��e!�,j�Ⱥ�ϖ��:�}���ևu�6-tP˭�a���"�:ZMzs��6�ѻc��-]_��
jdZ����Al�ȁ|h}���DX�&�S�Ȋ��[��rn���*L+��P�r��Vx_��� ^��Ԣ~<d;J���:��H�,�#��ʣ$��ΐ���=��s�o��M8�;a]쯺Դ�#�	z	x tV�t�!��y�?)�mfk���?ZEϔ����w�CA^��wQ��E~`b�ɶ�J�:CLwi�խ$�@�v�B�UBy�r��C<��-V{���Ź�7��g��2�<�-�!��ģ'Y�ʚa	d$@�X<T�;j�X��I��/�FJ�!K���VϺَ���%UF3��a*~���K:�����l,�D���*�נ������ "z�7u�vG1�翧�����7K�8f�c)��ň�c>�JI���!ށ���Ih8����ui�@G�;覛D���%3MF=Ǝ��j��Ԩ�$}Y�a�ѣdJdY`/B�Ծ�1�Ʌk)��T�G4�T%�,���K>Ƨ�l5u]t���MO��*ř�gY1S^ ����^��o�PD��04Vy9d��bH?���kaj��+D=���@�W�����'L9A�8+L.K/3FVd���B�].'x�x����(�{WQn�� O����c`�����R���)���*����cdc�a����E/,^�1 ��fc4�>5OF�Rz�`P%c�q����)7��t�M���?9��!2f�З�ob�?�v&E�n뎆�zsy":�g��IZ�G��u�����.c���`n�D��D �h,�da�:�jwK�;�	�� ;�Sx ����F�p?-���iQ��(�\�4gJLX�A��]0���Jszs)8�͋ �?������՝�\��$/dk�n� i��Sg���?�R5XB�����p��+�߻y�U��	aW(���b�A�jv�)�Ӥ5�l(![�n@/�w��#(�2GZ%��`C5���S����Vгwّvux�e��l�~QU\��s1ءU�"T?�H��m��vL�LAi*��ʉ�B���t�����u~�F�)�E���;!˰�������,D�M�;�;u�����; ��B���40�\�%9T�<o�.7��{��COؑE����9zQ�kϮ�G4lҏ�|�S�u���b��#�]�v�E�[2x�}�V�v��� *�A��\s~I3Jf�#�kG��	x�4�	h�G/�[���o��h-�bxj�O3.����];��STR���N�P:�n�	e�Lٯ��w��!&K����:�Zzn���ɖi8��u��W�H	�W����� ]r��n��D�y�͞�"�=��<��cԴv�A��;�����mt˗����Z��l5�kc�`8?:�M�wM+����o�E+�}�ow7���@�E���o�
%c�)�#�՞L���k����9�4�H�a��`�����v�3	+lX�����'�����qv���N�̈́P����\�(J���y�\�Һ����22���#=�'>��pa�_u�J!&�O�� ����OʚT?�#��iD�H��ѐ��cA@B�|hC���`�jT�雹H�;_����)��+�e��IS����wEp������q/*|�a�K+������0�;cӒ� 	��o���U��JZ���$���A��KM?p���m���X�f�<r������'��^)�����Ԁ��u�su\?�;XN'_;D �F�����h^'FxӨ`M 9�m�%�9�)��Vl׎v�~^��2�b7IQ�{�� еuv�vkQ�����Ӗ�	u�[�*l�QkWw���*m'#�k�xxÐ��v��c+� �/��̢<b⹪�t����p��/5�p?��5���?>V%��<]>��{�6;v��6�߷��c����!�mG�6�^�f��B41M�KkʥeaJ���;f"6 ��G௨�_�I�0�SJ�o��x�"	���T�xF'�`;~}�,o谦Н�W@ �C�z����m�m����9�!��z���H�L�X������?��F9R�w��� �?Iз�9^��eC��84�r�'��zX��g��@=L�8(R��iU�k�=1��{��1��+MQ���9HN�����Gv!�pTq[�����	���5|�t�^�u7��J>�>5O�0���f�+��
�_ߖO���(&f�` �st��}�8�*[�óGc2�E�{NAv}(Z�>kJQ�ʇ�$��.H�����'l��0e:�7�$��.{+F�P���:4C�&�sI�
�4k��h�(I;
Tķ��Z�%vv������ՈpD�ۅ#0±w
#.q�aF�|�nų�5)U���i�8�04W�?��gA�Mm���$Ƈ��tE�����˴Y$ �e�!�[�`W����j�z�+�=��k�Cň�^�����#���?i}�+��:p�1����eT�#0%���[EF��2���&�zz��0�h�K�&���[�|ݑ�׋��c@Tqw�Yo]�yApc2���`�Ӷ��m;*YA����Fe�Ul �cf~/�_8�U9S���Cin�Nh��kH߉.�i���L�_�ZI�uH��c^3�z�4=q+/� Vؾ���B��Q��ns���b��<��q�u�!��}.5|Z_��-�����+t��D�In�{Jheߌ�����Ӭ~_��f�H�$[��M�y��~ɗ��FD{QL)
�E� <���B�~��I�Ե�C��
WX����5w���&���rPs��T#a�Kg5@�2�hJ(���A��w�-i馼�7So؇*��>5tk�n.uY���n�J��'�q�� G�%[7���_M���-�ւ��Lx��D��e�ɒK�w!�a�e�A���!��>˨�˲�A�9V';I�x2f�ֶ=:�#�X�����`�ף�b��zG��	P����įH+NU)O@�kW;V��ⴀ6�T�#�&4�A��X��n5�6��@�*���<��U	���f�s{ս0��ٚ��k��4k�W~��Br�&��g[�33��wπ�)��&�����,��N�z`��.���÷�����wZ>(6e��q�}�y�,�9�L�i��מVkqF�bt7���F�w~�¬I�%p�L����k4����=��y��cE�D^�����>��3|
�ѹ���@���t)�WJ� ��L�u�� ��a�(��<A�Wz��s< ��>܀��G]Ubt =3���4�{x�L�g����>r��7��\q{ؖr	��� �)C@��
ۭ�Ԍq!�$����0�����Wxa�Y��4�V'�e����90�����p�6R�fj>��0su!��X��9rc}f��9 �1��-�K~C%lo%�Q��L��>�X�S0׉Yf�ģ`�I�"���Q�H|w�ā�u���@+�G[��uj��dm��"xC���@��_̍升>8@�j���pa�;
	��_PJ�6鴑��Qph�E����[�.���4�Z����Ǖ%��](�Zq����dw����B��e�e����8��O�eS{/�k����`<�/́]phc�`�m�e���U.O=F�F'�xz�=i����<����6h����E=��呔gyd��j�x����e��Z��ڽەFT܊$�)+�����N��rB�Iނ�:Dp��a(�C͊N�=���(���&s�ֳ��Mf���_bT�Yb�p=l��"�a-�di��ݹn{,|w��۪��-�r���t��w�<P���r^�ڕ7=�%ԝ i�8Y	�5"+�	@RϨX����T�i�!Jk�ZVHa6���h2-�z�m��7�{���CU;�N� Q.@�� �/V���F ������'ۮ6$���2���}\�V��J�Rp��I����!�is�o^b�H�y�<bl���˝c�C��z�	����;os =����Y�	��o�p��宋��x�	�
ƒ])���� Xp%E�Bj��_�&tM�T�t��gG�Y�)2n7��-�{KO(~fg�&Z���c��7GiNL�[�{m4��� �m
�/s���
�A�-�;&v��桜X���]ۖ���L�!W����k������Jv' ���@�"�alB���繩-���Q��d'��'�#����]���2�݁s���'�A���&7�Be1� �z�ǽ��E)�+x�LE ��A[�OO��� �;�1��#FBf�c�W@��%}��� `��Ss� �����ɸ��H�2َ'<�8��J�qE��Y��&`?�TlG�p�B�^ޚS�8J�s�'�ERW���+��p<� ��f	7��\���M��D��s;W}����`N�%�����>����JR,R���*�ԖwM�\�������D2U	�%gR÷�z�(Xi���Ơ2 >mJn��Θ��KBN��]&����WR>\=��Ęvwj)w��h�M��9"d5�tx��D�D���__G{�o?�C�@���\I@	L�� ��q��`{|mF��V���ބB���sKr��*Y��uYEi?�U1ρ��en��/jk�g���l�;�D�o!���jZ
nBg�ծ|a�o4�\�� �-���ԥx�����'ס�[+�E���+C�A���M�x|�(��gk��0�ܞV￸k�S!A��dA�(���q�o34��G�G�bc�	�R��Ɖ�iu���s����-V�@�u������a������,q<��W��C����\!��O~��g@Ol�m�v�N2�~CI6�{Z����4`�O�/-�boS�w�U��uF�4�N��}-O���8ˈt� ��n���m�Cz�w��;�w0n��?&������}�ey�����%�H�P�C��@!�s:�irQ!]ז�[r��-ЌY	�w�,g]9݈<`����烴Y����	T ��/���N�e��I�B-V9�m�é?�m�C9�H}amQ��CQ�bt���6O?E�D�D`��8�wG|{�,HyY�WQ��
>�����azA�@c�5ǟ���@_�r�-����1%�R�/�uDg�|4����R	ڿjE�S\�͛R]N_.Hw�KH?Z].��-�8��FC⁽�M�o�����D7�*&t��4�nS18��s��:��LO�vi�v�]��N�����<K��T�}X��Y ���=&V�T0K̲�7f0�� P���m��e��C��b��H4��P���wlL��W>'���0ܽ��w��ڹs1�����,�C|ǿ<��ה��7(no�.���:ެ�9\h�u�gg{<����x�J�b=���g6�U�y;��Io�����	x���d��ߨ3�鬴)�?:����ʗ��M�[���ufk��w��M��������c#q��Ie��uA���:`2��V����S����8�y����9�&7�k�*��s�w���&��c��u��>��0��t���פUN����> e,p��E�,�>�F0[7�}B���x���Cϲ��(Z{__���9A}�'��ۡ� � ��NGs�(��
B|�W2�SW�D_��\0^u)�w��Y��.����:|���THž&yW���0&x�w_n�E�~�T��R#O���t��e_�F�����a��_��(Qk�4W��H�3}ن���Y\�x�C�䀆�,[졟��n\d<���l�`"�.l��Ћ�_��$c#�O� Zo�v�W'�+�)Ho�Z���5�����>���Z�`h����E��*ݞc�ބ�s^E׭��6���H���6Z�ղm�ҋ̓SG��x����hV"��M��X�w���� ӓ�&cܝ;��i�
6�&�N�I|l�+¾�bY�8j�;�4��!?s],/f��3Y|E��_���[ω�(;
a���Ƶ3<H!�/�x����Q|g,hr@v!VR���k�}ou�mke���l~ҳS4\�����]o�f�d�-^�����O�!?c���zZ ��4���p�ŭ�L�LȞ����GI)����X_K3����h]��eln�"8���Ы���[�l�/s��Ԕ1�;
�� ~�Au깧C��"�8�Tq�|�;�<0�T�=�Y����_c_�%8��|��>��.%B�Ӎ������ԣ�t0��┃B��nܟ�����~�2`���N�J#��cȭ��t6�f��t�?��O�|��bf��y����M��و�&ʐt�i������Ҷ�o#��=��������J�ۍ�u�?�L[l�:���a��\�J;�㕰��D2�|�l7�c��2�/��|?^���dz&H�ښ>n��ayV)��ДZx��P�81.�+������4���~+u�Ԥ�3�ص�L\�+��P�:���ܒ�N�j,RV�o�E�#pZ��8z��Y������ˀv���W+����z=AIZH��A�v�
�����[���L�pc�+~f5�}�F��|���F��y� ��VIk���'� �[z7,��KL�������9a�?<L"E��4L�]��-����x�=���Ȕ��~�a]��'5�nD�;X�B64��/h��ϒ���ֺ��RK�"���U��y�h�^�gJ| p����H��j�޴��H��g7Qv$�M�_S&ĳ^MO9�C�V^�{�3�\�5�������������Ky����&�h�|iw��Jg�i��k7;^���q��e(e��
��;�y��Q@�q �;v$r�C6�6I�4>l��}�@Av�sx���j!̀9.Jѕ4K]����Qd�`q�4���X[pȩ��ݍ��s�V�#8a�����|�"�	��]b��U�W4�Qm#۝\xfue�e��}QŘ~�,Xh{�%M��k�Ԇ����I���i��{KTb`�/��u\��
�����M�D��7����a"�#���N�����⫉����#*]�Ņ�x��[Q�Ou#H	"h�b�=�ȍ��Ŏ�����Nkx����6>��5�!.A��O���f������=2>=_����-Q�Ɠ��v�UK�@���*I�j�,s����>��ܿ/s��	u4U���SMo>�D荛�,vK�{�ft���}�$-�"ɌSn���ZR��V0QPī�.���ݩ��d�~@�	w3�-A��q��M��Į3�!�E:�#�ļ��q���R�mјr�佔6�~�L�{H�n%�D�������V��)���/���=�p*;'!��#�W�|v�nWq�>A/�ڮ�����tʈ����+�	�djY��W�t-$�@�ɦ��p��<���OtYiJ��'����Vb��Y��B�\g��r�;�|�pB��]���Q���d�^u#K�H� �7�_��8(I~�n�'�,��;-nyw���c������'B�>5kJ����J4?�35����2��� (�T�J%�LS��S�;�6����ɨ��5�/����Q�����>lۤ�o^_�ڑ '���2"�����?Y�5MZ8�u��>�p�J�xP���� �U?��`� ��t
[#bxvA{Tk���VG<�)��"ݒ'���m=6g�ZR����j���DHB��}W95�db���+�!J�:�9��em6��x���cu��̲%���{+n)%Ê)��ҵ����ǰW*��9��́4�-�2Lxڼ��9�Q�mј&��f��������ʘ.,��m�A��Q�����=x��+�OoJx��<�J	v�"��-,j�|�����z*�FoQ6B��nbU��8��+���;'������x<���6v��*6�$n{X�c�E�)*���8�i���˿�y�S���PT2}L����:����g��G���{�,�30��]���,]21�]��9����ðR����x3 f��~��h�� 8x�~$�=
���_՟6��@����dÉ�)_�ҙ<��)ɑE,�?�z7����&�l��(}!����^�͵��L<I_aDu=�^'pmH1�7��}��fJq9������֥ߝ��D��fФ&A�y�غ�(��{��l֠�>1��=��Z>���w�9�{�Kߛ��(!�g��(��q2�ǔjӔ�0F,�ZQ}�ag��;Q� _�8���=A�-�ų��#̛�$�G�}�U�����- S��%ە�w�)�<��:W��
��Y�e�u�[�I�z�������D��*Bw�&�q�鳯ȉ�/C/�k��hc
�1)��J�%��jyt��kZ�$X�����K�����ɼC�D����?m���[���m�N��	诂R��w���÷��b��{��e�y�wW�F�w}�7m����*b,��Q�}׺*|WíM7j����Q�Y6Z�#^++����f�ѿ�^蕰oE��� �_�w2t���H`����V�w x:���^3�B�����t$�_�U��� �
�/��I�g��.�w�u	Y�jrz�����P%�����L		��qʻ��x��'g$n���/��>�q��T��.�������ke���@�QV�!��m���d�fw}Mt������K���ʿ����H\-Y�뫂vTk��h�&���@�y`��:�6o����Z^r؍G�(��x�}�8�P0
1�:Kl�����n�]߭�k�� �7<΄
��]6��M��Hl��U�=���;4Їɶ]�Yڱ�zy/h��q#�Z�l��$��M��V��W��I�\�e�aA���H;,x~�N2Aí�f�-c�
���W*TQ�)ߙ0s0����5o�����=��}A\�C�����(:w5] ŀ�`ِ�%o`[��'��Q�P�M}i�/���N�P*%�b�Z^���Sq1����B�����G��7%~4�c�u6}~�U���[/�6MM/���A�W5� U�`�U�j�)4)��[N�6�|?T�"�2�N�jO��"�:Fꠁ�w�W�͞�U������viG�5��P�e>��0}s�{�.�O����@����W)�7C� ��㒽̬�9��z8�MnHIh��h��8�����D&��Yr��s��#��ȱ�4=x �;&�d�Y�X�Iޕ,����9̚���gߞ�/�96����=`�A��I�m4#Ҽ����޺>V�M�:N�éV��<�f���4�퉲�)E�ئs�*=Gc��_W:�6+Q�k���4�'�x�C�{9_�v�bm$5��3���5vStBڮ��̕+L���.z�0�l���v[���c�n6�)�D��}p_�;k�U�2M�wh�2�uQ�N3�`]�Q5+��ۍ�ۚ�O�R�v�L��~��}Y�x��;��r7�ƫ_e�W����Uؐ�_��T>U�B����P�M�^�
)u�DU) J�������6����?�z�6� �=� sF,�1���m��A�x��S6��M��z!LM;�,���Jp���L����-��F1�E��۾�h�<�\�Ep8�=��LhۻJ<����y�F������#��ã����ޚ��r��|~t�diJى�u]�O�M�F�2�ᛒ�,9��HA!dg4Ϥ�7�����U�X6�������.�md�@2����6��b��V�X 7���c�!oWIPX�-����-�D�Hl�qO�����íC#%Y�U=��E���g���t�"�[�J�}�@��;�x;�5�S%F�OZ��$X���N�o��K�
����eI<y#�:����⇝�E-M��@�Ƹ��aR-�ZQ��G�NȖ؟�qσ�d����K$�DJc���ڇ2w����Pb/+^	S�P)�l9�g�w��20�,]v�t�ǌj�(�ڈ��k7�y�%�� m?�����Z=��Τ��o�>�a��s�!N�<��(����v���>�51 @�E�l���HA"�I���C20�YEu}����uU�B^מ���v���N}�#IW���]d��	����k�q �=�����'ONg��͝�W��0�79�gV��+�4�.dc �D�c�t��:yJ%���C�%Fx��?�)���R�Ao��U"D{ҙ�~���I������$�Dk>���mI�m��S�LkKG	�}=Xb�fزn{א���i%���:�D373�l_��w����y���UH&��7�?�Q�����|��yn�7���w��J��'h����P�͟.>�k��>���s5/��گ_�ӳ\k.'-��E�S�Rj��v��E^���E�hӨ���*�?so��%�0&���^J����'�fk@#e�%�Z4c���O�b����w�b���sX���!�6����w\�w�8��Y��3?G��+Օ�j���T>"D�P��g1;��K���U1>�ai_E�T4bw���X{�L��X��i����/<�$��p���x�Эg�p��?��2:wS|̾���@�&���8O��X�xw�7U��<6&�M���ik�/���N#��p��T���E�7�z0%�vޥ� �%���S:m�<���m1R�U0�����P����ݩ�◼�h�8Yb�:Q�sU��8���4�=-�)�Ћ�W�=��Pދvo�Aɇ.��6�v�/S�(���!��wI�o`��ŴP+��!��õџ��-�SD^�%ckb�P8	RP@��]Y�P|a�������(�s寈�}υ�-?��{zڤ4�K;�R_ȁOb�s�?�v���f�������z�B�Lb'T�
LR;���)L�����TU��&âS�9>�>��4��^������Z��5�	�)��İ@�a���\khB�~�Ks�󨇗)1uV(M��7�	��Ԉ�BK�"n���"�$�@	�b`?�G3�ʬ��o0�y7P�t�1��젦OT���;?��A�W�!�})�FC�Ay�+긊��n:+�D��f>�"�#�3s��_Y�D%�'M��ܰ-w�Ծ-24��)D�GI�-d�*�����Gn@����L��"��N8_-�����k���tuΦ�&P�ٗK����;R�"0�`2,�����ɘ�LÜ�uy�Uj�xs��wn(���]��������`�n/T���Q��&@a�JZV��'~.9%�j���y⤉аHKцC��o���	���
d��N���TD"�گ�!����O�KġN�����]4����s `���CPi�G*M�����ܑ��lc?� �x��V��_��5Jւ�\�O KEg�����[�S5n� U�!qrh�^M�%��4��-iG�(�8�[��1J��r��ui8��.��������*�c�5�kf��8���"�e�ʈϐO	2���	!�g�A[�� ^	�wr(}R��q���|k���SM�yf���Apw��-��0�k_Pk@�V����w��S�|�����N��-�A��t,���_��q����gK���0����x���z�xS�C\o؞���⭭'�zX�f��y�/.B�q(��.����X[wY�S�.�syg�ܫ�XuL���{N�}�����aB��v�����7^�0(����{���q�i����Bg�
�A��[���c�6$�������!�~O;�����+hlN�|
�y��b3�8I��j�,��cT��ׇdvӻ>���{s�b�eYUf����<BG?cD��+��>���R�Bu������f�
4�}T���Ia�Ị�,g�I��T�1���$�zXd�T��K��U0E�M��8�l��c�m�`�m�.�3�"�/�5c��p����)��8J��vA�ل�W��q�Oq�:�&Ib+o��;�s�JG��gO2+ʸ�P� ;^����S�E�Cx\��ڥ�UY1w?;�w���T���!:��\۸)��E�UD����*V&���s�·bifT����Wv.��O`1�3����E�[���/a�vpov���Me��$�ȇ�WwƅL�xĵ/e��;�rb��Ÿ�o�ͷ�d7���qȃ���[0����w�A�{O@��F=�ur�,-p6��ˊ���n�Z�PO_��;���q��+�`:� d�����͗���ngu8l��b��d�(�:p���2w�?��%|`�0Kf!��NQҩ煅[�یː!)$ä�oo��߱l݆OX��2j��2y3`��5,�4���C5$k�q���"��|Emx�U4�w'-V�	�o�~\|cII(I���|h'����	�s�ԽDy�-��AON +1��Y��nJVx��t�:��ـ���V:d�/۠��tRx�q�Fb\���ax�D2c�Ŧ���&�_���J�����7Z�y�y�\,H��u�!)�x($�p�B~yČ/��d͈���g������:��]���J�B���������V)��g�g��ɴ��%{���BK��&�`�J!ɍ���S"��${��ZB��C��f�łӬE�WJ/*��#k(�rO�{M@����)��ř�7M.zӸ��.�f ���¸�\xeZ�h\���`�r��vll��ҭʝ��
*�q_ό�gm�j��w5��g�2�PBW�@{�Z�p m��pAF��Q`�w�fc�r���I�#|����h���f\綢��&��دЎ>5��
�1�cy|�1�����P�NQ�ggT�����ا�ȈDT��{Lg�^I+���/�?����驈+���p��� �H�m�#�Ϸ�ҝ1qv��_������Z8GY$J1�8GmP-�Y�����K$�Å�~������9R�w�~�����	6,n���9zP*��(�j�{�#���[��ET��7���I��L���f����#��Z�2���Xf8����&'>��(q�1��w�|8�Y1GG���7:�Zë��;?G���2�����̜�����$���$�D��q�/r���Ɇ�pv$fT}�_�� ~�Y�o}������$�I���C���퐫���@%_yKp�*D�z15znJ��j�z�z�J1w�����5�Bc���|d�zF��q�p!�P��];�"D��헖��&z��������~��t���/8�
)a��)���O�]�"����]S�]�`��Bw������
l��~��-�!��k�Z�W����;h�x�3�l�Ic�BEYN���%���7���yxR8Bq{T��㺇s%Mq�nÉ��`��c?G�c�>o)3�g��E�I�y�ּ)�{X:�T�iI f_����~��Z����0==�#5���O{� 若���ZI�՗�B�n���U'P�3RG���/;��7C���G`Er���*{�r��J��0���=��G>��aL�VR�������ze�%���q�[iՆM"�U���s�=�����*����k����t~Dȉ�l����"%X}��/2v�x"q��S�|;�k=�C����5.Zln��7�Bk���E�RQ��A!?�L|�.|,u����B�	�#/�Ҧ�C]���t�B�Aّ��8�u#{���~����U�,������m �wB�v󱰺��Ls&�C��7�ֻ�}V�����_������U増So³`j���i_s�2��'�Z؀'�ۈѧ��v�@�llT<��l,?��I���p�^��x�z%1Z��r��~�UQX��v&'���+�0k|�m)��cu-L��-9���>����w�6�`�
��/�}zY���)>B��j罉r�CW�?�>����kE[� ����>�{(�Vx�*���.�g�#Gl��t�eH�3�o�.cz6z�Q�8b��^��8L�69�1��i�f���X�I"@�ݵE|?�=��9�7)�WOd���K8��甊b;���- ��@��4�z�����CZG�$z7Ŗ��=��.�ѝ�p�����Y
�5��t�*��'3,	�OR쌥���~���ࠊ`}|]��H�Y�����i�VJ�,�AK���B�2��R�MM��l��;lQ����P��t���b4I>���v-��{�8��wwo���du�#a&H�Gm�_l�� �d�tH՞�ܑ/<'�J�x"�Ҳn���6���ll����������`E�z\/���>���`��ן7�;R��q�S����-���x�*���z�{��th�i��ݲ�������/�K���4.U���d ��2�FŶ���N��Hb�M�;G�Ox��+Xb��0�9Qv� �)&U~R^�lI�d����kE�x�+�2Є����2E��V�|�������(�2����j7�����=�0W�	gW'�^�L��sk;��%ġ���[oɛ#o	w��va0��v��
���~���ݫT�&+�(V��a
��3,�}6d
�is��ro6����,rz��j�Su
}��9�_+���9Ӎ��� x/�IJ||�r��I���'���N4��z���vVJǲ29�N:�"}�aB�������>՗7i<I�5��ٓ�r����4�s��~G�D5��`%�H����J\s�!�ءn���R8�̇@��F����z�k�&P�`�C+�e9q�'���[Y�-�`\�{���צL�7��z�de"�`z�� 0��'�(,:F���$��f�M}��7��l�Z8j=t�"�~d◻��A��Z9�� ��MX�����^j��&�~Q-��y�[��=7ev��z����j�c}v>G�\L��`��WN��!��ϒ2fp��G��G�����7���d��W�r�#q�&z�����>�r��g�#]����f|�,�z�����qbH^>Á�>+��f'U
nS6�O�^��{�-����ü+Ăg9�)�L�>�!+�I~�<��C,�0���#��@2�+B��E����e�fc��2~�nO�	Ud�[�m�,E��EKb�kp``�q�S�΋���XD;ux̂�p�������2�O$c��hOoF��~���k��Ʉ>�����[~`$�V��ύz�2�ⱕ��K��'q��4�B�T����[���MW�O�7��ge����O�UT�t�̌8�I��}��Z��,$�"u$Ʀ����q��:�f�-5��|]/��|x_���c;���VN�V8���XuOz���/?��1CS�g|�&���{��M���ᵡ�4�h�50�&�F�A�~ JFBIDg���w�OC�aF����J���B��2��,,�1x�&<��ƙp��c��!AQ��;�J<���W��z��&�.��s��| ���n�o�����w�W s��EA�
�Z	��1�\�{>"�_���=�Թ�+�.f�2��%���du���{o4]���m��z�%gPmp��xU�(u=�9������ZѠ��j�� ��(WI�z/��=(Hb���iJ�_�IL	m�ZK�l����A*��N3nKx�9�B)@�~/^�K�(9[��U��0�s��#$�G��5˶?}�G�HR�sx陡��a��:#����q��X�'�e"�5�d�OY^վC�8�I�}S�Sb2Q�?��fgs������=�4�2{�0�b�
� �φ�2��c� �q�0���{r�p��h���^���wB�*O���|+șڰ	i���	�S�{MF�w��|/���!4�Ύ�\���j�<���+>xi�.�X�gj�����[��+�Fۼ�M�=�p�.���ղ��+f����57{!'���׆c�:���~aj$C�O�K5���M�ԗ<���IJ�~�Ak%���	�� �=����R <"xL����,4�=��O��ل���ՎS��s�N�َ��?�N�΂�i�H��\l���� 4���ev���|�4~n����uLL��L�A͟/<��i�!�~v�|
n�0���k�d����\�l8�JY��T�+v�hJ����%L�)���9?�DMa�P�/�k%�8����A���h�6?[��(����+���|�M�ƯA�F@�劽���;lW`�m�?�#	k2�W�_��'��@4ձ"歇��$F��+2?6��AU���[����Ql��r|��M�Imq*�n��6՝����b¾�:�]�>�
�r7�o�˚�\��xsSR�V���K���c:@�N�~>LS?���N����7���wF��s���l�����6���.V��ɂ�� �S|B��2��Я�����7��Y7.��knK@}|3�ު�qBs�qr���H�5 R�1�S
c��KA��|ھ6%��;<�0�{�LԋZs2��1���0��B��E�2�GO�\��d��S��uR��U�
:n{?���L�?xB�s��th�[�}}�>%dQ2�ܮ|{#�(0�n' ;��6�Դ�!�5��49-�J'{ڗk������;J+p��Dô���
������:�c,M��i�y�ʈ�q�]=g�D&鄥{_�! �F��֊��=�� ��>_H�mS�l�2i+tk��e�V�6�A��T|������)>I@��,쪄�h��%�ٲ�����l�י,���٪��H�q���({*�ʠ�FIi�ȩc���"�D�ezшm��Tk��kAQ�`[=�V�q�y�I�]�^���|!�8�]�00@)��L�8�N��� &��1U��D��WܶCᄧ��!�s����^.���H�����{��هG���	!^\S����H�x�W!�<X_�9����!�_�$Җ�`�(�.X��i�Ю]]���h}D
�!��M�i.(��i<(a\�c#�B�iL\z�<a��<�	��ƸY�=��9(BL��4�aF*�C5�gh�Q���2^���Dp.�>Q���p�~�XG�̂���GFc^�N������Z��,^�e�i�-
pZF�9�6��g�|GN�a�Q��b�Z��MR�����c]T�
K^5��㹺�ޠ�PYP��������\m�th<�v��"��xV
ali-rRװ���8�RE\��'��"b39���ߴ��� �Q��j7��␪:c4Eq�������*LF�(�U:@\�b��j�kd-�A�����*�㴩 #�$�� ��泹�5�fI�k�)c�H�Y��^s)!?�x����!�L2t܅��r�m�31W��^��l:���a�l��B����Q�j�i�8r�F������?��o0���Y
�?��'3GqM�s�֋PSw�e��˨~2�r� 7G�!bϜ�"\r��^H����ʧ
f��3��	�����IC^�Vy\�jR�|�����Ǳ�b9���u���{� �?:5h��GMőX���v
J�%<x��N��c��$��H�ѫ�j��6.`>XW��I�֚�*��Z۰�n�h�⬎�ȤG]l�v��wÈ伟DDV3%��<^�۠�6wO���R݂Ӱ��C��QF����p3_�Т��i����*���W�0�a"h�>�1��_����ag]ㅼ���M�X���b���F�RO{} �lN���['�\��X��O��i��b�;X���0ߘ��ڴҋ�r2�:Ǿ�"�:>Z+��E"�g>���8G�on'�u,4�< �L�6"�H��c��@���h&�EQrc�NA�v��+���k���N_7v��,lדF�5q�vV���j�#��M����H�߇n���C؜��=c� F�j^�B�m��V�-C�����Ɇ^������!_����4�c��ީ�q2�t��ǄF�S�ƣ��XOc%�00�YMxѓ���$�b�I���x?ZW��T)bQ�Ŕ_���휝� ?��5]�]֣�9���+?�����_�O�,O֔����)|�y�j4+伝�1@�-_�1����9`�B��c�j�������"�`ф�X�4�5�H��
�H�S�C�?�W� -�+���'����r��o�?*���!��h�SUt]�w��_�喼��c!26z	��Oe4���sW��Ьh*���8@�����m��?O7�i������~~��x�B\��o����o�X
]�q�QJG*�+�7=N6V����D�t������#�(�:��a8x>��UC�e �ĞQ��zX ��~E6w0D�;{�Z�h���#�r �,+������y�[�XEQ����~Zk�VI'����D3��������$�$��-Q�Sz^�+/ ϛ{^F�[o��b@���^o��{�8�>v|D�J�4`�Ȅ�X�R������}��7�j����_0��y�.*��������͉�](cQĚR�,�����ȁ���C	@���y���;���1<P�	A�uR�� ;`�"�S�+*"'@Ŀ��j�c/��iW��@�c��#���n���cH�Pؓ|>�����##���H��4�X�aX=t��;�0.�M�k5�0L�=n'������L���f�p2������U(�m` ��%F���c��av��5�|�ަK�w��h���}��K�A�Q������^p��_��{������Sm0n���لE!s%@���2JcE�R��Y�]�,X��I�yH�(��<���V�r���|��H`�Q@*'_��?��5���3����ڑ�"���o�k�M�DF�D�)��d�t%�{f��iH�5s$o�`����`
NR��b��Va-6�R���I���tvq)Ң�[���+����<�_wo�����ڎ����F���ObPW^$�˪R��\�T*��hɈG�)�!!E@��F�0].obwvxq\�MO0���zM����"��f��º�}�Ůꋎ3���S��&�uv�=$q��	���>������'��=��,8�EV�Ӣ����"-���;
���
�� ��q'���@ �IQ� �9�&�J���Z呌�[���>�7&�h�V��%g`r�� �$%���;Fs�����i���"S���`X���z�+���p"j�|\ H(#5�!��w��o^���;d����m^�P���/J۷^a��P�r�*d.��g)rX�P�]N����#%���/�(��kw�6�5 -C��T)S4���!ΐ�6��O��z�`9��5G�6�/�5=z��#�)e�/�i>%�ܘ� ���Qcx���N�*`�u�]'ξ۷+� W�k���K�1�CBd����޺ґ<�Ӂ��Kg��S����Ȫ���y���3��8�p�����	SOw���i(�5)��ͬ���,M^+�*�w��c�U�;ę��U߹?e��atB��a�n�h<�5�ï۔��� 5���w�T�g��i(��M���v�cc6�k="Q��j�t�ef#KL]����������:�J0N����<P��O��|��r��jQ3B���Z�4�>����6=�4�����^j��h7�Qѕ�;q?��*44
~���/l���1��~�;�zU���|F��J�oL�΄�U~��yY�h�(Zk�;ٔ,x�^��c2��O��m��֫|w�caPk7��:Ü� ��<nw46�hXQ��sU����hRIbH�~@�]�ݿ�<C��@�HR�z�A�"e&��v��Q�wx����V�
咣f.�zCr��������U��N2K�h۵��W2U%Ǌ��˺Y�8G���nsi�Vڴ ���mJ�BĨ���2��7\@\��!֛�>Y6%]l*�EI_����V��1H�%q~��A�t���ä��v0�"8�ź���m�6(2���=z%��Қ���!��k/�wh<ꥨ�`5�wKK�R+����w��Ŋ�RlW�����[��- \�?����-��j�#�p�K&��I�C^�w->�>p���uU�8v56��KS.���`߼F,>0	
k"��sT���pz��8��g�n��	r�P�z�gv���t�,p�ǥ����X*�'+��k,@`k>DG	�W��k-Pde���U̝���jb�bڐ>�&�n�C@���+|�-X8li���)J��f��϶��M�2c�;��崾1�T^X[�n��~��G5NV�G�@o!�����O�0[��Q�b�=�v֕�G}����xX���̜ EzL��)F��麳�,a5y%/�;��Q�y�Z����/�oL�E��mA��ȡ����Y}iP�����WRNE�0�Ũ��u��"%�_�g,ŋ�B�jJ�7�"v}���^'�+�4 ܯ0C/m����ƻ���gԽ�
�@Ui]k����yg{��<��Y*>���s>e�7p�,��W��a휋]?J�U�RQ ��| xy��]zӵ��x��{�K���)=
�s�D��R7�t����+�Yـ` 6?람����?�zlAY,��7��T��;T�+/kE��'�g�=�������������z���.r���M�&{7�Y8�P�0f�UQ={˯s�c�n�tΜ�
�<Zp�dpx���+Pn-���eM��Mg:+�c�ik������|:�bM�G��iٔ;��6�^C�1�V��G9U"�� �	�H�zZr�ǯYa揦�K\qܬ�>]�h�t
hA�D��4�nQ��n��Z<=�46�j�G�2��u ��P 󝷝���{�B1;���7�Rn�ܲ[����6�5���c]U�w��具�S� 
۠J�\�3 ��Z�Y_l��T����a��	3�6U�bv�z�K�>�\A�"�fC��+��^
��������ʱZ�s�.�@5rH��_}�
�[ƻ)兮��.U5AZ������,�1-7��;OT�K��a;W��n$�+���F��x��c���*bD���1Ys\��☧����Y�߸��XE�O�G�y@��_���1�Эhwdl����*[fB"K� x��k��$?��;�ex9dH�N�L�<����F����Y�w�w�U2����F���T�x�8���b�lY���K�E�	��l��08lv�L���wrLyy���X�%B$���,�S��"ΆuK�|
I�2��ѩ�z0�r��xR?Tf�8|J�}��hH�z��q�������b�J���V��0���� ,�����g�ϭ!O��\i�%%邑PEAǅh��g�oa97,-{��
ʛ;�Q2���F,�U�ozԢ�d���f��8���:�{]S� �~8�?U�;�L`7X{>w���f$_����?�Gr:���KIڅ����T�S�Ĺ���i�C��=�Ǭ7�&�Э�)�*���ȅ��� �����R�K���x�J�M`7
{UHr���J�T'!ők��Om�'�yd�g��w�!�q0@/��!g���Y��[�˹,����;�22N66I�>��ۿ�n��&�L��9�9�"���r(9��b���d%��<��r����tvp�>A+�Du<�����˽z�h�G$!S[6*q��h��j�y��T�N��Zϖ�M�E�j"I�V3m\�}���&�hWy.��~�6ZQ��3о@+�x%���4�:&��x�?�2������29g�͒����d�Ge�3P��h'���!�����uϋ�E��z�bA�OG�	�j#im3���U��y]jV\$IFmZ�����q���Xȧ��~���c鲟M�hg�h0�p��lHW����S�X�PAL�	nM�aYIVŒ�����s�������u���ϸ�J��flmܠ�0��c��7)�j�/Kl�)'��B:JM@�͵�Q�����+rX׋��s�H��UUY@a�ۻ�_@o��ĵr��ך[wQ��nB�7�f�>@ʮ����p���)E��Vu��>�|��dP����l.u?�8��/j�n�y�=��߆ `Y7�{��
de�W�+E��3�%� ʗ��T�j�v��dF��9 ���-%�	��ơ�x�Ype`�8��g��V�Vr϶��gg�m����ê�]�����3inY�R ,��2�19��l�4l���ρ5��lva���U>�|ǆh����=�axL�������[����RGt��ދ�"�B��6���$~����t	h�݈��j����͍l!ز�����������EO�~�
�
L�I���d����a[]L�T��|�����/�N{ӊ>ރt/�7�;p����V�;4 $~£�yu���5g��\����B�?�e���|���20���D��!� ��e|$hE�`k����\��دX����dI7�8gٹe�^�(��ff
f=��j�H΄H��p���B��^Si^pN�m�fE�l��㢋��ϛ�����h��c��8,�h$�!Um#F�%^��C��ׁ=�+���}�&5U�ј���J��/��/��XJ���}�tPA�%�����H(λ��'��Pɉ�;6A�k��b����'����E�<#u,ʏtJ'�iC��j�6<���O&�睛�i~���a�h�?�v,@�)0��?Wml׉�)��Ͻe����]�UH�	{�Ŷg����fՅ�׳/���GyV�-l��:�_�:�����E��u�y;^`A��Śh��q��%�lEC��i'�u�Ă�<b��8�nRvjr�@�'����0.)~�,<�R��}�M�!�+O[d=�6��'�/:��5��B��'q� �5�>ܡ�[�0�����`�I猟�*��6�Te�2�����U4�C���OW��A�!5K"��9��%e�4�((1��m8�k�p��T-�ʹ,ߵ�UL�6`���$��D�9��~I�8����XS����žL8�z���;����3��oM�v8����F~l��\e2�H���7oM ���0��LN�>z;Rg;�7�$YZ.>%���f%�S�S��C�,3X�W|b}I���EQ 1�t�ytaA1�Q�����I�ƛc�����;�֣(<��W�#Ov���N>��$��������#�ĠQv�J�B
�75���@���H������6���Ѱ��8 @��k>	������^�QX�Ǥ��[;�ГJ�_���&>���hNl|	3���.Ȁ�#A�pJ[2$e(h,5�|E�E#�ɕ+͗�~Ð�j_&uwp�y���H�m���/c�P�(^���*#����R�А������	SI��7����,fζ���,F;���w���i��#)ݪ=/PP�}ۦ�c���b�+#��|�Rf�Q#qF0�z9�D�^�ԟr����iu"�	���3$�9��F�M�Ƽ��n;m�I{��r�È �ؔG�8���鳏��8F�69�yн�gO����,A���o� L�:p yo�2]e���P,q�%����͵�T���%7X�����-�s2ꭥ�A�v��?�7��Cc������u��bZ��q}�\V9
ܪ�#��:�!�2�A4U�;���0�wbo!�ab\a-4��hNR�'q��>����x<WDr>�q�zc���=0���Mj��?��?t�<����>�؏��{�C� P�Y�*���"D���P���;H��x�sF0$�r+6y���������5z�������5�����uUF�/���ŏ�8����^ț�n l����`��_��*$��k��s�l�7�|%��xy&��[gW]&�)��p�~���'��e$(���s���40���
U�^��0���A9��������Υ��_x��,�a.h%�l]YT�̝�a��s  ���S/�J��\�;7H􃑃Z`=_g��
��SH-
�<$�zl��X�E	<�������O��Y6��h䤖9����p��9Ȏxq�?��pҌO�%Z�`��dl�����л��9����"��.ZF�R*GF�{l/�0�:`F����S,F�+�M#�tl�S���vY�񜗻�ȵI��~M�M$:�|�`�˲jf��Ɔ��IB��9]ݎ�J7л�_@��줼J0n�aL!�d�y��N�L�.�BِLqD%s}���An��)�
M`�r;U��:�9���Yi�0�#��8�%�D������S>Q^�Cr�詌�3�XWI��#@����J]��W��j��h��d\�_lk�+��i�k�Q�%�����6Њ��n0��̢`d�砖���K;��P̈́K}�4%�:��>�w��w��=�A%�& ѼhI��V3�?Ĥ����˫m�B������V2���J%�@�<��_<m�Ql�Η��(�w���(�|��I�m�ϙ�1_ߙ���H���y�p{���M#��ؖ]�y��d��J,F䩧���/�+��gRX�9m�]Û���7�:����/�ͧ���[^_�ƢK:F!�0ep۫n�
v����o�e��$���r�-��?�4_�S�P�D7C�R�9�ٻ�(5yh���5@d�=�._�#��. ��.* Ϲ��Ś���3F��8M��a!	v���Ҁ_�s��L�.����R��-�&�ASUT�f�#��,�I%��_�����[�dI2�B�%j��|0�Q$�>���{��E�����*ܣ1�KD�#^�����GW%n׳
Kq�U���S�}��Kϸ��p��U�����
��=J�c��������u5���=�!kO�iA�	��=3��t��\�$���
3�⁮�`0�i���s�`$+��A!|�b3��7rޒ�=��9SM�Q(�����R��h[�
%��3�}��`^pF��ck�~t%Z�(��?�4�L���ej e�06�΅�����c�����tgj�2)x�3ޡv�a,H 1xb
����%!����+�uu,
$oBg�
l��֋}�;d赝�ő�T�o�n���Z>�g3�ެ!1�A4��kC�b�v����ܡȥc���]�������ڰ�p���[SW<�t���v-����Z�|�կ:(��<O4�h5\�"�/c*[��c��reBϢ\��J�P���O��"p4�I��m����P�,0s���>�ѥj��	<����+���}E�����
l�4�]���>�����Y���t���ɮ�&��Z��ө�oR:��ye�i[
����c�����陈,.���(���ǿ��B�l��W��>����>\��H&nhD�'z��6�O��Fq�B(^l��qR	��b.�U")�e��{8�צ�k���is��Ѝ�B���&������¼G��*a"�F,�*Ćp.�t�D�M�%ƃ�OS� �=:h�khd��e�D��'������eb#�Szeq;�h��_gY ��;�,��잖��%=9��Ӻ$G���d/����8H�6�4:�:I����].!%�=�6��F��`$#��s�`�z�f���˺%��A���{f�C@3G�cnNE臊ǜ��9@�*�y,��tB���T���S-��'���IU��T,d�W)4܈���l�(�[Q�Tî\u�"��>��;K�MM�Hs��2c\7M�4k5������ɟ��'�G��5;-ԉ���s��>����Ǟ�kJ�~�������IϾ0ŀM��c	����2iζ6����O�a���va*��EZ�y�s��t�6v�����>^����L���-��B�o�ԓ�	D�BPѬ�ϑ�0�Ꞧ���{������
�ne���Y���v��?}mܐv;� k�&���@�54�1�`��&��2��JvP�|1��A<jg�./�O� K�C�����~ZFC9,ߍt�I���!Q�F�t�o��$��w�.�K��/��:T���5T�&L�@���T�^�`2L��8�dתE<$�g��%�����~cX0-����r�^	���;��y�<���/�p�E�#�J�ѣ�%����Ȧ��;O�N�5=���t+΄�U7ـ�p�E�\e���Ek�]Q���1%It���v3��&]˰�v��V9�y[���k��a ����:Q�~Y��j�6X,ꏚ�7'jT���k7M���!�~�ߝd����iڜ$<@v��4&���락΁[3��i!������^�5l{��,��[J�AH��y\3�}����LoZٌT�}�=�t�U.��k�OѶ$������[#(���F B��"�y�j$l����Н�#���g�qNʤ�H;����1њ&�N@�d/�gΝ����Ǐ��sOn��>��R�a;�^*�/�p�D����,j��EUlC�\�{����C
�b��F�k �r^3V��?��[@'��f�;�X�֊Y�V�� :Y�D��9��3P�6��կ9�>̽A����:���k�l��j���`��p�s��}��E�%��H���\>�B�O`[�^�j��O�5�A�,I'�s� �1�O���}�1��8Et�iN^K��b�>�]��$����'���e�I�$:%ܟ� ��d��D�����V_�fةQ}'^)�*��?���[xѯ�]P��$�H�"��+�M:�F��N���Pv2���7��4L���[[[�����tرS����r����HP�o�GkC��V��i^�J�k;�(���1�*��7M$/8�*a"�Y8}�yФ�F��%���0�p��B{��z��l]��� �z�*���Tu�/�6�ly�-�j
D��/~�*�d�0���k���h�Lȇ��.bڞY����?��:�/Z��j��Ȭ�P��(��3ߴm�g�؊�,*���R��3-�U��k_�n�ij�m�>��G�KQ�!6�X��A���G/,���x���4P��>�7�Jè\B�;�5Ч��}��93Zd�C�<X��'�oe�"�+GY�jF�o��k&�I#�-uL�_�K,'?�!<4Ps��;Ǝ��VQ;ȗ$��6k�
~���� up�_s�����=(ƷG$?��h{G�y�d��x�x���K%�	%Oe[@h�AT��>��JaI'�4�FR���p� ڬ���j�2o�&n�^���{I��o�=�}�.��qq*q>�l��J��8Q�~ x�|���������Rdp򵠄�nQD܈���:���� w"���Y�o4#�E5x���U�0�4�\���S ��jC�7�2E$���S-t|�eQN¥癉��zG�����%�0�|á��asl�U	W{��&� �����M���6��PC��+��wж��C8#���m�-n��\���:E�1��gO��(C��7E��i^6�OE��
q��.�s+?t�
5Q�qbu�I���}���Ɯ^��n�"�+N�w?��y��y>���9Sϯ��������M�S�v�r/xZ~�:��2�D�֛�="罁["I2��x��21�/�
�4 �kj�)�ʰ�ū�O-��镱N�dJ1,��B�s��v�DH?w!	��b�9�(��r�"�7} �k���;���Ҫ	Pr�C��W��Y�/9�g��>/����;�`�w(/��~��xx�����H��Ec�㤞��O��5�kZ��[���{cҕK���31�@��Y��(���s�]@���h 2ON�p�90�ơ�x����~A�GI�ȼΫ�܅dc"Bm�hE���.��� ���=�TR���v��ğQ-!��@B�)��;3l��o��g��*��G@�l��GO����v@�΢�Xv�(왊5)����˷��w�q9ݹ�:C8H�y��A�
j�K�M>�L��^�@=��D��u����Bl�)}�����{U�&׳�-6�6i,��[���Hи��!S^�M���٨��_|ޭH	fs�-�+�	�
9na���xX.�7E�e���y����G�� ���W�v�+�f
�����[��&�@�����P�	���s�R��9uF�����'m�?�pgMF�|ӟ^��.�{��b���(ˌ������ 'w�Ԯ+�h�V���UR�;�l���r������:"\�nQ��*M���GM���n�n�dniy@^F2ɃҰ�U��!Nt���WS�>߻H@1
@���5T�c.�W^pӦt\����8��u�(B�,ۆZ�u'��!5���w?�,�"���x��|k�@��ȟ�"������7��"�5Z@��h0��]��"\lhoԅl���ul%1}�[��1��^�ئ����`ȯ�u��C��6�dY���==��08�����|#ׂr�H׻�-W� ʆ�/:V�ք�g�om�2}�t�ߔq���U��@Y��)���CiO`�h�ߢ�uP"\�ǰk��3Q��*O�]����֞�hT�"��ʀ̳صRO~K����Z`����';�d�D�RV*tl��C7����p�v,�r�7SGFI��-�������"U���c2|�c5g�5C�7�JW���q)O8ѻ�`X5��������&뫣�G�W�8`2F�F�G���)H�����w7>?����rU���$a�.�^�]d6�����I�?�
�4�Y�����4�2�L��*�"Y�`Ü����h�TdhSm��O��,h��8�� -���n�i��4P�r������r��^���zÝ��cD��ܓ�t�}�2z�������2WZ�E��X�z����4��.}��=�t��R /+`���8��Y�ϐ������b�o��i���ޑ���K�f�s�ux �m��d���l{q�e��#E�~3���8�މZ+�J0hz�S�9~��i�f7���O�H��0[v���"I[|�YV"��s<@I��i�)��.�:�������E�ޯ+�������niUÄ�Fh��d����y�@b`$Ϝy}�N���?�U`?���6�뉪Fq.��!�eBug^�]L+��0\���ryT�+>��&^�.a:8��;��84d䍐�t����r�?�ݴ�<(�z�@��%,��*����F������U��&W����a}�D�0l��Wr���k�{��6�|��&�|��H�X Lq­B2.oI8L�D�]��7�4���e����g����]��a��.NԸEzr�5�/{�ܑ��!���j�9n�QX q��k��,�%�;� �?+�n=���5�b��FvG��Qĵ�$i ���q�_��\�f��'='���h�o玄֙'$d�{:{{��FhYG����-�>O�q(��s+C{�-�i-]J6]o�~��nv����CU�}�����>�z=��|�:���+�+F�Q��MT��h`ytC����>qW���î��L%��/�:��0��K����N(�9�Pp�WS��AҐ71f�����$��{Λ#����u�17`�Dr���|�v��
�#ER�
x3p�q�w�mo�0|$r�!��qaPG_Z�w^h��\��Z�W�(�Lx�������d�ƻc8~P3��4�Z�G��S������2�݁��/�k�6x��+�<�s��Z�^ǫ�3K���?*��m&/d2�9��T9�AG����E*���;�}ɕ�� �S��p�Ue�m��4���&C�h�Z&)��\I�\���n	�^�Ka$)�\��=!:���d�@���`���A�����7 �ݕ��2��	�k���rQu�u2m¯=F��U��sr�Mu-���Gj��IqJ>pQ��?�`�*�6��$�-��u��Ͻ�ݥC��{���X;���T�n����z�8��#mv]�b�`�����~��Ŭƿ��I��%!c�@G�/��t]M���r�C/ؙ��[��F R$�w�!h,��u?
���ۗO�@�g{l	�Rb����{*�{��Ͷ��+��"���7ƾ�W���Ѣ�!$�̼���wj!�ذLamWe#��-�|_��Y+���u��L��e%�ȂY��5�
�/IZJ�x�V�0�5�?�G\�[V8~⅌�dǈH}5M��o����?����Ϻ#|N����IMvj��gГi�m,��6(_�7�P�F��A)�IfD3�sn$沃�>$;.���B�Z��UƳ��y^ÄN����;@���|�h�ϐmGs1�0!�3�7C}6�E<���c��n{�Ov4?h�<��a3���x�|.��#:{���Zxv	&QA��i4�'�\#��XJƬ�a��-�
��$2qO��m������ƹ��������nK͙R�a�uQ���G�O��pê��Ά�0�"|�@���ǉ��ڄ�ʥˀ�Zu�#���a]����������?�Be���W�@�݂���~C`�js�ȷYZ�@��j�|�Z���!-'19��3�DW��J�F]yҰ̜u��PG���� c�}�\W"8+z�X��,�!-}����r25i�U]����X3-Iٙ��i��1N�9��vN��-�>z:Q����e��#)�S���ep�+qG�x#Gh�ĝD\�ٲ��L��b�im�"D���b
;�)����Ӿ��p�¼�_�q��������Ke�H(^�Cf�smQ���Ǣ
,������k=��Ǌ�3�e3�7Q#8��k����T���	��.$��Щ3)�����F��~gP�C����#cʶ2v���Pz�ⶐΗY�#�.�0ˈB��\5��[ݼN�^�	�����6��L�wE%JO��#j�������d��8/�u��B��ims�NvIa�Ӷ+�;(�cToM�T���hq́tu�f���V��!���ixC(��<��Z_c/��][�<��pEs����2����j��pl�]=������ G�W��;�W�1�!���N��(���;�U �.,^s���gt�\iڝ��2�?k�<?�f�37����v�x���rŞ��ɡ龍�j8�G�?hB]W������D�^@ץ�8�o!.�s#�]]��ئ��L"��_�Ѡ���3��P�}��z�)_g^#���Ѡ����(-)wC$KN3\0����/��Q��4�{Z�n'���\{/M���e;	�63)��tW���y�P�D�A�h��4���0L���%^l��5d��Ta-�&Z~J�	:��\�9Ä�fkb���OG��vG���k^�L9�5�F�J������EoJ�d��̉�u�ޭv�P��>i����.=2d��Y��}�0aF�a�BLzzf���e[]�Zt"QI`��.E���I�����������-�u��p�Ĺ�E�!1S18\�w��6�V�n�j�4�]~
G���S��5���f��J@����J�E�Z6�y���o�b�y8�'E�)1�&_�'�6ȹ8�-�Ȼ��Ap�S�;��Ebh˨����]z���¤�z������8� oW��4Ie2*99g1\<���o�Z+��ϩ��>ݷ���LT"f�>޽z��I��〾��Wc�bP��0�6`9������t%�6��|#�n&pN����I����lz�j���1ʍ^|&�g'Aí_��3����%�"��P^�.�ac�ȑs�`a�/{����J�Op��|K&���]����N����Lw�a�)��DBl��	�y:ؒ&���i,����d���G�#��z�n�#@�J�i����Dǖe��d����A{��j\6��{
i��Sb̔r���dß����/��4 3G�Jo�A!Ͷ���Wq"'$�4�en�/�"ϖ�	)|�C|Y�N��������,�����m�@��}wT�M�#�xJh�>m��uv#�D.h!0��1\�ҝ��ZI�/�6�����v���1�>ɜnxiy�>��e$J�pi�֑��J����}�ᖌ���x��*�����KU��w������v���k@�Zt:���U_�q"~v4�>��?ڼ�4�PЧ���>�wzk���?8(�o[�}��Hm�p��!f>��+�x��bAIW-����B$쫤5;�'X5��`+,zO(���]��; #��Eԧ�9\�� ���u�$��U��q�΢��Ѝ53������^�K�HH�RT�J�O��-D�m(��-�%��닁9:��.6i���o&�i�x�Z�3
9U�&��<|�:6�s��SQI�>�����]6'� ��6+3	�@ۊz
���r�3; �?3��U���.c�V|(xt|��v�|M�H�G9^�5�tۣ�%���3�����Fh���R�,���s6�z~�����)c��G�ۦ߶MC3��	;ҧ{��4kK��&�	f)�w�����>4����V:�L#=�mL%�:ٖh�X����܂��q�h�+��ݦ���V�O�5 �N��+���x+,��=Yep���vy�%���T�� �*��;����bvJ�����]��Ȁ��q.:��lb�H����Gx�&qQ�d]M�^�d���[]�S����_�M�eX(_��3M�xd��o	������Y��A��s#�q"�T����4Z��V����fl�c?�ź"�K��E����䓑3EA"�d�SWX�lz�0m�t��NO=�-`<g�Q��B���f����=]�LI�#��΀�X��r�+��сb�~�����\��"}A�&3)T�v�${$EHk��TGaPm��L3�.��gK)X�Tc0r��ˣ>瓄�?Y"�Ϣ�~�q��P5{f�u��[������+Wu�*��c�=2U^�kv	cq�K�0Jރ��N��G�����+����ٶ��7]f��0���E"�B�"��.7Q}�`ӓz�����n|�����o\�h؄IW>e#�Ɔ8r1�&MXۃ(q���-�z��<w/�±��QදYg�!���QsZ�U}%,0*�V�yP��GCP�1���~�m�T��Oܑ�7T�w27��/LM����2�����m�ϕ��2��f#�h��枨�s�{t]�{%��0ܝT/�12�Ǝ��;"�-$mfVh��q<	���>!�S�q���NG���(�bK�I�jz*��ąG��U�y0F9��K�SP	������9��lhP����D�o%��؉�~���4|�k��<�.�3B�~�a̺n��U��aj�"�¿�)��q*�-7��I�~r�U��mKXk\��맨����\��p�$���)��O��>X[ ��G|���1�����?��#�ʮ�h�%�wLР��^{^���xlc�N7x�u���ڃ��U!%�F���%4��ԛq�.��A��D�-d7G�.�L]���:|?Rڐ:�-і�+ۖ2�S�LF,�gG3��p��n�'�","��A�7�2ՎT�i������5}��o��3 ����G�QT �i͒!�Q4@�x��6�\��]_MU�]۰��_ɽ��8[�a��f孮E��΅�����y�w���n���n%+�������f�YI7��xgS$8D�,zp�d��2�B���UtQ�K�ϠQm7=����q���K�6C©�b�Hɨ���˟�e�@Q���R5N�拯p��F�,G_�}������a{��r� J�1(��ܾ�L,�9��9V7h�ߵ;�]��֙�!B�̘?<8a�^s��G햧~0N�ɢ��,i��0�����"�[�k0s�GB�SS0DF�:����Ľ�=��_j��址���P#O�W�_��7H��f�K���R�0����\s8O�L|w.�"��3�c�8%mkU�5�`ȉs9k������2v����@Bǉ���a�8���>pI�D7xy���h�@�;�
�l=G�C�QT�{�z�Q5���84;z}��p��|H������3Js�Io�09�����z~Od��k&$�α��yc�C,��CM&�c+�����CsA�c� ���½���y_�R�4������CC���"�C������+|[�|��z4�n%ԯ����_�DOHC6��|HmU��k&%I�@j��X������!2����g�7�#۰���}�̐�W K�����p"�Gِ�m����@����*���v7���?�z+I�A�'�;J�5�暶؂�!��gll~���C!^7m�_��K�8���G*��gMP�y��Q$*���9�u�����D[�-�l��*rPzv���7H��a,?�q-��С���C��h8��p��ю�ϪZ�?�aZ6���yQ~%���N���:�/XՉ@���qH"EHɆxa��j۵�H'�o��aa��������~�]F8f��(9��f�K��e2і9�#����3��Ԅ�3 o�S��k�`�vS�9��s���nK��z�9}� �6y�*����UsY}��3}�v��ݑ�����6��P��'�zG�֤��u�
e�1��XΑy �O�HWd?��U0�V�D)����s]��������|�k�0^ F���D' �_���}P|i�7Iw�n왺'U+���I����b��+2Z�c�"�#��0'�򎰐-�idS��/�I��V�"Pk��X�-�Mz�Y�w#l=�+�	��dU<ՙ����'Ca��ӝ[�L��W}��l7\��A�d {��}��Q8b/�z�ߙ��]��ƑF��a�-��G$��@��yb�"J�o`����fC3jJ�����¹"�.6<�.y�X��~�)͋G6��jF ��
�-4�5T�Un��?z��@����8�V�dju0&H��[P����mIh�}Rv��]�mh��s�(\�6��aUye!�G���1bԋ:s[�P}�������Ѷ��e�͂�r�m���:��u*ޣ��9%S2�heٶs��C�`B{�N���t`��Kf�r,D#�N����x]��dX�KH��U��� Ҋ3�:��8e�g����j�jSd�t�d�w#C��䧑ے�)s�|��5�1� �͢2�D�Y�?�г�wf�f&l�pΑp�Uz��AvLK�vg�֪/N���2e����Qu&9�2�������39�H��l�%{|���V�(Z]��7�����?��������
53�� n��4%KF��h�~>.��(���盵�䢟g-$�����dj�_*�����t[���G�s���	���%�"��4+��F�������f7�Z�A���(nc�A�<F�E�Qv[��$������cP�����J=�$�z�K=/��h,�l��X���J6+8�������ƨ9rGM�υʭv�g���7>B����!h���Eus�M�D��i<&R������+r�;E�� �ak���(U�uш� a�K=����
�nݓ�$�֗��x��q�	�	J����vO������:�d�;�k�5��]��Gq��Ę����Ejǘe����!Zk~�g�:>��]A3)��f���W��f5�����
�����O��աP`( :7q��߻�b{/Q�[z�x	�L����K��0�� c�o�8]ί��io��7�y�"����Y_K�%5q�o����Gdn��hv��G��}�0>��D��v4-��fdY��e$�-�����SGe����4�����iў�	�G|���>+I�gZ�&�]]��a��o��z֮�O��v�j`NyE�	\�l70�F�۹��|ս�Y�ۨ������������6�b��sV�<����{���N��u�D�xY��\���R'�繛F��d�L���AZj~c,)u{���d�ݶ���zb�H�7��z�uMbC4�c{sӐ���G���İ����d���I�n]n��(�ˮ�X������67Uׯ!�Y(���n����6��+f�����*>���T5ڍ�b�z��1�+ˍ^���r��'��L V�cEPv�L�6�:��4�	ƛ���r�6yQ�N@�t��|��$%�>�1F����D:�j�q���v����� ������'C�vw9�>ѱ�%��>D�Pt�4[K=~��lxàMi�|_��3����VR\iT*��V����(qǑ��E�;?6{0��#���2�1քvb�U�����D�C�P��'�#�ڟO?����z��Z7� /8�4�a��J����uL��3_#56�����;
z��^�{6ѥ��2�ޓ������4טhCD�'���lE4�<
F&eW
o���J����Z��vo$�l<E)7��l��y�RUl��.�Y�����6�u��+�*\���!]�)��
x�E�]Ay}�O�c��_{$у���t��hl%ӵ���A	����*�A�#J���T9����R*Fx�0�$N����1�"��B$���u�&*	mE��55��	ӌ�pڨ�%ᶠ����~����6�0���\�ٛ[,I�z��W��~���=��/�������KX4�0S����#���sUʌ���'�zBы�����f����}�Qe��4У#�����!Zm����M���=����������-T�ñ�;(��ɝ?Y����1���V��+6�m��F�`�C�E��$��A�C��Д`�wz�"}s�����<I	�_���7O��)�����uOn��-;%1Pl^���Ж��@jrݵڦ�1N��1T�V2�ac�	J3C���� `L����\�|z�`4��̅N(;C^d��������JT�	�/l�C���q�V��^"����f�ݖ��^j�5Z�gGv�!_�;W9��H~��]�xe������"��V�&5Z��ݩ�&�Ys��kA<�.a��*� s��(I��v�(���4t���)!��� ��'�+��^cc<�a��Ix�	�������덋�?����R:p--��T��!�z�B�)"�W5"T\�F]�ŕ�;A ���l��
W��T%��A1֠�z2�j=�v�'�USաiE�P��f� ���&cf�W�&��p�!j^��Pz�M����-Q~�d����*�
φ��yzOouo�|ղ1�g�A]�z��������Ո�鎸.����ﻍq�s�6�$��NoʛG~DH/�G��Ě+f5���m��W�]1Z��g��B�ɥ$E
���k���/[������>܎��w�JZ޻��d���!:��r�\4C&���'Ei��Ԕlи�َ�g|"���ŏ�KxcfQ�M�_��/B��dSۤ+��D��1��8�G�46�%�jz�D�	�Z>���j[%�g��@�7p�9�����ó� �y]A2���SR2C���h8��'ʵ<���'�[%ݐ�\aE�`�k���M���m^�j3��G\�G����V,��$
�7��.G�O�9��\����
�g�F�g���v��3�Ǉ���'�FO	�d��Q��7=n� %��� ��L��zTE(����˔kM�ւ��|/Ƹ�O�*�#��`mϙ$:�0/ekQ`��%*�@ZY�SL]��L�f�M,O)�Ϣ�5aҜ�ꡗW�7*��r,r�4jT�ɻǪ~�V�qj���;�e!�9c���I��߻,�[5a@E��� '/���UH�Y2�(����ְ=GO�Ü�����̥�	�e�>�<�m�Q�U�	���sڰkP�o�8X����<�[1���~#`�������[r����<�#��m�WxJ.[m�s������ԅ��XF ��ԉ��+�J�7��e}hz���Y����tV3�|U����Ǳ$#U����������Pʁ1�-�.Nƺ"�㜪�>�C�)���ZJ�l��n.�P�B ����\�-�'�~ƥ��٠-�}g�r�����;�,��=���?�S�)C�p�=�zw��|����n)������b	c��'�֑}M�ix�����V�F!�Y�:i��G�L˶�d<T�mu�	K���B9S�<��$}}�*Fm�!g��d"E,���Z3����g���b��P���pN4��~x\��C��~���@d�@��z�[��6�Wn��wf��I�߾�X)�Oۗ�����=v��Z�-�P�b$�|cr�萞U��}�(^�מ\q|�w�~V��W6�tz�Lo#�f/���!�"]9����2_F6:�/<�u�N��Żن�c>K����tV|�a,;��+�sj����@�@.�r��s�+�5�q����T�|�{��8�T|,�&��\l��bD3��U�z/<Ƨm�7(��WX���f��6h��A=Ӥ=KJ�����.�̪ո��=��p�m���	y�wN[��_������i�t��/�!��"w'����v<���l���5����O�F��s���-�G��TH�5��5(�KʪD�8�8��+z�x��OtV��Sj6?*�Ra�!��?0�
��ьy�S��<i�P��i�M����43-�S�5 �6�ݡɄ�bq~#
�ѴD�\s�c����B��\���2�~�*�˧�|Ƥj�*�M��8�C8�b>9r�s	J���p���Ĕ�<q=3�`Y@-�`���2��B:pYG}K�0o8���8MjH`��/k�x��</�I"��#��s
�<,l�� =% �zD�X��_��i���T�9�1���˩��,���#N�Yi�F,vL{���9����}{�e���k���	9s)b�+�[_bd8?Hs�4�DΎ���@���s�q|�9�tRʭS��\� t�&��.��T�y�B7#}� mW�ݮ����H���U=K�Ϙ�S�i�}���4�A��"x�d����{��ݠ�1M`�s�A�U,B��^A����KƧ�J��2�?���i����
8~ћ���&��E�]��.�3l�����Ɲ�~��x�(�̏	��k�Y�0F��L�zS��rmQχV(�~����׾s->*��WC�5�6LM[vVp��M��kT���o�S]��PB��+�d�"�w��!��pu#��iZ���ͮ����]_@-�xL���=b�I�y�0DXT�+_�Zp�[�u�W�U�bR�9��Xa*<��}���j��mc?��i;3���)��#2��QnI^6�w&�z5��5f6}GZ�Ob�쟗@m��
lm��L{�1��}�aL��Y:Jh.;�+}�E]�!��^�[Bt�V�>]�t?U]~�#$[(k���4��%��~��L�w�U����}/i:l��*�MgJ��, �oܮİ�~i��1[$����^�SE��ܼ�;]�@�3����������Nv��p�@�?���=Y�C���ՙps&�|K8���yGp>0�c�a�ێ���U��"���q�.h�y������J���������t%������ܽCR1��,��b9{���ܤU�0�RJOhF栧2��E��p�b���B�\0'���������m��˗o�G��Ό�!����`�o�L+�2N%&���W�Ws?�+6܋u��X�GZ'ڟ9](�ğp�����1c��8f�B}?X�2��T�%�K�2�lQ�L{���Oe�Į��U�0*�����"�+QDUТ0��}J��E�7�%'��f,� �z%-�l^��z�u�䃻��W�ثUF{y?�5וtG4>�{V"a�擎1��t��v/kH�؂+{lF���W��r���sZ�xE�j�:�o0:҃��"jm%M���Ș��菡���G��j,�n9<~Jv�
�sm�A��#'2h*�b��L���"|C��[��E7�y�C#_ ��f��~�6lB�}+��m�����3bm.y��-��%җ>9�J,"�)�[��4o5�Y�̊�Rm�hj)���
�0�紨}�m��J�n���ň�(��I�m�.�Zr��8HjEgТS�y��Ct�k��m�R�y<S=�,�${u��&�\G8��j�R���DS_DZS�`�y.}#���զ�խ
W��<K){���
^�VE=&ӛ�:蚜�'��N�&z1md�.�҄�8P��7
i���{�`0un�I���:>�v�jw��ۈ���a��O�(�@�E��'�:���2k$o�GQ��Eu@�ـ��, p�Im.�3�w�Wجx�u�\�d�~ͅb��!1�������6p�%�u~�n�?�į����,KvP5ʭ��Kw�'O�n�������,�`yc���nۑ��B;jt$Un��d ����|��)G��'b��J�M1���m<��cw�ݤ!�cY48���i�ӕ":F�H��ID���M�՘ ����[����m&ł�UNK@T�T��IU2 s�n%�B.z`4��d'��a.��I�����ޯni���x� -�1�P�VF�O��'[NWgą���^U+��1�Æ0�	��,q�|�~���~��uF�yO���i5�W���E�(���k!>�S�X��m�2gJ�,�N�����~�M��r�s�;��K'���-۝֠��|evȜ�A��V'oD�Ÿ���8��� ��!���&�"<��-,2��?�]�]6�}�z�y�HF��;�� ˿U��)��B��Ik�i-e|���Z��s���k28���%:�ո�
ߞ�����r`X�~�ij��rs�#FO��i=\T��9��]�i.Z 4yC6e�_��K���Ya�#��&犼+�Z�.����m��"�scO5�]}Z@��;)�5{�1�`��/����9�H�>��j4k�Bw*𲸧�I�p_t����1�ڦQ4X���6_M��|���6���[f$�kn���Գ���ؤd�2��y�q��|�S���/��G���o��+���zJQ���%SV>B�A���:���H�u�a7�#�!a��a���v��a�_�\"t������Q��sm7T��.�<$�ǸzE����thO�Il�P/m��hè�ibku�8�����˖5'~���@}'5S����>�)�����wi����V��D1���?5��x��1Ҕ�?���`��5H_���|܊�X�EBoֳ͛�1餼�	�����G�����d|�]Q篃UnmE����d��A����AΚ��\���3n �ʷ(�E`�A�V�S`)���fݷc+v���(�U6�\�slix���4��Y,�/~�*b�cG+�����;��n����@{�T� �-����wR��Ǎe������c���#ߩ�F��k*P}%�� ��ן��P3�K�ZـP�yr�h�٪�����?��1��S�{T }���ibt:=�v^^u��Ŧ	\��|�
q��t���j6_���c'*���k�����F�_�� �уr�z L��g�q��q&
��5� q�Q˜����Q�8X��xUЩ�]M����sUո���tK�+|��G|����� �`uU@ه\�4�=�+�Q����^���-LJ~,���"����˻a[��,b����=�������0s	�{9�==̼���#�nV�3���׬�(V2 �i�P����;���͟ф4�[U4�RJ���O�����%Vs��?oG�����R; ��bz����N <��æ�l�Ӆ�EI��W�h�28gY��K+�M;Wxs�Z��.-��kN�%�I�F�PT��R_w�Ob�Fpoew�#}7[�Mh'[^��72ȗ@��]O��������Q��o�3�ዖ:������Kq��>R*Tꈝ{�֕�7T�hɜ�';��1fW���ѷ�{�@��o�C� ~�m�^u)B�_�-�L���r�͡��_a*��k4�..�d|�I}�.��%(t��p�"Q��fkl�����n}6}�ee�������A1&��/Z>��f�!��Y�"`���f�ǥ s:������`O�'*�\i���ZKWM��{0�mM��q�M7�I��!L9d�����n'O� T�0g�?�V�4��2S���F/�ظ,*��S�&L]x������q�ٶ��k��Iͯ@�s�h��$"k!W�s�sT�@.;{ m�������̾�p���9��?k��U��Wt*Sh�{��/���U�:NG���u���*m)��Y��)=Ꮍ}���d�S{늸���P���cz{�����͝@��������������#�\�~bR�5���} �����>�����,��`x3����H�&���"�)�ļq�&Ix�V��w9{2?ҝw�?�r��U�/��=�
����6��٩K�d������Q��8q.��[�o)z���)�W����X�/�ō�Y�M��`�qկK���X�b0q{wt	}�(z��2���}@��U�h��R
�JsB��o��y첚D7��)Lv9��y�BC6������m�Ѩ������ϛ�|J�x,����n�7����/�-�4k�6}t���CD�	u�=_��{�ֹ��ey1i��)$�%���"k�z�綷8L���H)�9�ҦF��0��	�%-3_cN ?$��L����n�9E�W��hu)�U�ܴ��.ȁp"�Lo;A�]=/��ݬF��6�q˳�n�t�r��z(_�QC��Z��9YP�*��if������x�,VBSZ���<з�`���%.��M_�s�^��	��T�,�|��<@��w�/��i�5����{�:T�`S�(gjU�C..�A�0lA���s����sD�@�j7�]�J*vA,�Ā1��I�˚�g�}4s<Pv�Y���ܠ�����哕I�[A�>�
�U��@VҼo�N(h�5-:��o�P���}��]5�@�[jo��f9�M��]���Tڸí^~}zw�{F��EKߍ���n� �7 �����+�l��-�PZ���k��Җ�i	>�P����h�[n,����L���*s�%�r-q	c����?��ۋ�� ܶSLa�_r�� �M�.hp��ġ:6��wF �!.���U�����yB͇0�Dk<��}�H}�@�|�j����rQu��m�̪�o��)����v�	�6�8$$|O��ɷ�Z,���� 2�"�l��c9Ƀ)����F%�{�i�ө�ȸK7"�i/���|9Ș��f��z�#��b��4�WUD�����^�	���,/����FpI�,�[�_�Z3��6ͬ\`m2�w��00�x���zK�2�K����ZR�@=-$�b���3R;;%�E�G<t��Ё��%5$�����x_9�aD��+?��=c�Z��f�7��=Ǭkh�(ڞچ�ʎ�S�:ܞ�k�aw`9ee�V`M:,"�D �'|��c�~��*�&����T�׍ဃ6�۩Rc.�oylUnI֌��d��)�'�s�N͑@x�n�Y�D���lH��[B�AFY�؜ˎ7��Wg�׾~����Kѧ�5����kC<O�U:������y�Z*�"� L�\tc�4m%�����Q\�����t_��Oto��� l�}�[Q+p�pZ�3
��lXQ~7�����K#̖a���Hp�1~��O�w���-��C�5��k�������.����4u��=ŀj�n;����Mg�ګ����~72�A�F9�ɶtpN<�UlZ��օ;�L�6��t��C7>�i��ͭ�nxH�ȑ����~<P�t��j�R�gI�`!'�� 4;�N��۰
�A�rB�������/vX\v�%�'�nܢ��!Ҵ��t���9��?��3�,�]R*]�gA������1��)��*_DhƸ�ºT)=�'U��*�4o��a��:�����lUU]�ω�:��>k�61�Z{orKзS���	i�r��� p�k�ܲ$Ư�F�.�@-�1_H�
̝�j��E�`�N��	aw&�|�T��?alF�?�e���1\<�>g7ܖ��������.�c�D�T,�:����Cy�.Ū�hH��zג�� � �]UR��J�����"�!�a��r�yw�ࠎ���v�C��ٕ��%����mv���tU��R8�%[��=4�$8?y���=֓�<ʲ�J@�	�'��\3�y4�7+�=����2�w����?SrQ�����^AU׀����a��qC��K�Q9�ø�,Xz�9�[w,�^���4�V�`Hd�e!�~f�������z��{MiS���K�Fc���DʢEU�t%N	����y�sP&��Ҕ6���.8𻆄�+���S]f�0cNUv�9�Rctb��aL����>�ݭ̈s�l�T H�?�7�RO�M�֚���|�;�8
�RA�*c��B�y��0���6̓�=&����(�mi-�0Ԏ��3���E8h��.��u��@�n������.�W���1�\Q��ssu��C~��x�1j�zD1�,��-I�~�$�k#_�L��X�|�3��g|V�W�N��_Rz��Υ�M�L2�&i-�eΧ�X��b�#�N�	X�aM��T��9�V���8"X��9�-�-N7�6ls<3��=�����O��`�o �!HcL�P��	j��;#'y���4h}B�c3�^��t0^�a����g��}��\�x�A��M���/�L�oN���_�Liv�y���jZ�LL�����{�G�b���L�V�nKǿ�������	�v��2[ �Q��7�����΢�ك��5%��%�^��� ђ�o*�;�>�ʶtn�Q5��>?L�� S;?����9K6��Z~��m�����u��@&+��T�������q�\)�g:b��G���I����j@)�{$���rĠ��kr��?����y� Y�s�C1o�Z3܉(&|͍��5"J׮>A�4[t�25��~6����ނ���GK�����-�D�7���,�[���*�{w������]t���q8�&֚�I��U�J�T�0֊n��6[r�[�Q%����V�|%&���2z�`�^�2�R�����:�f�����³5W@�9��?_Usx�m� ��-W�kP��G/�u�y;TŖ$��r��}�}D"L�z1:�����;�����eR&�+�J����_g��ѕwc؜4Wĕe������mD�Q��=w����`YH�����<ӎ�ri�mB��5�..�U"$�;�v���}����BKdt?.rZ��ND�T1�!U�.%F2:J>����5��=p�!��L���ɦ�K�=z�*R9��,�n� J�RK�m�%��h��]�k�M����'�F��I�o�2ԛ���f+��L�<S�`��G+��|G
��^d�HC!�]�$��}׋[�fw�Ѣ�?���|��5��eX�����~ь�?������V9�����oN��E"�����,��e���AڷHK���$�%���>����"U)�h�a�������/3��W��rqڔN�i����[�n?.�A�Q>�:�[���O\�'��dDO�Hԕ��}%�L*�zu��m��P+�az�.�2�G��dTn�Ă�݈%��p�o�Zu��#�U]ұ 2�C��]�Uv��(�r���uc��W"�:���ˊ�NY��Oh2��7"P��=eg��f/^����ҹ/gQ�]�x�n>w"W2Ӯ�招�J�|X,����{1�e9Ņ�r�p����r���K�f%v7�B�����z�	�$��%�x~j�/�3���=8:�3y�`���A�ˬ.N;���07OpU	��L��C������8�.'��5I�ۇ*ƙ����=
�i�*�6ct�'|@�7u�@�_�hn�;��z��2�@5M��*zE�����	?�a3m�9Q�K�vĿ�E)W3��^ӵ���9�g
ZW���Bd:�]]l��38���u&�`Y�ߢ��G�gx �ʃ�m�&�,D\�z�r���NJf¤?5��1��
M㒟��L���x��#�y�x�#�F�
��T;R�������` �EH��'�œH�u�ۜ���X%��e��a�:���?׭�$sA��$45G��"�cN�\�Rq�5�R<\]@���{J��F��	��&�$/#' �ɘ�e~3zX��1Y�Vu����u�`�-��JZڛ�K�2q��_�?w։N��yY�������T����ܦgr��su-��v��BA�)4�x�ME(��j*\�����g2gZ��n�3.IE�C�ݭBC
��d���o���f��� �X����Y�P<�3�����]V��8�ES��Fz�bV��.%�_ݷê<��SM�4�m��qܓ݋��^�Q�D\���2��O���3�0�{lp���e�d�곫�Hv�8+��ڌaP�H	VOmu�j�<V7��z_��_!�;����ڙ�зZuR��@~h`��Lv�+�o�0����^5с�ΓB�0pyֈ-�(�x���b�Ɠk��vn�p]_�FQ��t�w򼕙������L�RKk�>��Y%��?�J�tA�~�7)寊�& t�p�����&85�8I�,����&�&��6ņ0�]I�g�~���]	l)��爚(k��:J|A-3��4�o�9��9l�2�I�ޣ}��j3�� �ɬg��q�m�M��\���]��l�(��A�x�k���LCRb����be\�V�F� #Q|xjb�'HU�bTI�.�b
/��)�^��`�X����w��j!�EU�b�����N7s��^Y� ��w=d�~�yW.��F�%�@��I��Tu�jG��N��b��Q���tC���vXEմ���F�wYf#��.{TY)E� �W3����G����Y��?�wр��l�+%/G�e��u��@c����-/�Q��J��=�	B�s
<,�?5g>�h��s@�S�-Wc`�,=����hmb�T�+U�㑭c�+F�����6�=�]�Ni�2����"B{K�w!�B�$;|����ԍ�"�>�����*ײ�ҧ��������ͦ�_*�Cm$0[C���lb�fؘ�5��'��-/4�,�������͜bh��~��ӽց����]��3e}��/�|
]-?�k5"���b�d>S�1q��~M"m�o�vc��J{6��q��Y�;�
���9���׮X����u����g��`{\�7 ���A�Բt��a's,M?��O�po���n_��v�]w��	Ō*m��z�F�QDJ57m���q�O�@�M�����VDX���f�K�.��G�ْ������Gi	���j�a|��!R���bs����6�T:-�\ Ɯ+\������T�i7�3yuh�M�V���	��r'do��p���`�2z����˙��g*Q�D~�@�z�dЭsXL��ң���JxF�i�p&��@ܜ�?����╃�5m�����\_A(�(AU��$/`E�jx@�
�!Zpm�/d��d�� ]�W�o� U��\��2�jq	kK��KY��_�r�6�����Tߧ�Z��s^�I~�� d�H�E��n,�����%)EB�F�D]L�h9A�ʼR�:Ў�6˒ ��'N���%
Ρ��$���E{B�,�L��̇����k�	�h�.�r_�j���t�z�c9%��]����{�˹7�>;	��E�s!8*韍��Bm�:��[���O�W	��=fI�M��0�-�g�+>�M�S��M��D���<\�R+��>��/V��m��H�� ��%t+��9<M�9���M�Hl/�W�v�k���	�Z��0O&ވ��'d1�U�E�4v	���jðWQ�f��w�e!���8b涖\ƹ� ��J� �5£i�9NKߒ���|m������VB�zax�}��B�����.d5�&εRN���s6[`3��|�"�j�ü*u�Ai������v,��V�s�\ͯ�>^�\V��� BrG��� [)��x$ρL{��&�M͎�x�Z�����ouu�t�/ ��s��6�~ӮI�*`��D�5��a%������&�_�xg���a���`l��cg�f
�wRq�=�� (k�XC������4ǋ{N���]�K���#f����9]r��D�P��f{�f��h��� ��m���b�:/���߱m[ �xC��dH��$�� ���F��3��<͛c��<�ۈ�*�A����+V�/�#؞0�~