��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>%��}w�K�P
����$<�0�E��CO��Gg�&�1�c#Lw�D:q�ٻ�2.��+O�m���@��8,���Ҋ/����t��'� o���A�ذA�@�Չ���|�𨛜U&����Z`�.F_8��D������>gE�}_��Œ�&�9L�Eݨ�Wƴ]v��8�۾/u�!�����|l��"�j�y9�����`]`�	�5�f�4R��.�[v��R�TOICQ�y)���9���	�<�0��Y�xX�H�^�������<�EEȆ���]_ã�� ,UɌ�/��ad.��1,k�ЎI��͙�7L�#�a�'����_e�4��ݶ�!)0�B�����>-�G�]��Z�.	U�R`�Q�f���U���L��L��ѫc8��Kzb��^����$;��J�þao �������e��b�3�ӑ榏,($NM��E�?��Zl,_tg�|� ��
�ҩ Qn����Ui�E�C�~W|*�g��H����.Y�ށ0��9�g��!l2�Ó���>�k!��������A�C)%�M�񸳛%�@\ݨ���jU��6~���`�Bw�z�}0V��us=���L_�c�VF�YZ��Y�|�MRK0��:8C�d5:�0����w�q�?^ ����u�m�Сf��)�(<��4�h�CU44O9�ZR� Ⴎ�Ψ��Μ���1
� DI���)ۯR'���u�BI�����($��Kb?~���8X�U�o�$�1��58Pdh���'�G����Ų����xr1����Eb>�ڌ-Z}�,/3��9�F�,sL��n�V�a���` w2j�oOY/�+g������[~�M��<d��R��9I�{���:>�����+�6G���ʖ��ѭ#h|�qTw+v�����K��9��dK,J[�O~N�ݲ���5f�Uw���u�An!%&��sX������7��X.xtx�M�����g�H��(�4�G+TE�򩒦�0Jn�.�����_�Q�Q
-�o:�M�2A�D&�iڍû�H�}������:3;fy�����L�$�
3���W�{�"kz_����nX3�]�b0!eb�&�.p<�{�22�q��b�������|$�H�q��G$m�ܧ������NG����##>M�R#����K��'ٽ#��Mҧ˹J��viMtU*$��a��ʸ�Пe=Z�5(rA;�Qf�����ס�4���ӟ@\�"�q���󔐍%6�N���a��j(A�tĻR5Z�GW�����!.�:Tg�QAd���(+nGL�A��k��\����CnPL����;�,�ph���;ڻ��g�}.������>�Z����7UMZ���>X�z{k�Q�� JԀ|/^�3(�n+���+-:ˎs5&p�#����=�cb:��\��p�y\��AA,_Sz$��\r\�:KTa��&���f�4�R8��oVWElRIP���;�t���d�NN�0��h�ƅ��[/mq}jD�=��Z>�X�E.�QW�I�H�0�mlx'�S��x-� :qƭ��\w
&�;�%x_8:��}��;0���$I�M$����K �׈3��&ǣ�eYen���.�@�!�?��Gɱ�ڜ���cC�����*��r����tH��Q�𳡾�:�����)�l黎ܛ_q��"����U�y|&Yjd�h���<W�d,
�<��,,Q��!�Nǰm��Hv����\��f�囦KX`��.�����Ǩm/��H��=��G<P���ʣåc�o�w��j���3��"�l*��Hb	�:D���|'��}j �CԚ���������dL�B].�D/�������<�Ӵ9n+���{��AV�.�g���<;�� ���3�P.��lqs�؍��A/�p
�N_vXv�#�;]w���7*�+�'(�'
ZJ����A]1hncK4!uQ�luz�e�����16f��s!q����@���dIB��z=?�^�p:[�8#j0�����u�(,4p�֒̲�͑,7)�y(��s��y�����[]�<�e?�7��4���q�8�s��G�xF��i>�>�b�N�~�*Զ-2����>�:W��4���c�-��L��C�v�����^h�Y)"��9[Yj����x9O)���L2�T �ے7o��on4�T���ܦ�jm�g��E����q�j�]�|�Y+�-�R9�����~��d,羓I}>��ߎ|����%A���w��7�k��c��Z/z��:r w�S��+R.�zu�����U�Ia,��y]���X�'B�/���� ��D��5��3��Q��*�,�$_x}�KfT�jZT&L{\M��d?��{��v��w�LU��`0��O�x���0F�'f�/1o��fK�_�}���B�o���	q�qq�wu!���Uۙ~;�B��Amv��u
S��>����%i�$�[�=�+�q��In0��8�Oz$�
�f�"g�T9��/ �v��H��I�!�2���I8�t���T���ka0#�-9����_����L�=�@��&��1�L�����;T���"��E� ����Z�=�:C��	F'�+�X�l�H)���(�G��M?�aR�z�@����-�;N��gCf�X�:����jFgG�>���'t2�*�r�`��>�ɸ��n��+㶽Pӭ����,|��?כ/�j C�P����Y=1�i19YVK��v��u���Z7�'d ����WB	i�ƌ�u���t0$0$�� _���샛���H)�<�����v6��Z��ȫ�<+�H^��=8��529:l����1���V/sLǰ� .���r���f�^ �z�w�Nlrf1��A0W*f�2�����(aV�׿�)td�j�Q�}P@���k�eFi,�&[���LG�`��)h�s��m��!D%��Y{��o�*z�W�wu/��@F�R9�%�܂�ޙ�9�>%M����Z�uf�<��2���~����~���<)v��̫��,��n[��ShR�Q⬴�	�Z�^��m�rz�!űG��"���~4�R1�
m:�yk�4���X�?b�B�
���e���_�3�)*vQ��]=Q��L�b�o���H�pQ#RXF`����~��d�>b������P���Z�3�|.�9u^B��o�%;˛�	 ���=�`�Жx��>��k��'*d���g�U`@D2#��S* ����?t�ɐx�>b��'���"��}ig�8thyǦ�����UG��C)s�ܮs���"dr6���n5tMS������i��-�v$]��9�y�?��ġ(Q�?uo�-�,����{=h�����P�ӻ@'�w^�Z������=N�ý��B��������Ul+K��A,M�`U�7#/ҡ"��lW���$����AeL��UQ�w��5 �mJYj$a�`�Y���\4$g���l�GNIwe���ZF��VD���u8���-��]g� ��n˼�KsAF�6�k��0$�ڶ�;8��V��.Khp
��a��\ae�}m�0�vX\����ŏ�`��gf �d�OC}�!�i���4AͲ4{���)�mS���Bi	�UE�M�1�im+wfv@�?q����jéYb�p"�Or�S�'i*B�[��ji�
Gi_���YQ��W���pWˠ[{>�����?�TRB0j�:��u�iF���B��>�|=Ĵ!ͯ����(`C���25<g]r)�>�R�qG%��x��A��G?҄�E�e1_��x(au������@�_s.�<���<)@��w���M�v?���`DP�{_f���̍Xk�L�ΰ�񏵺�*����ff�?�a�$�k���T�ʌQ��2����i��X��=�wP1���h=��s ��3���t��7m'-O"œ]��c,�A7YJ]t��x�(m�~���o��2 �_mn���um�	�IFY��/X(Tcq��x��#"%�'b�e%�,�.ݟo��X��#H�x)$~��eR����g�a�n���Ԭ
n2���-Գ������h1���%-I��<g�bO�XQ_j������]�#�X�r���q��K�>���N�E�
	�eVc�HWRy�O7��hE�Z
���M �?�A�`��jk.�?�B�Z�Q����ęe�Y��8���;4[L�g��Mf"w��v�Ĳ[].�.m-K�I"���2�ms,�wD!�WC-�G?�G��&ت`6�1^pj�����:�p2��e��bQ�:����c�ʃw�l��@3��P(������kV<XI�"�iUҹ�k��z�{��SZ��Q�k�j��aI¯ŵ�dS����_^6������jm*9lx�(��F�:i��k�w��x�����
KѠr�Y�Vg�"�Tț����K��@*5�?3��례�a��C�d��ӈ>4�M]��M�%�8�4�[Em��T� �A��s��`Nc�[k9�Kv��
����T&i(����6<�4b@eK��4}-���o{��z,�o��ϻ�G�������}� \,,:B�����I1�T��E�i{�:h�a�(�C�WMa�d�I���O�L���|\&˗�|@Z��Y��_{�w穘Z��kB�3&��)�W��5����Q�J� ���c���oT4n�4�ŐbZ�D��A(����y�4-B�Nq\B8�J��%��2���<�Ӡ��2���Ã�t�1b� �K*�n �ה���U�w�ɕ)g|��?�^���$���P9��f�Fے�LI�9�J���x=��I1�|N"��_���(�v�D�p�q����͇��Z,���V�h��w���P�Qi6Q����䯁V�d��J��E�X]��[�Z��x�WVdܓ>C���?5 '7Y��#l������������W�����k����;�\�L���/0p�D[��M�������5���H��cြ��hڒP��bW狽$��<v=W�U �Y�NZx{EZt�M�������ȳd����bg�5��B擴�����$�� 2��1�1r����X���(��|`S��,�E���e��p���
��u��$jn������M�>����-_�όL܂��cV������˱�U�)�^�8���ŝ�=��� ��3Y%!0��^�s���wx<��`�[�Y��L��E��*�,���4Z�X�J�]{)*�]@}g2-+���?x��N3.��Y[yH���oįxC�;��/��m��{�����I�۲�os�T]��~�9~��]�h��S̇<��%���k����.�kěϲx�ly�ENϩo�6i�';�c��$\����֡=D(�E�@���Z�4�~�oֻ��nă�WWr����_��qk4�|��1�i�&�&ē;�Տ��3�ȑ����;��m�E�;*�	<L�<�5a<w�!C+{��F��Ç��~`�K� Zinө[�&���wŶg��'q|Ǭ��/���R$�}�t_�07��S��|8������J\���|��^�+tKק0�Ě�Ԓ�m�j=�xb�R$)���_%f��\��2�n��+�	�$W`�e^8MehN�z������ B��fc��m�����F*�%���Sn.Y*�K�=2�Gя%����Mު�r`H�=�����'�kW�Nt]��`�ҳ~-�z����&���B��T�3eN�@��g�4�+��6Y�gh�8�� �H)�i?��F�ٺm �#�z'������(���!s�(	�J�=[���g�y��Y�d��X���Duw� ��$hX�'�����f,�.Iq����H�ӿq�@��lH�=m?7U'�d,�˽.�Hn��
���u���e�3��)�;�Z�d�W�Y�U�-��J�_j�E�O�|��cj,����0�	��@��}���5ɽ1�%80`g�����Jx9�0���}9�;3����ɐ㐨n�tگ�����<b�K�A�`װ�f�~Ұ�33f,y�x�]�,�3��bѐ�0n�4����z��,VS�\��Ӿ٤.�z'�����ul�A}�P5��(�rU������n��a�ȕ�p<�wDN4���CI[�[Àe֔;Ck-�4z~��w�3��Gă?��4m�:\:WYb�W��D���Q=�h6й�yћ������ H��t���hu�]S�ӽ�� '��`����`t׎���4��ׅ �iݙ�V,~<����Uf�֌�ۋ����Ȓ�	�"KF�cv�j<!=2��c��������@�J5YA�l���u&;��������{����IHLs��1|�Ғ͘�*�[4
��F��Lx��C���FSt�������s�ۑ�B��5�x�׵�B�N����fiM���������c;m�tEr^�J%x��	I�f�.H�i�

�?>�P(kqRwW؝,�=��5��`{3��6��{*�!��35D�����%�i����\�^�M��J���Y�+��t1�s ��W��V���9�Y�����'v��݊�ǃ�$XZb�̋z�X�����MԴ��ڲ��eD�����F��v�%�
Ȕ%���;)�Y٤/�n�_(��E�Y~����r��~(���fA����J���� �r[�T���u�i�e$��u������p���<��[܏��f�wZ�(~��>߀��	o� w�V @ Aߎ��l2���ɠ��a�V5nk�e&�M��y��pQm��ЅJ{FM*=A��d��9��ؿ
��.0�nfs��v$�<���1��������p��s�vhײc�D�=�oRdUX�C�0�.=�.D����B�����W�S4gw�vBӼ�aq���1Q���촴��# YO�)���������KiS;��vK�����zZnӏIpa��s2b���I�%��e(����Q5�"Յx��e뒄�eD�C2.Q���O8NC��(�֞`H����ten3L�P	Lp�Yc!��ޯ����@���''�o��y��2f���=�I�A/yaD�pO�����A��P����M��?>���8E�uSBKέ�>����9 n���U�?��4��k��^�2��B���ri�7g��B{������G� ��(5+Bs�����T��a��R&���eEԓAu����8����`⍥E`��<"l,��Wއ|�&Z�͗Hx`����J=�t�W�gßSy�+�ٜg���a�OG5��(���t�E�d;n[�J����@ ��^�b�(%�na{o���ؗW0A���W�GjB9��m������@��28(�y���4�{�B�*H�^�
T�)�� j����]�*'�>2�s�	�������ŷ$p�9��|3EQ~�u�#�\���rr�B��-g��=��d���8��ٟ?�N��	�ʇA�e�:h��~�Ƀ?��!	��-"^CFtUݗ��&ڷ4q�_h`(��ߦ�ƚ� �W�v"�p�H]�8���7X��IG*��Zt�ܚ��MאnU�����<�ked�<:Po@��z�
���>�"����;N<�,��	Q�,��d#�<��)�����CV6�O�{q������r$R�l󆭬!�� Lq�����/1��Ro'��h�Z7c�S�&G��r�F�5J�>��AR�?�R�;�F�9�P�x�[���6�ɍ��P�h�?AG�C��9���_	�ǍX�c�(/��)��eN%.ˑ�7A]#�QE�`e�����:�xKM�1aBl�oNs�2)�w8������Å��b�⧎h o$'�) ����d.A�齎8��s�U*f���Fừ�7�H���&s��Ti��m�>��c,����1a0�.���~?�T'����z�	�'���}�Ou���l^<�w�l�Q��1`�s��=܎�W.U�2~]c���Z�~1�/&>|�e��d2�6��/�y�=4�& ��|�3]�����Tg�T�}��֣!f^��������8B'M�
�u��|(�iAf8��c����]���-�#=n|�G�˧R���-��w/���4s�SK����»+�sE؛��YD�(�0s�ծ��� ����A��u=p���� �j��U5RH����h5�X��=�(~$g!�NB��P�&�Z��5�3�ݜ�jY�� �3=J8D��M1���n�u3�@��M���ҷT��VB>�Ҭ�s�H�j�Vߗ���V?�ph�&���f�'�`��o<�(
�A�}i��;%�Fҟ�	� �p�5v�'c��?L3��Wjs���.��:O�u�+����;O=��'���ɝ�[H�5B�#c�H�#�h#�{���B���������J���\�5pnp\ҩ�M�\?�N�壳�����.d���Dn���4,��#&��>� 9�+q@�.�h^����̎�B���R͎�Y��3p~���֝�{Bu��ƕ�� ��W���e��_���5ܭ��<��>��L�������	ߎ7����,aH@�-���z���}�㚂zn�-w��*e �A��NCܥ��/ 2���J'E����4�[�����ڕ�d	��=�=��V������9�0`���u��
娥z�'݂<�X�]��XA!wc$�����Rd'K:d���I��p�A��tB�*bCQ)5��d���֮<6%񲍛n�E,X���P|�^���*0s�.)� 
=G�a�6l�i+��P�5�Xk���3S(Z���8T�9�ˡ��GY��iP<�6�D7<Fsi������y�"�ah�.e$���Oh���d6��	vc*d���;@!�-%���r���PUK���V�����ڮ�w��zv�+���x�ǌ�VS]e|�6*rP��*��Jژ��ЁB�28�y�]e����_k�D���#�W�d�
G&�A�xU�^ w�J�:ϧ/C2�k�7��!fc,Li���H�;��D�4#�"�1�b;q���Ά���T\3�Mz�েb���8}ʌ�g�ծ�4.�
�lV(�``&f=`�1���W|���C�,�!��x���i�Z����n1�	�CB˳F�7�	�/��#4�j#g~A�O���gi����Ʃ���aI�q_�bjƟ��[;yB !▽)�Խ���TP��u-S�t���)�F"�Z�(�! �vh�~}��4�:�x�Y���-�#� l<��@���0�E|��z��1"R]\u�7��Je������[s���l���ֹ�C����`42�	�B����0~y�ݳ{+J�l �(���v�rCh-�	���L�XǑ6�L���W7/�~ْ (����4�%h<�R_�R�/<��G�=�ޯ�!բ�T�N����r*\^8���2<~�n׃#zN~U����A>���g�>�,!�a��\e��GA�ޡ���W�Ȧ���}3�,mՓJ��@҂m�������F,����v��Y��OT��
Ϝާd����_|�{J¦s~o�����C��Le�[�x		]T�]���0
}�N(*�1�S��SCl��VV}ȳ������%J��/��Q��+R��}��O�ił�Z<{S�~�g���e{|1��������q@!�2k��	�Me���W�ļo�*�t�&�w�
�^���_�����m�YZ��Q]
�U�Z���(��bׅ�@���1M�����!��[i�z/������?�`<ԛ��1�1�p�.�[Εz�7�y��E��β8�����!~Q��Z��H#p$�` �lc���T�8��I�.��O-��ޤg�SR}�[ ��ؑi��c��N�@&���1� �@^m�^��Kw�ox;�@O[#�&��/7N��4sl �D��r%|��0��w�A�@�Y�T��Q���N�#���@����jj(�������[��z�Rz(����J�2���$�1����C�o2��݋�w���a����1ڴ�J��9��IG`���y�*y1����CO�,�gC�\�\͠d<S��09(;7;w��%.][ڵ�挛B�x���]\�3X^�;�R~�er��A�ף\�E@C�;6/ �H��2ZuZPv��*�]G5~Cͷ�L����c+�iڂ�I�ntڔ�^F���ҩa�KB�4����z�]*/;�����䥬��E���@��J9�����T	�Ss�w?+F���{�j}�u��3�~�:�u�i�=#h�H��~)f��iِ*V�TL�Y�v'O3�ɞMq�(^����.|G��f��Ƀ �Cg��k����y�|��(/�����|2�f����aw�f�T�v�q|����y�\'gIß���{h��2	d�k��LW�Yz�fx��]y�e���v�l���(j+MHg�ү��N�/��b7���1S۟lN�xm�O�e5R�f�cА�n����v�'N���RT��
d{&Jfŋ�
�g�%���a�����d���Y�Pl�k�>�N��e(":�(H��QK�獿6���,H�+����f�=�(6c@l�e�  ����4f�b��%y����`��O�E\��^�����'f�d!R���~��˳����t�6�+�Y�"j�n=�Q&��'"Ps� yLP.$�k�E�%/�f���W�}��t�6.��C��y��X�pd��u餂����+�8b�OLjQ�`_�x�������4��Z[p}�%�� �*���_�M�G��B"y���~�d�11,�������C�h�SG�9;fp��ӣװf�����1�g� 2k�9ǣ��zv"�=�'Q�fl�0��ov��0��C�"�O[F�~�Y�>x����tjiE��	�N�G�^��=�5vF�P�7-�~"֕V�emx�
��70�P�Xg�ME)`8���Ƒ�?���x�j�Ii�؊BeV�D�0F��2�j��Y� ����3O����>��Yơҝ	�٭�_\�$o���W_S5r�u�dk���;��]�#�����W}���ց�-ҕ���)H�x>�s��-�5��NɳV_�t/+ٷL��f7�s�<C�F���C�p���|��HiI�0R�>��u��ws{�E��qX�¾�'�l��������?OT����r��V���{��;YE�z6��g���W��"u![4`���F��TvK%66SmđkF��0�U��No����g�n�E��C�A����+Hk�֎�찴�3�ᷓ����B��ɰ�Hs�{�K뿞@��r�I�R7�3���-Ψۥ������,����6?,�-��t ��dpo	o��Ϯ>��!�H��'�J