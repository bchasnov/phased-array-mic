��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|�L��58b�Y��u�o�>�ER�')u��0�>��^s����(�����vÍ?�X0i�!$��{��$�qu��q�9�aQ֖2�}42�� b���ml�"#����v���������d�=�I'v��~�W���Rx�!�ǒZ�Ln��f������9٣�n͛h�K`�z�o���d�Ϡ܃�������b���1��#o�gNt.0fF&��d����3��{_�l*��X)�<�I}x�p5D�����- h g�b��5bl6���6^�����:�7��[8�ꕕ���p[���C)ŏf�7	��9-j����D�BE���>��X�6
ʹe�P@���g{�V�;<� .^�<�.�@2��x,.�]�7[Fq	R�af�	$�E���ʿ�[����$.�;�b�y-Μ�3���1��ϻm���va�\l�2�7��Z����$//�b�H/x�~*����7�s�q�=�آ�����)�B�'����܇K)"gVk���r>�(��ϕipmP��X>nS��J9אI��
['Cy��+n�]lޭ�hi� �?UO~��n�`@]��\����ya��<��Ir��ŵ1j�vO��v
5�k_zO��	Zy]���<��i�sU.���j����Fe�ٮ����$~����{Q����wp6mC�8 �]
;ĩ�K�暚+e%G�r����Q
�ٗ�k���7�W߰��mt��[M�5(�WZ+ْ�(¬��H�D�D6�O~;yt�mԠb�X�n�w~��T숕\��Ivoo[����j>�P6v���^:��w�M�{:�	�Rm����~}�7�9�S˃w��hH���k�ěolzK�,�sT�r�m�#It�MG@�Oђɽ�����=c��c!P��; iu<~�{ʟ��)l����x*�=�	�B���5��fXR��K�B�� �$aciGE1}t���t�@��+q]G��`x�Q�*J<vנ����x3���G�����B#K��LJ<9�ȶP1���M{,E��J�8�`��xԇ�Jl�K�(T�s�(���'�Q�ruMy�w�	�y��Ы�M����9�4�'bm�c������A�܅:��o܍'X���ܿ�冷���ey>Y<
5�E$���iN�|k>pGcV�BNb������cc�d��o��7Ҩ���#H5j�ܮxM ���2���%�p��I��.o!�Ѳ`�8�h@SS=Et�Xw�>o�^H���Id�C"bq�
��!WR�u�9�6�z�����{�ާ�V�x⠗���Ԟ�9���~_#U��X�m���f0΢Z�ó����Zԙ��Œr���>� $��gM�����_�J W�I)D|�ڑ��� Ų�GT��DJ��p�k�u㫐T���q
���/͌��Y��;�\�5l'�}a�(n���K���kM��~�l��2m��ٱ>�KA�J��<q��{��RV|����� ���|�2��
v�c
z��'���BZ`���*X؈�㥃��ą:i2�C��z�I,zo�ݵ�)��J��uً�؏ՂB3N�|�G��X6�0/~�I���0>�×� �*V���~��~�,3:�1$A`A;Y'W4�pU�܅aR���,���]�#����W�[�h�҄��}�zܬ�5��348���
����Ә~Џ�#6�NVNe��y]Ӳ��9��R��IP|Oኗڻr�ˏyF�ct=��=��r��;��e���+�xo襒����J<x;�@���a�¨�+�$�xΙ���ZB�Ϸط��\�)�=D�9D�ioy�8�Ὃ 	� ����ſ�>��Q�OA�p�h���8�FY�J%pnmy���ؘ-�9=���KO����[�o������B�׳�^=A7Ȉ��R�ۡ��o4޵���U�#� ZS	�^0��>5���zԗ�SF�!�d�7�Y��/�,�t���Z:T�,��U,{I�����R�e	EL�8���{'�
�
|�_�"R=Nc%��y�Ҽ�B��2 J��Q���y�wݙާ�1k���	�N�c��^����yU �ٹ�i�3��}��R@��!��J��M���:%�΋i���ST��.0g��m〿�}6;<6X@w��,z!r^w���|c=���Ԣ8����%0@�����Ө͎D����&c.V� c�g���R�kQ�`+=6�
�2vp,�2�{�%�� ��]a���#P����M��A9 �:.gx9SP�2�,�v�_�<?��Tv��&(�<,`Y�������W8�>+lI����*6F� ŧ���o�mx��3��G��@��q�]����|:�84�����"���JY6,��o;e���,��HU�$5���[�?DsH�B��R���^_f@��"�hQ�P%~�Ac2�|�)ѯ$
���R��=d�(�`.f��%�O��pNdׇM7��ֶ�[�h�Kŀ��i�൝��1ҫ_�2�֩�N��~�K[����!ڌ�f'�%�!Dҹ;w+|y�Q��`t������T�O�ћ�K#�Bhqrн6�^cSk�xՑ#���z~wi2���j$t�u�0���r#��K����]8��v����7�u���#SqF����>X�@8�iޡ���0'o>wh6�[��Šs�}5V�`(���x��Z6�Ed��^X��&�����
�h4=��+�ח�g������XH8����}�E����ȗ�rk,�T5��H���F5�t(���	��uל�2�^��"�{~f��}�=�.M��6���x�M�Y�l�R�S�I:1��+TW|(�35dk��,WEY&2��c�k�A�lm��I&�|*��W��t8��2JF"BQ �����F~��i��`�᪝���zײ�dڀ����/��zf��[ϸY2�lA�fa������;�y�Ղ�9Rt��J�e�����C�<cݏGN�� ��~k������v���w{Dh���z҄��#����w6q%���� ��k�J=���C�t�ߏx~,�,�t����/u�CZ�W�:"��:An˗�<r�#��p���i��z/���$-��]͕�
,V��.�j�[&5^ȏY����F���q�я��r'��4P�*WdX򭝃д��q$�%F�� �\/bœB��ʉ���1L��%~��p+)Zf��|>��vC��]գ�RN��������`&�ө��<Tn����~N�B��gN���p��5���^܌�xrM�~�Yv暤����*. @����?)S��
� 8pg�+HΫSe�����3ަSMM��@
q3���m�S����!J��(=U�ϱ�t�@�IbkrN�Ae�k�+n*e�4a<j�:��,���܂��ϝ�ʃJ���s4�l