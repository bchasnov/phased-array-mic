��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|p�n�U�4���]dkf[��cXOT-�\�������GƟ���M� ��SƵ֣�߽�Jl�q^�2�@8'P(�6$�5�s�t���=|���-~-)_�k]�t�'�@�5��e^ ��ᖨ���L�$��&���п"��A=D-�tNS���U8��a���v�e�Ԡi]
q�M����z�@�����������^Y*���K��غu%�%y�V�_u�Y8�$��o� J���S}��e��L�{B[
]�Q�'�lR�f[����&p3�ȏ�l��&_j��d�i��1 ��RR�G4�z�4Q{��6�G�� w���
��;p��)�]:M����d�Br�Q�˖��{~G4.]�ñ���{6ӳkL�8=+e������︎���V����÷U�� s��T��H_F#[�s���*ˉ c ���f�-f&Fޝ5�v�F91�Si~+t���茝s#
��hݝϫyj�j9@;gC�v��>�7�
�ŢD��K�!� ���+۬9��|��-���p#���*3�Qȗ��v�D�/G�����Ͷ�!P��í���چ-����R�M��}ՠ�tHTr�e�<�nGv�ę=f0(��$���G���d�\��&l�U��N��2F���}�>��0ߡ5F
x_AB$�<��ў?u2{7���K���"BN�=�g`��5���Ӿ�� �����v����	�ؤ��Cj�[_�ݨ|s�{�}���0�p�J9���)���Wx۰9�>�Հ~<����(����2#E��g'P�E>W�I"�I�Վ^tZ&/�B��s�5r�<n���C=O�4vM2�SN �Z�4�&�I"�AH�^3`}~
��Q�Ia3�́�謷�-ϒvzĵH��y&����D�~��p0V�2i��S6�v�?FnP
.j+��Fy!�x!D���0RS1�fշ��o��&>(/w��؜�"������Ҍ#離�� �qw����K<��p�Fz� �e�EF�i��t�P;��	242V{���ˣ►ep��6vVd}C��P��D��'.phrC��X�1ܗ�/ ��`��<!.�!̊��,��R���\������d�2��������w�j<�����	�$/"�����{YԉS���N���P4	v��o�h5�㯢�4f�V����|�"�,}CM+�p%�6*���I��}�O/�����y�?3%c_uol��O�`sHh�6�Z��
׃�'P�~ѹD��!��!3A�u�ʙ�_�Jڟcƚ}J�/Vp��R�&.�,\�خQ�"�XP8y3����H���sCciX�z�A�q\9_:^L���6Yf��7��76q_�"J<&]<(;���v��T#�^��r��TJ;t�Tn��|����.�J�w�������h0��I��	��*:����}J��g�����n�ʙ�$KZ�b$�7F�TH��*|�k#h��RD����̕S����6�%��x��o�������m+�]�?܂��0�~@��2��>��7}�?��_��Z/�43>�e����0�{̔��� ���@��W
}��z������'p��
b�Dz�SB!��$��"�y�ԅ��i�1��)�N���v�?��ٝ�{�/�}/%���X���	�8w.�0���XG=���w:�Y$���y��f�_�IuȜq��I�ؑ�l9n5n�

�L�X�ډ~�g�� Y�I78OFx�J{����gG����}�u�6�t�2�Xb�& �<D~���]%^���4�C�ϼ6�|*���z9�.�Z�����54]����2r�'�
0Y�ĩ[ ���F)�{S�ӆK�ɼ��ToYf2�9����tkB5��@�s��8�	��n̦��'E��(pAG����-+z��Ɠ>2:X�i>�L�/B�G�3f1Ƃp� ��9צB��YZ�䕔���+a�;G�#��\*[>!��d~a����ϧ#K����w����,$�K��k�0��=��?�3��R%੎+}�������ڻL`�D�:YE7�Gm\�27bGE5:NIt!
���J����3]�Vu!��4�H+��G~��2��3#M�׺� �� �^d�/W�@���(��L�N��a���0)��xNt�;'}�rʟ+T��޻(����ӝ#��e-�����I���0�d��,���=n��0�A�^�i�_Ve��%@D.��� �w�9
�"�.��8c(��H���2Ezv�tݻb6�ė��/u6]��Y;����}T�a��,�����H�$!�k$�z�����D�hk����<����A��ի���!�̊�C����K�ysM�y.�iƁE�4>��5S{Q�$
%�{Y�{.J���~�H��B���?� �����.�	�F�Gx����m]4���+�F4Yك=���h
���t�Ҥ0ik�0b��2u`= {uvB��,�H�U�OEͭ��h��0�񆞒EU�a1��n]������[H�q�4'���uHAm�^T7e�Txy����d��|Xy8�/��V�5u�V�
C���aj�+ݓ��q6�������{��xې�Q���M�~�,���c��ǷH���?��D��`��*��-؞�r��{�ӺK"�ܸ~����x|$|K�������0���Nd @�xv��F���3�1�H~��}{���rQ�R����q�����o�������bS#�>�ŋ�O�8�Al8s3�8�3��j\|.耚2�O�f�i��́1�\weq�~ Yw$d�y��������v�Ʃp1E�8ĦY�̓��.qjE�78��t�l{�I�#+O@N�y���]F7��H8Ƽ�4IK�]%��d��b����9��r��M��UuoϿ_g��0ׯ�p��J\��c`�wXk�	9��\a��pJ�f2� ���b�[LJE�~w|`������qE_�I��ha�����pR&(������3�fRH���k����]�|f���_� -`�&���>����4��%Y'�#s��W�]�,Kv�Ԥu���l�
8q��ځm���k�+�z���ʍo�[>d|�KJm6�\^���ڼr�"�⬌�����m��x��w)	����Z-7}��3|�T֢G��	х؜��0�� �&��:��w�U�Dn����w�cF�;,rA,�Vn������Rng	I��M��9�����tWU�M���M'#�ӛ
ە*J��8繞���3�[P7�<D�M���
���7sx��
�&���U�[|m<�n�n��yY�S!o��=����d
�$�h�6[_��$[�ri�,�i��Q\�䄂��� ���ݩ͐�
y;����9�n�y�1��C�{�9H�����'�<&ɲa4?�M�f��/"3����PK|IR�%
��<��F56�h�탖5�9F����U��'��	�#¦�4�R#��Ǌ�/��{<:ݟ���W�b�]+7>�P�!�Y�= ���N�/L:�*Sυ�k]����0�c��-$}��(UN�"�7��X��6Nc��1�P���Y֍�:�KE�^Ы���,���5V���Љ]�������Ζ�Ul�R'��Q{���s���#�{nw��t�yåy��wTb��KM�
v����Iϭz����x��u/2M
D�9\���K�vX�����,9x���M^j>�5��'/L2��N�c�&�C�#ɨG�q.��yխ|g�ГHܽ�IC-;N�B��C��	�:7�?�vj�z�5��0%�X�;& P-5[u�v�)'HE����h���Axq��M�\2A�dW�8Q]Yf$I����=�f�KU"�הQ�2@��w�¦ up�(ܾ������+"#m��I����\��MR]5EtƮ�kZ��-��5����	>��趃����I��^E2��Zg�M�Yͮ8����&��Q����?�st��F�ق>�Uu��7�Ki� ��7�I=��� �n�{ջ:����!�R��!���\���[�q����
�x��+in&>���0�Op��9����eڗ�m��#��5MwN.bj㫸	t2���,�B+��Io�s����r:�mHژ�٤,�y�m��}k��Q�ď�_o7ʻ���,>���|z�}Ļ#{5�b��Fi{&�F߾.z����̀���)�cm="�w������z�����4x�OX5�᧙���LAGid���L$�A{�-B�Kg�_yT���y/0Up\am}��� *�k�Wϭ�6�m�i�[]�����t4��'��g'�����`ߙ���%G߶
ˊӊCd��╩3����,k�lf��8����)v��>�Y9֥A�툼�=���GTү��|i5,�f7����g�g���%=C���Q�S�g�z����"�����w�%��f�#Ҽ�3�o5�����߱�*�y]
mI}�ЇY��ԅ���Ȧ.�>b���ظ���Y��S�U�٦O�����>m����뺄��� z�ï�awo��~'�,q:���Ib�6@�ܹ�ܺ��rđ�.pu�o�Y��x~e2
@.9��y���������z��d�}��N�< ��3��mV���<U���j����B�͘]v����ٰ�e0�/�A~q������C��J��`����1��Ҭj�n�ϙ��* 6> 5DS�hϧy8^n�����A���̔��w��
���u;'�/q}����:-d�6��?ρ8�`F�{TIu�_6�辛�Rq������x�NjSJ,�tK�&�Ik�Md�p쒼R�qE��m8
0����L_Z(``y��xR<F	9�-)�bfӢ���W�������'�*�}��+�#�n_��Y�l�s�� .g�R�*�5�� K�	t��|i��y�
�	�9+�N�mx���1���ᕆ��j�zF��Y\{�'Y���r�b	`ק��
�M�5���;�C"T�r$��/����#����[YZ�������۸]M�0��Ih+U[�\
��7�KХ�|kJ�}��?3�0������i�d �g�v��mG��!���b],�9͢�K:p����R69! ���uoJ�)�y��4�s��ͳ![�]�8����ś�q�0��޺��/�z��~RD`E��"9�B-'V5����Mi	G)`����1S��Ryۀ�KFH&8�v(\"H�2�h�@�a4^V�StGGy_���i�nT�������7ӯ��<��R�kֵ�W�nᙫzy�jK�c�*�������#>�=U¥C��>y���0&Y���!p�p w�k�O��*:)� �Oh�q{��>)(�Ju�n�ed�R�e�t�u{B#�'�^Ev��I�bdS�a~n�uQ��)!���+���\�'�Jf��+D��S�5��%�6�#�z��܄)��;�d+��5���(	w��?/c��)_V5P�����&������<�P����n�g���+ܿ���{��j�����J'���̓E�{t5�a��ݣ�
�ғJ���/�sv*��v�5k�O�e��W�pWAu9d���u��5`�7r��x���ı�q��Tr4iU��Y�0Q�MO��1\��	;��Ynx7�p�tʿ�lr�A6���)f/F�EÌ,Q�ʰ�qݳ	����fLC){�_^�u�ٟߤ@z��=�o�b[d�LE�k�oD�,�Ɍ�8��y�������-�?P�za
Q������g#�)P�F8iNsX�l�T�D==��.�q}Q���.�~?�F�F�<D	�\����a	-�P��@y�C�pWZ���cb�*G�L��f�|?ID��5Z����2Z��:G6~���g(_]rf��I3�y����h�Wn�����;�L'cR�I�r�ZV���?���P �=9m�۷�e�wq&r�G7�/��ǲ����X]�2;�a�����-�>�[���}A=4�4�t�J�<!��*g@�v���rԾf���`b5�k�f>����-��'�K��M�V}^�ghr�|+��̸;�������u��P���9!/C~�	*��X�x0�&Զ�(Z��
^氮R&�4�*�l�� �TУ���)��P��CR*g�٣�K#α�.���U��M�g�qU�7���ev?��T��\���\T�=H��x"_���DPB�?����e7T���'6�b�L���Ʃ�����xV�N�)ˁTG߄ (��K&<��J����7͉�$}���q@%ڽCN��� yZM'kepϸ���U�D�2�#����ߓ���@瀲R���������b�$�WT،\�s�	xxĥ���b�7�T(�u��CY8��"����pe}
9Jiط'�����>�;�\���t7_�SŐ����ۋj�i�����op�JIˎ��
˸(+^L���D!*[]����?3��|ݻZ�`4S�m�f
����O�9�1��xi���Kv����5,M}zy2m�˳��U��>G������*'�<\�R
��7�����[����\� �DQ@��$�n���ŋ����8�۸,��H<w}�5&{#<0qͱ���
<���}>nt�ˎ��6P����wid�0V��t�k@�����6�F���5�߻Ʊm�3�ϡ�)�FT����F��W���I��}��XcdtJcڏ����Us=M&�]� Ks�=G�����MNT�l�<힏�*��n��w]BV�9}J[Efm�uKQ|.�3��E�_w�����\�����f�:�-ͧ~�3��!�8-�|�n�:1��B�4�x�ub�4Pw�)P�-I��6i�$e���������ih��\�u�6�u�J��z(UE�����h+�G�d�=�����aPR����V�d���*�9�<-����_z��9���~�w�P�\G��x9�o�/A>��ʐ��Ѐ��~�E������
�BX��51G���ND([��#��.���61�FE�c�۱"�S3Y�H�P��:�C�3���f%���Kgd�J��'њBwK���I�Y���s�����`~ty�
�߯<`�E��7��\[�/�,��2��T�7��w"Ay�TD+x���!��\�"���T�E�����9������6�R� ẋ\���I���D��":���L�]/`� �}N�d��"j�T"2��ۻ��hW��s��$��5�j{��LM_���-��C���'��	�Z=-tw�7�� ?:��^kJ�]�M����b(�\C�<�n0��7ۆ:��2!��:�/�O춫�¤ѩ��+2�?�3��Jg��8�~�b��3&�1��*�)7�^Ê]_�Ҝ�У)�G9�����������4/��;e��.^RB^�"�"��*g
�ў�sP �BT,�?o��P�6XFك=6���Ǧçb$��s�x(�ef� &����<F�l��WV�*s��}��'CA�uVȏ_��a��%!����ߞ��Y�C�9���)�g�M����r��rw�k��$7����M��9�5ڱz;��i���`	l-a'm�����F�(�c��3D�,)٤:����z-��ڤ=j�kUZE����i��B�6����{�����;�҃�~�C��}y��w�͆FINZo�8�1Q�������4��-���5�iI��f����$عr�4Y�����;��tD�N�J�ro7�G�U����7C�)�|.�4����e�P[^�=ٝ��n��~ԙ�&��)i{�ï�����}W�(�b\�c���2�ù�v�B�=���=Z�fh����x�A�zAט�[�?$�k�'c�A�e���^����ݥ��}���K���w��H����{���3{M����:&�!�ծ:xO��p��1�_�bؓ�a���A~�<��K���. ��2�9
���Ie!��O�DH��!���ZOZ�����Q�$���ڧ߻����M��lh�ƣ@~�uh~|H��!����K��x�Q��u�h�0�wG����|M�W���ҕVJ��58Ɖ8��=�/���<[�ԦB�fR�طSVϝ&��7L1^.��X�I���� 7�l��[k��l�M�)Ds���{7���0�qH���6��#�o� �-�jX��nuH���y��t�C�Y�|�2��W�>�e��[���~`t3/�������v����h���W���9�+��M��b���Y�h������ A}�ę�.=ը��}�	�BI���b$٢��1�2�;G�V�O.���YX�%(�y}y"h�d�vv�������3C�<o�UO��`I��+l%<Cl��R����`W�$ۨ
S�!f4��Je��;d��˘�h���DR`���R��򹰻��ؑG��L�}(Z��\���!�����ͼwJ��؇�sj����b��Lҳ�:��������5F��#����$�ɕ����6S�!g�� ���N1�����Nk��������Rzz0�"#����G+6����T<�TZ�=�J,������X~��B��U��B{rJiV<O�H�Q����'mb�\�|Xڹ#t�~�
L��;��'Z��({UkD�=�!��;Wg�e+��~9�\/��W*: ��A&��$P{�9��R�^�9�+~�]a�{�.JB��W7���W)e����JW���P��F������vDϫ�$��J9J�k�8%i���*���"ك������J�~zծ;QM�R[oi��>p�d�9��J^!"؉����fnfh�==�\^�9����		�Q~�X��׾�Fz7)a����g���Lr#Ǘ�W�Ef�8���;�>>.Zi���#پ���_�S�5�.�w0�����t����}��*Ѧ=fO$��+;���Kd�b� �ܣ�hlܣ0�Ϝ�N?&����lgPu�Z���OG�0d�,+%�:w�"���Ǿqvsat��Jqgt6B`��\o
$J��73�ݽ��i&nNOD\5���o�]S3	MP��A	�S�jw'�(�-�DTZ���d\�"�g�����7�,�D��j�.�����ҿ�0i�J	;(��o�'��3��C�r�)f}2�����F�i��$�=��)��͜�7���kv�s��Rr�p�X�jENW͍~�L;4\+�4CP�2�����|�����y�����"TJ^W��;�5�[��s����H�[�i���u�{'O�^��$��=�f{����~�8d�Q��$跍�������$����j��*�	rm�?CPf��>�9��uE�.'�9�.������+2=h���[��w�\�"������SR��� ؝����o?��=�Z �9!rz�S�cD�*j�2�V3�%=�/j��yW$����R�
m��{>%KV�Qn���6H��CS7��	��:R�V1��>��H�](����fT�$-m��+�ǹG3F�;���A;u�d/����O�T�>SY"�^�G�:{���6��6����]���독�uv�#ޔ 4*�^��uơ A��~
� 	o��Ck���0<�r� B.�ϱfy�K;R`z�Oco߂��C"1�	zB+��U��>��K֎�	X�!���&2�[�]��ۥC�M��#P ^c��?,V�2����8�m��j|�0�C��y���jЅ��7)2@b�u{e��;R�l�r��:ުՂ�W�MTG�aH�����tH��{|a��[@bi�w���X�8�fCT���eL�)D�����u�"���1���w��ߣ�Ld2�� �1�ž�;Bh�N/G�>��0�z��"�'2��K,0�}l����\��~Bv�O�*�ov('(.YYqK�L�`��(Df(P�3����_�x�]H�N�s��"?�gǐ�����\����ݶ��,��r��=�=�*�j���ѽ��G�>��!椳������m:�>�����k�?���E����*S��}^$�A,����fp�mLb�>aA,4��*xLNo}IH�P߯�˅s��vS�;WB�I�eϷ��q�B�r��t���K	�G��/�|V�(���;I��ӛtg���C�lʺM��6�_��n�|�q��4��(���A�c��UH%�Y󷡂��UσQb���G�>�wW:�(uzA�m%����:�A��ڕ݃hU4A���+�g%���0�:�1h�@0��MŢPE�h��d�W�F�ݫ4�*��Pޖ8\y��0���u�� CQ_ދ��j~�e���)���>��?����.#^�кc����5�[<�������=�3����S`Ha�to��qk�*���w3޴T;T����]�0Fj��V�S/ѓ}b0e�*�=g�����,R��U	=��vJRy��^BGB��XW�@�����8�C}RIk}�0�����?V��,����y�0�P!���
n.W�͎�𥉑jVd[�ۈ�V0���1�"�y������f<�q�!>����".���F�8�i��%�~�I�͔_Ea��ھF?oJ�S;O����BG��R����Ӵ�s�Y���\�Ղغ�׋�$�/��X��l��wy�z|���//>,�g1�S�=�δ@�)�����E�8��!�nb-!cq�����j�ع�!o�zBt�3����K%����q�	d���:و�)`8jE��tf�e��9�A/��4_��[�v��%oz����W���R߀T�~?�i��Kڼpo���I7[�b���'Ɗ�� *э��Y����c�H�r'��ڦ��
 ��N����J�����̻n�!�{��q['^rUT?��&+(�ɜ{��)�n>ߐ�E�9�p]����b�Ì1^"�}0<&��ʽH	hr�X��@�B|�v,�AC-�98=��" 3��XGL?� ����2w���ټ����?,b�'��`�9��s�����K���.,����-��HOv'�K�V��c,��,%�'+<��J9
�9���K`�ub^�fޓ�e����v��o��g���݌?��@G∛���_��q�����-b�q{>�5��8M������ phJ�3�-��d!��;������a���/~ou��%���Ʒ����d�c�]� t�pKLGu��y�d�;OyAuH6��$	� ��H;��h�z%���~�>�2�"�H�1�	yKd���
u�֞?��ÀH�H����N_�#/s¸%�bRӭE9��L��խ����1���7`�xr���郃�b�n����M���v]�7��$v}|�����-�Y����U��M%5a+�����cO�Vbd���Of��߬'��T�^�+lh#M5�`U�j��z������䯋$�v]��4��{���>�3��>������&HP�I�0� ���θx]�%�#!y߱����b�N�����gθ'�e!EL�au����p|Q��cj�n-1��]9����8_�2���s�Rc�p�_A)&�ޘ���'�4�0K���ǬG��DF>���:"��;��b��.wՆ�وVѮ�	��%�|	����L˯��x��0�k��E��31pr�%8ݧ*�T.q^]�er��.����p6.c�Y��&wVp����M�R�4َ�E(���ؾT�G�R5���M���][�����N��=���������$T���{�_˫��K?_�s�*�u�(Eǀ��WR�n?Z�&�T�/��̫Jfr!䣃���(�B�;���T	�N'��i>�\Pwa�Vf��~^(��_:�s�~0*ؾÍ���A��­�ƭ����;�>����#{��5r���i
{�sYvo���o<�_$��:9z��-2i�T��k�J���Znr��b*�O�=��1�q����J���"e�C!B�-ڸ��L��uWBϣ�/z��v� �[V�п���m=�,*%-�!��4]d���!���� e�r�-��o��B��Α�Q����k'#�qQu�E���(�@M?yО�5d	�����B�
�>�f���{��<K���B"�LMO�js�&�=ﮖK ��8�YF��51��Ϲ�c%�&j�:�H`��G [�W�R��qZz9�bLn���[\�Yv�'���k�.�d���V %�h%
uX�5�|����J[vU���1����I��>����keT"?�ЊB���1���C��r��!9h�m
>� &�*�&�Z�e�=� �0G��Ly}�@��n��N��4���V���`������c[LH`���1���!?ƈA0Nf�#W �А�qĝN����^��kO&&;\(��@]�;͊W_QC�Z�x�u'JJ������rMUXMOWu(j?���'�dɏ�*���& �8�#��?�?����Q���7,��홚��If	^�J4��d��y�^��f�8S�)��{�yٽ�$0��[�A]�3,�7�Sb�����%XCv�+hq��g�ٿ�*�<�A�����q�ׄ�<�d����]P�'����)TJ�&�ë#_��0L�}���&G�ӑi��������[�p�����޺��2rM f`��p�vcj��E��k��D����M2A���]���D�1�_A�7?(R)%o�;�����$��*s���,����PC����Nދ�尸u�]��2��g�h��v"�lS�x��|~�����A�
M�-v|#8�,yϽ�']$�?���������W�J�@�T���_�
�!�@͗�eX��K�(TV�8i�1�7R���?g4�;�Ȏ&]@�K�>�4yi��'��fc�#9�e 7:p��l��9y&7���P른o���A�9�;�P�jmKIfM�N�²��#�zڬU�&���n�۰�o��pBܩ�����v}��rN|S���s&�5�9o?(]��	E��mK� ����[L��Ά���U�?I7�8r�����A�s��S�3�� ��<�-rE�_m��� �i���Զ�I�hH�ta����%����`�\=��`�XI[A�]�O���o�,�0��M�J�2��	�ݭ��:��bF����Ì.Z��̡�ϵ��|P
Z �G���a����T�=�ۀ��-$d�F!��׋�t]˘x;e_x����\���͆��c�b� A�4��q+��A%�
S>Uwb��̶c�&�x�먹�gOi���p�U|U#d�ue����}�7(���OI�>�L��n����{ũO� �Bnf�h�2��D�:�d\1>c��/XԿ �m�Ջ��|c�������1:�} ]���~Ư��Ę��6�z��ҿ���U�,���Gw��*����5nb��D�u�o����5Ϝ1�a.��U]p�T�m����ϙ���4��g�.�Y�w�U���8�E=pv����*���g{	՛^��s��)s��`��ZNO[H9���_����+���*��O@ᐡ!�M�� �GCi���I.t0�@+�{�J'�E��1���V�1���K����o����aܠ���`mz(�.>�OL,�Ēc��͑"�����ˠ�؞ꍛ$�����������n�6�ܯѡO+&�bA�"���Ao���W8�0Z��~�)����N��OM!��u�wE�wX�7�_��"4�yx��7�%ܭ��e�����5��/���f3�}A��.�Q���P��E,���n�)�-�+��(}�q͗�T�ʻ��7�E�4wbT�v��f�jì"4du��~4�	��o)`���'̯nG��N�F� ��lc;���@����?.cI�PwSs�m�@��rCA���D���'�5Sw��П�x?0�/�F SP����mg���,�P�բ��6�E2��S�<���D��cϾZ���p�\u�S� ����j�t��*O���_�Ž��VHe;m�x�\Fa��ȑu=����� �Ce�����k7�)[�*B<^6�{
g����5�����ҷvfa�3�/ː�0z%������
��g�+��d->f������9��
5��Of𰢒N�.L$pפ�\W��7;�IEb�Y�M���myًu�2s�㕤 ���
 �u�rٙ�
����� "�h&��8CV�I��8�D$ܮT���cA��5'�^y���Fjg)zi�^f}q�dɫq<˸d��kC��+���xoa_c�Xi���X�:n��Q�N��k@q\SE�Yd�Q�Ö��xDVe��0�{z�g�Y� ɂƤ���Z~{��Am�ۦ�׳{A�Ԟ�:r�{�-n�C��	\�@LQ�W��ق`fP|__�d#4��)	IJ�f�
�w%kD�@��N����<䢑Ҁ<���]���uN�Q������%)`�$�d�/ հh�
cݴ�<�ǟĚţ.��H:$o�:'F�2�<�J(/���h�)�2��vo��f���N������E�)wh\r��]F{�*���\�ۂ�������E�8��=n͝���Oqa�ΩDꗨ�\CE���|��8�L��}�.a1�׭w0��#��44b�8ֶw��yYF�iUe�X�@��%�q��d�L���0�T��ݙo�.7S�_��[..�l�x�u	S6#���"Ҿ�a���`B⓶31r_%C�ܔ��b��b���!��z�K�rO��(�\����Gٶ�4_�BĊ����>)��|����u�y��H,0�V����w�Ѣ�>'���4x��\��d��0YW�o�poŔ݅�(�KdDW[�T�s&��b��_�bD����+��r��w�GXm�x�� u6�����`�<���	@YpL���q+�7/��v�p���>J��� D�зs.�vn*+�K�ǐK�xVFP�B[��n)��UMhP��������晖��L��D����8����tfq��0m�k7��K36�~�F�� ��]��SkZ�[�����o���k�R����`G������}�pe!@l�l]ƻc�{ꌡ�,��#��@��e	T@�"'�5J]� [�h:���?����#Zs'�DH�6��N��}��)e#�@�|�'����i �� ��{o�[�B���qvi9����bhI��\����%��������tIw	�5|G��-�#���3�ص.wmk�9 �\R��F(�7�(��@�^��f�<uF1~�f,���|2j�,��?��	��qʢl��Y���Lm������PG������`6`�����XE7SY���~�I���_����x�m�5Δ�BR7ᝇO����}p:�a�ҵ-�ڿ*�m	u�s�㯞�(%N1f��>{sX#]�?Y%`<��d�\��_�Һ�
��29�a5�teZW� B9ϏfF��~� tG@�/�8}����j�.5o�x��{u�7 !�F&�l�!��Lo�M�����w�-M��lP�i"&d! Ý��qbr����`*�*L����T�[��6��^��l�p���A1v�8��tJ�E��-J��,*�p�9\���4�P�^�@>o����s0a��m_�*��
H�������{��W0��?$�e�-a^$����u��oU��g�#l��܀�?��į�s �)@/{z+߿^�2��c�4!+��ِJS]����̧p+�_U�O/�����8�,�ȥ�q��8G����P�WQ~�@��ڮ���A؈dS��8�q\�@��?"�+��8{UA?��Q@M�&ĕ�O�\c*A8�e�nƇ�Mލ��-�}Ѯc�#���SW0�1���:����O aq�K��p3:��U�f�[���d���"��ם�F�
XrG��)1��Sݰ�s�Q�yWǫ�Y���rm�i�w�NW���V�r�7�]`.X��q�>��%�?Pة��W�����7&��� .��4��Pf�)�?6y,�_KH����I���f%�3��L�L0�%$����6�˩M�?�dex]�>�,d�<Uz�c������(���}ތ�B�(\	ŝv�\�~z� O��4l�VЖ>qt���5A�BZ��8F��׏No9�{c���dpU��Ek��g�zk���Vd�}�u� ;��ڙy�".�ed1J�u �i��Zt��+eZ�8qC7U�@�ď��ݛ�|d��H2��Tbj3"q#Ĵz;M�O(bp�(���3�ܼ+sZ���%�����oiK$_�����>6����׷h���L`s��J���� �NX%�@�ʱʣȢ;�1�5{ѓU7�-Ȭ|2c��4�Ȟ�Jv��;Ƌj�o�*���s�L�����"�n�!�����J̷��NPL?�Q�M{	oP��	.��&/cv�l���7��P��y"���5�0�S�'Im��f�p�}-b�p6�&�b�Р꺐��z���u�N�""׶Yܻ	��*���v�︒��T�(8��ZK+ιd��O��2  6_8z��(�A���LG��c��9a@�h��xO��r�h.(X�3�x��SW��Qξ�S�ѯ�6FC�������w��U&�&��mh�h-m.���gGa7x���!��j�)$��#�*�;�>�u��Q{f�!�ܥV�.�K֛:\ �k���<��E=�r#4أc>����P�h�A��@�ʸ�?a�-V�,��e� ҙj�y ��k�i��b�1='mO��D�+V�q�<����Li���tbO�1�9m�7\��H!l4�h��q�� '�^S
�"ѷ/}Fou����8|g�w���E-���E�J:p �קL5��"~�#���y�
u�}W#n�,
EU�����OJ�TJ�ޥ�]\:��6VD��}R�	�0��'�\���lO�G�lyG�L�1+�+E�+ѵ���p�G^�i�q���(`�ԩd:�����Ŵ_p��m	������������?�Ck�	EC�*�������UKKV�,q��\ƚ)$��)|h���n C����R��,Q6����{�8�P�*��#0��?1�Z�fL��Mݑs��M���m!��d����PDlP'(�\��d2�J-����I�T��R�v[Ȥ{�6�O��F�I���n��4%po�1�߳�M�[Fe�*ޣ@�A	���W���,ס��]�Z�5��r��Ԉ"YR��"Zn��E�Y����O��Z������`c��s~�����R�Z���p��?����G�q�]_�y5�C����5����WǊ�ߵ��|)��v���ǆ�E���3���;/���}�~'0�C��@�|�4N���h:�,�er�sS!�k�2%�~�f�c����K�gW�Ŏ(y�hq{tY�?X�T:��=�s~֌-$�}��xz�����$�շ�U���S4�:�9LA�� lw�t~�ĭ?R���go�&�����0�l���*��U��LB
�	�(-=|M?���w�'�^��|4N�O��OV���}r��8h�
�^4�`��޴M���j��y��N�'�����m sT��`ʏ=xH�Mt�*�J4%mK�n��-���3��#τ�٭j�{OOP�M+T+���������7B-�%X~�]�N��������G<�[k7��$&
����	��P��@��n�^[��z�C5�k�]�h0Ԙ[�,r�*@o"&�>��~�^"<w�#
B���U�m4��zs��1+��2o��4/�Ļ�������mw�U-m`*������>��!jl��"����@�W�M��Y@�Џ��3x��U����E�*��qV�������N	}!���ى��gb�;}��P�-AO� �ݬk�S�5HXv|�bf�1$�)G�dSNF�:�6S@ڛ��v�<B�����@[~�	2���qDJ��w�q�˵9��Î\��{7�1q��SYއ��h6�5�A5]&֍Ǳ%	��B_%��d���f�c-�����wc��g��? �J�͜�_�n���|����Q2��cWm���I*�a�%1�3��K� eN��w��'(��Ҫ��2�Q|���-1��Ԥ.�X�0�Y�qeP��"�.���m�緸-�����?j�F��f�Yi�����l�XB��!��P`AZ~�H��n�#G#H��L��d��:�P��d������l��5���q "*�Ht(��*��逷�⤀�M�8~?�k����J�(I��_b��L��������������_Z�96�5UT�ʐj���A Of1��
�ߝ߿z
�6��%�anG�j��Cy3��py-L���Bs.����ԑ�50t�`	�虁������e��a"��bθg�aF>��R>�Q���-��y���.J���m�<����5��G5%3W����/�e\�)zy4�4o�Տ%;�qQ��hȕ�+� <?�UVo�nABwVo�^����m˚@}h�U���;Jxp]ƌ����*���p��GY�;}�.O�qb�#�?����W^�{=�8����Y���OR@dN�gkh�������>K�N����A)�E��/�hK�LY㐢|���d��;!��i]m����`��"N&�,eFh���,o�gyx_��=��|",I"~�p#�ځ� Q�p�܇a�zy^� OG� � �;&�5�;�T�P����0�^+�=;]�0CS��0^5�h��$�U(*�_k��x��@:l���nU�2_U�i
)5=��@�dw/c:1��aɝ10��������<�Ԕ#{�7?!�yR>e2�̛��2��G��K�X�=���o 9�����p^�S�NB�L�B\K��Y���&+�P	�kŶ��@[z�D���~������<e�j~¬��^*�7V�-�'2Մ�쯭���������R�E���9�}%(��,YP�%�HV�Re�}�QXʚIE���ј���q�l��?����CE��/��_�w���:�����M/k.�"��$_�̆,y2�mt.��K��#a-]��1)`�1&�J�2 r���Ј���)C���m��ӎ�LS-b[g�:`��?6I*Qz`.~�Y�C4����5����\�%��)o�a���4)x���9�ڵ@򲫈_�}|)V�2�K�(\�JhV<x77� !wO�P4z1�S����q�ƫ�!	Z0���S�#��/��[����x�������A�nFb�^>�p��u���.����rF�4�$�Rn�?��%6W*pc�2u����ҿ��/�y@�d�ZpDO���B�� (�s4;��dxM뷠^����P\�4�r��P�y� ���txZ�&�7�f�KX���+��,Tyw<&*]�6��<
Y�e𭜞
P�ir�R����k���&k��g�'��`�I���lX	A�k�zڗ�A�|������h_Z��U<�fg\3�H�����X�Ny_�n9C tYI�_y�M��X	R�v�����ۆ�#��oN�̨2Y^�����2o&�H�H\��1_����	j�׃�Z4�g�0��uJ}�M;�e�$�n�=���X� �U�J%���V�-i���?~�gZ�c�4��l���kmGx \Zv Y����u���[Q͟\�����b/�^^������UMnjc�>	���I{��ۻ�K5�v �#/�aDJ��G:{��(�<�|�5�`!��xb��������B���~���As��|ޢ@��j��L]�s���:+��o(v��1�<i���4�^��b$��HT�G��7J	��:�^�t������cD�����`뗞��:���a^4n�/-g�e'騮(�ފ���f�G�g���I ���^$J�A*9�>ϲ.赁�!��I$=�*�P�f�x,=*t�/����{p�HW��`�Ũo<{C�Oَ�8��6�[�������ڒV��1�.�Z��a���y�:������z�l�c�?���i�9$U��1�F���<\����_�C�\p�X-��]1��������w�f��$�,�N�V�Qd�}�����-%�ןWH:e& X-�o9�X�>�|@����hKƇqvvg
'<��i�Ng��<D�H�{�N��|5��Vx."�Z�!�!ƆTϜ�9V�]�{��uU�LV�7+�[��������D�`n[1�T���H�S�I�Pv���]rʰ��bbQOЧ�Rb��W��K���-��m�1���jf�٧�(/��Rj�`3b�2�[��^ G۷�p*��d����m�E_y���W�*�?��h\�	���`�VC���>�	ȝ��|��y�����1P��s}�I]zYEL�~��B����-�l稶\)4vr� C|����Z˽��4�N�w���
{@ۅH�m���$Z�'��i����]�ɴE��"�j�'d�<�	Q��KalCw)��QP�Aר�hF�b��S�un�~�p=j?N1�.l�K�L��"O���M\������O�Q�α��G�
�J�tuh¸e����˺�k��>���ֻ��I�Ή9���נ	F̄L�
 � � l{����[D�abe�=�? ���l���]���A�	�/�Ͽ�ӹC��!7��z�帮"��J�������,����?��4�|Y��1TJ;���#��A��VX���=�(cԋ
U'���(z��7�����,5��%R0�AU�0�kF�< �(�i#�LhG���C
�K�;�Ϭ�� �W�l������e�9��gF��S���MT�"{���Do��I�
}h0p.��Wݢ^�J��7i�I��$�[����\�9�}>�`���-;Pf`�I��p듡�yWa"�L�_���6�\��v��'�#��%�����C���{D�ǛKd��ڌ}��� htx���7�Is�s��|*�g�,�m�P�����!��L�:������eM�L��) �~~��l�'+E�c��o�7��4/��z_�s���$��0�_�����	ee.�B0�{)�σ����SpF����B�����ߟ�Ԝ� ��Ȥ��赙����&��&����\h���e�J�n�Ep$��79>�qe��cC�r7�~F��9V�k�]��L�kDa�lDk,ŉ�6=l6a,�h�['h�`��2�C֡�`�Y��n��ȩS1X"�9:W�	�HV�}�����7�xS��S�̷Ws3�;tk�A�`���J�$�#f+�R�XZ��mZ�k�5�hР��7�,5�`�t{�9է>�T�.�le�:��&Jk���Z�� �.�~�+�F����m�*=���2���B��S�É����K�O0=��Q�_I�$�����o�����W�}'�=���j@��n-�<�	,i{r<:o>8�lֽ�d�z=R�[q���-m�ʚ�f�ìA��<Yd�2R*�8�z��l6 XO~@�x;"�{T�����������;�\�<:�k����D�I[ df�n�?�ł��)��aY�x�:��?+!)��
�4��b�l:0`v�J<��0)�V  E�:��5%�y������R�#� �P�����xZ����L$ �<����+{1@>�ׯ=�w�Wo�*QeeIp���Z�$�[����(n5�&ZO�����Ģ�݇A��8�98�W�,�3��T5�	�}��Kr{{��r(�� hgkR�����.�YΨ�6�@�[{����޽��Y㼂��{� �BGl�Od9���A$�)�B��@N������C��m᳭=��l?t��|���f�I.��x<��lW��ۦ� �[��r������6����/}h���KxU8Q��n���{�T=)^����gl��Z�y�+�.M�d4��՟n˵���1�e~U6�Vhk�����g�ޑ���@�fpkse�U7��1t�yO�?�0j*��Ϸfn���=򷶺k�u������G�z��v|����m�@̭`.��0�)q�n����I�=�!m�}�"���c]��bEts�6��;]k�l�,]�bW��	���T��0�M�h�ߤ��c
�>p����Ph����n� fA����uR.KR�s��+��s)D�E�d5l��ͦ������[Y�v���$�\���o�!��'�Z��Ӏw;� 	9yoi?�.�$�H0-mb�:��giP� ��*��9�˴������/��ܵ�_5�5IM�]�U�����x:C�u4Sָ��Ԋ ��;	�7M��u
�a��W��x�[��c��z��;���B_���Y�N���(��� �";]Z �h�����*�`
������{����k���Cc(.� V��� �L�oG�3@|���3��U"����j�[E
pC	a�D�U�m!<��?�;�*l��N�\;,�Jn�:
5���S��X���^Dߗk� ��\N��
S��r�#gߪ@\�66Ӵ\��ZG���bG���_�nD6��"*N�Y|GB�,UkX+�/�6���|��Q��yw�$A �`���m^�q��m;��e���c��w7������_cO]���lb�:��+�6�����b�lĩg"��Ȱ�o9�-/�oǥ}c��������0�χ��Iܥ�Ђޖ���L��!(澨2���/^�M���a�.�����d�[�L����zR��sI��侟�,,��[[!#AN���i�c.G*ǐo'�p�+�i ��m���`���C�*�*�����g߂e�/lG0rѷ�ڎDAk��g� �m������40�h�-I#4U�s��s��t�od�f+�-�dh�u�d������^73??���UIF�i�(�ަú�+/T��-����8 3�d�4��� O��q1B=OΈ�ȲT��p����v�V���21m*��n5��I�zl�زܾQ9�� -Ù��H�&xS�t�&Fx	�tq�V��=9=Wuo���{A��G~��ݿ��@�Y���EW�gt��kvo!�/��a%�A��Q*���/�t��S#�8��*ϼ�8W0�R�����k���u�d���סB����]�����a�B�~��_!b�~��u}�ūT��M��l� >j[�ȳ�x�mo�|`����<�v�*'�<�d%����州�io؞M{r�=�;�ҋ����7�wS�-�o qi����c*�s1q�I\��Ŧ���t@B�F��-��wa&5YR����&t����[��H*�]�I?���D}��xÊN�׫lƟ��+ʕ&����]0�KBhJ�Ă��+M{$�V�`N������)�/��x�υ�gC�yh3d--q.�ΠC@�/�~�:�����D%}� T��i��o�����:��귶@��V�R�A�D��?k��]��d��
_I*	I��U�@qD'Q
�ΥQK�� 0?�'ߡ��w/R��