��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,��.��̡�+P�FuX��d-��N��$%�I߽7>wN����u�]��j��ܹ�Ucל�|�=í[~��k�5�P�ؐ��T�5�����#�p"&�l�z�Fr&b6��,���Fԟ�Z�_�X�;���93	�����Ǘ�M�~���٘�2�c�D��������f� 3łߥ:ա�;kv��ތ(�}��r�{|�Z�LP�����!�Y{������I��܊7Է^f�L5�:�	�͎������W&��b��wD���Jݎ�IK��et��1���Lt�:��6�Ui�;F�o��!b��\#�Z��k!�Y�#Ao��U.H����Ƈ'U������0JN�]�[�萙��5��!M���@gb�t2�<���#H���p��Z~�5�;�k`:]�@9��!�}��\��'9:���Xz���r�٫�{�$4ʄb���V�]S6�$����3��\���e~�b��cu�ӃU#Z�T~��8�]~R$|�:v��E���Q��4���G����l���>�I{8����[�>�NVf���˕7ǲXQ.�4Ę������K����<���V�����L&w�g30���owu���ױ���y�K�ȪP�����5쐖�ױ�qV�����蜀o�0^�egb����ŕ4��`�1�7�+���A�,����1c��B�M������e��WW1��e)�m"}$VzF���,���E��a%�����$��=��Q����so���SrqҨ�����II/Zlo$aN�)�,�&�o�����*��j¿�wP���QDФ2�"J�1�I���?�sW�k�����v�*���[o�����֐!��*��5�W,�|�A|�)N�(�7}�ԋ�%Kݕ[��<��h� ��v�7qV��+x!b��MMLIS��}{[���.���Uds]?/ucG$��e���Z[�s��N��#���Cwϳ��r����]��lm�u�l��c�mG��0�i��,�C;�-�WW��|�ځ���Q�8d�N�%��~�/<�'h��]�m 	�:�W!�7�k�|-�*Фxg�
�J��lf�,� X	7X-<fa�2I�+�Z�i�����Q����Í�B��4���Q£y\��.z�C�֛��1xI͞U�ʹ�-K�CK�6�q��d`�h�-�t��Z�V�21h�����i�5�'�
�9z�׮G��.���Ց!~��VS\�3xВC����/�yvI�E���T>��׽*eK�k2�臔b�=b/�He;Z���i��f�1�
-�D�9������-�k���Ց�������)p�Mj$��;�!\φ`���-gn/u<Bf8����fLy�e�P�:OG������Θ�]�%`n>�,l��p�rM��(�:#R�/�E���Y�z?� �"Xc}��������zy�F�,q�����'�B_�:<����]��Wj|N�{�R�/Np��+ql��f�x�:?@T�M��� �:�Ơi�qî���?. �Q�p'6�h�<ǅGW �{@q� <�3٤���PE����/��J34�NP�P�c�u���,Z:�5^)}�E�,?�\Y*w+�j�vib:���A�q�2M���m����}sk/ː�`�Exm*N^��v=q�.��c�W��R��ZyS6��'��)���M%��ܨ��^<g��s�܋��G+g�|t:7�%�X?�r�����b[�\����*�5�tŃ4ZY�����0�*���IV�st��gC���҅zrL&O[L��n:h���Ő�"ٹP�)M��1@��g�\���ƌ��	PT�ј
������������A�x����C"�+�Z�^��;���4+�"�����>Jʅ�i<R=�op�/�\����&�	��Պ>�
D��O�Gi7J��p1@)d��uO�6�I��n��}���j���c�9�Q�sKTI���0�':�u=�j�|H
��ll矸V�|/�*�~Y��jHa��0 Z�Q	��/H�����4����w�S��c���lF ��� ������5�!��m�`d�}ಚXw�I:��0f�#�D����q?7$��a�v�I-Ί�rBf���@�����X�JuU+��9�|������i�L�8S<a/}�h4N�����:1����:��&�'Hr���F($�>z �����`1^l	���N��隞���j��m����DB�[��MH3�A��[N�k�M��X���D ,�8�5�15�E-���1��/5�u�䣻���͵����{m"M������:���!q=�J���J�j'n�;��y�i��k�=[R����#(��9|�yZЇ�SXƳ���v��:�y��\�"�
c.�j��p�_z�ǐ�$!�F2�0"!O�G@[��|˶Ch�́�|<}��������br� ������q ����>L�##����eg���FV�h_wc����A�wۦS*��� �����ۉ�w=tƱ˭8C�gPf��Siv[ԛ�u�0� ��