��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����Mڨ��˳0]��?l
�4�!�ߦ����"�p8"	~��kB�J)��NbM�L��\jO��#y��r�3wA�y�}�S�{�����X�.m�lM(��R�g������B�*�NV�X-?����$��$�3�s�`;��y�@�u�ߗA�R�|�Ԝ�+�)]f��������҅i[^�"[��t��00��6�ĔR�*[�]�V�t���9�c%kz�Q��*N�| ea�z ��@������mU���h�$}���~�k��'C ��� Z���>J����ׯ,�'��3@akCc�U�U��?��a	6S��K󊀧uh���Z��&���9�+�)�b�В���ɀ�t�]z[��z�/`� !g�!*��P�����I�<V�� /o"�����@�g柅˳���.���5����9�i��)�!Ҏ���f8�vh�3�Z��ZC�:3Ϲ@�+��&�Ư���	��������Ϋ< �����"�����!b�'G����Z�!�R�l��Ã���3�����y���H�>����/{���?R%|��n6���gJ�2!b/ΧW�}�/FM��%����� ǜBk{�.�-�ّWz�*J`����'29�05�J�NYŪԚ��N�F2���������q��y�-Y�	����D�0���7��%��,�-.�O,P�y�w	�	�JT6'�Z�Ҟ���4��\��י����Ə��g��y��E��q�"�ӊ��N���H��`����=l�r�Ed�tP\��� �c�G�����/�('�'˷5����+��3]ʸ�:xõ|D,"���V�d�@��^Nm�D�dK�+l����E�ȟ��_��O�՟	����ȢM�6��������U�²��;偐&r�+����q���_j/�/3Ew�?'�Y���7ϓ,4���W�X�`]���eop�B����nIN�_K�����+�-�J��^��8��c�.)��+eR\_�-�/��?���}��@�|�VBp�zq�4���tsT������wPφ�(�,/��3�3~����]4�_x}����M��t,�Wv,�,�t����#���ιXz�^U��#|n���q��LlW�'_�@aQ�Ѽ��Սu�7�q��"�u$��NɌ;����B>:�?���3�
��uk�iz���u��`����sK^��b�ɦ�����u��8�@g�!0�U�p3PR��O�����=8��֠����a��~	���j��LX�)'֭^���ց6f�\T��@:�EޔR�J��՛�)h<�2G߹w٪�}�&�niԩ�������R��0x�;�-�:��\z�`^�7�zH7�W�!�~����Xe��+�#Z����3	�鸵;F�N6-?�@%��ݸ\�1�S��R��b�e��
�Z�w	�8[YA��X��.kڪ�������q�@
*�qT`�I�f�8����cAC�-��gу�Wi�h-���9��	�0��!�TN fE���<�G���{�5;�<q�NĨ(1�f*麗dQu0�AH]��WU�x����#�!^8Db�])E��L�U�D���y�2<�T����~9�u�3!c��w<�#���f�Q`ۡ7Q�SX�Ujd���OX���n�+�K��OX����.����׮�#��v�!w(�j�o>��]�D�TBV�2�� �4�y�QDN��W���$%���w�4	A���V=�.Vl�bH���#�r�p��y��zp��
-��.�����ڢ��Ң�����ENm[��Eo�`#��
4���r_��+��ff�y�2�X1���T�Ҡ��ҫ��V)���6�64�g�&G�`gY�=��o��w�켫\�\|0�^��Sث���w:�F"w������F���e��_��$ȸVA���y1��X8h��L$�px��')�rq���3�%��sĐh+�����p^*��=���{���~��Q���^_��L����
��Ytȳ^������ �6�6C: vJ� 8_�,.�}�j�pXޯ���o	:�[՗�-��hL.\Q��2Ny��\@�=�f��[Đ���#�ApW�0x��4^1İ�C����P��J4�iA�����y��&_�_h��ץ�~B�Y���fa_����M�j8�a��1�o^ֻ�)�]���˃��א+
���g���/�5kT��s�y����k~�����*�'�@M)��b2�F��X� .�o���:��D�DX�M$��l����KeC�����!}#� �'�u?$[ފrT ����#?{�.���ò�������{�֚2z�^쎼��#T�~[i꧔jw�jq��NSr}�f��_���P��h�����\���a��@�(�X�(rތ{D��-���)�MRсl5�֕��d������]Fio�?+�'���,oE7�l*N�