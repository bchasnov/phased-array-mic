��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�uwC�5�b ��ϴ�	+�
Ct� "�J~���z����<
�����'k�z��ߵ,d�.��Z�Ӝ��2�x$ҟdL��h��ʔf��#
����;�;m�ȋ��[F��E� &'{=u�3jg�b�)��LA�u/5{<	��������
|z��ok��n��kJ*CAw��� ��T*��1?]�Ʊ��!��p�Ӟ�3�8*-��(�lg�p#���-�C���ӽ�Μ�I`o��hI����(�����Y%:I̓��؀w�4��]��NL?�yP<�] �WX����M���:�C=Q7��L����C��`�Ӻ,Yk2��;��K����U䐶Sƪ���)
^[���M[�aW������>�$�q�S��.�:W��ϲ���k�?<:�nH��w��.�/ �RyЋ��Q���传�	��p�ۊnMrߗ��Hb)�ǚ���=#Y�U���zI�Z���6p�3��9j�aG�_zt�~���I��HLb�6[��B&4��d�B[��n�n��$���~r8Ú,_���x�V3{�D�nf�D�j����ZV.|dd�<�}w�M|��.����q�G#�_S?���sւ�)��Z��M�e�� ��Ah�2ES5
ƍ���O�T����	<����94j��t�Nd����t�S��jz�Z>K�1%���A:OP��6(���2�.q�e�(Y����w W���&qY���D=�j��886��֞8b��^cd0[��kޡ4=�OV�@v,�j�"ǂ���f���$��Cy2�VL$���j�:�g�V���j��b:�$��k
[̰�(�a|wcs'�����8�.R��-D��@yd^L�P��L�-d��7��L&Rn\VZ�ĥ���nG���z�[ �D��]���,���$�Eg:��i]3[ARC���t�8L֨s�+��$�"y�[�q'Ǌ����%��^Z*zg4a��<��A�j\q���� �JK �|9�W�ia�bY
$�q �B���|]���釶,�ꎤ���۰�۶q�7,�����Ȏ{Ӽـ��
U�+؋�H�&i�[�Ћu{���d�.���4�Hٔ�?��%G2� ��M|��u��5�����۴
��w��7��f%E��P���s���L�t"���/'He˥�r�BH���f�G�}�M���Y��:�#S\:j�C�JN���ʏ��:B�3�Hd�^��suR�[65����,��ݬq��WŽ%���@��/T��"��e��t�eX�9I4������jA��`�Rl�q�?�������bp��^GVU����Gښ�*Gi�~H��_�
Ff�c�'����鵨�r��N�#5��|�W��h�	���������x):A�|uj+�-l܂%�h(�cJ(����gC�d��^���y��ֹ�C�d`	���eC��Ay(۾���>��~@ua0�}�)�#_7"Dr.>~��xPˢS�m�O������\��:mh^#z��m&�xc�Қ�#����b{�˴���GǓ[%��-�#���H��n�^$��c[ʑG��8"x���?��A<;ʶDs�Ɖ��� �`"q
��]=�Tá�޽�l����XL��h�����vϼ���jś)������Q!#��lJ��p�.u�}/q�7��f
"�z��H���K�$�ט+m�y�kZ�xp��1<����@>�Y� ����G㽌1 �]d�G��-�����*��^��M~m_���dO�U�l�BԘZ,��j�$�Q���]�T���YVF�@'���=�S��R�`�3,��2!��i�~k�«\�~��2a*�-]��ۅ��!<J4���K�ᆇ���3��]v
 ��xx�����b�j�k�����'1R�Y����Y��`�05Z���#��?֩7Sj� 93_�.zs������Y����c� �p�"�g~��u�Q��c�2�<Hۧ��2���"�qz%����Fa!m�@�5-�e�+V4��K�lvF��o����烕G�DS�z��V�^;�F��j���K�I��B���/�0@���Oo�/������*ݏ� �(��S��ī��	dv�8>�t�d�Z�%;7r���L�-w��ygg�!��KW$S�|T`�̸���dv{���u�:�l�<)��Rx�-��6�.-_ÅQ���ߘX��کG��0�K���w7��T�*
0��1xcxc�6_�R�!�X�r&X�V��9Km�!r �π����!�����À|�t���E������m�;N�f���8+ �ĩ"��1T��p�2��)5gXb|��g�Vc�=0'N{��D���)�%r�8j���no@�� A�0?��Y<�P�P�\��q�8��?�Y���#��.v��F`>.���H���xkU���9���jd�	�;�㴚� ��S���H�ߙ(y|)̣Y��}���x���k��C��9�:���.��`�Mͪҧ��5S�P4[�if��=:���{n}0d <� z�0������d�ˢ.�:3�\�&�gt���g�q�?�J=:A�� y�P&ѣQ�I������㞱��:A��F��>pD̯'[�y��I�Z�6�`�F	��TbB'Q3#

f׹ᶗ�v8�Sĕ��E�����{��޵���
Q���өMN�8i��p�U�O�dq~�k�
kҹ��f�'[ފ^-|ȣzPN�3b^��˳�{��LEӻ(���d;>p�r3��G�"ގ3�M�: ��LӦ6y��h{]�9��G����	�3�Z#Ł���������=|Ş�G>�z�:�C����>f��PZβX�
�G-E��	'=
.��e����s���h�:}��J y����Q� ���*���o�G6�r��W�%���L��� �߾�W�w%�����!\�3�))q�y���6�b�������O۷�BpT����h�!��s����U��[�h��[�W��pWwmf�{�W�6��3wv�����^(`e
>}�0?�r���\�N��LX�_*]��;QQNr�H�j����Fz��H�8~!%�Om�
��>���-`-��T٨�$�^��a��O���:#�w�)�T�=���Y�:�4�v�V� ��)�օ�r�Z���&��i�\mZ���BN.�Z�֓�]Vh7��������Fk���.�?��Z@p�,�1��}�x�������5��
�ν��0ݠ���[*�<eL�4��r��vڼ���K�Wc�~��������C��v�&����'�qo��I��IL�ıby�j!���V�߉��o:�@g��
.ם8>o�Ʉ"T���X�w�+0o~[��"�vU5�bc;�Ý�S�Y�K畴K�����4M��u�/�*��
?�� Њ��O'�S�s��<��'�K
��rW��O��cjW���B���.}�4�ݤn�{�bN��:; ����9���ni�"uK��k��9ޕSx�@�a��}�pXl=�չ�,����B~�	&����b���$͕:�؂ٷ�
դ�e�OAA�DA���[�|�I]�=�n�=16����b����Æg/����:�_qw�6��{|�����<9���*�<�I�ߵ#'���L�W�iy{�K[�|T&�HEԁ�B+�)��������EY�n�v�+��BW���"&�]m^��� � #�Q�Yj���d`<ջ�PD�j4ǎqm�i� qG�L
���K��<$�W@ҽے�h���Ň��m�;o])�%W}�&Y�S��}��%6W����|�Q,�Y�5~�O9��l�h��oD�����߅��"����z�這 �+W�"p�tw���Xs.A��� 3F��.P����2����<�t|??6+��� QUYc_����N8K8֤t\�T9��E�R�&������/6��-6I��d����#Acv߽�{�T�I�Ҳf�L�1.o�5w�vŃ/K����P��Fx��t����f3'��=gD��
`�ʉ�o]p��d{��!D}�+@;R,�IKFW%���B��h�Gs��'���4͔��+u\v�?� �n�����R)�֎̻��g��L�i&�Ԃf"n�i��~�1��d�������v��+	�s�U�!��RV$/+�5��&�"W����䫢zC��я�7���`�a�/�1ˍؽ��z���t$͇�RrP +x���F�A1Y�f!�g�1�	�@�UU�0ʅc����3	wc458��ڡ��da�&�򲺲w����� ���ͫ�Y�PR`5�Ϛ1w���������u�QF������_�(l=U¤��x�'[�K&mVWq`���,"fD�<A�iY���6k��+�,p���.�Ǜ���o[e���}�Hz��_���:�p��������X!r�b/#x/{��ۢ�CZE��\����<qm�TC/_6�ɽ
��r3ӧ<g實����[�p����E��F�/W4�i�)X�,f����n�^����NR%�~b��0/ӥzN�%I�	�?UN���o ��y�6�L$/8���"�O)��d��@��Lc�GCR�bZ�E&@�"i��H�O+s�M?�}PQ鉔C���:���"]r%��!+�X�e�R4����f�F�&�]�7�������)� ����]��p�F�;�%����A�Wz�C�3s(�&J:���yR3��h띵mJڲ5�h��+�EJ���ר�6W�]�	G)HB"�m�8u|�P	GYfeԎ
�T��o���^qPq"z{���"�B����G	o���r��i�ލqGR��/�*���A����),���+����Ѯ�P��_������=�j7��n�C<���c���_��Z��6�ק(t����e��y�����M�V��khj��n�h�HӰ^��(ډ<*P��'�L�J�:߱��i��O=԰��O�3`S�]w�����3�(�5�;<M��P�:�y��L�q+R�#lэ�<��g�,tl�3AX�8:�Q._$��Lۙ<|�e~i�YYQ9����}�0Fq6�Q�C�')��`|
��6�JS#���^�Ɍ�pj@,�xX��+T�l�]�a�C<>6�����/��Ň(YY�1�vn�o��nv����ݚ��V��};vT	s��`5cpWB͐T�h������zi$�v�nz�^Y��w�$G#S�	�ӿiib���9ʔ91�uϭ��I�BT��]NQ�xLz,��O��}��k�~[tu>>�Q���)�x����`d@�tS�:j+���q���a"����ǥUٴ���?X5�\:�+���z��s�fb|Y�u�2ǂ�X~gɸQ׮��� ��S׏��E��2�68��2Q�ҟ�9�l �;�	A��w��N'D`Z�����&(�����xf��*��o�;d�"p��E�K��W;�C�q�(��S|>	I>f�YԆ$y���t2N���h�ܦ����`��
;� ō�����U�<w��;��E
�"��H9k�KŴ|e�� ]����ݧ�;D�p+�^��_�O�C
�w�4�Cx#+ }~*iMkR5}.��V������&\��e�0�ٟ��8,`"y\D���+`�&�'q�bc�e��ٽĵ)���Ǖ�]��M��%cy �)M���)e�\QG��9BSk:�����32�X���Ii`���>��]p7����>DZ��&��5m#���O�c�OD�>�.͍��AF�;C^���9�y��47�].�JxeYmŪp�A0�mK����%�)ND�2���=�)���U���>Ic�6F��g/]Y�}�^�;:HfĹ����
�4�j\P�&�)E�Ά6~�ŨWB�߽ l�ͬ  �X���%���́�n��
��v+���ߧ�ʓ��z"�y��%�J�{�iE_�-˰?.�"Pg�$Fj���e#]���v��8�Ҋ����:�=�L��A&?}�#7ԭ1��`���	Z8`)5"�q�kO@j������*M���ݟ���Y��EυD��݆�A�_�,zRC͍"a=�>]��������4Y�|/� z)�?�C�'��T�Ӡ�{����d7���/�1���녆�-�1�M]�udx�V�	�:�{�ȪD`��ꮸ�-y�Q���O"N)����TP�����i��i!\��8���Yv�$�\�0��T�2d�+�H�ؚ��[�S�n���������U}����O���e9�����Ǐ(f�L��ˡ�-�ɐI��g�s���!���������]-�(}����+ǆ�?[��*�n�c���8�,��xt]_r���;���~������a�[^�����>�8_F�V�uS4�͸[��R��[��]^�c֨P%�PH>F��@��3�CɌ��t	\�Q�s|8�t0A!p�b���v�����yy��,~ ���S�Nu��LA/��e	�M���ݩ<I�$4�k������i�����b�"/k��,���6|�F�-(*��(���1�[c�٤�b�&mx9�Y[3XMP�V��/�S�K������Hx�7�����㞇��v�4�J�n�΋S�k��$đ�*u��_���"�[~��tXd��咥��p���p�Zm�������h`��̤�'�쐫Ѫ�"y�)�Z��TK�kSN`�ҕ��Y���\.-��9�Q Z��z
�������/R�Y��Z* ���~ub�ΟEֻ[��%�ޮ�v�,��2��@��HER%�<5s=��W;��ap��8�0�4,9]-�˯h3�������w��Pˡ�H��}�6.Hu%�����<��Vv���b�$䬥�՘J�]�Dxޝ4������k���m���#���tϱ����V�Я�.�}�]a\��ǯi��(R0�H1ʏk�;�+����)BOG�B�"����)�l�X�H�(Qh��r��+���f"������8ȕ 5���&��F*�n�$��H\!@�˘Ҧ��7
��)1�b%Sah����*�Z�&�?��[����+����OW��b��q�s�����}��6�T�4-�mq�y	�⋊�Cwc��r-�ư�8�򀘵̖�������_��HE)�is�$�`�6_�υ~�Ժ�ovŞ�MO ��i�Joc���<�W8�� �ٱڻM݌�1��e�e��|�<�ȫ����%<�*��gAf���hI���NI��?$�n��p �:(�ŢC�����)n��`�Ղ5�T�v~x���?a��c�k`+Ȥ��џ����P9
1�xmk*�=j)D�V�Y!ûJ�.�L,�Z��]wG�t&Ga�w���Wӕ^�G�����5�'r'�����Z���^V���o�U�B��'�t�2���e>,H����t�r|5pT�m�8�; ��oC�~��|
�/�U��ƞt���!I���0v~p��̷�B=�7�fm�w:�H.f��u��K��%s�<��z:�̟a��郎&�ݝ���+x�+��l|cb��~fد���v�7��\�1t/(G(�捂G�(����-�6�K�E_g�u�돉�?�hw��5���u����5ڄ����{s��@2ݝ���E�[��_���JtQ=W�g���bZ �z�����"������� hȄ���"��n��-��ܦ��e���u���F�����K����8cF�^���UnE�����1m�D��J@M����_g1����ۀ��,�4�/�%<l���c�-,���1X��GG�P�&�<	���\�y���,�RK�S�QQ�����yB]�X+�L�gK�o��~.k�*CI�=`��FX@��psP�M�+�쾗A_�{9�\�1���FM��mG*�7(���[�|tU:|��&�,]!;#h���' GM�02^��W�x#lWN~%D�5/ �s
t��B�E`�,|qv}Ɗ�>���[�.I�q�}��J��I��^n劣�zP=X�F>R��P�r۩oԱ|yn��I?T}��L�T��9��IaB���h���Ѷ1&RO���t������Wq�B�8�-����@�;!��
0[���������X���֗�B�ڇ��]M��^A}��'���b(�@�uM��	�SJe�Ǟݪh;%�6��2�U��
6���\t�A���G0pV��]�\Q���1ZPT���.�l�'�Т�E�u������`��+Y�Ӽ�j1�	���=�j ��K���M/@��۾��u�y��x-��Q��[6Q�s�µU����:0!�m�k�F�m{כ�-�T��~T�!w�x�(<6e�LR`>�.�}�sV������ʀ��L���T�-��z"����r����@b�<�U�\����"��[�"�x��N�� ��Մ@+\��}�{s�v�j�9-��S`�/_�:0:��L|�A��Rp��.W�v�AN�q/r��N��Vv����.r���gI嘠�;=�]b��<>A���yϦ��&�Z��;v��*���R+j$n�Y�y���{@�l�������z�br�2�l&���D^v�3�a���"�������1�♏��?���=���˗�U�5-�b ��y(��l���F�<�R>������aU����b����u|��6���ۚJ�>��D���2�v/�֡���c�Yf�-պ&í��lA+�s��yo��ROw�脩X�*�7f��������
��=����`
O1c4���c�U#;_����8}.��ng	o8G�D�~�C��V��r'�*�w��	�	��2�fTq4�F[X�A?��e9�u��5o���#���kV�n�F� sZo	�q#�7?����P��`��?=�ʜ��r@#�������؇�?�y�#�\�VB�J���*�!���%�*�ۍ�]PG�-��n��r2�~}o���b���XCyJ~�
lh���G�l�Cۙ
&�?=��sڜ�@�g呙,���x�ٻ�eL���},��?���k��ʮ��-�Y?�V�<z^�{_U$���t�I��ld�c1F?)'Jp�qAx��k ��c�#��
�_����U*��+�l��Kbq�<CJ1p=k�������g�j��Zt}��J��]�N���<M�_��v�Z`j'pӎC����G=ǂV�*n"��I�-=� �rX�aA<s�>���N/٪��	-��o]��<ބ�K��^�����dXw��v�ܻ�x��Q�Js�ӯ�'޹S�o�bcGn�!1�yb���N�m{��S�*��偋�U�y��W����!�4HiLlBJ�\tN9��?�t���cr?��v̆��{�{�ƆU�\ܜsF����>)]��,��!V�M2N��ʋ��%�Q.3){��
%��Z�S�
ă�T�ղw)��Ơu�R�d�P���dK��ⲛ4Ъ�W�s����F.��/X���r�z����P�h�|C(��4+˅H�h��>�s���?*;�ͼB�քϪ��e��F7O�-t9�j/�%��m�Y�d���n%�0�HÇ��CDw��8nzׁ���_�:��P�W.5�O�6o�1ܡ���A�Z����%�I�>���*`�b����tO�A#���1t�_7!�[�"8M��ُ:3_����	�%[8���?t�d�sPY �D��7*�o��aS"���@�۴̤B�����0:ωB�q.agM�(�J�e��V+]s�)X��ĉ$�s�ؕ�3�h��È��ʃ������g�D@���1���nm�,a�[k"��	3Jˁ�	hpԣ�?3ŋ�z���'(��夛i���TӍ�f�|�`��	�t���T;E�3j�;X�C��>S!^k(�m�����4��h���	�~�O���N�GS����W��S�	?�B���ƌ�WOk���g�������G˗	�i-�J��>oEs���tE�K�VR	|������W��F��'q����R,�Ύb�	�/"x�PXB@
}-q�β����ȫf�����#�X�L`��f����`A�ɱ[��WW�����ݫ�Y҃������v����ϧl��U؉��n#��p G�e�kI\ט���+���s6�q(]����K`��[���cH��O����l�NC�f�' �f?�tw��?�D�vU���я�@���@�@uN�\�����0L	2ˌjK��,�'7�8cI5���濜�u3�Q����ฅ��nw�?�oy�f1 X<�m꒑7ʪ���sʙ�h�
d���i"�VN�Q�hp@���T�?�u6�̮6�e�xKY �=�쀫LϷ�=��А`����:T,L']�U�`7o-Yʑ�c!����fεv=�7���k��g����
��gAϠKk���껽��s��p�R�2�UO��~�<�N�}�y�#���{�#Y�A�*'ĩ������y�vNV��v9L����u���Z"7۫�6��?^?û�w�@��$��;otI�)�*k?�6	!W���Y.��oY`m�d�H3�
A��8��O���2b��a��9��I}��2�tq����"}��.`��V�����r�&T�f(���$� �L���Xx����0��#�nR���˙a�'��'=�	�ث��/_EgD�lp�RUA��3�'���;��x�����m�=�����Ȕ +�5� ��N��&2@�k���-�`��c�����Ka���{��2���=oArj>&��憼3\|� �k��]G�ЦO �Do�M�>;j�C��v��3�SZ����Ąf�{��H������k�wJX��XΙ�������-�֕�q��>�w�k��F�HcB��v����MƄ��]�W���Kд��W��ޛi�Y�A�d� x�.ލ�xe��/�{7�5���ݝ��~TU������N��~��D��7���7,oͩ�@��4���	@뿝��m8�`j�7� N��w���b_��y�`�5��N7��=l�a~k�H�L����_�-zh����o���;������w��+����k	��n��@\Q!Sq�)ODm R
�bf�O_ǈ$,%J��]j�L8����{� \��Pj�]8�5>D�r�LH��q9��|�i�*5�i��^�yN�sU=S��8�))��ۧ�?�+��j\ۣ)��Ĝa��(��_�Ħ��D����W����3��.��Ua���Ќ��B\����*T���qPy�n6�^&y�h�����P��D�/�v�'�ǭK��h�I�7K�
�����ԛO�_�Cm��I�n��A�)_���t���:Xe�eH������K{�oln��ڿL�c)��Q)����t\/.�«Л��+��I�m>���m�,�l�K΃��Ry��c+S&��g8�х�1X�TԘ?P�����ʣ]�I�G%���#�;��̺�2�<%sgk B�x)|��Z5:z)��R>�k�j�>��0{�9����ߒMz�S�	�9S�Ϥy����>�0���1_� j��~�F�{Sķ�}��r�w-/�-��#S'�<���Y�V�$���|~i�#�I�2���S:w�Qx��Eq�c�K�\!^&��E���N��5,$����ϛO#��F1H�� ��6:V��j���!�/_��Ը�J���Rח*Ɔ��9���?����f����d]�*]��R!���O����7o�o���48!|�Ĥ�EC`��q�v���s�F��P۳/r(!$U���D��O���sa
(aKӲ[~u.���mҹJ����=���T���.��o�4�3|T!F	��p� ؆e9�-�b�ۂ#H� Z�h������W�'{�C���1qNܥ&��EF�� vn��,�����Λ�Q@�Ӥ��ĩ��J�Z�% �D�త4�J����i�kFtn��Z����������3ś����z9�����I���� �%���H�\S��K򾲉E6~�0Ө�B��C�K�6U�kK��L4��mI�R\�T��w6��rw\X�m���+|*u�sm�eu"w�J¦]RP������0:����ҵN�㮯��b ̥���&����<�S��,��w�3����dLk6���"�*�I�8�&	�<�0{�`Sɾ�p%�`�����|����x��W�08�G�Yr�*�-��{�4�m��)rR2���R~���>�����t�-X8p�pgJ�"��Ӓ��"���O]�<��d1�/,sD��L�����ػ$���_��*���u�nS:+$�#����K�Ff�#p�z#镅��p?T~��*|>;�ZHrV�[���![����u|_)W �����W��0����|dX���P�ۿSQ���:Eס�=^��Z���&�>�?;�C��w"�Z��0f��g�������w���CV��N�/t�����F����o�ņO����4�W����4�ϥ��s���:E	�� �A�_�<�@S�e��s����O!�����(S�&�a�0T�2O�-uU�3t�u�2pd�կ^�(���
�6(P�I\~���Hw��bjJ�C���c�c&���:��D�D.>�r6��µr PoE�?��,Wے�/�7�����)Q,�?A���%�}?��pE�._�������If�[�nB�`f�̉��6����ͳ�	n�|z�O#�%n:!"����0����T��f�ti����+���x�li����솗R�v2�?�&Ӂ+ۺ�~���T9��%��\�������������u~}"���s0	��)����������N�����Ҡ�$���u�AU����&�Pb��l��᠁�Ee�4
��:m\�����S
�>��n]W�Q���
^O�y�l���6JF���*��qLN��\=�WMHTT��k7�چj���ֳ`�8^ī�<�����Df�U��s���'쯪�B�Ű�ů��i��~���ӎ����.��.1?ڞ:�)_7;�f����U��� G��������@�BT�������A@[�VP?��q�2�-}/�>�Is{UD�j���,Rqi^�7ݱ��x�\�8np�k��71KҢqh	�#M�)����H{�(�w���:	���>�`l���S�R���li#�=��A�p�8�]Y���ݽ*�m�\I|[�H�3�E�&��"Q��m	�uª�G�x1�E��E��U^��=)�%+�m^�o�"0�ƒ���:�4��;��j�5�	2'���m&������4X5�����3�)�.m�Y+�f <�b�o����
6w�Z�!%c��e�c�����ɀ,͵�~!4p���j�,&�y��� �O���Ð)�L�3��BV�wL����	�ŋň�y��B%&k$Yq?-�*>�
���Ɉ��+��M@�+-U?K�aS������F��V���D�n*I�W �@�U��z�p�N$�d9BX��>��?�/!�J)U�$N��[�PkF cȘ:�1�\�w1ɞ�����Os��|�,!� ß^yV����L(M�j2����'��4/�l�;��n�n;��u��꘤*��.���iA����D�@»ST����'�3:%-[A��'�7u��(B�Q���%��׷��I~_�Psg/����EX�YK=��p*������u�3K���TI|�ǵ��h{%���,�j,l���������kӺeq��<�HR��\�(&��m:��x���w��5��<u��)�f���%8Bm���*t�k���6�2sϱ؅�,E� �Vn:1@��|���,����4d�auw��&�Vt:E��g�X\aV!@��S�erB��C,�F
� �>�wU�e)�eP`�cрx�����?
2x����q�ɑ�#5���m`5*[p;���>��gL���}+���_�?X-'�N��%��:�P��nԕYC�����@�K&��?�9$���)�Uw�6�9�����
�ӿ'W�Osf��sf�Άi���̙q��cA�q
K�w� E9\�62�=C�zd�.�{��[QdX�`�0����.��a�DwEE����d<rѓ�����c06����w��o4~Ռ7	��=�{+�Q���Do�R]
�kW�VsV��t�.�F}��+zN��;�-���8�r�}x���� ��'m)M��-�T$�����?�Y�Yt ȴ�2��t�}�qs6��p�1��N��ǋ���\�|�߿Yi~\X,��l��r�H,y�Y�}\W7e{=�� ��߬�$S�**��U���\���'[�Y�l�iG�6&�jk�Sf�mYH��qF��S����x�EN�D�,� �P�Sz�@\�z
�lG"�c;@�?��g<I4��ͣ-EgF��@����`��6��/�ٝs���8ry�Vv���j���k&�s��:k+���`ԑ���W=[4���T��Z%C��s�4�{�c��������m'���9�lXw��s�rΫ~��<�@+�g���º�g�r���^"��۵�_�s"0HGТQC�Z,���m��,���	堪�0����WGb�p9BP��sz��jj,e�Э[k�'�HÄU�!H>�b�Bi�jp�Wp4y�(�f��s�.
G {!�_��O���)`p�ߝ�bMUR����Z �A�Ye?�dJ3K�u�8=�o@����MQ�iq���"Fv< �S��ec6��9*�땢XN·�'��]���*X]�!lӉ�n՜7ډⷉv���!�1qU��m���3!���C��ִ�H�������_1&'�/D�4�9��
5�A�4��Q�.���>��?^:�q�1�ܳxf!�J�eBml�˕���`�0x�|b��hv\֑9F"�͕�=�ǦEy=��	�$�&�D�C
 �@S��

g�҉��/9uR�`NҺ	����0|&6 �����2��}E��!h(*�G��g�)��3A?H�dP�#�L1m�SW�M[	��x�'ߤ4�٬�����G�8Ol��&f�� ���=T�$e|���Fs��һ����w[)��7���^���L���X�B�O������F���;F�}�N#�Q����C��j�jW�#�u ��6ݲ�a:I����p�N���*�Ϸ�����ݞRY��@rk��7>ۡ$7�{�F���}֬��|�ݓ�y&�]z�A��v6��'� ��\�S0<��}�� 7i8�Q��/.P(�G�����԰9��:Gk�atg����6�`e������FJ���8�����}�y3�ppet]�`��:\q��ω+l
����u��l����z*��ٙKV"��/Q��eҜ�0���[�e��8"m����<��ʢ���0�S�u�]V?����@��*[��#��\��]٬~�_QƓ҆��"+�[W���}�uj����$�%��O\��iFd{�e0 XYN����������`�4q����. �;�%cz�dHl�m�?���s7'r� �����&�JV���V��O��0F����pCݰy����)�b��ʛ��*�G�Z4�u�#����ZYz�<_����� ��S��8�z�i�e� ��V )0��L������d�Xl����R��4A���;��[B�M�D���1�ǼԞ {��x�N�Q����6)�>�kՅ{�藑U�s�r�`"
<}�]�����T�WQ��F��L2���n����=.�e'2�n|�E�zvuqػ4t��z����lS���m_F����u]Yï���q���^�4�ձkc=A�������7��޴�[��я�9)���Άs��e)ƍ�=�#��(���-Hp��z����ᨈ�{1Ig#�$�.�k���x��܆�0y̯�����(�m`��_�S�IL탅_�F��2��vѝؚ��H@�x�d^ݠ���&�y��<
VF}�g}��R�����t�S�?�zf��W��p��gnX�G9I�V�-:o�y\o�Ka��͑�uT0)
�7���w6�60�`���q��䋖��Wp�>��{K�����Ia����k�?�e6"�y��pgKL���*�����+?[E�Q�]�_O�����HdV��~���V�5�}z��K�c��N�G��r�rL^�Qz�@�[2���n^�Wޕ_���w�n27��u�F�d��i4�/��5>Q��2�seM�eN̑9��vV�Bb�'���i4#E-�a!�s�,	���@XF�:p�����`WR�9���ʰÔ�3jWx�e��om����e�+����7��y�
Cz��3W��r�r�3��]��r�A�.���-�ӷYGF�Up��
�+������v[��\-!���K�Z�=�+S�^��KJ5�-:��刎��S�	W��Mm"�_��g�֣�8PѲj���d0C�*l�)v*�k����\�������H)��E"���_�^�L���\	�G�%��\XP�p��"=g�\%�(�/��[bU�[�$#�ٜZ��A�-�w������$p���ۭ@�.��jX`�/���>�R�����j���͖|���[���3�A7
�O.jp0c"��=�=]-�^����>��r�'��g}m0��J�҄���b��D�a�� g�Y���-LQ,��xn��J���m|�4Q�eX׃�I�����:��y�8���s"c\{#ճ�e<�k��t��]�s��L����V�U��l�����0c��7���w|T��+�Ơ<�s��x��`a�;�땆7X`Gz��d�4��4���31C��و���ʂG�n��0���^�k`�f������k�h�R����a`["��R#X����v_Sa��w��x�s@p{��v��(�%��C'gt�<��cз����r����7H|�a��YV���'e�����9��pW���,�|����"�B�"`�I�Ө�{�����	,�M�Ձ��Yb�?iZ�DhT��$���a8���O��n�J���B��d^@��6�ma�
*�	���c���$`Ka*�*N8ω����~PJ0�]e�X�v3��������'��#�T^�x5�����".Ě��tRu��+��4����մ1�Y�="�t깝;_<���i�� .�륟<'�F�E� ����N�����y�y�;�$u��2Ō߉�>�F���B4󐉵�i�BK��"lט�7v������|��\�_�f?{�u��	, �V8�ݩ]�@����;:�?��0���@�E^���Ȫ��Mc�	 ��Eܗe�����K��27M^@�C�֪��!�����]"�j�
��g�ר圎:@�Sb5�}Ĩ��.Ո)�e`��sTԋDsi�q+'wW�Ō��/�5+JD���[�88n)�K�A�(�5Hd�~%�C}X��Ob�$`kY�r3u��xY�q���j�78R��0L�D��t��3xʵs�
�9o�@��ws��w�3R�x�D�M��h|j�鬂LM^��~�^�F� �����jB�k�[�t�	J��8Ҫ��%T�᝕f�Q>j˞�<z��p�����'e����s���&�$�ٙuFԞn�Ǯv���S`�wϽS5���S�!�>�W����x�;{E'�V��ʴ@�͔^dPK��ן��Wv��2q�U=0�q�H��nE������ئ�៬(��*S���B�M�hU�p?3��(��)�B���pJ���
*�����I.���i�Dڕ��
��qܡ�g9Y?ʗPFXO�7�L����aE~g�_��m��a����b?��<X�2�$$g�]�C���$/^�"�T�M�$�
/I��.ձ��z*jmF���An'��7��ǯ��:����6��6�V��ܱ1g�]�'���IM_��w5��F\�Ȟ1,;���*�*�syVS�Ӊ.��s����C������X�I~��剬�6hp�
J�IV�|�g�*�m�#�HƆ��k�q��A����R��p2Qq	mO��Lw1��b�:����ߟ-���V�كԔ;��ө����>DG3��	P�����'R#^6�/'2������e�X�Ե�@ �p཈��x�Yf�AB�Oơ��`2 �@ױ�{�6�h�I`R�}����Z1Ӛ��U1;Y��v�k¹x�\<�fYxE1,�h�������vM�ߠ�8��_�*	��$��Hr�#b/4�(����ѱn����ߧia���^�K�x��ūQf�*
	�6b�#�������	g� �|5�f>��j\N&��,����C��E�_���(���cF��8����%�7Z��z��h16q��/]zz�Di��N�%�i̯X6,��%���_�~�����T�<��l�3��u�~u��J�a.S9���a-���-1'���jxC�-��e!��������w7}y��1٢ݯ�Y2�k�C��o�u��3�q�˸��Q�nlR-z0�*�*OTB�Zl��u;GV�
����B�H��VpP�˵[�W���I#�1ﳑMG�����/s�.(m��D̦4����4D�>+cj�!����E�g�eFf6K���,(�c�ÙO����n�c����Jy���P�lof�4��������$��"�]��R⪌}a2��yG�k
�|Q��(��Sʟ��rzhDx ����-�A�M��͔�Ϝ2Ơ��E��x�<�o�`�[�F&�-��.T:B���6G�6D2�Qh��|!Vo��Z_r�t"�w�Սzq��$�R�Piz�R�w���P�HO1��@��ڝ'��@�P���\�/>��yq��6���^�� }{��&�`� ��񋪾 ��ߨ���R�9��:5�7C���1�� ������l��:w`�������5�l`1;�X����Fhg9a�"ʡ8�,d�z�gV���1���L�_��5����gz�/_s���6+'D�-Ź	ַ�ڄR�[����nqO�G|���V�\�J��<p�y��TH��U�K�]Z����X�56��1U,A��`�+'�~׮Y5�ѓЀ�g�.Q:��̧�_zE�����ڼ�n�u:�)�*����U��#<7dh�0# I9A
�6��\�j�3A m�m�.|u��X���Dnl�d�<�U6���na{���zѦl`��Z�y����:�Jlf���l���c?��K'�=��;F0�#�0��o�}��B2�Ow��elV[p�O�+�ٳ6�Q���X3����B����W�k/?�n8(�!юH���������j;)�Q�-	Mґ�!� �8m藽��$�/g�{:�U̇"]��G���L�P�
�aH��J�Ny���=�l]��+�Ĥ������9SM����vu-�Mu�(��qeI�4���^DD�oepV9�x#�puS��O|��4�$a�{�/�do3^�'���$�Mꩱ}��J/�L��So�{����=_儣]N���׀�oi9�O^�H_�lu�k���V;�r�X��I�d%�	<nv�_�g�FL	��=��d���Z�0������Χ2�f����Μ.a���}�C̑41!зMe�tG1��Xhkz� -�*j��y.�N[��(R�6@�&L���� \�I�0�RQ{��f�8�^�`�8͘V���^g�^X��>xoj����sh3�nߑz�S�y�_%py�������ڵ�?D��6�G#4g��1�ű�7���׋��̛f۠�y��r�@c|�����}�,@��ыle�UQ�*j�&D�m&�8j�Y�ͧWUF���~m�{�/�v���r�;u��ۣ�Bl��M��
d�A��Tb{`8��g$pQ�?|�nkQ����L���Z�
*����﫲z��+[Q��4�����x'�x=��ih��(̟���_tF�b=	�ͪ�ou�G��wY���W�%�2�#q��4eo@���N�pV�Plf��"�10%z���yЂ#�T AF��h�ǘ�ʆ�����l��t����l�dl�k��.�^!�a��*���KX�%2��%$毞�nMe�ǔZm> b(��T�Quj~ ���c"=��o���fŶY"���$�%�eT���y���&��'�R�﷈Z��hH�wʧ��YW1�!�_M{��� �t��t@Yl�v'���wՍa����C��΃y�iW����ȶUq�I�B������q���w�Ɍ���J���v�������Z���v�� ����a ��(���ķ�|q�����U���[��#8w�	��<�1�J���#w|���J�Oe� �e����`�|$�#P��fC�S��E+G��[më��a³�\3��D;���B\���W(r�H-���� D�䋵�}&�e�ll�a�$ �����������ev�G�Gc��ݞPwBR�QaQ2G��dQ�+{�)̓6�����H(�J9�oH��I?��2CY���i�;�=I�8�C�<�*�΢D��e�nmgb�+`�7����6�v~��#y;lT�ao|L��
y�O�����Ǵ���n(��;/�kg������vZ�:����7��a�A�a���ji�w��F�F�ϻ�&��#)̲��ƻ����LH鬫*B�`��n�˫�Π���q͸���E)�8��N�1���Ս���ܘ�_H�-��p�;hbh��x��g�\�^��򊞳o��tO����Būw��u?^q&����1�- Q��U��!�6#�(�I��yy��Y?�ec�JG����)�)����f^3�4�wX�k�a��@�]�!��e'�y���k~o�L{��L�{��,t����( ��XF^��B�Al�K֌�X-Cc���#���m��_}%�d�$Y#�k{�y̤���FqR��ݟ���!�J�����Y��-Oѭ}0���c���Y�j�j1b�Kդoh�%���G��O ��`/���{G̻[�}�L��+�4��ک�G`���1>����Yq!)�v�W�:�Թ��K���������I�CRp�mע��'Ҷ���S�Tg VQŋ]U�l�G�M/p����V\�P-?T��]s`����?�z���W7X!��:��O�LA0��ZŊ[�|�����5�^.XÈ������_fÁer���Z�S���50*���@���wR�������ڟ����=�c�W��9Ki�4����D�ØEinEkF{I%b�i+��,���G| 4ҡ�^g��jwO�Z����o�5�2�xm�i� �O\Rg��sBͬ^�Ҹ��W��δn%!��LZ�E��Hb3#N%L��2�j|��H_�1P��7[�yz�@�AB���@�@}U��|��%WQ�
�[���6�R���9��I�Y���Z�vxa�0<�*��P5y��D(��q����_ %��;�1�X��j��4�V����q��Q/��W5a�l�=���7`�B<7"�h�¹�V͠4��n�q���/:T�iGG|�����A����U⪬���!f�]Dy����l�>3�yR�M��Z-��y�#��E|d�圻�3��
Bϙ�3�����%�Z�TWq�k�� �����P�~%��)���`��%�P]wbj��CC����H�F��0���UP����	=8n���%HR�����.���-k2i�Gu!��w���'����%�U���(ۻĦtI:���b&=rO5�h�D�m��L�W���%���ش"~>C�]��%hi�,�1T�o�~:`�,���F����֝#�Iu7G3��k���:S�	�U���v�_��,E2RGVP�]�����f���DR���^��H%�XT��tҝ �����4�F�
E��ze��15�X�RF.b����\��^y,�{�Q�a�DQ'�]�3⭞���iQ�_��׷w;�q2���:l\�0!�����J��]D*�!�l�t�X�{Oo&G��Y�dH�|"E���(��z�l�&	5p���Q�������yQ{έ���*��fĬ��:{NZ�7��>x��tn6h'�����v�|�/L��x=�c��6$elk��#{И��{&4փ����qS��x��,||�{��
�S�ccX,�E�.G�	Ȗ��f�c��J9��|
�����e?	�,��������g�H*�j5�@�n$a+K��O�]`n�qC0����(y1@:khKV����jW����S�#��8���؝�`��Q���s��>0PG*,Q��1��{`3`ĉt[y��K�^��\��vz�SV��R���X3��஡3�n�**G��L#
���l#�����Z/��d������\4G3L+����!r�g�:�mA��e�1���:{���n.��*�#�+�+o��lgl����z!"F���<JIg�D"���/�2u(ve��!3ed:�~Ld�u���DSF�7Y����*]�/���e<�Y��2�g�E'l��X�dk ���@�J��لN��ճ�Hԃ�r:-��M=��ʐ�����v1��L؈+����F�ߙ#4�wqW7�a?����+�*I7�]<7*���%�r�]Ե⌬~����{�����#�iN����<�vw�� |e �gG���9��Tj�ĺ�Q�+����ܦ�uz��. ��vuΓ��&�읩B�\s����2��4Ǿ�l��H��|��`����B�,v��F�����+�Ե�h��4��W�j��@GP��笽�e-�IM�����Kk�q�^l�{���'q�C�����Ꮃ��OLd���rapL�f�A���
|;@�`���RZ��4�#�x:5�ÆV��*��Y���qX4ܓ�7�'ڳ�9���ba���D�x�es��^�h���-|x��sZݏ�����Vͤ�=
��?�K���٨X��BL*��P.��0L����3�ˀ�!J�)r`�K��-����cKÒ3>�8zn%Cy����g5{r�,�!�Cul[���6��YTc+�ag��I��JB�7|���j,8"ef��c�5ǘJA��q�@J#s2��n�_�u���e���0�;���d�P)V;C���[��3��@`�1��ɸ��K����T����k=�������!ܳuٛdi�m��g\�j���P�U�{qC�wF�t�q%��_�Is���|p���Q����K����|�س�߿Dd9�<���C �ؚ��j��^��=��mm����hg�'h�(�60�y��*-�EI���?y;H���8�Wl{%������XeW>�!x��!^�0�a{�h*��&�SɄ_�Ζ{��s�0&vD�Y{��@y�N�GC<ND�����j��G6�w�"Kʠ�<m���v?��`����� 3�o��t� {U��dIX""<��cB�8�C6�	bhW�k���ۉ���f&�w:M(��]��X��k9Թdi^��n>l����6KM� ��G�ۘEl7F��Z��<;�R���#G,
҉ၗR��ۏa�f?Nf�<�6�g��;v�s����%�5��q��Ǒ̦��{3��"�{=�P�N����e*�x�4�gܽ��vU�Z��U�����&n�E?ѣ�hk/*��Q�x�@ͬz2����5�/QC�e.š#7Jbz*2-�ߠ_�ʯ����Si.�t����fO�h�h��V� �����ї�4L��+�V�P�Lp�/:\�,��b���!�G뇅j�S��K�G�M��/͝����n�t�6���̦��Q�l����L�L�	��9���ɬT�m<�5��f�Ee����Ƣc�2cR�>�=�˟��������ڈ5+5����Ԇ���K|�(6@W����<�&Yʖ�� e���qu���G���G�?Ҝ�?�J��#"-�8Gz]��8o0�T����c��U��ǜ�g�oNWS�ߑ����.rط֯�Z�nc��z��>>��/�r�"z����� ���Z$�P $]�PtG[ٛ�#܅u����ݙ�G��k�*v�<��^ �}��l�n�e�?���7�"�$��o4c�c�m�w1�:�7Z��@� �6N���5 h�ʉ���5��S��U�|[�"4�[ J�z�G��qY�I|Q��N���fw`�B����#���y�¡[\G�U[>�6GA��K�[�x�	b��C~�b)�A����#cS�BLm�R'~ɩ�dט"�X��؛�Ɛ���ѻ3��=��=�S�hdh���]0^����C6��Z�inf�g<�7�R	��/�U^έл�g��QT�U�m[`�p}گ�3]�2���$'�`{1Ta��H`�Ԇ )r�wF���<O;ͱ�EV����(�,#'�kᾌF��մ>�MY����Gdkh�s �j`�F�O
D��X|4F����dE�9�_f�ڳ0���!�t�G�`ѹRȨ��r�t���њB��
y��c�!���� ��Ȉ_Z�b�����{]�=��)>�[.�l���՘��:[1��L��"B��b���ap�>���s���-����z�dR��4݃��8�pO���� ��za�Qi9�Ij
z�I��S͌�·muɟ�j�#V `��d��#4���!�7g.�^�ߒ��f] I�3=�J"���	��#[��Q�lc5�tH�b�47���)��y�K�6v7}Lk}�F�����#�����ߑ�|
���lGO�0�xu��E�rV;��H���3E���w�fgV�ϟ~~	('8��2?f����#j*�,���j�?�z���o�})�6#��&��֒����8�j��KN�g��3t� b��g'uFſi�{.m�e],^��9�a�Y�jP������t-�:{��3~�H)��	b)lk�-��5�1�V U%|�Q� ��!ϋA~�Y�]��<�,���O��^�,tN�-%뜪v%~#�BVM���G�{l�t�8tw��O���] �q.Bo���Δ�� ��������Q��.ϝ5Nx[_Eb8�+�i�JP����ٍ0��c�#��c	�M�j�6B��/�~��t�J��n�1_ c�`�m90q֫5*���!��i�]���g&3�&����^��#�Z��y9(w��N �\,��v��(+�ª'6�}��m_7�#H���&5G-ϚF���n��U��� ��5��`�Jx�L����oV�Z��� u=5�����`�mUK�E9B�U@ڸ��eT��u��$�y��O򵃻4�LÖ�.2�8�Y18�\�q��h"��k)az�K/:��[��<��]���e��I�ˏ|S�xc�]�y�h;ر�?]F�m���(�����7�̭U6�r.&�4�
����G�[Om��0�����C��[���"��3�9
ڋ���Z3PՓǚB_�jJg�mS��,�%e듶��h��mL`�L4���D�X$��K��Z�GJ">?���
>x�0˨ >a=G�/[(�K�?���X��A�ܭ�V�8n��
w���urM� ���"�+6�K,����D�V�*�b� ,�|Œ<I�m0I��	�������Nߡ�������L�>��]��Xj	�.�Ň+h����j1D9��N��_R�S��$[�:0������~���*�M�^��g������ui�.����6ᒔy��,u��E����5-��R+}�dho�{��>����l��Ռ8�
��p��䠱��e�õ��{@�d�����+�9�)�5Z�~�J�ߥ8�;��v)Cy�q9'��q��ѝB�gqc����ᆝgb���l��f�f�. �*�:B��LA���6�s���9Y�݃R�Ը+�	da���_N�N�B.x�d��^��+&ɤm�o^�-�o���B�R��l@bFDu|�Wm���I`l�| ��u\�Fu~���p|��ص�h��0绻���fv9]ZhIN�>�?�9U�WPD��O�����D��T/$10�^��"��j���^n0����/1�!�������Y*�+ Cܠ�z%�슩��Fΰ2晡K>F�v(��-tn���gS�m���[n�}���G���G�&�$~�y^A��w(���)3R�����ê]uI��M�%�ؤҝG�rc�]��ElGA�K��S�Ⱥ�J8�V�f��I	�vQq>+���=ޑq�>J�����g���.�7���G���%�u���s���ޡ\��0�2l��Tv˞�5�d�C���IOld���e�b�V_G�쇘D�����(��=���;��`�u����#�.)�?ʶ�XE�I����z"8�ͣʩ|;���| _u�(�Ρ������<�Ġ��i��F����}dc������<�����?c�ۆ�Im�C'�]���n�8�si.�LM�����}:�b�\��T���!���vi��z$�%ꐬ��k�nJ����
8�_�p��w=S��4v��O8�Q��ly��§>�I���I�p�!S6uG�g�@�g.��F{t ��)w�}v�.ĉ!��_��6����BgWu�|O���}"AQ�9��W=��U�L��6U7{N�?_����XP��i<�Y��,���'\�T��V��q6�y��c]ܵSji!��q�g[�|���kU5΢nAZq�n����Z���W�8�+�kwُE�@��v����b��}?������>>PGɖ~�����v%���tٖ�r9���J5�`�V���G[��t�7]6�в?��jms��!qU��,Yo�(�I�%�%�~�h�r�>��G�M��,�zZ�6I2�_�ȥ5��
��UO���W��I��Z��������� k���}O��pU��tK��81i}��œs\�I4S�T����-���2u=��(Wmf�(]�p��C������*�}`:�;"�e"`���KdI�^7��:�,P^Ms���jN��&�
}�c���Vq���^rTw�ɣ'�ʩ�!5�\{�.Ӧ��2�A� ǐ��q:�,��z�Z�����]�)\q���}�&�2�S�ܹ�y�9l�#_�\ �����,�X��NVs��sϋM�n��ze��"�v�͠Hw7�a��,�� g�+(�1`�-t-��橶��~5���xMe�_�e�L:���6�D̟R\�Fq�T���5u�5�!x�� ��P��N_zG#c|��@��z���R��<�_����"[)��Oa��y�$�'��$��T��7���X>���x����Uc��# ��?�=(��s�("��\sy�hM�yq0If�8}v/�\�O��<�����"�}�=���Q��_�z�"�5��pA�����0�%V��,��MB�T��=On���u��)��g!]�s����Qa���o��N�p`fj\}uA?k3�Є�U<aM��d��C��(����O����aY�1e�R#}4�c��xnS�2��稪@o���yxL��!�3��m:�u�}�jU�+{�D/�rAl�i�l��w��b�qo�)˻�$],��x#րu`�n�%�v��� ��&��!� %�U�$1C�^���	�Qb|R,�S��Vv%�x2ซ-�f�V��5����S�cﹼ��g������K���@�&oQI)%s}�<����	�I�1S�����]��u� l͙n������
Zg�Cd��D%?�L���puB[�ي�h�, �*�KO�1�G�_]�Il��iB���J�fE��h���«84�����$K��s8�L@��q��w؏54P6�QQ�Ψ��o��T�A�Q�]�q�S�;p�NV�Pa�D���# ]��G��lc�W9�\����Z^g��@��!�x��g-�F�=��4�)����ct��M2������%-6��p�*���4�Q2���	�i�F�����~��aw��;vd+�����n��c+�14���G�/�v�A��%�R�Il�a7V�#q&��	n=Eð'] ��7��k�\�4��nB����Y:�1 C���4�x�S�D~�]���Q��.���[�-WR��=U`�(;.����)N
L�НR7Yw��6�D��P��H*!��`30^��b��5�iC�W�A�?�;��<9�dC�+�]�u�K�V�Zn\	�����A���Ֆ.��cإa���p�/����։��֚��=s�2ֆ=��0{�`ɞ��$*&���	a)���V��}T~�͡��L�d�:%��j5�0D<2��������p���"!ͺ�w��2a������x�7l��r'����.��.f5{+UVd����km���� �s���цV1��\pp�Q�̀�9�t�>�",�Q+bl�$r�V� %'�E䙄���۴C�	��2H$�l���v����y�=�=PH8���X(qȎ�����w�Lj�|�6�1���꽮�,?�#�7�ؚL?��o+�2�nfy/�W��������!k�
.^
t{~�,�W� .7`Zq(�z	��z^L*���8%���� Ơ����Aأ��j�1K�A*M �Z�S����������-��H����A)����A:��"A-JDoHx�{I��S͟�Ss���d	p�mqO5X&	&@g�h[�Xy�g�z�-B�Ǜ�5:��
�FƯM��7���u��L<�'!�� ��aV/����㋊悤���'eܑIh�$��_�����#<�Y=�E`$�6�gz��Z%l	#��]fr�]Pf/@���m��R���
��]�<6�X^߾v���������aZtc"㕋�����]:�f�qW�Z|E)�z!=P���X�.����
@��^~}/��݇vq(�/pw�8�յ�|�������(y��c϶�;�#U�j�+ʁ�����x�.�?F��O64�ﲱ8}��3��J���n6�K�g\�_һ��&ЂpvV����yZ��ꐘ�����R�4��V7dq�,�MG��I�b1��&���7ꚃ�8@I�d�v�8�r��>(��o��Yl�v]�}�͚�Ӈ2��j��U:r��|��L�o�b�w��O ��8����q[�cP�c��ʇ���4����8�a����z0z��ˏ9(ka���c��Uwl/��#��G�W��h`z�5��DZ�沛?�I�)�`n�i[~2����$�v4J>�p���?�ovg���<�V�նǷiʞL{i$/r3݂���Y�p��6�.Y@�{2����=��J��7̘�y�@0���U$�e\'��=����STF�'�?���ME�� ������)�w�!"�a4]6 d���M<�B�e�U7Ϳ�ti�X�{.۞�}�7KNLSmt*EVd�2�Fy����|��k�yh:V���vt<�eO��������L��,��#� m�`������Ⳅ�oόv�-p1J����몗�1S��K��B���	��l�b�ש��:N|�ͨg:ٟ���T�yK[�����[���_�#��&E�B�L7{�1)R��˰�T�7�!q�����+?m���������N����4�g�,���IG�!�A ��W�"1M"���l�5'j>�j"�6���A�P��Eee��i�h͌G�>a�J���g�S��o{����"�| � 0!UJ<}s	[�h���p�_�'�n�h���U�9����@U������q]P�U�A=��J���H��N5ѷ���e�-f!�
+o���~��#��~��Lb�I���Ku�ğ��&���;~�q[Ijr���L�l����J�K3��F��C��s�w�� �ւ�Ql	��.K"_�k8�%�m�Gv����7�T��F�
�O�'�lvP!@�W1%6.��݄�i$5ܫq��f һ�t`�p9^�E�$�Q��|��Qh�����a^ذR���2{ي�5����O��N���ĕ<��;8�}'~�tU���4貘��]�������A�t?:x���2w%w��P&�Ꝉ�8�zmҍr�gY	�kR_�v@��%�j��Oam<@[�rr'ѢN���+�(byf�`����P���N~<�h� �@�y��� ����<�ݢ)j���=iY��eD�/pHN	�y)>!��]<�l�e(���ׂ&��}��(z^�Ǭ����2'����룷?s� ]#�L�	�L0u���<rؕ&�'D��T����yNT}��ۥ�y��F[mKĪ�5������ƌV���҉CP*`>0����ͧa	}kL�����f�c��+'����?��s�{��6�]d���pV��fWDg��2�O�Oo$P>-���y��6�c�����Ea;�.(��6h���K���B�.K��8z��Į�3����6��!ݵ��d���@z�Rb��5G3���X,P�wGV�:L���RX��0{d��?jU��(�w1����J'�e5zRջ�W�Ǎd�RdW��\I>��NQ"wpOé��_��a;+�$��&cIꟅi�z2?���� w��ʑ��j���ɢ�����%�� Zu�4@�D�~����|���MI3?&v�������::XM����8H�E_�+���L��٠e��g�3k:���e�*nbkmJ��p��/������8��'*B["��(
���.ˉI@�@[��z�a�O��ռu�-�Q�z���]YpSf��X�妊�>�M`c����:!23�}X��"��I�D(��_R�\hJ�G�f�EX���w��:�܋��<͙�/t��kŬWf[���>(�o�m��@��a�Rnu�� �FB�z��������V�)���4������J�e�=�E��8��ۣ|��y��m9ے����b��ȌaC�;g�7-�������/�g$�4�N��C���`.8���CÍ�cDj�s샳L�9N ����{5�3�[�2�A�IYsɥ-࢝���Ł;�zx��GR����Hb�8���yc�����^L.���VL��r�w��)�Q���5����U���&���Ԇ'�LRn���h�+�v�Ϲ|��&ٜs��ѧ�\R���i�,���ʢ�n��d��6��C����up6"��֗�
)�R�G2<:ʇ�nMZV%<��Br�����:r�u� r%A�v���ZS��%����-�U-�a"G�f�b��"Z�oq��\������d+w�|�0�٫0�ڲl����� ��� �z�b����6�y�c��.�R���5v�1��M�sS�k�m�?xq��i}���J�K�c�.��	��6ȳt�7/�߁G�>��RX���L|��;)��hAg�]V��،5�)".>�7 )�������='U�s����v\�գ����f�>j�ͤ���U����̎hE�W??b�<9 8'a�2��'���Z���E���h�`���Q�P3���6r�2���1H�B���!����oZ`�����?�^m�yS���[e�ո��]�|���l�gM҂x~�۔R����Y2��</�c���C-wX�s���J�d7o�����Mbu\=��F�֗ٚ��F!�A����J�dW!~�1׍G���d�����%���p��9���t1���>IDe0:9'i�Iu�R��JeL��=�ؤ�(����!�`ڶY�i/�*��J��H&[���-�j�^��BXES��L6y0��ӟNي2�P�,�d��y*!���l\Yܥ�\8��L��8~h��FcE=_B���=c4DLA9��)�?������ॸ.~,��	��x%Ԭ�gY�Ʋ�v(�}�U�͏nM�tp�� �\����"&؊�=&�HX*�'�BRs����X�;���D�_�^��������f���3�,�i3�����oq}@�<�X�~�p�z
$U�0oX��OD�d�i���۶ǿ��\���ӛ'YD�Ũ~��[�n���7��O�5��͙��F�y��ڨ�tۃ◡�9�ѺQh5M݄�v���0|)|�%FE�<��?�>�j�!���NH+�ݪײ8��`���>qچ7�殇*���vom�Kĝ�?��PuH&��������Z��5�}�d��L� 6���Ԑ)�<�܋�k"��E�0���RdL��or݄a�*�����v-�i<M��M~?[DF�4#<�����
�.>!��Z��#r@�Z%ul�����E�ܽq&���3X��f;��"Jӭ��
Z�2�.J��d��e���8f�aM��M��Q�M�w%r�횏������7jEO>��<|3b�W�� ��?:q�����+�t$�_��h�_��\�^�F'Y��W3��W��On��~>��w�!�9���\0�����b�,6ci����|�	����C�����V��r%��Un�ZO�����|L��	L ��������v�6�IQ`�~L�a�۱fX��]h<��W��:���L��3�Q6)��-���=$���X�G�+I�ı�;�!^��5�l���FI�&<h�"�t[]��{� �6f��3&�����&�H"4��$|~�ocUˁ鐫.1���K�L��¹�ep-���
���X��Q���-߉���,��#L���̤>0`:�X� :똙q<fp�� g>�$_Ϊ޻�'8_�H��D��P�Ć�u�K����K�)"����Ȼ�ۘ(fJ�b?���0���l�<D/��3����g����x1��!���_���(�,��99A LSK�i@�P'vg���z���^�W�`�m5r�yp�-�>)ܕw�����A�-��ԛ���7T�;̒��]}�y;Ldie��:�cKD��1[��4�3��H��?�ɇ,�#],>��U���3j�5��
Ze{5�g���o�Ĉ>
��V���5�!aН~��$ �eZ{�1�-�f���B�-��3�B�N���AY�Ā2��j�he
\Fȋ�J\HNp�q���{2�2I��B�������i�'љԟ����.��}��u``����0��ܱ���eiO��I!&�0�/!��� ��dh��qVH����`�z�ʇM��e��Cя��*[l��Q~�華2��9R&L�
&�]?_��C|
�V�T�^�)s���K��\<��'�[�M%w�#7��6�)���IS��aZ`f>dG��,����s��p����">4�2S�t���0<��>-��@�ɓ�'��f�L��z�~�ǁܔRݚ
�0b��2��{�{�ļ^���]>Z1�Ѐ�c�zu��c����p@�9�7��w���;�Yo2z��(�%������xi��EcC�b{I.��s�xç�Ü#�����T�r��;(^�;B'x�o��2U��#}<���X�=��f�xD4�>BH�酭`�AÄ����	F�hZz0:�ym��լ�:S�K��г�Xa�u/�4-�\k[�"��s���߻�F�D�!��q��J��g'�� �!�9��y��t��S�P���8Q�+E��Vf?���옓���
]�i���H1��v���*��,�ʝ�=e�͇��4����(^5��K���]�[7T� ��G������|w�Q�5R�Ф��1P�'va[cc>�5��Fr��a3kJ�j��s?�э��Ƶ[��=G;�L˲�tq���W�Ҫ��ԛ䀧�DA�y�B�������	����~D|�ӊ_����v4�P4l9�M�L��C�4E��ʹ��S�{34�.�)I��Ŷ�N�i6ݴ��d��݅"�Β\�Z�3qtS���TF�=�������>F_Os��:��4����bU��[#΍�!�����e���:#2��F��
)��D��J��Ԉ&5P���P˳�j�� 6Z��6�+$��ѫ�cM��0�(��݀+T(�c�_�Z���A�۴�6���_��K6�Ìa�ƅ�����7j���F?�E%W4ӗ^dr��9������������a'���!u�����קU���㨬g�\���?�]M�c���� �����8���d��r�e_����jH�euvc<�,��ꑉl�
	��w%@�PA��~ �сV���W,��s-�姅T�� .�Z?���]B�0��dҗ|�
���P�7�F����@�m�tqyШ�gǋT��BI~t�X��T�w	�X���#X���!f����.�(K���p�Q�Wb^��ᜁ�=�#���xZʓ��Z���L�y��}I���i%x�Z�m ����(�H����R��4dQ�X`;�!���b� ��˭�*[��-��d��$��h9w��w_ >gX�e�����p�r�b�$�ym�Nc��mz�(\��)�G$|���3%"͝ �5�qܲ��,	�}���(��Ն���OC�w�ԇWE�xe�'9���M�4�KB�e$Y��e��b��ԔI�f�GL���U��^ <�a�F�V�C�ϱ⩬��WiW�Ⱥ]S�|�~� �Te��N���Oj�rI=�u����8_�&Cu��U�e���j�|���G`}c��+�04��J��Ҽ�m��R|�� ��S�w��2ą����Gx��-�}�`�`��N�2;���K�'���"��PAС�e��1�i9R
�őrP��ppZT��c����	-�� b�� ������Y��qI'M�8�S��^�1ȼ�L�]����Bn��A.����+l/�U��FЋ�I��c'!�y�D���c:6o��0���[�G<��z#�[���b:��L����I�ƕb�գ5-�ʓ�(V%����d�"Le����z�#S鶳l�n�1�`�$_���26Ⱥ&9ߏM�u�&F��g��E�f]t`Q��ܞO���]��;vG�=�AtQ"��QD���د8�:�v����@��4d3��S�}; ֑*a�Z9�G��'��Y�Y���EŲo��Hsi��v��S������	&�GRZ�E]�[�Ǡ|�	�	a�+��KЇ�Wy��.���R�
5����$� ��r��à��U��o4����fc�8�f��1���*�>�E�b78�k+�0��^��n%������ԍ�:-���C�Tvz��:�Dz�i�)�g8o�6��L�\$)�v<����Z�#���s*!��-������e���w���-f�EȋvgN�A��+���y	j��a7�:L�Az���4/� @���AO�]ޒ���Җ�vlX^+��8��b�*�2hj���ŬZ��\6X��B{d�+��ĉ����:�+�1��p�B�p3���a.��s�oz�ߢ��?�p�!H�Ң��*;�
8����W���������>*��fM���l{e*�!�Sakʼvc|.�\= ef:�6�3 ���S�tEe6ZP���x敾���-��6��ݝJ6IN��۔ٺ�?�	����V�%g�VJx�S\��R���$lD��L:��'�4�����'08)�Z�ᐆaOqS
�4;%���l�a��rﴻ����)V�?���L�q��m�u( *OoV�|�gW.w��>���O�R�d�����i���ޖ�'���R�y���h�a��on3w~�D��rW��J��*��Gsq���F�%�D�$���@V̑�PH+Kv��k���Dˡ�'�x������q���V���N�U
N�PBÏ$��]���k��#h*튏��p�n�<�Uj���t��c����@��wEBm�p�_R����k��dN��Y=��]J�h#�q`�3)�)�>��34�r���~ޗ��Q���a[C���!�W��H�	ޅ����4����^��(�����i�/%z5���F-�EF�(����Ծ���m�ws���d&����mZ�((��*��+���c�t����y�A#�蛍rs��$к��׽�d�R�:�tm<ǭ �x�$U�4������6�L�����"�E��(�&�~�4�LI�^����K���M�i�%��&��
���I�*��/=h�3�d��ˑn�j����������;��-�"	�Qo�G��,�|�*�m�3;)�T�>�M3$ζ;7G�Z�0��CB6I�A2�;��!<қ�>�8��dRl�۪Ƃ	O��:+:҃l3�4���#Y�4�O�aU`TN�a�m��ƝD�e9��!�d�k6{��R�c�P�x�a:~{f_��UMG���?�+M��I63��˘�#��7/eT(ҍ���Lf��%/Ocߗ'��bj�3�/��E�r�,*o��/3��` ���lK��m=F
��4Ë��?�S�6B�Yo�v&D�E�X�<�"����NO�|�wM�H	�(Sg����lEhY�_�"�\�D����ǧ�x[v��_G�iO�c�%��JU�y�N�ڦ O�7�% Co��A�_�f��Cg �;Y�[GșW��`+��<]�/ȓ���������}��maJ���z�%��c<��>)���ps�x��a:����{T,_vۉ��S�v �P;�ahP�>��jiwg�U[�yx�0�K=���X$>��l|�c��s�v�x��u[ha��H�ޒ��/��[Fz{3̂v�k���X�
�)m!ԭ<y� ��m
s�ն"]84b�������๓�z�e��u�J� �V �W-�(�|+~�{��ݍ��36�\ՒضX�Mߥ�,yCL�(��:���K`~o�� _��K�	ĩj�M6Z��i.�ى��j
�o�����x��gM����ͤ���(�lf�~	ؾcz��`v�j��5�S,F���{:\j����?XN��`)q��߭a�7cF�3�:�fZ7]�_(-�ٞ�i��N�z%,�;�k ǔ�w�zk̩��G����Y>���!�:���p�X@e�sl��N9:� Kߟ0��l�����{�`�n�=-Tq�y�N�ꉠT�ѦnK�$�6���
{p [�9�(O�x����~�{�!,���Ξ�'�}�J�]S��,��R,��\3�~50�?H�H�̋�2!�*�$�9*��9-M�ۥ�j��GM�+Ԑ��s��X�C�f8����X�C���u/>U0)��fXyu��6/c���E)mn�+^�#0Fy＾Uf��H��:�W�2�����Ή�O�P��� �o�0�����^�L>[5��'�C�-�f�{Q
����;=�#o�X.��6_J���W]�'�t.���X��..i�{e|���;���Y�R/G�f�$�d�'6U]:6[
�	�+N�梷fA)jq���s�)�Ҙ����^H�FI�ȵs��-R[%y{��߂]&tqh�K��a� �m�����	'�t:U�^�>��H�u���r4a�-�2�v�xs��4�o�kw�%��n5jU~e��t*�URrm�X��N"��S�H�Ij��{ҷ�����xiĊߊg�?_#׷��`��� �i{�ky��,��9��>�v��W-��2a��F�\��/1��&�QkF�>�\�q�e-� m��NGV& W��A^>��]���6���+�����Cn4��$�+TZ�;M�Ek�8�M�tfW�L�g"�[[uS�ڷ-𠵽���<&(��66꟔�\�u��O<�$龎��^s�dN�����
�%T�#*J'��q�K��ָ���EX�h;l��,@ZJ��G�#+�gf�W�c����[�����@L��H����
��I7D+���f��~�bT�B�R�!OVzYH֚��D7�2�z�������w��@{qPJ�M�1G�y)��J0�}��骻N>Ⱦ�7t��T��A ��R��K��&�X�Q�8>r��G�#-H��$qp�̒)��d2��3���|.S6PV?K�F��
>�I�_���2�dM�Zv�f�TnD]�E���Wt���S	m��<E�H���覚�j{ܛ��R."�/Z�U���#?��c^'�3��������G��Scb��j�Nŗb�[_|���|3&��|w쑹
Y�>��%�b&��`K�(F�8h�:��߆?�={�-"��l�h(�!:;�c�ڂ���U,���|<Mv��W�e+\�j�L g�	{"\�TF�K֛ *���<v��-�42���"���Vte���n�%}����?����!S���h{lܯF������)졙�ԛk��K����R�28Ĵ�
���������{7��_�����	GH�=�C@��̥���zn�����Yϭ���������G��у1���p�;�eLM{T研�P#�A�Dk.k����4�p��<M�ʢ�|b#j�<����-hÞ��.O'��Ȑ��v'a�8�Wi3>sĞ���F��&�����Q��z-``&���a��P+�e���,�z����oRf-h5������g@V��i��ir�Vz	���$,�,6�ıE�;-���؈HN��w�nN灒����)��]�@�:Ԁ}>��.�����Si���(R��!<4ɓAH�SK�	����V`�&������ZP4��}�ҠW��{�g!܄��^VZ�E+�/�u�8��Y������P=hl��$�vzY{ �6��P�s��\uO�i�`R_и{��Gֈٲy�������21��T���/��.��H�n�����60����t��w���66�Oɬ�F&~�z��b��aAܔ��f](��U���7)���ca���%����� }0p�5�'�4�0�e��N����$��t5j���x=�f��)�Bރ[Sn�5��{�������T��ک(��`�j���WC2�wy����W���6v �g����k`�e��xk8�;�Ȭ���59�vd�%�����\r5��0����2@}dgN���滻FP��x}�s��N����"�N*.�7r�P������n�|,g�IG$/�P�ۖ���KO/�LW%����Y�d�_�${�4m�B�G"{ю��zi�����B���~n�(%Ps�J&��2q��A��Z�d�z�.�XF�?���t�Ka�bE2%�Aj8D`�,�צ��G3��_�X{�w��-�d/c �;o8�X������j�c9��Ç6��V={x�%�{:(�f��-0�<e�1�;<5�|�k���^S�&�o����b*��ߵ����F��c��P��L'IHL=#��]�����2��oe�fi�����,6زr�tY#Uv�Ib���. ���m��=���O�yI(���^lN��/u��uS���jt�0{����̠X�7���o~շ�L�~"�H�pb�t~0������:��吘��}����Z�����X�;(��Tȵ|�OU���s���\��i�ȄC����U