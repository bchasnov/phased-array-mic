��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\����q�?��e�I8�b�Ǽ$��"����ׯ1�V0���6��80���ݍ�F'��$
�����d��,
g���S�X��7v��]����ݷ���*���������snlQ��S���P �� m��f�cR���dVjg3#m�����(���m����)bƗ�cԧ�� �O0��m�N���QG�: */��/��;���E��{�H*M�*��/	KU=!��ޢ�H�����}����S���Po��_�gd�l>��'��0e�k��yM�`����3u����S��0�/�Zg3��y��B>��ֱ	=�����<VF�k�=߿'�B��Լ��뿜m�2d��L�2��tX���j�a̎���o���rʓ�]0]�b����O�hA��H� $�*�LT1Ac���. ��u���5h.��Y�N���WY$iL�����d�\<�yA��$�p��Ob����Oޤ���HÐ�$��UI#�R��Wʈ)H�q�V)�b}���?�9?E @��wD�p���7g"�����ngI��,o�� z�M5w}2a��u!t�p�
�V)��LNoOr�Xt�o ��X>sO���%�{(��΀ꍄ��+�,0�%O<8�!���7�bt���w�!I�0=�)�����3�J��I���>�t�gd`ʔ���/�\]���d�5F�x�z��ʅ�Ԙ�����RF�P_��.c�!u��#E5����f��XAzCJ����%ضi����=>�v�P�:���$`�.�b��I����ڝ�GI�o\"���o͊�#M.�G%2* L	�s����<� ɼ�.[G�D��+`(.岎�z��o��4�貹i�ӄC/��ΚJs�Q(9Oϣ�7��JOE�b'�3E"���<����b�rU�(���%`�f���f�fK�I�Fr����;*[��x�Ⴢm}쒕�<������Uo?I��Ub�L
�2���-1���Rq1T���td8t��a�g�y�>!�n7�G>"(�G�Du��q:��w9��v�_h	�j����SnM2�z7�L�>KQ�v���	=.H=pa�7�Ώ�����<�������W�P�O*��m�>�/K]c���J~{�1Aڵ���E
�!�\�F�-�O*8[2���av��A��A�Ӟ�Z� ր�6��ӥ�Q����!o����m��9P̩�}�J���%Fd���Dc�O�O����4��,\��� Ã���
W�8Eݶ�ۖ�����P��(��i7m[Д��T+��n�x��u%��ޙt튘����Z���)�8M�[���f���r`d��*&]l���D����}�5��if8���
��On��B%x𼁲&�E=�pZ�b�7�t˄�reG�4�h~DrbQM�շ���Z]�e@xX��x�O��Wr(�"���&�����Ǒ<cI�*�Z��Y��v1��\ɓ�-̀�j%��ʞ���mQVMM]�=g�	,����~mPއnZ�����	K�w�a�.b��~X�\Pn�	�,B�k}�N{D���ame柴��P��:}{�o4��9�ւFHނ��ӂ�FӠ��p�X�+\�M�&�����Z�s� /�C87N8p�}����"�;�e��}�}g���JL+޸U~�no�v�+RQ�cٳ��M�I��YL����¶2�&Җҋ6�+��o���`V�Ɵ�q91,��卓�CɎs�[K����6ΤA��0]M'2��aO���Q\��<l��p�Ԁ=Ɠ����	��q����������G۱��j�$&F9�G�p`�}���*׏�]C~A�'E��CAa�~A�H3wz��6o���Z�[BB��q����\n�V��q$3�!��l]|�Hȶ0�I<�!�64o��\�c�����6����%Ʋ��\�	���'�f�ui�E��;��G�e��PF�Ay\�[���s+qw��Ae��;���a�}�e�
�NLFAJ�K�}|��X���Y⎥�C�&~�'���J<�K���X��-Nêf�dX�&��sAÖ�HNQ�rN�V(9@³6���>�?����F+ّ��$��bÙ��lIe������.�|,4F�&/{�[�}�L�[��t5�[C���B�J�M����VO�
�}Hj�L;K�Ĩ��\
�q��B#d)~y��Ў���W&� %�0�YJ�-W����A8rɅX �
���wzDo�`��b��uC�*W�c@+�*^�q��5
'qTH��vF�6t�?J�kq�{���?�<ҷ>;.מ֡�<a$pU������a�HM��ea9�|u^q:��Z:�/�Q�u#��ˮ�h����J��w@̎+�)gL [�������Q��Tj
<����ؕd��@��V��*ak��,�t�-hI�t��e͙�������V�`30P�5��������:\�H��]���Ζ%~縵~�-J>7/�TҐ��ZeV�k���"�opՊR���8�C`��3�"�����Ț��2�?y�U��o��D)����K֔���Y�U};mw�G�����P*��w�EKa����hu��L nms���i��D���{T��m�����I�g�#B�pU���@'�c�9�r�{� ��*�[IWjW�ӡ�$<6��28�{�4�����{�o6��_S����.]�����=�W�ܪ-���%����L�S	ـEyT�&�����I��(�����p��c�k�L�S��&Jϟ�<~��?#(O�[
��r�m8�I!P���}�,܄+;�2�*ҍ��4B:���`��4ehC��B�"�;Ӭ;�)�_Wn��/`��wA~�9���>\�ύD2�Գ��cFs͹�	�Z����ඎԞ;���Hp{�G�[�x_E�����SE���J�y��v����4���V<IJ�Z�c�'��iR�A��Ii1��/J�=��I(���WLB��a�%�ә
pR�.�f�gID@��ų��:��Y�M~�<b�r(dQ�l�i!V�#5�3j�]^{��}�/X�C�Et .��%�jc�B���1S� ���apwN.&L�����zf�>����z��(N�{x���C�]�"�(�	�(!⍳�<d{j���%�Ӎʈ��	 ���.]�l�Sw�������_R��瞲�a92Ъ�M�]�^�iD��-�ζ�[�(A��+V��������ܝS@�O��/��q��0�D��s��
~�����}��~�ʌ�`��VS����גyf��S{�	Hto��n��,��p�g1IMU�H7����@���)��,E�Ǧ���>¬>ב�zңA3���&;3�Q����QIy���X~��R���@�o��N� 9Mo��L{��l��C��z����>Ų�#ZHPs�|�6w���)O�j�e�f�l��釧���&+�\�C����2B�wx�: �S�sc�l��j�ǩ���R�7`�A���E�^ȻO��(��J�41�c�O����ʀ[�39Dz���$wcҼ�!؀h���Ք�m��*��e�!��y��ߞFd�X���J��`��M�����^d|.�M`y垇$Pxi!g���g�A���&S�� ��`��>*\w�j�@ğ�Y����;<��:S�M��,������AJ́U�I���f�:�C�d� ����y�*v�O\�Le�;8R�4V�$��I��.a�a���p!�v=��R�ه[L��M�f#�z]�p^�V�zA��Eӛ����9+h�C��V5��Ϙ8Y�m��D�cOl�����2�h�w'K�|<���<y$�k����H������@�57*���3@9�(�!���ŧH�L�\�E�oz��IU�<}��v])ɟ69*�Pe���/5�������v�dґ�/\d�~>����!З���5K7�$_��Ɋ�.��嫠G\��hq��a{���
�Q�o�����S�+����R�U:��7��ƙ��jc���4F��LV$��;����ZV�����C�C����e���ϷI|y	����<�ʴ����>��c)!��{���ɋY)	�"��jlʣ��51yD�'$��B��SУ�k�-V֘~<0q�����cs(�旭^�����wos �0a(B���pL/=�N�I��&�E���(�S�!�g����C(뎽�;�M�*J���6=�%�����U�=תs��mI�4�k�stbF�z�9�y��ř�E��A��q�
c�.W��
]��4H=���6�߅�ok�<���p&sa�#��50���_���'^u�TJ�E�r�݀��;�÷Q��]�Rz���c|^E��>Ȅ��X�?��V�H}�
�T�t���J�咶8�M�B�V���F)�\B��)�
WD�A˦9.��(����c���v��
F
��糫���%�,<�P7���d��m�������w��&O {���Ҽ����ϲ==ޤr�������X��g��&�[�$k�H�FU�n�^P�[���DkR%!�?=,�$��O��K�w�$|xw}
�y�Vݡ�<���;����5`d���k9�e\��3z�l���7���������������m��ی7��BJ|fȶ5���351|6���K6��p6(,�b*�F�Oy��7�vp���Pr`�Ji�^60�q���Hμ�r��7*�9cF�AJ�����Ժ��S_��~��0���GڽY;vP~j_&���1�]~ri����(�r���h[f���̀� ww���Kr�����v�Z�x��Z��� 6�~�`�m�!&��F$^`�����/���;9�ڶ�f.K
߽���� ����l��ɦz�,���^-��|0i��-���7������1�I��ʬ��}R��^߾!�|�Ik�R�>���ʎ��f��>)���(F�,壮-��B�+%D�������I:��-Yr�r��'�b��#h��Q����]
;������ĉ{rPF:QjKjU2���{�u��,�1�%�O�Ɍa�
����ˁ4�`�iʢ�X�|a��J�cA@a�~�K�Y�AͧN��noo��:�4}3cb1��M�������W���i�?��_�mS�C����gR���Aymk*��P�?�t�kL����?��B�x x���ف��jR����%* y�u�SH`���`Ƃ�I���=��PF�J�qw3s& O��d? 6������X�W�h�I!~��R�-�bC���e �St�i!��p��9�a?��>�����#���\uɐ����{�'K��j�al�i��-��Fa~��:*M�nC���jWz�J��
���r���Eѓ��8<��2R���&�C��f9�k�7P��4M2��p }�BL�B'�~x��{f�H�٤	����"��s����{I��4�Fo�K��p��:�����d~�Һ}]�d���P�g�*�@f�zҸ��_���B�|6@�Ŧ��dxF+Un��t���f�)�M�� �wo�~I��,��Y�3]5��d1E�8	 �.�NK�	[Z�q�[�&�����\�w�Ղכk7ڳpE��S
�A\ V�"ۉk]���D����zFH�TB!�x�YN�9-%Xnǣ���1�����q@�&3%�q5hΫLB���(��^�i�%hg<�����ɳ.0���S-i�:�6�a��ˮz"�mR�=L5�Y�ǿ�`�k��-v8�9@^\��~&�i����R�j>���ݰk�E!����Q�I���:�':��H�O���L��s�脡@����ۀX׽[v�Q�d#�3i��K�E�|1N�����Y&7����$}�L�ͧG���������ʒ���0��T;x�5Y���D��o�	u���l�Q�t^�Oխ%�2{���,�r�d��a��� #[���F��s����{��@+���jz�ȼ��v�F�����'�����dc�I��c�U?0:��T�=<�n9v�uN�T������ʴTo�>�ty���Z!~��	�?B�Ȏ���;�4v��xzY	�k������
���h�=X���!6 m
ڝ�D�(��-�_z^���:����E���E�W�}�cIq���f�Ud�^��U�[�Ka��]N�a���E)���e[�*��"�����<B�l�%� �Nj|��O���ʑ�f�5�׾�Q�˴�/� �mN�9��BQNՋ|�;w:�K��y��j�z���Uۮ'5p ާk�͈��o�h����<e$�g/���OA3������?�E ���6���[:-KoV�;�B��)�9'$��;5'捑����vЄr��7�S�1%������{�6yB9v���̽���Su>A�qo��}�Iٵ&�y*R8�o�t������z�����|�g��OȬ���H&�� n����"еGӇ�,&�i��vvq�Mx�_��T��l��8I����}�De����i��ܤ��Vʙ��m=�7i\��[�?�u��3Pm2��y�	��YY�&��fS =�wL�R��	VԄ���(n�fC���=g�Gwɉ�{	�[e�,� ���}��l��@A���G��Id�۠�:��=玏���c�J�O0��7K��hPH�b�񁬴��~��CY�:;�1/ZmsPZo�Y���Y	3={��y��������ےR:e޹45lv�ĜDQ��m��F<R�����3L;�ãGE�3Jr)�˶T­x3��+�rk��$B{&��I�c��MR�]W�⚑����(K������FP2��"���kۧ���"���p��a�$�4�B;H6+}�Mf�������(���a��i��t׵
TkԄB~���>y�K��3�@r/ʪ��!�-6��!�a���T�=-A۝4��.� '����5٭�W�3��9wB2�(�4�i����ʵ��=�0�2��W���h�vO������b*+�TI��*����. u/����8�����]5����Л�1���g�K����̐���o��v�{��T�EJ_B=^0il,���'��tx�gsq���:[��x4w����݈B;���B����h��E���l'��|�!!��������E�N�3�Z|���������;V���Ǆ������B�tfא�����`�-���1H}7���=7�k
S��U�)NG!�����o\⷏�x����w������:Pi���J���b=��i���(� q	�B���ӝz�VE
I5�i,Q�n�?���`A	�^�j�fܰ�JU�^X���D�|��?^��&��$�=���/Մ����̲���ޞ��3ѫ�G,�yG-��m6����x�#K��J��Wk���o��\�#����ޣaz���~�bTբ����;�zV	8zz�5��r��}�8r#h���Y�I@ >Q7��:1F!BE������>F�{���}c�vb�����0ݬ����)����4�PC������$3�A����E��ڔ�=D`^L�
8��o��c�ZW�08�V�^������O���u���e�m�i�9�!��\0��F�П�*\���	Պ�7���o1���(/l�w�.��'���h��;s��ee��G���DTE-� �����3Bs]/�����8Y'�k�e��6�@��A;S>yH^�8���]Ye��\�m��"�/�aP�9�V�+��a��;^��� g`��G�y>��:n鲩�i�
?����̏
~�6�oNz��\�\K6�_IQ�]���ϡ��M	��%�&����G��]*�g��z|l9,&M���gJC<�������A����E��\Ya���k��&��x��QU���	!Oc�= �I=�\��B�4*|���#��fJH�T��?{̨��F�E�ce��)>BWzO�1���)����1�p����f��r�ޢ�
ٽ�z:܌#��/�y�����:1t�r @"�=���w���K�}�cB���[����s{fm(ك[�'
A�\����xW\FdB]c�vt�#wS�a�}�9{4�ߔkAShq7��K3�i��dO�Z<�f'�T��VZIq7Ľ�t��Siډ[g?a�n�C�0`4pe�  u���e�:bQC�c���(i]]V�01pY��4j ��n�
&ӧ[��'���#��[��Fw�YIB�x�ȸ��5΍��{l��k�(>�@���ݻ���^1|�ۂ�%Ԇr{�@�G�m��Q���S.=`�ޯ�kX����!�.nF��-M↉����^����Q��s��~0���/Q0�`V��p�t����貕�xr��#��Yؑ�p��B�V�QO����nn�P�yg;Rh���5�B��7�ı����g�6�^��$ä�ɏH��H[,]VzS�_�����c(���/@(@����a	v��{�7�����4� ��#E�{m�6�o@��5���g�."ՙh�Rf�4w�"�j"յ����n�0���"M��S=��E=�^�}���3�C(|����[��/�n.
\9�Θ�H�=��N�(^7��q6��~���b�I�Ʈ/�V��e�d��\%OBO[��Rn����ځ5�0�d �S�޾o*���s�d���"�f)����93�1'�}{�PGX�u�Z���s��y��4^%�)��>��ظ'w���/8P�1iy������Ћ` �6��*�ُ�+��>�ykv�1O���5RG�PK-%��0;���$��/��{��Ц��wn֭;[��C�iV/��iA� ����sۺ�d�n���C^<v&�A���Z�ڗЌ8��;�"�u�0dO�<��=�����2�+��w�5T-v ��0���.��}�d#G"v)�ve���{�Jo��3ׯ.�����<�8�
��lb�0D����_�c.xq&9���r�(5�R�b�A�oikdt��tQA�q��I�2�6�<�C�[G��೨�a�g'3�Ej>�zm~CFF;Jڌ��6r�k���i2��L�7�A꣩�-EHOO��̅�Ƅ��@�]oVIf;��Ari �(`J6��J����}������f�Qk6'�w�Q�:Oc�����U�*q�L��x)y��<�:��A��u��Y\�f5�b_��q�p��#Ui&]hp���R��b�FG�R��ƌ|@C�	�I����2����/i�D0-�D\�"���X�x�ygtK01�I[a<����f��
�ɠ@������ͤ��oaWh��/D������"����mC�d<9���3������#J�e���>�M����R	�@�5Df��z%��w���F���'���~ q�"�d4X�F�w:�SO��{�O�Qj4ىZ��[�ر,�h�ޜ�v�s�u[�@L.Rz�w����(��wdoWƎ2�ͦ�ǮB�/�jU��r9�Y٠��Q<ޅ�pMT<z
(��?�j�T�*A)]a�j�[��ggU�n�F+x��8�u���;�p�t��-1�G`<
�kl�*�� 7T�;�6�i�f���n�h��g�-���^�m��a�b�+�=�f�y>VM̜`��f�X76߃�M�_��1?��q�C��6�Ũ���C_DL}���Yc���\�l{��}�n��(q��k�̜,O�2�{�[p�i5�x����.�\j��$��)��P�0o�*���Y��TO>���ꟍ9�hā_+�_y��3a�����C������ug:��![1}i��^������^�l�	�e�4�����d�\��+����E���]���h�覗M�[�f:)��;�����]�K�C��v�"�D*�3[��A����62�����2s�y()_��N�sԤz*����6C��Kf��`���t�V�ޯ�,����T$4�(JIe
3ÓE�>`Ni�@����q C��J�5�'Hƻ ��u!�٭ڏ)@��A1�Z������=���y����3%a{C N�o(�4�🡾]̽��}�ɚ��v��b�B��3NQ���1�+l�a".~��i4�W��>�z�/h��T���|]�s'<!�6�;:�"�LYY�&V�X,�%�=,D����t�M�6�28���ҾgD�����7�Z>���X�	���<C|Y-�`iZ$޽�o�����m~��W���P��R�ͺ��`����{��};�J�|�+\�P;��"Nάjn�D �` Ϡe�Z޴X��a���0�|vϞ�HdÿDq]��0K��7G���q��m���sixun�[>�(,�����$V٣.kʀ�}��ؗ�x�N@o�%�Ztv4�5��Dk~5�Z���B؊O$��#�U1K.��#`uC�F�B��(��S��\�vy/�pڟ�Ѵ!�����-L�u��.��J�C�+�*�XAs&��/PȾ�&¸Z�bu�w�8�[X�3���p��z����|�[��� ��{fWLР%�.����V�kI���WY8魪���H�ɣ��:�k��ʫ�G��	5�/@��:����<2�:�z�:����k+Mh��Z��47� sf��٬�nA�X��� ]��Y��ƑH������"¿V�yvi�N ��(�]�Q[�i�,J���'}�YV>�A+W9�¯H �-�L�z�}������p�_T�!&��:�j��nv�� ��l#��F�bk�~m\ޕ��q�<��Rk�xF�j� ��Y�Y��wE{7�DEX�K Xc=�Zi(���~-�{�_�eL��,��˅��R�m��I<�ܑ%ΒD!�}��]Y��)�{댕H�2�ątI�lLb�7�}��w�=&������������R=�=�s�C�v<oH��8 �����L�� ;g�;H�����l�Mf0ki��&���41�ޔ7�#��L�v�U{23./`��M�B�ql5}X�(r�u�����z�F��T�p`�@FX��L��6т�O}��M-�k8��ds�\O��"�~�k�5��bI^��sJ[N���0�;�e$U6�K�ViȠ�%M�:.ĉ.�bym��G&�M$�lY��\U2a�]^lb:���n�W��-[g��^0��B�2�-��i��SF��rɿ��I�%A�\o	50zT��q�QI���ӎGpE��ς���k�M�2��{N������m�.�8��fY.�5�O�1�bV\�s�Y:@��~:}�l��\h56�0�k�^m]����'<�+��#��B\��'��0�t��}�L�� m��$-*jc�Đ
�8���J�1�A���þ ��W��ndX뱶�ElN�8^�5�f����tr\a�+>놃5�s�'rw�����q��g.�#�*�w)�v�F�]���@�w��%H�(u�ޡq]ɑYqY�c�TN}�|�S(��ɍ/ �oa��X�bol}��?�y +��������g�d2q�\3��JP�g~�eBRi���%��[h�ܒߝW?MȏT�.Z����ۭI ~�Ǎ �_���9��ڱ��H��Iw�{ *a
�*��Lh���S;���~��<x�RA�ТscF�pA~�@Y-��Q���ۃ�Z9]Z��Bd�ȳ���?E<3�#�E�UÛ8:�[�����	?_ �$=�%)�K�ج���>#L?bΩj!A��`����w��<G�3׵v�_�s5av���7z ��>��/�
}�c?�쪞Cw�ZQ�U�x��YPZWq�<,�Vb�-�1.7�B�`���f��-"+=W:��'�1�۹�f����j��vIЃ��,$&B�#�Je%���<ä�M0�\[�'R:])g@�F�i8�q*$��d�\��2�G�s}����V�=AA;�`���f4�8�iF����~bNܾ����X����ħ�W^���x{-�3�:�|���h�،���ܣ�B�S�h�R��H���ڐ(B���GgU�H�x�������K��T�W��\1/���fkޮ��g:�Z[���?��K��a%Da>Ŷ	�ȒPy�M6�>(u\ڜ�O���;Q��b���a`h�cc����+5��U�<+�#w뻩'�Qf�zw�ճ��V��I&ɐy�|'�Ь\R(?*���!�4�M�Wf�������3����"�%��Z�|��)��!ck���B��)Զ�.<��^���5rT�\0���L�.�7A��|�jNa?Z>��UE | �1�_?�*�A�q:2�-�>���w[;��#��͹ϗ��X�@�Xr�eWG�~��:Ί�x�{yWB��[q8)���9~�ܤFM��Q������e�V������P��&�]_�+�v��	�_E�,u�r�Y%@~z�����vvv�AmpYt�1�sY��o�,٬��mWj|���+�W��<���v$v$�G&�g�e�ZN^�$l�D���Q�˔��g�S�A��&�n�G�+c�b��J%��s��p��;��'A��m�~;AN2�����+�*�2�r�T:\�2���������P�`�0@�NN^E:��v"�1\߀?	sM�,��W^�	)�N�?���3�(U̎ZBQ��xw
�u��;'*�|(|��'�5`�4��1��h��y�t�,?X��^Ɇ��v��1$6��I8�1�*��I>�6#X�ɗ�x�aD��-����m���,[�{^�o��BE�}�u I���)�yp~"L�e�	0�BX�E���*y^����ol��dУ���Ţ��������Jv�2 һl��ߐ����x���jĹ�B#��K��9���{\�\.�U�6'���o������.`š��g�X�o%�w1mn���+�L���|,T�]Q�e�G���g[K�c)�)+�a���	��aנ��]�\�"��:��ZwS7y<��LHA�����ʄi�ז�2��		���	��r'��8���n�� V��4=��j���f$�_u"c)�Q����MGs�0�D�Xo���yh���k��%l��|c�+z���`} e�p��?{PC\�-��&~���^�H��T����h���Ɠ��7�KqK9RT��x�M;�����ڔ��'��tkZq�+����$�t]xvii�%��|~����k���[X��ٽY�76�p�nqV�Gњ
��å��񓊉�ڂ��7V��ΔS��=R��k�Q�EՒ���+	B��'i`0�.�zc0^<�SE��Y�v$��o69|�-��0a���:^��<�����#���4D��I�F
�A�������tє�i��r�R������:�êju��ҏ�����uy�n��&V:l����!�E?�_�x��˒Feֱ�hZ������o���8��.<���N����e���ZHKqXk�Y�y4��)��^��㶣��Cn!��n����U(�@�[���zm�E���h�`�C�d^��[��	�k(���k��C��Il��U�!r}N׃]7 b��J�sL��LL� g([O��P���]����͎u�J�7B�d�ת6U�I�z�e��y��m0�EM��oP��ۇ���W6��.q�:jf�(�b,"�x��,㿋l2��1L������Z9b�Q/O���o>��%���m)�4*?����u['�Vʇ\&��y�l>@t�4�.�c�9�A/������X/nϾT��2?tW�^��%�hK=֞�b
-P
�3Cdz�����{Jwio�G���3"�3x�(�H��!�^�| ΋���e-..�6;��X�=p�¦^×��.����ԃ��#?��Z'\d/��rO�=���#z�?���I��]�s� +[ظ\�p�rL������%�pkIZUyl҅�����DC�Uh.��"�r)��v=R���+;Zf�=c�B��=�X���*��YԑiF��K�� ���$o��?�`��fMYj�.������Ƅ|e~�iH�Da�?�AB�C�_0������c�2�a�����L*f�RU�@�=O�\5�Ǹ��3�Yk����OЯ���D�zz[�ɀt� K�vn�d�'���aA@jZ�n��ag��P�I�a��<�Ӻ�N�!ٵܡ�y^�V/���6�|Ym���0��&���o5����]y� ��F�2�?�X��r�!^�[�)ȿ�(��?�q�)��b� ���˞C	���n���ęZ&� ��0��'�}K7��
� $Ѭ6�i��T6qL���LA3P��@����TĆs��dG٦����AG0:7�8vٻv�^i�_�o��L�Ay@��1ϑVYӓ2��ky\�S��ď�s��~aQ^�t  $�]�X�E�����Į��rԐb��W���ʾ�O�s)��Vk��@8%��ם���D|�����>��JH�FB�$��(x�W�Um������@�X�h��,1O	5��1P#c�h56���W�'%�6���E7� ���/.���Ǐ~��oE>[]�#3�w��[]W*�;��,ή���V$'a	�4��X4`@�� 0b����@�懢Vb<�ǜ��qwɡ.���/t��i:X3�TE��)0�;{��)[5�Z�������!�Z[�󸄃\W�lU�4x��Mc�jǮ|��h��wj�O�2�LwY�`��*[�hS�y��R"<]�Ѱ��^���C-Pk:��젷{9�6���5w�'�s�җqF�m	�j�-�珛�t�4�B�O[}�m:O�Pj�.�k��m�&\�ExՉ�Θ9W�s�~V���^H�.�[.Dc1��b�oZP���w`������D���LH$�A�UM�}v�36��`;z��@�6�$��K�x�n  PY�c*�R�Y�x��]��Y
�xmrֻ|z>�t4<��
,]���ڿ��XLU��@��F��:�:�|�p���|f�6 �9j�f2�tݯ`IGp.o���N	�����eތ�C@�K���D.@rR6�ȭ}��Py<�P>������%����A[[V�O�C Dڡ���X��������3��45�j��&sL�um�.a��g��p��d� 
Z�2쉬 YHQA�ۦ;�� a7j�+	�[�՚r;#�9�9q*����+n3����Ӛ�;2;ǵy�|�-�۔�By�;~�0]T/j�ӏ�9�ۛ$Sa�n��|�ḇ<'�*w�$�p���-��f�̳�g�,r��v@X[R\y{����	�͘�.p�=K�a@I6�No(�N�z�`PD�O����'ÿ���� :��iao�ʐ��Ŧ��&H7�F���a��ｋ�^>���tt�����v��G)K%j�I�y��Bb˶��ǡv"#�z{�j�2��*ۏ
(x+o� R���vH=�?��Tg����GB�{�̵�j�ߗ��l��:u�tW~6܁�[z�'6����5v)�{�3g߁[�A��e��;tܦ�tTZ��D���J��$8V�<�p ɍ#*˭�OCE*�<ӊ�iD"u'�����F���U{��� �AM�R�q���x��!�qtu�)-"F��|��[�����|�SW��)@u�o蕖4	A#�Q���7�۳��9�M�(D���\�Ƈ�f�~N\`ilb�>�sZ*��J�kFJN�G`����~(��e��������/Ի)y�����
���_���	,�ǙI�c�v���sa�D����Z,NbX���w�k�.�Z�V۔�`����U6��}� ۜ���5�~жp!I�ܝz@��n\c�Fa�)�ֈaU~�9�6Y��J�a��<���u�B����ȀƐ*ɯv�p�e.��6��#���[��4���v:u\L� ��S$e뎦5���ͩq��(a[h?�rd��� �I%�g�����ѯ<���O-.�~e�����+B����o&O�Rl����~�(b�u[�ɇY�g+f����^\�d�j���u�ݝ��n�+�u��no�H��/C޶ e�B2��lR`I�(6�&2VpH�w�,a|��� Z�]�L/TO"��@ҟ���6q &��@�*-�����=05��b�1Y`��Lk`4�@b
�>��_�!4'��^��r�4 ܍U�Ad�5��V�����d��ħn(倳�0Y�m��z.7�ߤ,�h�����ni���.�_+���jeg��r���Z���H���8�K�H����\�I�:�ZN�"S3���+��,L�g�F�ee��
�������� k0��>dK=N��T�x�%�?q�'�L��l����?�M7pH��JR~����GyG�F�W���L��x[Q��ٹ\������>�7STo��٘�<��S���Cӭh;������k�{�T��H�;�}E�D�!y�)M����9�����Z��O����:!z�]_r\���\WdC�B9�r��̻�+��������F�$��%Cu�����<4w6UC�Ur�v)���(t��_�{O~��띪�nS��{��>mo�v%�L�*��֌�������Ef	��J�X{�� �q�5�	�S�I�Z���13���W�I�M�՞L������p�9��\IN��lvp��n(�_��4RP��-İyUj�o��OZO�HBS[k�g���9>a�������Tg�n�-$3�G⺩��,r(j9ޑ����Q��sT8K�H���p����~%z����S�`��䎢��`���!�g2��ԥ���Nܧ�꼪l�q��w�q]m�U	go����`M���F�')}��mJRQ�;�;-�~#`|�hC�Ti\O���X�٬�����2�y���F���Ѥ�4�z�_�T��;����{4K�Vy�3\�a�Z�l�c�.����r�:rl�Ĵw���?#�$��$co%������_�N��Jqד��g���j�]��u1A+�Kka���G�p�mRz��.rJ�8�P�>c���W�%!��^�װŎ>�!N�MRA���u'��b�C�1`OFU8i;5��A�<<.��_\V,1C�V*��)���� �����H��7�<2S(�L���-�U��l*����*�h��/mG��/��OWN��ӽ���KdPfZB(E��K�-�u=F�{;y�2dBS������ͧls��W�ާ�Ky2Z����ry��MFܟ�R�(JL��z�ߵ*��A���Q$���P����}��O�9���.d��=�>QĊ����>.�}&�SD`�0Ă�f1�㠶d�mUs\_Ki�����2n�� PвG�?�5��L):�Q�p�E����r��Y�o]��xq������'5>o�V�6^/- zg�폩�mo4�?�-WL�	&)��'3�T���%����fZX���e������@<��l����ǐ4~%��ܦR���a�y�)��}�|�V�H�i���[d���d�@���[���F����O�5�E��6�'_
��,�럄��3�����x��N]YO�`GX�a��H����GrHv<����PU�+	�s��PjW�ơLa�-��u{�u���b/)عRx�����;�o�1ܿWa9�zAͻ��7L.ݯ�j���gcw��]��u� em/�,���Il�� Dq�%j���npXlFMM���s���QIT�UM��������2N����t��T� _�[k(���L����]Nza��<��p�(i�,?���̐j�z��3�*L�Ά�!�c�Ȉl�W��,1�9�&��?�1��U�A9� ���?���j�p�9UCЅd��\�$�yXt�ځ�W"�����83�̘�' @q�e���\����{"��ߗd�����ߓЇ��e�!1Хh�	�2�誚W�jt�[$,���>�����]�tND�Wp<m��a�bD��d��q,>�Ow�F��������yC	��F��`Z^�8-����|_ �v��=\$�W5���x8.8ǙnBB�����2�Fњ����,szK�e��E=C��/�<�Ub��c|Z��RYp5m����̌X�������D|�!��Dψ�j,�����'�����������=x�;ڕ.<�%�8�Ŗ8�:�+%7��+,�.����w�2�s�u����S�ԐNz\c���B�f'n^c�mc� ��oOw��R�J��ݑZ��!��V.O}y8�q���5�ԇ�X^��7��xÉQ���H���}�m�QI�J`�̈́k�j&����i�����99�D�����1s��?�۹6�S�G�^��f���,��.�k\��˩F���8�n��p���L������N6zAJ"L%V�h�O�z}�*���w�>��'��
���u�(��e�~���U�M��E6�4�K���+��Œ�����b"���,Ճ w,>6f	ֹ�Z�D�H[^�.m?}���c�J�V�|���V�("�Ob4&�� [}����S)��$����%��x�)5p�d,y���ᅶ�̧��T�l���t�Y&+^ן�^-�Ѷ����|��v%�M�xoen��=t��#�p_p	NO/�Z܂�Z��<�-BXq��s�\�jE��������j�m��຃;�Y=��Y�B�UxZ��� ��&�N��FL���^g��+��8�J��Ʒ+o�9�[T�tM:�b1]���}rC�1X���Jګ��l���	��+>��Ǿ�q���w�p�jU�)ea���{}���Y8�h�O�g-�V���66�v��k:�$Q-��'L�F���5#�!W�#tLҎ�`�^y�Y\�]���u������|�y�i���ɅI��OqQ���:��M��Y �8���Jc��k�*)`�ʷ���+�+]��>�[55��<�)�
+wr�����Mm����/��QH�����F�e#��)�$?��',�O�0��F"���*�+_:���6:����Ƈ�>������,���3ِ�<����r�N�[�~f���2b�7I�MZ�d���{�!��Y�r��Z�y���
m>5b�KvD�G�[T��X�����0��l�B�6�s��������B��œ2�T
!���k��t2��fE0)�7-5��5��ɡ���	���	�aSɌ���s�R�=C��,K/xv�0k��n�~�X@��'^]�]>%\�~��`�҄H�U1����U��Fe�2�`YB@X���\��H*�3�����
X���X� B^��Mciy7�~�0w��m��&;%�g���ح����é�+}���{�?7�{G��(�O��%��|�`جE�ZH�Ʃ@֮sv��DCi���k'O���n���^�G� �g��aB��sC��f�%47��9�s7�s��2-)~�#����ê0˭ �AYq�jN*�K�L�~+]�3h'���h%�D������w���s���ҍ�`��Cd����Y�md��]�đ�����#d-9`���^�W��.�����63kK��7�~�)n�xϺԭ��.��~�e�F^r+���= �t<��N� �<�6֦0;�E�f1|$=�ĸ�d횜���J�$�vs�q�?�k���?�
Waj��a鼟�n� �g���u�hJ���x ����ۘС&��P�@!e%đrc	a��u�/����:����L"QP�G;S��>�>�7��� u�j�]�(��g8�����T�2&�`apX���ٕ� �㭌q��x+���l�B͏g�w�B[C�e��%v��GN�ZbMCԥA�-��lP�*�whjU���V��>�I�oof6T�Q#��0-� =��/[�}�<7m��b=�.F\�|D��}t��.��;��q��#�O�`�d��r�� <�p��Y��5��RE6ܜ�;^#Y����^x���C[AupW7^�����l6esQ����5m��
4awU��:�x�_�C�:6�
�w�������S%�Y;wnW��1ӿ9�Eҡ���8��|�,.�'zXG�K��2&u�$��	}7}��X��R��W7k3"y#�mQX�����N�*�]�k0Y��C��U�IC����^���ĥ?�8�Z�A��Ȉ��}���k�CSa�<�R�؋?�����26ʍTX&M��C57�S�QdT]�9��C��n�l�c��ц~�f<E ������n�#�s�aO�Cn�glR�"��Yݸ7!����-݄a9u�,�&`1�-���'��!?�w��ڨ���v�|���9��t;��z�U.W�����S�z3���#D�L���ڄMM���+ݮ)R\�D�����m�]�oo�գ��\�2�m�\����3��1Nv��E�	�����J�=���{���S�����"��P1�<���'�hx+0}�Z��[�$s)c4��������'NS9��	 ��@������:>i��[�ّ��_Q��.�@��	�	f��̢��5�G�9��K%~�c13O��&S�񠡪�m�4�m�ҍ��T�A(//F�΄�1�H�͡����� �ԅa,gZa�]eTg��z�eߙ�� Ne@�����/$U���}��/���(�{P��ۋG��1F��8BFZ���X�
��jZD���ǁ�T0�Z�T�%[��ߐ}�ҬÉj�6��������L0�D'�:�f����n/����|@�D��X��{(F�*8,/'!$��]�m2ܝ���E��O��X�W2Y&)��@����z���x�]����u�*t~o'�=c� �'�ad��r��d�NV�<9=�D�p{��Iy4Oe@�e������w�Û�dρ��mڅ��Bu'���3t����$U��Qֶ|��ߑ��Ӣ���]m���먪�������~���F�B
�G�tv�#R3�ƴ9XtƘ���3UO�4�I3�K�S?�IQum���5B�̹�#6E�a���_?z�zK���G��Z���ݧ-�B͐j���K;HM�pu�o奊$8���a�w� ?E�
����L�����O�E0#'��Nl��u2r�<���D��V4�!��D���h1�G:��K��[�Ӄ�2����ւܵ��]��S����%���r@��eI�ΚO�������4�YS�1�����i��Qш�0��GY�"��ʕ��Xc?�;3�JiP�_|����<U�Fpf�}Q,�ԕaz���Ij��⑒;u�>cj�|�q��^���k�m��Z���]p(ֽ�h�0{�tn'��:9.�m�c��Y��T��<^����R�0Xu㮶�#k?���ٳ=�'�9@��m�\,`��j�A6�1��	?�Ԙ�ֈ�ᥲyuy⋔�Kǰ �5r�z����?t�b@U�-��{�sN�yp�
_����d���$����$��Y�O+����|�_�X����Ҙ򾙲k�N[�Lr?��O6s����4`�/%���l�ern$=�+8U��3S�/?�8殰�ЭyN )\�q��;�����ӣ���:����Y����/$5�F�ލ)�&tIzvP��5���n�-}��4qv!�Z+b�?b�� ���������=�iK�b��{��9��!`����	�kv-�u'9�(�a9�r�HC}�L1]��(��$�֠�Al"6�-٩.�Ơ#��
��ֲ�J�œe�jS�����-�$E�t���q(m��� @p�����i4�#IΙ)G�f[����ƍ..��F������8_�8!f_r	6�hZ�/�8�zt��lb�QD�5.���̵3�����ɮ�.���̿aa4��$�bZ���bl�����^v9���t���@����14��:�
A^�a���/�����!G.�Ec��'d���vZ�V�O���x���p�ק[�ؙw�[Cc�ýػ����;r��z�cQ�T:d�uO@�&rų��� 5��8���4KD'��N8� 75��/k���}�\��*�D/%�]8V�0�P�~N@�I�U&���1��b�Ft��N�X�v@�P�������ȒEz�"��;��M�c���2�P�lj�� �v���Q���}S~��f�bʪ<V�ʨ(\�;\���@˂{�#S�"�]�*���pn����1'!�'��"�iO���{F�
I�ɯJ�g�C9W��ZJZ�=�� ��N?���X��!��!��蝦�ꚿ7ٛTّ??�s�S�a�;��G[T��82��zQDR���! �� ��Y��$(���$z��=��*���T�7���d ����[��?�No���f���O��$�O�m���\�}����O_a�ai�h+�N�w(�D�Y5��O����M��%�f�r��[��G�ܒqO���m��+�d5P[QK��V��_v���.I����YXLq���Z6o�/����~ۨ>��������wn8c�+ǝ�V$�6 �v��[Kڏ?�ك�#[����,�ɸM)"�������{�S�-��eL��d#��>�Q1k�������*���(��m����&���# �������qabq��X�{�3�"�S��EE
��ථ%l�V|~����P4���z��pW�^��22g3�o5����_VGP{mL����wl�Ke@M�>��U]��5����.�04B*�]��bnP%��~�>�������#���"8;����I��6�6�ب*εw��uY��R$�v��U��N�xj&�3^�M`�a�=�c7
BZ�Mw�����F�,�ͻU��Ĉxv,�j-��f�F~w�����Ѱ�ۉF�}�����К��ɤ��c�5A���@I��{6I��<�Vp8��P�0�%v��
��8\{]f�t�߲v�N��z^�
pC��/�y
��+s�B��>�{ɯ��N��c~�)����9p�������(�<D���w��>��u��Ng$���"��X��x��=��/>���� ��g"X�|���Y�;}��n}����v	��8�g�FE6A���*r�1�S�<�$�d`�Ya{{���ΩT��l8c����%�\i5<������c��rq�uV�qYG��VJ\ݚ��:q{�<0`�CT߳��P�A��+L��,G�O�eeVԖ�MJN3�# [	���,rs�&�uq#C�Ӄ����_߆o( p�#�:&�?�Ըl��Z�-wW���-���깋��9��|n�Pf�A��3C�c���O6��c��8`���|N�U�!���'������}��{e��y��ډ���|rJ�1o�6{�	D���k�3���	m.�4/��Ӱ�*����h�)���N�&H��J�`j�����c�6�^8FځN�7���g	� Z>�^���Nք'��X�P�3�-�j{(��0�Q�6s��̒���#�n�D�ļ�f?�wy댛QF"��@L�qK���&��G�+%�6���RP����S{�$�"<�T�4 �?S��&�ۖ��#�_�m�d� ��GM����:�nT��q6����f�~�"a�k�Ц������6�c����������o�f�KΥZ�e,�y�����g|���
U�Oq��ƃ����⑲�6T���Ch����k��(wr��j������O�a���D=���26b�Rg=��4-=��R�>��9�Q��6I��o�M��sw��'l�*��)�K{�����m�П�;�mq^r�۫�� o������x@P'�&7\�A5j]#�mO�t���1~I~������k��z�;y3����@�W�t��͏א��+z���Y;��l�pv�׋.�}߆��~Y
ነ��[p��J��C$s�LY(<��-u�%W��_��� M�s�L�{Y�"�oP������5~Mz���MO�"��{�$>xWPk�E|�C��z�W7��H��ϑu{�Ã���	���t���~^�`��$J���iWf0䢰_|�wͫW�z�l��	ke�v���bÕ @�|�ZIu���h!#W pHϵ�"����� ��۴d]I�F�O ���F��%M��r���@��Y�!(�}h�⍯�3�6�P������j-�][�������Qec��d�����+�<5��h����������o�(E���;�:�՘��(��}��<�W<��Nz!��̝8��2y�Ã�k�+	�L��L�%M�b��?�5�P����cY�����n��>��K�A�'�W�.i������q�s1UÐ�A�fYX����_?�[N����L�&��U���V����,��C��"2#���	
�!�5N���mIi)h9��x����d�-�RZ��ߞ���<���r���T�6�����{�'S� )�؀�B�-�Ŧ�9_B	fy7����R��Rq�M��#��Q6�(�e�ې�M{��Xi�O!(*��|��ah�!����	k�y��֐� �e�/_�RMlnR��  ˯����i��̾Sٿ���GP��r�O��	�[����i�_N�C����U���p|g�E�ס�1���~x��k�{��T'ޯS��h|�.Ke����]J �8>��wd:<r���#7͢6�rx����������Q7�s�V�`�;��E� S�
c������o��*����i�͸p����6�y$Cnr:���ɬ��b?���e9�2PapO�Co(# �g���xD���̷�&/�s!�i�U���ޤ�BQ��'��W�=�����[a%����[�̈K"�`h cڔ$W�%��v欘��+�j�P�$�%b[����,e=?�jF�>��j��ƼNV���7���,��5��^��׷fK���2����� ���NЊ�f�f�i�t�Q������Ev�b
�.���ZA�ZoK��ҋu�����;�{q���~�^K����@j�����Q	�p -�v��(=����j�#��]&�w�_������d�^x�����#P��/ڠԭ8��m�v+�X��}?}O:�MF1�![qbQU{w��>���-�J�;O���G��Ô	VCs1o����*;@"�:t���x�1�ŗ �1��n#����m�ˊ�hp߮��)����ѭ_mU�!��8���٩�\=�ju��4n/1����1g( ��DI�e�7���;��e?nmQ/\��e�4QW�j�r��Z��v��}��M��J��4��'*'���C�:ߕ��t���c��B�nm	\xu���Z[|`����ҵr"q�h*�UR�����Ij�t"��a�%0i�5SI��|�;ⶼ=�i�A�����l�ڬ�/ c��b	װy�ѪpƓ�KE.+�%ڙ���1nx�5��)�9bRV0�I����=R��`�V�R�ʔ��I�c5�^Ywr8��V��-[�7�6,�S0}��.v�ȳo�ya��C��/�4��lQ���f�9ɀ���+���Щ���am��U_ĊV�7h���]#�Afq����Z� o��C�ܢ1O&�tT�]�R�>s���u��J��\��X����2�%�NY�h��U`���*`��]	�?FD)����z��|D�H��k���A�j�#:χ>~�I�'����>�#�sl�����2��s'�5N����D,���(�'�bY�S�>�����
YIZ"&Ă�6��Mj��^6r��*�]�_ 56S�ֲ^�Jͷbɺ��߿7��������$C��7�:��a�_��9m���k1��u�k��r#q\�5�Z����ѣ§3����c����,�K��1�V4r��qT�w�b�&@5�dZ����B�I����L��ׂcO�i�|�~�^�c3.R;������΋��e�T�M��Tr��*r=��\3�����D{&���Mg!�]&xZ��ƿ��o�^���q��J�BV*���f�}�&������[�sñ��qj�QR�q�7��4o�9���`^#�9����L�?��>�yZ��.� ^l���a�c����`�Et���;jT2�N+�;$ªZ��E�������@�.������俾6�ପm3"����v���)����!�t�ۮ��[�
�y�#��|�`�mWV8���=�̧��=v�a|��kl�[$XI���}xl���>��m_�� &ۡ҉����3�4���(�_<��A#��Y�9cK��0�g�P��p>������RE:��+98�H�Et��ad�_��SG���:�-���z��2M��k���1�G[��ݯa/�r�b_���@���.�����z"L3�@�%��	ޣ����6{�^뷏�R��d��pVB(!o���]P�T9��]�v����z�u�q����,��D���Q��q�\�R�C<ouT�1����/�����s�+.��;��Pr�SE�e�]�Ao+�J�| �������ʵ������t/�o)/�_���eF-Z�ܧ-7��i������.�iG���d��`���4T5�Q�|�����ů;n*�ܔ�?.{+{�h�#i(DlCA��Iɖ�p5�ѓ˭yIg���-t\�����BH�Q�N�r��g	�,�F�ݧ���`�X���Nh�ܾ]p�;�@�s���r��������D��H��G �A��F�jޙߌ�G]q�E��!MÍ�� {z�l��v|��ӄI���&m��1�+4�ܨ�eQm�;e��V��F��YI�1;���rL6��}�;=4ʈ�[�
x�%�L�k�ܦjPE�*Z F�Hg�����_�d]�AlP��=`E�S�����Eߢ=֤!}o��t)#��l�d>�_!����U!��k�K���zJY\�j��.�y�>7�L�;�Bf�>���oNw�E+�G�l�<�:�9�j��v�0�eOs��d e9EF�w�C:'�g�˅�$�_���_�qf;��s��Qoh��6�(oyݝO��o����z�#=��z�S�t(�؝���C`+m5�3}}��џ��-l�-�é��,V�� ����fjD}Ɲ����g��5(�ir�s��g��,ڔǖ���d��j����*A��/sg�ދO{:M0<!lԮ�}]P�	ĸՎɖ�Eڶ/C��wv������:���y�辳�YJ��/fj��I��Q���/BC�ZZ��^��w�6Է�G:��\7/~<eμ��E[�H�iv�BZ�I����t�䇒��f-k���e���'�e�*�6^{�l�
Q+�U���U�B�-P��;�[I�ă	��`g�ƵN�F��xXp�4i'ʘ��$���r��\�^�=�T���
nr�31�3N㊶>�AO�GV3i^L��ϝ��oh\> qrf{��	���j��~$�C(�[���qkH켞��?�K!�T�ieS^�Y~0�k�I��.#ܔ���}� Ň�2*ɐ��AK1y��Ɨ6�GQ���~'a-Ʋ�r9�m9G)�D��{��Qc��Ӹ�`�R��5RƳL�R	i�]�
�ķ���y�5�%�����X?�G����]�Edg3Md�R�#��2�mp��xI�$�С�0��)aί�Y�j�t\��+��Ia%�ob��հ$Oi�룛M����0��2��
]��t�e`�/
�PI�dK�L�X[����a�,��e(� �Cm�`�[xY��1��p������B&m�_N3h�s9�� ���*(Pu�\�d��z�w)�?���A2
4!Z����z-!p�c��z�A0]s]P*J�d$���(�9�g,C�/Eϫ���k�c����M�u�y�?>7��ٚ���t��u�\�����y��V����%#�'w1������L6�?�7V���(���9�E�uv��ì�äJDT����qO��S�&�*��f%���%5��3��ҳ�:�FދÄHnʽ�S/]S��7�U0=o|�h⽀�r<���^��`�7���x��~DR�;���N���V�u�d�����|̑1�ٻQUh�B4!�FИ_�� B��3�H��*f�$�Q4�9y�{��Ӻ^lLa�����m�Gbx+�A��n��S��3�Zb=`�Ck*�6a�A�?5`�H��.�<���i`�M���P�
c�nTF�i:�>�/�7;���{�I�FLf�����	���lO���)�~�B,A��Q6�ַ��P���gL�H��MC��p\Dt���<"��d�(����I���x���0����)���ɵ��)n�M�I�I�s/T�!���)_I�I��i��_x�9ud������~W6���:Cko���û�o�E(�:$)��B>4#�)�K��Q��gH�VN���Cu�hR��5hw���je��/�U��d���
�0Tϋ��qQ|h�������'x���En4k�Q���&�S#ߛ�t
x�ĸ��3}��-W��	Ro�	�T�?�R�&���?K��D�d����@9����	U㔌�,I/����I؍#;�݆����%=9��#�;��]�yl�p��Jb�������t�x�C@aZ��ag�G�O 𭾗~j���Gt��T�t ��W��#�\ڀD^U.�pl0�M��j��7ί��Y�xv4 �8�
�c%��������{�!��(�S��uW�azf��d���t���Z�k���A�b������K.��P�׆�b�HԂ�<n΃�35���xR��ogX k6h@@k�f|��+֭]�}���Ƌ���\�h�����#F�N�|�#	���&.�!��'ժ���?��z`����sI{e.�[�y1��Dk4e�&X8�����\���k��_��e��uE�&j3	���K$�m;s�#�P�����e�~beB����ʓ��K^�d{��$�ݡ ��
v�W�лq�ₔl�T�q��;o�y��lO�*d\|��" ���ӧ	QL��h�	�W���vm�|��kv��0܏b%iÅj�V��(������M8Ix�܃��¼G���C{�.���o7t8���� �M��Y���E��X�n�O�_��Oi��?�t<�BwZj�Y�{6
��,k�._�@hT���C�Y��?b���^^QO���Ll/26sY�����}G����{�ym�n�)�-e���yx�DƏNK]�f��T�c��JŰ�1y]K,�k}ɋuz��%���<����J��~9}�|Ԏ���چ��Fv4r?r sɡ<�=��E�%'+5����O�j���磨��y'`[J��e�x|g���s��ǹ1��
�_�L4])���h�-(f�dZ�ۗ!O���ȸ&Z��Ż*p���$>w�a8�PI�� ca_�e�������2�iG��
[�D��_�W�b���eE�|J��`{9ǌ*R��瞣�`;�	�A��w�a`O�fVm���l�ŧ]��(�/�$����.��c��t�/�7��=.K�b��{����	n�uCV��'�Ɗ�:�އ��ݚ��Q�6}�v�H��lV4�S^����b�y���GxŐ�����<:w$X�����Gd�LC�
	��J�Й���o~v0Ҍ���q2#a��I�������h��P�s��r��B���CN��ۏ�3��@�yb�A�OpE/b+&0l�+�YؑX������?qe��[�G���ĝu��u ���g���q�T-�����1����,F��9�P��8J�L�@�nU�5�B�v5�,����,�S^.`���؜8J`�׽@V��~��&7q�TA��ls+d�4���^����͚���x��*q���l�����{4�͌���`�&V����|�S��ňd����-D��y
�ݾ+�+R�;���1:Aّ�h�z��>.+`�H*�H��]��mUj�N>8��
{.<�S��f�i�qs�6�04�Ԓ���Ũ2��Z�*ȫ�}Sõ��Q�&\���;�ü
l06"����m����N��OZ0&U��bUOm	��g���f��C��cŕfY`<��s[��7��h�&=���6���l�usC� ��Z�>�d���C4��a�"OB9B�־bbdQ�;�k�mCtQ���,��0��wF=y��x�:�������Â��:�l��)���z�)p%)CGrZ�T�R7�E���[���$�vO`�ׅ�1'��AKX3B���)�3(l�7��/�%��Dm���9���_.��&U:p��҃O�^�>�-�2����;�l�k�n��C���z��~ݸ̺��)�`����)$�Z���然b&#a$��~���� T_>6�}��S��D�d@�P����:�_z_�Bx'�"�6�X�ˮ���D	�\�`f��k���ׄ�'�~���6C�gǑ������vI�ǂ�u��Q o�<�RX7�f1רR����d���]��֓P
�{���@,`�W�q�����b^+c�4>Z�}�my���HCƤ���_B�U$Kj��N�Y�E{���YS+�_ҕ8(���PR��u~�	�_ �$�
�B,�TD��M����Sy���]Q�ڑ���|��t4+7ɞɏB2��BRt~:�q���w٫�c�d�Wrh@�v���"C#'���S�c�xҜ�Ŝ+�Gۘj�9���	; ߩ�s�Us���Y�3蘛=`0qg��0Wc��R��~�;�Rrx�$
Tک��1�|�ٷ�j]��d���u���C	ߑ�m����f��.p��#��"��4�h�%�3�ϊz��i;�+zwغ���:���������8���b��n�k���脠��z�XQ��-��6�E�"�ޗ�M�$uc�; �m\f��5�I���D��(-��ʪg�6�� aB@�uˬF�&�Z�����>��k�!�xw��+h3��@�u�p"���Dx����R��k�RI�nH�g��)`I���ȝȶ�4[A>#~5�S�	�
�|�:p���g�ʝ�p�Z��4.�R��O���[��=Yq۸�O3� c<�̇�y�|�)��!�I:�R���#�2�Ռ0��vp��O���<f[ga��LQ\�,���� E]��$aH|��S #�
#:��Dm�TڎK�z]m y03�f��#;�>��p?� ���Dvqv�"M7�V�6	!�%!�v)���^�(ˉ����\�Yu�2AP�
9E�Hu��A��41l����m,��� cE�6�`��pBE�ճ����@��s/V� �R�_�7���A�2vJf�����B6~��󊴂�H�&kH���k�DSL�a|9�&>`�8��f�[��*!�h��^�i�EI[���X���w�7�ĭ��^#{oC"�.r����|Q�[X_gy��*Y�j���|�vIf�mG<99�<7����W
H���i�au�Y�+���˞�#n���v#f�bLqǲ�J�L{���������U�g�x�E��vJ{�m�fd�{� ��b��Ly5\��ٙ��h�X��f:=�ˮ<���É���<m��M�j�:�IY�b�����t�=	d��6��y�L3veST�>$��%�c�:�D��LR�`�W+*F���S��:�6+�;�/�$�:� ���6<�:7ۿ�ҟ�?z�xeP��jiBm7���I,������s2��P)Iǧ��^X\ol|�h��Z��TQ����"܊��®�K@��ϓG��rn��V���O��Sg�^^H�А;�8⣍�'n5x�p[��ቪ�#Z�I�����4{3�iz6l�վ� ǒE؍�+t`^�1�"<?)�`!
��'��N���j�ڢ�"%�S��2�K� 56y�0�i0�ư��{2��Ѿ��i}�Y�َ��"4��Kf���ba�3قu1�]�Is9x��ތ��h�n��Ȫ�C�9rP���2,8ktcx�v$U�=<������,x�ٸ,g�!���}=�K�r�������/���j)���${���~�aA�A�zA��y�tIi�1D�����S����J��hd�D��
�؆����g/��5΋�	���i�V�<�1��j��{5����n�R�4���oܷh���U���uI8�S�)����r)-�g2Ĩ��4|�$�M1ԣ���GVt���-7@;t�k�3�JVe1�qm��=9��W�8VU��[�����c�C�s��c��9^�7�o�۝L�8��D2l!dSO�	�e`!G=��W���B�Ύ�$�r U�.�'�p��h�F7���
�]�qsI4)!6����á6�"���dd=����T��c�Es֯��'�}��"8���h;3-3f�Gl2���g	u�aDBl�?�Ic�M�&��۲��p�p�lVX��|.��K*�ZgV�o�P����bvZ_��[���� 9��~��u@�ۂ�Fۣe�}c.N�$5n{B�����-�@
��o�^�k+��a�HE��z�,�R��]
�8�&c�Sa?�M�S!H�M!y��yB�3����$��3;H�nr/Б�*��>�/>�[4��D�B��]a���{vA�4���:�%^�������D"�[4[��P �|�v�Ц�j�/ֈ��o��8��ӭ��ƾ��-θ��Iɚ��~Y5:9Biӭ#�$Ru�j�w|�Uy�'>`���఑i�أ�枿HD��t�.rYJ��Dh]ąv��2��nJ�CZ_LG�Õ/3���P2�1#��A؁�|��K<{9��$�Է������L�]�t��V6�6e�:9ZxSY����h�4	./{#�/L���[j4����5�� �� �ϐ�&�Pw��Y?�չ�}i^��p��{��!cJ��q8���Nw����V�Orjy�,Xj�#+��#d�>�Ɩ���;ɯ|����S9P���Ę.�-ڨ|`�ta�����)u���]�-p��&�%͑��}:�'53�Dc�����he
@�^6�ڝ�Sr��(qķکh(xd[��zm�o�������_��`,�Қ�(�/�ӻ,ܡ|3O�������dYLپ������ ��-�xPD��d�g'*�+�XF4�*���|71��>��$9��!x�byz�U�{��/�a7㔩��ɂk��-�Tކh�z��9����f��~Tr��r<��߳Ӻ���d�~k�l���L����_~G=l���y����0�����:��>�X#�eQs))�#�<�i�Vdm��*�6u�U˜��/6G����:($�'�%���4�h���w}��?)��V�]�Q�y���M��~ >��������4F�(��!�#N����,+�	�����&Zg�D9?@���q�u������'��7����f�0���IX�B��y&�)+}d迢)H/�?N	��<b�R��k������,��v�{�Ux�q�� $FKiJ|������k�uf�>��®�㡬q�)D���6���A���T'/����qzq:?�������S��)�uY2	ع��M~w_R�ڽ 9��� �kD����bw�������'�f0���d�q�~y��W��	��?����=�[h�PS8-������{PH���Y`���������$�[WL�����co�.�F2�a�%+�L2��а9����2�9V(w0�xgfX�,��S�&�#WE@qp&$���/�����Ϻ�v���B�mgVouH�|e���tˎ�:��:�����I�RQj�O����&ږGA˨�:�me�0G��,��m[�=�0�Q�Q�6���c_v�RV��v�8�>|�\V�9�N����&��A�����{szt�~/o~���P���ޠ`���"�ļpHOP��'����\*z.S������fOR%=�#�p�ST�	6ig�ODt>��1��]���b�C�ĭ�1�H�8ؙ#����Z�!6
����\J�C;^T�Y[y.��e�6N��*_�3�
�خs�ʣ��������x�)ALu�j� ��,X��� ��ݚ�H|��{����0%M)>�f�2;t\E�����]�o�R��,�	7�������wk��|��:g |���L���g}��O�n�qf����0���(�\���b�a'��D��.��y�DMI����$�/�����JŔ����!3Y��`G�����^�t�Q��L���"ܿ?����>4��<�Z��`�͡�n*���g-2����b	t�@��Q(U?c�H��_��򕝰B�ݔ���kB��p���?�,;ͧ�{�|��܇z2���[��0i6p,)�����ub�r�q���7ߩ��;�T�fi";�����k��A<?� �?���NHIZ�'�+������q��2N��t�"H���{�;��͂_2�*��~��2����%B����-��JEXA͉���?���LY�@����˸�m�F��1� ��,���~y�J��	�}#�]�{p����܏&���B1�&@\}��M���į>;JZ7u^� �=��@M�'�A+lo5��ZVS�rґ2�,�DT`�BbJg�g^�ʆ��Sk��K�\B�/-��i��b���1c~�dݬS���2~�<�gށ.�{��H>q���I`�w��= �L��ܼH�����>yP1s�����YQ��ډ6]��~�EW_�+�U[T�pѩ��jo{�Ӎ��W�Ux�قeH�nj��"�����R�_e��%j��p
�'�~�^�(���m���N���,�щG�p���|Xo?��p��s�=)M�d�
��}`�L�)�pK�������*���6/�D�����ed	�ALԓc*M��L�V�^�D�f\�i+&��C\��H�s���˴����4���08GSI"ܳ>=p�c�)M��&�.q,nSv��N1���{��$
 1���)I�5�.����YRf@�SoŐ��=��6�-�H�"���	/2'O�J�;2�ϙ��+�/.{�{���U�~��a���xGL@�ږ��#�ĉ�ؗ��Q<�9u�r�,��:�M�:p�J�Q[v9��lN� �x|$�$�1�e9qa4�\G��D=��,�gE�?�w��h�˷��0T+[��9��c^��UE�]Y�()�����a����np�)IتE�мQ�E5+Up̰_��4(Y-M��̮�;&0샣�TS�����-}p�tV��{���yK�Ͷ>66�����綞�3�7+k��]���Z}�W*H^�O��W���2<�	7����.k^�t��-Z�R�Z�s`7��/�_M����t�a@���>?���\�1��+��"�V��zC�� q�}�<T�(Yq��L1/����"��  ����QO"�Z.@��Qț�0�����&�k�������g��2PY+�����_ C��g�I�3Rd�3fE�0��;�m�۪�5ĸH� 
&\�9���`C8�MX��@EY��N���:1k�O�%���K�lJv���i���$�O���ɱɶ�Ͱ8���Y�N�x���3'�(�F�&�̼��e� ��V"�.^QߑZt�귵�PN�u���=��9���j��.9q�\[���������Y��/˚�Y5ŗ�������uPԨ�'����:��T>�'�榥��G��sAk(HLn!�bx&���5����Z�x��V�v�4w��X3fe�.X҇$�����(�u6� ^\wA�Vo�9��a������L�"�U��d�Z7bK>�=�M��l<��e�_t��,����	��xK5��b�CL��.��q�K!�jЍ��9[�Y�$��1̙�-%�Q�@.�s�ȓ
r2��#�oӄ�@,
�sx�;e1��V�E��5�G��C��1��~���Фya���XAJ�����
쌯�9wA�z����ۜ�Lc�~�胘�(TpCam<���c1�~��Xp	�숅�bQ��9�@%2[W��@������{���ťJ0�i��:h�(�s�g�j��á�d\?�O dy�8�Ӝ�%�bI8�`���r����6��#Ɏ�  ��f��.F���51��O����q4]���!X�6�;ޡS��h�#:�^V��j&)v���T�Ҫ�)H	�"*p ��5�S�����*��3pW�,�ߔ�^��d�AX�����������+��(��x4����S3�ս^����B8�;U҄�,�T'��S����;.p$S���c.���f�}fO�j�C���=�*_����������_��-T��sx���f��L�����̏k����Q�䏅��9���C�%��\e�~�qĔ	xi�OJn���Z#: [»o[���Mo�f��������-ς�����<N�3#�W׶���C[�54o�Y�S�-��� ��-A�.�����i��eE���`L;���3T(��xN�MZ~�cd�
��E
�!�u�>w��f�z����N���N�U>Ik�����.�[�R�%a莰48ulj���d������w�����Z�1������
��4Xj|Mh�*��N�z�
3_���bP�3?3��.��,�m��p�����<��J��60���:��Fh4�ݍl���#���SJٰ�E��v�&4xb[(L�fO�~���e�	w��;(���[�� �A�4^O����$�gq���d�a���G�|0���&��J�����s��ɿ�H��4�G�m����H�(y%7�G�͍��ӞjZ��鳫�a/�*Tű� n��Ru[�����V^�����{;�����#L;�~U��5����=��?&ʺV���^��n�˩������4X��M����Y���ӑaovL�7(Ɵ��mà|��.�!M]PY��Ƽ����K�.���9�L��m��D�4a�pI�ޙ����ZL��>���1֩Q^A������j�q>Ĵ�r������/�;�Xm���x�!M���'���o�N�98{+�9+�N��^�",�W������y��ON�,c"+�9f���f�+�V��nn�x.5<�:�3����C ����u�.I��V��y�h$^9�8<o���a���P��[�6tY<|й6ts��]�x6�dk���d�Z�j��]�ɇH�^~�jz��P+Y`��7�:$ҲO�|)c����!O�8�8�/��b�kr�D�
D��032/�i����L���@	A�Q`�D�:v�^�x�T6֝�Lf�����ƍ�J�*��5Y�+Rp��g:����,*�R�nY�)���E=u~�0��.��c�\@���*���`���=if�o�A���T򕯓�n#����Rn?1߶��i��`H���GS�bWs�tNV��4YHb��̱�Y��_����M��р}q���EfT��{F;Hj��iѻ�8t��
�VM��́���KF���-����f��t�'R�\ԛr���������LZ�2�u�!��NL ��2/cKb2/d>�����~S6��W��B��3Z��4�ƚ���Q��T�
���:�q�`���	:],m}ֿhX��K�I��W�����¯dʺ��]o�r�N�5/��a
z�T���E�S�<B�?�W0ԉ����G�2�ug�6��46k���e
�]�L �pZ<���XD���=��[���ϡ��3h�~����%:mx؏��{b�4#}"Э��ݰ�qA��*�%�49��W��2'�r��e1f@�1X�Ż�Q���I9��9[	]��@�s@�Є��[�Gu���.���/����Z�̌�g�(��(P}&�9k��DO������ �Toy�E�Y�W\�>�T[M�6L��VhO�N���
��qO0G�{?��L�j��2���+D�v�b)(�6�h}?{!���=̆����ڦ!"̲L��r��Yμ�Ғ�:���p;g����-�n�F9�#�[D*�����<J�s��u�	'��I�,����ܱ�C���.��|U[�����~��W���J�3JW�p�y����\��g���.m��`9��]���e�o�N?�_d���2�&d��`nW�q�[�33��{�`���Y�y�AG��?�Xe3�6I�OH$v���U�Y&��	�A%8C��
��k����#�_��pE�ٷ)x�/���/k�w�"�uvCZ�ե�'l�(��e���@��ʥi�X�̓}�M�q���*�M��nk�T0gy�^>;��ȵ��ۗ��=��Wh�$+S�A���HDlV�����J��6V�!.8e�N���樘y�t�Q�S��kqc��R33v�SI��V�ճ ���:��m�RKa�;x����l=�4Y�g:�|���O�b`D�鈤�}9��a3��۟����?lˢqB����`c}�|�UB�>���vk���O|�jM J��u���s�1X��~ۭ<���fw�g3���˹]�/s0��yB?�"Y�
��q?y#�j�I�M;����&�˟k�@/-��B��z���4#�_�I!Ԉ��h9�礛��|���$w7Ex���F0�Z�h�h����q4D����y@o)$�&
������CKNF�F�����G(S�ޮ���
�<e���&��D�φ��0�T(�`�Xe��|�P���c\{�}(&�J��^���(+��y�`N[�&���
�+G����o��u5���r��܍ukޣ�z��bc�S)+ߐfe%���=U��XB3J�k�j�i> @�b	�А��m:��Yq�8�c�&&�6�U�懜�ƾ�9_�&[Va����<��/A�����0��kr�pu�3�C�'���L�K[���r�)Z�3�F#'S�z��ݿâhί,d�$-�F�I����y)iE.�\Q3O9��,��A�vfl��=LQka����f������	�<c��(`��8���Ţ4��2Lƒ?�[��@Z�Ui�P"�|�<�+��"y�ٞ-�)���ae����o&�]SOkۡ7��L����<�S �"h�&q~BE[4���ݹ�e��|�c�D���?]�{"?#�������GƜ(NL���ѻ�s�;��4�43Tݪ7X�j	uf�� G�E$h���#r�=���]B[�"���%�A�ۅ��9��U�<|�I��r�����̇�i����c�4V&�v�z�P�2K�m���i�n>�Lj�h]3T�˔Sc��Z�3��خ�<�Ԇ�&ti���6;d���<'�| s�X1?��?dC~獇K��	/O
,\�˻j�)�%I�c�i����޺ӫ$"PV
��Q�<���&���ؑ&�oD�j+�`b*笀����������>�����i"e�w	���%���N��Yf��ft�IV	�Oz:Πw�g��.j�g~w� '��j�88B��NS�MS�τ
G�|�=�yl��ŉ�X��
�mN�~��H�������{~�K�KcF#��3�e4| ��5/�!���XޗK��_�$��|�1��G�b����.`C��1�p��Oz�ea�l{%��U��^cm���}�S<�n�x�dm�̷�8��~z�WC�W++�&�m-ƲO,5G�X��Ɋq�>.�Tl�+ F�Y�� �O}Oy��h4�3�#���o�FƧ;C������b`N�({�3�8����ŵ����\A���?v�w��e�C%���2N��6`l�Kbn���㩽�>qFyǌ�B�4������޷�o�@�`P�R0�'��?X���k3�M;�I�꼮�lP��&�	��k�\yxlG3U���0!��;p	�b�~ �����>�obOp� -��/
J�E�+5�����9U��z��ކ�)S,�lCsV<���k��l�#F���,�H��gyX��N�ǒk�Q�:�[�8��S]�~�d��k���o�����7f��Ӳ���.5���>|,y(UQ'%�%�7�]��dT�ͨ��}vC�N�8�X f3��^�����AY���o^C�Uz�~Z�yx��R��7K�m	X&v�]+���/D=�m�%:ERaZ��K5nbci�;,"/>����C>�?��=����^eK�Q�%�m�1I�w�\
�:��DѰ��98g'*�VT�;�{朻�!��8����,����BH����ڡ����2��n��׏s|��S/R냪�[����ތ���ⲿ���?������$Q���z�#qm���[��2���6Ȃ_E�мD��ϟ�ބhITe�y�#�Ȝ'���Ͷ���gv)
�~|$�_�ޚT�l�L�vA9�@בG��6L����2VZ���0��h?N|�=�C>���	�A��J��a�c�q$�7#eMϵ)2wf�M�da�9�,�3��>�z+Q�\���K��~w�a�d[�r�;�$m�$ׂG�*�D�_� �]���هwA͛#���l���U*��D�v�8j塙ɤ9����"����;���ees?�{~����*�������0�p��D�C��F�@��Q�^���S�Q�἟�&�[�Z0�t�ږ�L�K�R �>�A_��A����J��jS:�{u<��'�^k��vn��'�XY�=C�����S�?��ԚJ�8�C�Ի��p��PG���ws>d!MR��!$x�����q��Nڸ�s �Φ���	�$"�@�&�)��Z�(�@�c�rN1�o<2�$�����I����`�2�K�J`�e��y�35��ۄ+Ӂ��vL
�c�4�U��P��q�,�%�%���^bǧj���/�u��b���ew��t�4b��6�����Ӣ50v6Ljd&��q=Ⱦ~�ԏYGSB03�7�g����7��u 3��qvW�U���K��8����|�K���xM�z��`!sg�#��]�V��[��h��׆x#jD���7��Y��]O�d����|̚��ܥ�`-�h�&��,����񇚿 B.�E�R�K@�T��c�/�l<��'S������w���[��@� Mu�A���?%�����i�� ����I��r�H��Z/Ij�f��&�{5dʚ8fy;�.��[��D�R��h�Z�i�u@IW��RcP�K|8ӏ�5��;�z�+%��@�8��`�dg�6�ky��!{��o�3�]��xަN��V&	`@p����X�-��^��ӓ���HX*"���%�=�{�ɿ�d;�"�Z�L��ܠi�+g�nTX�d���!Y�P�x����'�L�#�f�a2��kT/�I�?v;�G�)HV]��9�Y�}�̌ v��4*������
!ӭ'�V:�$���'v팼(���mܧH�BtK��Ҵ3�*������/ ً�/�K?�s��\d�>D�ݼ��3�?�KsiM�$3녊����L9lzOU~O5%w۠uR��"+�� ��P���I�/�U�|����J��j.�cq�3�P�;����5v��ɄO��ģ���m��$[��W�$��V�XetL˒v�X�8�d������O��n�����W�Y��M�0^kKĪ^S[�f�������Lm�w�� E]����Fa��*��75(�f�h#kS��SO�6�ւ)��3`f���	B*	��(�Ic���/l�#ޟ$�P>`�۲��q�ֹ������޾T·��|�f���_�-E^~0I2��� v���B& %ч\N�s����=ub�@���A��C�Q4&�f��՞��b:���~��P�O���#��ȃ=%��R�_����}�7Wt;?�t�����H~�~�.uP(����ˀ͉Q�����mv�Qṋ��\��OD�*p5m������I >���oWn��}�s��m�?��K�_;�n�����Th���٥�jA�g��U�������s+z�y�A�6�B]��҆"ލ~�D���X��-ŏ��;���T���2����T�YN$��	�'A6N	� ��t�.�>=KAp��x��`�=ۦ�	PVd	lqtqFs��X�C����h�}�ze� Է@��jۑ��?���s�@3�E�g���I [M�ؗ���8�Aq�+���+�6�4T�b.f�F�j8W��BOOg)?v�x,�U+ߝ^F��w!j�+��U��Y
p��ܻ]b��Sg����Կ��d�H�K�}�G0є��zp����TĤğ"w�1~�%�=�"ky��P�Y
�<�_�3�K�[#��dg#҈��c�b��Wt��Kz�:a�RR�H�q�ͲW��*e�!�Bq�7H���B�������)�!z�X���ٮ�o���$,��
oH��~�ZC��,36@����S&�v�������A!?�Y��a��nT)�8%��zK��\�� Uɑ�y�1���7U�(:�{�H��l���-��A��0��[t���VRE�Q��2T!)��鏪L�����Z+�@oj��PK��h�_v]3=��Oei$؋�&��1�����l!C��*�˃Ce�8E�ݠ.F�~p��O���]�`}���@�^<~�Id�R)�e����Hw�,׆�[��4]�~��j��w�l�)��R<OԲH��^e�*L~�o��[�|%^����&Y����*R騗m�K��Y��| d'�r3E��p�v�6���gW��y�.7��g!�P���|)'��e{�F��E����F��L�>��xdv���翨��:��`v�@z�O��	�W��y�b�l�[^���
y�6�BJ�1��y''P�L��"`>N�:�Tݾ�&�g|Y*yX�xJ*U�ߴ�f,fh��H��n�4�����괌�)�8
u�La_���-��p߲�M�Y �V�ʬ"ܑ.�V~�IБ�	ԁ!��;u����ԓ�Y�5���K�3_8�ж� �K>�+`�2��g0�au�
4@�!�]�b�e�x��M؇��Rr_ �g�.����~V���#_��BG�)�x������Z\�6IG�=��5���^A�H+�F6�6�B�u�\z��ːw�����3�\�������b�N��H_/��@`���J�(3'fMt
�=i�U����2���o9��r��(��Cʺ��2PD�'��vR�oR�RR�/#���%!_�����?��+���d�l�T��Y��>�fJC�㸫0��꤇<�";w�`�Z gtd�֨WC���X@9G��IF�e�02,K���)��R�k�Z�����b��u7(5��׮��;�oƢ���a-�$�����?��l��)��'aJO��^�gÃ�7����"�Ϸ�;�|Xo'UR�E�T-�/ک�Ӗ�� �#�ݝ�`1W�b��d�}�.�ܲ��֗���2���b��:���2z���M�h}�-�n�Un�+���T�p�@'MV�g��S.n�_Gw�6U�s�6B�6 r�lY��B�����ՓG�U�t�G�0q�ǡ�41a�"͑���(��9��g�w��%��3>T��_��ꓣ9�|��:Y�m>��@��,����B7I&v(���n3۫}��C!���1E�(c3L��|��7���g���¯[⭴�`x�A���E�>A"�g{�d�g�F��D�#K�W�}`n�*���o�}Z�<�-�	� �`2�m�����]<V�YN�8p8���������������w���;P���I_d��c�K&���{�Q��ԺdC��'`5k����U�Z��t{'�a��5i=}�ͤgx�I5�F/�g[	��"I��t�AeTdU�����*b���Pvo����4�����~B[Փ���*�b���z%	|QF1�cbf�>��$�E�֗�TI�U�5Ĩ>���̳�(��lfj�z�U�:�i���znז"�fm/w8����A��a��%����M�������S2&�"Ƴ�ذ�w$M��Z�AG�C1JI$)fmtN�z�ef/�Z��U'���IזE�S�@��X���lv0w?�ц��于����d�>�(;����SGh�O������'��y�[6�0	��xj��;�"I	l���9DJԗ6N��8#+�x@,p�4�*w�|Ͳ�ۉ��`��� �+� N{2h~�z6Kܺ���� �+�'JD�I&�4�t�5��ϠK1���-���+���`p��XƦ�2����z���K�R�k}�0����a�LbP�
���@���U��˥@��j�FE9�!^�M��]�@D$2�옷���X;��a�#�����y��5($*{����iϦ\��=�ޣa8x3��/d�`�P�6"���l�#tc@�uE* ���͘J'�N�H;�+7�t�=<z����  MBd�,j���Ƅ���Rl0��Pؾ�t���Jq!�89�:y[���,I�8o�O��>l+�n^wBn����K
�{bV�yl3o�g��8�
Ӱ22e�U��mgǽ~�UW	vh#�ǉр�H�U,����E��c�F�+��a0q�Ew)�$�XI� ����߂�@�<�� ��-b��!T��èdأ%����%t8F,o�Ng��c���2�����V���+��k�9�%H��$~��KA9�N#������)Qǆ���H�H@�Y�Z�/������9,����T3��١T�fɍ�z������@[)��T�Юx�!"��#��=I=4!�,������*�����x��Ҋ��O���Jd�{��.҃�;�@:�GnYӋ^��T�>� t�U5�S�o7%E?���TW��/<����a��A��]b�R�\s�uvt�<�����~�qɟ�[�0(��!Ϳj�߆�N�Qr��S�)�tj٧���DA.�$!?\�F,��7�+�Dn�jeҝ��޾}�dň����p%F���S�hpy�u��^���9�(���^�j�wٸdOð�S	��h#��k;H̙L�����7�"�~c��$-�溏�&��t����r��-��L��8��L3����y������L�J+�����Cv�G�R�?+plkF�ϛ/|���d�@VG�����n՚�;��EW�a����h�j�]��ޯIi�S`҅��������&Հ��¥���vu'Ѥ7���Ʌ^l�B?����6��˗׿[)O`d��@v��-s��6#��ik����i%�M[2�Z��Qn�����$~A��R��g&��Z��f��"�2�oߗ�}Z5�4a&dO����jk�y��F�X ��!f�lbO+��{Ǳ� ���~-f�3��\�&�)L���&�%��#�W0i>�x��Ê[�w��m�r;&x�͜t���Q�']�2���Vu(����˭7�^vF����;�\�j�>��.�s��ÚL�� �6?u�c2������	�2�&U�q�07g�>ql�<Au�y���w1�o�9�(�D��I�eRO��m&��0��9��`�
>`�#�n�����4͹o̘�x���K�E�PUu؁�0�P<����Pc��_:�v��瘖�O�� %�d+
b�k���Q IQ�5y[�F��Ԟ}IrJ���o�FP�޻Ա�J#p��$��O,���T�rti�2R����"��r߿����j��j��'	����1L���Ҽm�v{��0����V��k�q{�翁��f�A��Ը��d���>f&�o�����p�~���N����t�%�<@����q���)%-A''F�<���y9�u����c�<V��݃$�l{��UC:����WV`hAu��u./=������n��_,�%��<O\^��xf�0������} ��7ʼ"V$����f�tq�0éQ����_���˜`��M-�G��� �����"�&c� �. $5JM5d�m�} �W{�i'�F�Q����%�ݢ����aئ�z�DfR����D,�r��Iة�y��a8�kd�[Ġ0�������D
�k8�K$��O����;m�ǉ[�8�7�Aj4�����r��M�a��i��N�NosL�� �
6`��A-���[��Ơ@���3Ko(`Wo��������l*��v��u�m� �'w=B4K��+�;�U��zfi���k�3l���,� й�-������<�##�iw��e'�8G�nw����s	; ��C�,
Kݱ�n>�s�K�N��kF:��Oh��S��*��>`�#&q|O>�_C ����-o�ZcJx��N�0�ȸ.�O�4�l�`oi�)@_���*ģ��=9����}q����� ����L}��(��4y����[erk�[�`�[6�6�����q�5�k�{в�Q����]��t�k����#zQ8���(K�8� ��\QGԶn9��O��@�qB1�5�����������a���`��OY,MG,�7��A����C���w5�R�9~L���brrJC��-����v����݆�[�k[��9�[Ԃ��ya��k��V[�<��ds^wo9�xg��V]O-�>}��C�+�fQ�\~	N�6�EV�a*�{�f��W8��A�a�s�;g�W����Hq��z�6�͕���XY,�z ��c�o~�$��ܚ�ր�ڌ�mdMb���.�\i�Y?��#����gG�/]�$�1�mۇ�ș�i6Q��[0m�QZ�F'2�n�7����� U�g��`R1*"qs7��3�:��CzG����� Ƃ�NVA	��{�Fh(f�ˇ�����m�1 V����v�1�4���~�$m�̼<�,���К�y�+���ES@L�t򱯈����o�r���:�\1B���dk��H����XFSB���t�q"�,
V`�����h�$�"t�,4�D8a�2i�"���':n#<ϖ$�����繺2�{�:)��>�ay�01�L������*� |�׻�H>�%��T�a�d�26?�� ~Ͻ]�}���L����tG��H��/ϥ��n��/S��>�8�x�e���2J�Z�ʐE�(�e�Rr��� e}���YF�*j�9�G�B���5Ri�����t*}#S<�u�{����v��漃���[��΢&W�:�kJo��6f��q~.�W��K��������y�6�?���6�-͍����e�8?c�X��4�� ,엛��
��h�GMsV$5�P�X
Yx�Ӵ|��&��w-�*����p �j�1m+�������`���������g����x��ŀ?�*�'�g��Y��������/���3_+���� GytI��7͔��F���7O��������+c8��s6�J�G��T_>�f�@��.����	=
`i�,�-��U����^��ȿ����*��X�"�ys�
��C8���s���K-�cR����oē>��	�K{B���"���{>)�.(y�W��T��Twa� �7$�v�]��I�^&��+�%����N������H�{�E����EZ��טڃ���$/��|��}lU��uM�: 2��^��׀�����Ŗ>��z����C��|:|����A_ڤ�ժϱt������CA��8��,���fOt��TE���j�m�����u�����z
ݽ�R�H���ŷ��1]
4����W��/5óov_-�q�>�:���4��fP�4�f-Z���j�K�,���]9�wR@���K����bE�3��O]a�s@�߁� �M��ͣ�B�Sƹ]�w���3N�G�� ^|�(dn����wv��g�,;�*��|Q�!G�a��cc4@+�t��2��2;']�A
�����	f�����ҫ�k�����\_؊U�叚��i��u�+qH%�l馀P�c�N�����M��+`-q���m�׷�����	N���׶���K��aD�4J��іo�j.�}�=s޺sWi�I0ŗf���lf�Uq��dý�=�n�q��m/g��M-��݆���ȵf[݋����O�菵�g�<.�ߘ��I�W�6�S��{�V���u��L#P;S���	�6�����0n��p�:����Β���:��g�&�lli��|O.)np� ;����3^�&��2o�i�g�Y��@O}
�J��"�t_:#|qk~c�.ˑ�_^SH�����}��X	�=���p`gw��j��ZnO��`Ų��w� -,C�9��U#n�2N���bz'B�q8φV6֌�Ք����rR��G��Q���u�$�_�` 1E<���~�v�DmT�ƼR㴊���vjȋ���ܸ.y��֒��+Cwt�ô�EV{��W�n�s#ӝ��qB�S6z���.7}�]Ҙ��S_.�wҁzq�����cA_�"tw'�z�h�2�ク�0q�铰o�Yt�i�6�f���D�s#n��;�i+�g�f�@�����p|�r��^rȕ�3��W�2�m�!�C��OV0V˓��t�=���X�Շ���ޣ��)��G����:{������ԆN;�dȿE�������a���ґ���Q�K�~q\��Aae�\�ʻ����Б�C\�rR��{~�����~�z����
���M1%8�����1�aRdjtm/ۑȴ�Ǖ��wn�a\a�J]���K���P��XؕD��|_WL�;���]~� }�S��l�Z�������@��r���9{�4�o�H=���I�8�A��'���ߦ� �S�P�T
�3o���y��<�<U?N�~]F2�6��
Ļ-��Sm+ԁw��5���n#X;KA`�"�m���3�cXX�s�2��m���(H����ۗ�'�{m#ei:��5��'\�>�,�z��b�k����u�� :�F)��a��6�P�q�c^�=�^�w;i�� (ϥ����.����˹����ℎ[��#ͷ]��	�s���?o�^�^CXcZ�R$o9�֮���+�[3+m	�W�ڊ��7!o�X�怼�ݐP=[���HV��`�%_x����f������/��MZ&��G��V%K����j��Ǩ��\*�K>�a�]��=�P��G?u<�כ'��m&��� .�A��t�p#i0�Ul�f�!?�z�D�k�JG
�R���բ��?�Cn�A���t��-�$�W���b�ߡ��T���1��g/�����8��[ݳ,b�O���#2�!��e2ڜf��Ke'����#H��*6YI���a������4%�ҫ&�45*`>li��R�)��+~�4�\����������������4]���Zq+C�}�����e|RKx���[F�c:�~�8*K<��L@���_�5�[qqUL[�"�L�B���d���J�R������nXn�T���e�W J�q-T�lNWbN�����4D��d�FH�SX��J�Y�6��!/��@�aD�)�!qa�$V�H��B��K�˺W�\��[Rx)���';1�v��l������$q�՜�N1JlΩ��6OA��C�'p����)���Y�Q�U�IW�ٕ���[1�G�;���Fr숮uC��� s�b��sH��i�����x.�w��_⾓��s�O�yEV�0��.F��38Q��F��'[up�=kSq�xy����UV�©|�4�m�;��H�q�hƅ�+�_�g�� ��,����A��Ӧn��ﬗ���F��x��B�D��g_ l��8!k ��JW?��Vǖ��A�B���ъ��A����M�*��q�����$l�wFs@�;����1���%֐�Y�V�#�/@ЋG��޽�)D}�r�pU:��Xpi!��W����U ���q9��U������Xؤ�t;(N}��Ի���}ʬ��O$��0_�-���16z�.�K�J0������^�V�e�R���X�̣?�U�l�F��K�Ά�U�j5��3Q�L=�Ő9P"�A=G���R�[,D>��-ʩu�'X	�zq��z'+�L�x��
����x�Ȓ�c���m���H�n�kH[Rз`�`�k؁�_�L$�EnK�����ſ�!��2V������w�x����T]<'a-V��;8��B�*H�Y�&����d��^�x¯��W)#N,����~U$KS*��$=ΐ�	`Z/;AZ5lɛY*�L u�^, 㩩>��˂��n�.��z+XS@'<�#���.Uћ�fW��Q,rW��"��=�@u5�v����Kn~P+�d~t\zM��\�b����Z�Iw-M�/B� �/���k�%]��1�ݑ�Ai�9=+���`^S�g|�S��">�ԛVD�3�U���2����=�̬�r։v|�t�#�����m�L9X�t$�����7�B�Lh)�'�ӏ-8X:���4���Z<8K�V�����T���Q��+=rӏY�`bS(�S֤7	m���9,\-A�K|�0��"��������	֪�T< ��<���P�t�����?���]�~�-���lV��6ǲK���B�� q��`ִbw�5���cAP@�#q3�W],�w�z���g�$I�������1PZm�+��UU��V�u@����,������,��3�z\&��}vHb.��ReѢ���^
[х{00R���P���2��T3+��՗n�\��I�ׇ[%e"m�BkOg�Z�P��p�E[�v�񎉚�#z(M�Q��Q�ctO�(d�/A�=�chd�_Dg?�Gܺ�޿����{l�Akj��'k�*�qջ�xYCQ���K���)E��~:�*L�hO�q�[�Wk��e�m�v�`�d(]�@X3י3+}w�~OLa��+Kb!�U�,���T���5�v!�g�诚Y�vrG0U�+<:V
-�Sn�C0�l�'�;Gm�,G��e�.�0�M��0����6�}��3�N�����^�|�D+J/�lc�͙��k�y$�z�i�lަ�����N�(���$ƪd������,s��؃\b�[cj�l~�F����J��2���k�e�$�RhwP���6�4I�يA��o?�ӊ��:��Z��pP�
��WV������Ǽf�M\XjA��U�z�+�����#�\���!�5��	E\���� @��{ͳ��f�������\�R�SAݔ�cG%0օMR_SKJ]FY�4��4�)�y���O6b9%�����c�`���e~j0���]���I���K�EVw�&�lN���l/b��̆YR}�1��e>�!BH���'��nN���2Ddq��+�z�}a�r��(�4��,ɮ�k�Sm�R��Z�b�D�	N�<�~
�t:c�U��B���>�/�0��RŲ��)FV���/�a{�.�?f�l�����Dw Hȕg� 5��lbi �����|�W�����V��Y%	o�w�|y�{��{�Xa�����Щ������6�@S$�
�*Q�F� ot*5ko8��4��vb�8��ld�D���o|�7f�5A�j��n
�?��q�0��75����J�a���; sD��zS�;�Q�����c���Uz��"H�k�y�Q�3 ���*KS�Ġ�1,�	D�A䋄�6��9/l~�Qu���زTK�	���^��v���$��8�Mo_!��%9�	 3��03 ��ph́lݻQ�O#~���x��{�M5���8=U2\,���A�~o,A�Հ8	���<��a"Q�NH OZ��9���u
H�.M��πC�����N�ER�a~�^?��~���q�ׅe&ΐ�Й���a�@{,���uH�uE�{YD���#�]I�9�-Hϛz��,�n	��{Ӛ��`x/�0���!<I���@�'��c�x�}�q��T!�đ1ؽ�Z^�E����	��φ�b��d�2㿣&�$ف�L� qжhE�ӌ�͉��t�1M��j1��̝��������WW �o����	N�	`����~Í����=��j}uz��F�=���]DS��i�}0�y�=��!]���=@c[�=1��@��MѴd��>�G�t�j��/������Fw�՘E/�� �3���r�������l���G�(��檯�`t�/��Z����-B2[m���N?�hu@��}NV��`�ŵlK~��_�j%pY��G�M��5��깝�1@ae�\�N�
d�?]���<h��7��JL�}��%cQ�,[)c��3?�F8�p�Se��xS�w��cC�U����+��^�5���2�P��L�dJ&�R9N��d�*M!�j�>�g9x��І�.Í�U��m6�-��?;�����E$-��x�*��ί(فN��B�Lx�B�΢@K�B�#�窖�#��{5~��}�$5꾼d�#�T��v�\��m&������rϋ8��;�T�?W�����Hd�2̐|Ȣ��oD���mҴ�{�jD�k�o�7��h�K��O�#��D��wy ��̢zm�}+6Q��T)Y��;*]�3�>r%�����N��+�$�^gt��m4%N�v��e}X	������':s���}FcJ������4 zr��\	�FyL(�Iy`�mN/*P�a���h�Z�oF Z�\{>���C�Gr���LG���`�vJZ#^�eę(�ȟ�70����=D���y����z�ZN?ܗ��Ñ�-�m��)cI�3pй\H�?s��:i��$gE 0z A��qR��x`�z���;]6!�WZ912��׭��g�MJ��=5� �4p�M�A��? �ҟm(�H�ůL��^��=[����7L?���%�2)�_~?���|��;�rN�P,�md�F���y��-Tx�+�5	�N0����s�N����f��ix�V$��)�B�ׄ�2��0�0��%�YY�?Z��;[y��P�C�bF�	�Hg�2)�J��:�L� ��BǗ�Kn>����hr��� ���/0�yy1�^2�.����\,MPm���ôDa϶vtTi{bn��xh���B�����z�l�;.�N�d%�N�ʄ�۹���Q`�e�j��M� 5�	��#�
2ܔ�Ɍ�S9�5����~{7n<�t���<j���ve�Y����	�L#�Ð�@*Ӥ��c��� �l�y���wbd�ڟ/�_`5�@� ��k��/òQ(]�a��(���=,�IW/5�����"\|�0����S��ϱ��5L6��Ǡ��*e�D,�F!^�H�!ߺ�	�z*�h����spd���þH��G9,�(U���\�l���e���|�#�C�#	�1��4��o�>z{uDV�%6�k�aC@U��a���(,��0	�� �u��5Ȍ(��W �� Z*A,ڦœW[ZnF���fqZA|s$A7�G�AU��͘k2}�CS�������2E1V��CQ&�4:���'}�ib�9&��:��ZC��jT�K���������b�A�h���������Ҡ�C�T���<���} �u���geV`
���}&f����8�z�-�]319ۗ�7K��o�������?{1��'o��F����C�y�[H�,9(�sų�r ���.�$�1�~x�Rߞ���&�y���În�zٶ>zR��A+ٹq��q:j^��.:��N�R�G��@u08�k��p��ƅ}��_(h���ʜ�8���,��0� �)�1�g����?��9�{�|��������?�R:�11܂�Њ�tݡ�3�_So5�[9��sLl3�W�2�0ua�p� ̈^��r��1�D�i|ʑw�i��q�h��N� ��b���-�!j�屌C�k�Yt,=^�$fOS�o��(�c$����W�qjz�g�s?${�w�`$�=PL�������s]y�ZK��Qm�� ч�S��P�(c����N�7@E��f4"rM5�}�>�����&/+���LS�㸘�����mL]�9R�2�G�&?�#������m�� �ILGн�j|b�UH�� +�x����W�D)hn,Z':�:�����O\<��[��z��"� i�������|[(w�g��AHS gf<�DeO�����HHu��1��9u~:E�E0���]Dl�������|%Q2�L���2�)���
+��_,�!�//��J{�WeLZF�:� V��Y(�>Z�E�X��k[(mP}r紽��F���G���������� �o��S����t��#�l����%�)�b�"�����v��*�eS;ؘ��rY����r�{������X�V"�[�r����sH�m�h�<�	�NR+���\�]u��Nɦ�\��C�m�*� I��#�_�fT]v!ka�m�����ÊX����+nh*&d��dJ���M$DY�qY0�X\w�K�!�|Y�+X'�m��5�cs�3�bL!�/|)���#�ܨ����dBiMw��@�z�g0<(�	h��p.�<�Q�jk�~�vյ/ �>�a��/�������"�?R(��G�Fœ����yx���#G��l掋:˾�,�C�V#�穩�<e�ፓ�W���}<EQ�2�S�������wYI�z�_�s��y�h�Ng�r� $�K����䃰=sR�<����c���-o���H:�"��o�1@�!����:>��M]F���W�B�H�&� _*w�3e[#[��&@X2s�W^6��������{�罊�}�����c0�۽+;���)fݒ)�p���+�m�5����1K��oq�R�5GV�Z�S@\m3
.Ց@>��_�qp�[�5�S������Ĉ�-o*-|�Ef�̜<G��a8��2ǻ�L�YdԷ��:�HA���}*)�ã5'�0a��L�'o�Ϧr?��>]$k�[pm��7r�0����u:Yd �mrZ=�+4�s]����hv>,�6V�Q����l�qۭɽ�6�FJ��-������ݪ1����j�I��(������7,k�1����{�9�0b@�n�6�w�2̍!�K��M��P��5�>��o��E��( �Ә�UD�i�H�A�İ�����"�av�wE3�K���� ���:�HҤY�C��O`�6�KN�}Ko����֩+�sNn���2ʊ.�������Q:����pex Vr7%��J���Wr��t�_@�����&Q�/�V�SP܀��YĹ������7`$�D��3����U��^n0�%�{�&� �!��kJ\w�goL�vkx:�]Z֪N(��Gg
�5�L�@����-qߏ��ZTa�n�1��Z��.4�Q��2��TO!�����ۤwC��'ќ��$N�(V1g��s�$�l+"�~q�2ǘxIJu�U�Efg����ӵ
�y�h��v9�mo����Q�w�Lp��V��B�����Eb7lX�ʕ��b��WQ ��������M�<�����a�YI� �>7�xH����`}5�w��:ő��m#����%�N�n�7��sFҙf�:�k�4�/@�iQh�$Mr�O6�����!N������ێ&E���}�{G���!ɣ��v�����BE�̶s3�C ���(�&���_<��K�+�}ҢY]�bC_�f�?�A��L�'�)�ߚ8��Юs��C3�^��䤫���j�$�t���	 ��"|�qMtf���Wg�Fz5�fJ��M�c0�� 
��.E~���U�>ɠ��1�7�����@Y!2\s�mj*sU�?DĨ�9�WmV��)�R����oI��Ö�椼̡�%*�2!"��5��@M�:� |1ܠ%�n�J���X�$�oL}%���UE�s�7�n5W|�X�8L�|y�2�{Q7(y.b�u21֥��+����Y+��o��Ycv���&�l��!_�W1iDƣ$��JD�W��ؘ!R�kc6꭬ᇭ��%~�YMb�xXg嫵dš�(�d���1�&�#C���{R�����:�I��(���������AԴu���!8п�!I�:�?�^�p�Jƃ�4	�R`�&�.���F�9ȇ�@����������%�]/����;ND�B��ӫ�4ʥ�����&��./0���*�Wb,O/�����>u,�w�;���m4L�#�P����;��6���ti��]P��oD�H R���jBU,����ԟ���c~��[��s���cLW��Φ["q>t7L	��N>���	:�h��a����6�"֚���.�@MI�ڟ�������S���0b���5�+q]y�0QA�+���F��!GH�a�Û�����ugv}s��-�$��(7���u^ӹ|
��&�E��C<�F��P^�ڂ�,1�G���P� �o}b�Pc�o\���xX{��3hg�W�D%o�2d�,�ꃏ���_�����F��cF��7�]��"F�I��P[wÅ>P-6^��1=�!���ƟJ]eɻk}�ֵD�ɣ��d[���Fo� 9��	\MZ�-76C*��!�����䢣�=��R����@�|bo���	װ�$�qpiC��y�`�Q?B<k�7��n�3��X����F�b��γ���B�s����Q���Ş.��6�EIvqBl��]�G�*�(�혭��vI��y�����)뒜�bb��m9�E��I�K�)5�Tl�G��ڤ[qH1�>���%K�
�X/O���l��.���� �K�悸r�[40�uH=����_��-'@kI�utIǵ���k��@*�x��C�|��2H$��H9Eɂ(��L>5G��F���N6�U��( #��ti�|�3S#�v�^Wq��:M��V�cHRA���T���O���o��-?\���;����=���`id�K�f��
���@�nJ��7�dH�S|jp��Xj��a1;�z4��<���8����^l	���G�����u'4����E���s���2+���nPu*_�uU��_CqM��(�cd19�q��񸅁�� Ȯ2W�1���rMp�BZ�'oq�����Ä^�:WʂZ@��Mh8�F	UE{�k�\&<P�(f�c�b+rvi�r�1rw<��i#�����ް��iZ���#��/��vv���z�D/�R�&�v�(݋�= �`��H�7�0Gi��*z�GvzP���]���Dq����}������<ihel�4�3�,�#������&��=|MWY��ʸ�a2�D���M��U���,��.�<&�T-5%���9)*�'?c8�b��E ��o4,!�U�+�1վZHy���ٗ&��k� X��|�@`�ύ��K�4�yہc_\��D��,�!�]#�`�:��rz�N-�lN�$�@�B�J����&��5�cJS)��h��5:r��7���4t�1�8@���1dd3xw��&���۴����x뷮�J��?�t��O	���C�2Y3)$ >�.�k=qC��V�iJ/�5�ZXu�!�5c��>�!�j�]�~�T1�b|�W���m��Hc��(&�R6���TΦ5
�,�������d��`t�D�7�˃�)�X��{`������d�Y�l�����[�4Yv|����� T^�dV����l-��XuGyּTX��oO�2*UXk������{��!�˅iѢn~)["�fk�^:2���6���A�|���������X�e$�8���Cd��V~�M���
����L.�z�¯Ư4����k@�N$u��8׬Iׁ[W��f`������ *}��%����-�j(TBHi�������w��i�ѫ/���H&�=��ә��p��s�'6�f�*��F���z\�D���&J�o������4�i{��£����xQ���p�y�Z�fJ�yqF>�/��#�݀v+��9k�VH���XA�Vk�&@/-q^�A̜��U�N��M�~����py�5�0�f(Ә}��M&5���Y�����b�V�C�eT+�"&��#
/X$�Ϛ�Q-�,~$r j�vw���'�g&�J��˰���(�����h�_	�.��]֝��"uT�,��(ߦ�ʋW�m��	�L��$7�5�j����/M-e��h��@�S:�P>z{�j��������NZ��?�S}L	�_:�T�{?0�u��jbm�I��/?�4�5*�tT�_.���X�<A�t�`�R���h�O��di�h��4�c��h$Ǜ.�]K�.쨡���z��{�g<Ð��f�`lt�!޾��)3t�t�R�1F�\ �cgn1�-Fܾ��[ˎj8z5�W&1=�R�Q����Z�%�>zgR��#" �C����2C�8��~�ް�"S���dA��m�5�����ln��U�s%��\���=o��Sj*�L��*Ԝ��1��|��R9�氳w�:{�@����� �y���h
���k�\gl��yu�v�ς~�SZ*:��!hb�?�;��'5Cl���Rr���nJ{m4'{��%"Iz���à��!��xpt�=R�c��.���H<�>�
9D�l���~��߇����y�8;1��~�z7�J;�m�ɋ�&�t�
����ۍ<�%�Y���p�6�x�����߫�Lv	�q2R��G��BS[m��4�h�4F��������N2T�N����7�o�F<w�~I����]���.o#�A�{�#5��e���$�h-��P�툔8��4&h��H�鴻.M�P�*���{I�����W
����I�0�����@���G\������5��O<�,Jws8�����i�i���l4{?�f�1�'����1�%��6��H�Wj������Vo�Hd:�	���mTNV�L�yF���( �F/@"���ۅ斝xp�ٻ�+���3��pTSI�d�FH(
��61g�2�I�d��5�^�a�A"�k[ ��_�l����:�.��aZ�E&�P7�?��F�0�zwH�>ͷ������8�v��D���#x�1W&B8��at�ű�Ml��hc�`�{��Ί�0ߚM^\�����z粇u!ŧh�u�tQ���n[����[���F�|p�<�������e�1is.J=�o^EQ������I�j\P.���)�"';*i��.�5Ռ�wz���Z�y� ���Ƈ���(5�a#�
�y���8Nn&�Mk��z�4��1�Y�\y�o� �˂tY|���G;�_I�����]�-ʖ�)���CU�/�j�?tV��j3���Iw���	���>�6�	A��R!%q�=sԘJ}$O_t��Z˓���'�Ae^Y퉠���I�o����{�7�K4�)���YE��Na����g���4�kB�l{=ĄD1�����<.�/՚]��֏��b�[��?��(�qZ��l����8����\h�95������y��<���d����i��"?)���*� +���0grD�@��F��W#�CN�O/O�����AX��c*�`��J>�2�������@����1��'�?�i̮������v"S�g��DaN�����"��cz��H�O$nf~'�39����3m}���\
|��Ħ"��`H���jx^������@��@�#t�h�]�v�_���XaxkP��\�ڍ=�%:���t��9�Aq>�5��X�ca��ud�$��n{���yn����C�փ`L����S�`�&��ա*>�@0Mlh#��Ӆ%�1�}� �G.����ڥ����l !-,[�$l�P�虀���1���.Ϣ�m�SƐa��v�8�>����EXb�P�
�i4}�����C0�������ہkM�]5A���k#�Tt�$Bb��`DJ��׼.N��Z��)CA��0�K�<��a\���0y�����0��D~����s�S�S�kؙ�\��"̭���-��3A��X�'d>mbh�nI=VT �5m�-������A�F�X��5��+vIޙ�D.}#������#���{���޳-��R�yٿ������I�G.Z&���Y�j}!��Fu��+��u�Te;@5'G%���(��������!��S�`��,U�i���
����Gc'����
�b��}�&R�P�ȶ�'�s�i�"�n5~�䕿�N2:�C��5�!��Ac��f�&.
p~�JT�-��ʝk	��	APVc�	��/�@����p��{\�-��!�濍{^Ou�}8h���~�������Y*�	��	)8�f��{pU�᷌o��v���ڲ>o�.��k�*�u$^6yM��f13{E��d
���}�ͣ=Sb��Ø��M�a��ԋ�5��s�3�GNdU~ ޛyU�j+T/y���n�A6���ЃD�ϗ߮SEF���k�H�c�5.X�B�����0$�5��#��l��l8�g�F�8�L=�C*�d�=U�Mŀ6=���"�ْ?�{{:>��
�e�;�e�z�|��,�[�+������u�8'�y�ATT��b��B���n($�L'6k��H��B��m�'�?
v�� ek��11W���#\$��Bە(>��)��L�/*ڡEH��y�Oм8�@�RJ��31^�
S˫��?��[�e�¶s5a����(is�������*����م��;�o��̑wg��9�L������� #��ĪǶ6�i�C=��"���r�ӟ��8��qA�R�c���kU��)�m)Jh����3������PfK���M�"���n�3����X���v�X�H[J��z���E�]�B��P�a1(QoCdxt������C�y2��4w�Av��b�%�#䄚Y�Ud3�ֻM���݅<Z;2��a���ͥ��*Z��Rڛ!N�.�m9B�'6#ek�6W���ͷ�J���������	 b�lܼ�3��[����Y@^�as���.��(P���Ǎ>HC�;���"��i� ���%2%L�Gہ�OF+.Z��2b���Gّ�g�Am�~��G�s�W;yфF߂ع<'��\PqUYO	 �2
���B�;�$r� pΏ4/�9,���:z�EB�Ƽ���b7�cַ�.+OGC���Ī 效��S���6o�v���r.�,1D�VLi���S���z�^�:f#�T ��1�t�2���EPp¨��,Q=ߗ��A煠�貳�2k���TM�Ӷ�s���/J���4ų�k=l�����X[���'n������Ix:���"R~6�����3ٹ\�jY�
�J�I�8g��|wT��3Q��5��\s��<�9 yB����Go=<4싌�h=X5��!�#-Sʹ��0��W�|�#�ƎN�����U��uw�Nk�>�������i�-�i������`��U�Éj�r�����p��(�s榶�dq!��RȺ�Z"�����7(e��P���1a)
Z��%m���iH;�3�sͭ��lu����q}��-�SmA���`�������^�^>I�j�0Pg��f�����
�U���>F�:M ��o�6$�B�B7�@ Z@�7��R�|F�Af8����3/442ro@y�3,+��<�6i(��1��C�o%ٰu�/׷f�B�l���vt��Q��v�k���r��n���!H`�o��l�qj��V�ϸ����폕ڬc���k�訂-�ӥ=P����=%��^����v����v�����&����Vm�j��B�_��' �^6��o!W*[8���S��F}�<iZ�Ԫ�#��B�h���&H��"�ڙPe ,��/ ��0�f�?z�tA����b��*��k�L�9��Y��4����X���wj�t�3�M�(Pra�}|�M�kPBH���O'.�Йt�#�}{~�+BW�s��U�g��M�8��Y�b�:��	P����q� �lCL�,2'G_����-���I���e��鿮[_��^�3R�H W��<�^�R>h���I��	[ϫ�H�{�Wa��HY���7T��H�/�ZC�@�8�%��5o�����ԇ-�M�-�|��=�ߔqw8h�Ax_�:+��I�c����+<���SY��)\�c~�"����<�s�1�c(�'kx�vnTa�����/�C�qX�c��ߣ�b���%]m��.kDl�`���^���-��z��
��B��<Z���v�N=�1~B/��A�@��hb�&�8�b�P0�W�ϰ�Rrt�[�̍o���T�:㬰@��i�����j{{�/rY��1��*���'�φAK��w�zy֑*_ψ�uΓg�ow&O�f*� X�j�l�^�,�bT_fk�j����������}�Q�n"�u��S�?\6qp�}�\�&`z���l���A�5_m����A@�}��!64����8|���uWC����b�fV���c��QF���σ$6��"�zw��↽
�.�Be6.�9I"rq�5)��@�q��������.�S�uo	v� ��Յ]x������"!��a�O�v�Q��  2�މ�#�i���t�qdU��I9��T !����LVX���d�3R�K�[���,Ī߸��}B�X�6R
�t�&v'x��ݐT��RF�9����F��&�|�O��^z��ӕ�M	f|����R�T�¹��oP��܀ PQy���4=������:�YAɚb�)�J����g�z�o����ቂ)��wTc��H-�Ԥ�n�c���V�=����N$���x!P�ď��-�*�b�EZ�6�`r[�5UN�{#��8Rj�"x����Bu���̽v$�^�#�8��L2�3�/I?7�%��ӥ��C�y��j����֍4Y�n���Q5[���g��M�A1��q�VgM�BT=D�<�Y���
��� !V�<�������}�\���I*�8^@��xm!��Zcb���=�Z�,`��bTT��+�����ruƓ�����C ����SvX����W�}�aSg��z�S���̇�-�Ǜ� ���Y9�M���#v���a~��Ζ%"�2C�Ae���t�g�������S��#]�Z/�������T��	��7k�53�|b���l��9�zL�D�����ZA��[�v��h�"{�q]���d&)���5���oq�On��y��q�σ��P+4�����HL��;��`�O�����������~���79���J2��;s8�����=�U��P�x��Zl�7=��d⨽�\�Ԁ�x�J߸�?�ࢯ��@sCb#����m�! "-�Č�v�}¯�~��_�asy����
����7�x��:2n�Sy@o�p���:q%]��~��j2m�!؉v��)�N!.��L�M�L��� ����хk]��UD�4��b�%��?�[>kB���a�9\N�=ǩ3I���놸���yyM<K�e6�'�R<���[Bq��Ι� ��F2�`���/{�CԺyC 3���k3�0*t�ٵ)�M��M�A�U|l��ħ��J�̪#�� F�|g���q�C<^�����k�j�M���Pa�0�gż�)$���a�tX7:ǋ�b�bD�/"Ր5&�|��1kn��%�[�^M���`n
N��͘��L[.]R���w75�ɸ��ڬ�?��� C�����9�/4�!�@{�Қ����,��X�B�M>�m32��h���3�p�M:��r�%��7��X,��0I��ڢ�����;�l�XZ�mk�;�ڻ��2Qz��j8E�L���t\?ш��bx���F}����p�JLG�/O�6kY�t�ب��D�E|�h5z�g�F������&sN��x�j�{�w�xo�8އ��9��a��ݙ����E�QI�'(���5�A�Krx6Ͼ��u�d#���z� �QY��n�C�N�J~d�T� �������~�R����I�\%;g�X��пi�t\X���T�`�#m��7��)�'�Tm���|�9�>Jy���($tp��m�羕
�V�. �wx����v���_ؖ�˶O�D˙���p	 :��Z�$vs�9c;}�yc�޿b������'�<"垿���:L5���_�Kh�~.!k�;n �Ρ��(r,tx��^��>���nw�_�^{M��f��t���ʳ�1�埆�$��қ�̜�o/����4��豒|��
�C�SK�8��h|N�w��-���<!���5��>��7Qb�m�ҡ��H�D}�����0�_1fm6t&�d�ߡ����\~��;ni�-}p�`NH���Cۈ����?�J��#�!�03���g�	-��"�;"���}3U͊	YOr�D���3���!�G�����e�V���+��S�u����M�{���>	����;m\B����rr����H�-%�iu����	���_���e�����K�a�-�~�^��:I�?\�#���Ü,���!�|�*�s5��^ ��&gc�D�Z��@l�T����N_�i<L����):���-���#{K?,R������"�dT�2�+���u�j�r�̺;�?_*�[��#_(��z`2ֽќ�~�z�2��S�q�)ڳ��c�ڬ���(P�L�C$�ǄǱ�v7G�p�9�V,�CI�n�'Bg��%딟��>p�E,�ڶ��x����p�>7ӈ�~vvᄛ����k�S24�;6LDG�2z[�R�!�����m����W��:B�lq����e8�9C�&��z��4�,V8#n��w�q�6������������ғܔ��|���s�D�C���ϚR*� �Pj��Qv�p��G�LԱ����YӜƹ�]�V�HSF�;�9�r�X>-]�0͊��7�g�3}�.�7�m��?v�5Q��ո#pX�׈���=��*�	!ꍃ�x���Y���u��i��c�E?����ÿ: 
�}'V�6�YFz��,:n�e۪Qi�}�m{����?䖝�X���v|ߘ/������yd2�'�����7�+�Wg�j�,e��H3��gxP�	�iD.�ꖾ2h���LbJi/��!z0(�E����-�7�Hy��@��ٟ�I �G-<5�4�X+�y�;@��*	\��aK�	q�e���"V�%2�v1�	��j[��y���Ǫf��?�#aM��T�?�M
|j�{�7�an�-��!����k��Qx�4��gb��r�$�h�3PJ\!Ws�S��_8@�Y��3���b�z!�2`����+))�����,G�����&��>�s�<��_�#nyC��-����B����|F���L�C
�����H��(0��"��"0�ǫ��1xѦJ`�o3�
�	k��y��+���Ԡ�6!HXB�4"��@ �RK(��x�Υ��=XT}�����y~+4�҂�!1Ď;����(f�$į������*2&��p�<�9=�Egk9�K�nl��B](�O�������[��{���(�4�Q�L�]^A��3>�yG��N�)��LJs<����Az-��������-L���_����M 8��ٸ녵�/k�������`�V#Ӆ5TC�q�V��s�>YT�T�9�h��T�"�)�`_�i��zoa���˄�kw^&=�
`��(cI�g.�b����4$RG��[&��>.[Bh��u�zׁ�ݶ^݇�����;�\��&q|�;�
�Y~=[L*��eP�kdp�ʜ��>�H�"/0�]!%ߨ|���H�))�tm�-�	��d�b1'E$<%�s�-[��/Pa���z8��j.���X�c3��U�\$�d��}��OgI�"�om��,����Z��[g�h��L�W��^:��+�n�!W��n�`g^��z�@!z�`ZѮ���Df4`��Qp�j�p��:��X�t�o���Kח?��{�`p�~����~�;"51.E�/�<���FՋ����O~�'j��u�@�V�]K���?�ybǡ��e�ɧ�ֽK�E�"'�w��=ƈ�V����5@HƬ����3���2k��0�O����ܫ�b�,Sx�fިz�RqLb���������2��u`�_ָ���;벃�-�3i�xW�\�Y �Jq�=�A)�^g�8]g��GR�I�Ǆ�؅?�X�j��v��O��Ҧ6�ق^O�H�d[�B�ؘ.~'���r��⋢��Q[�'j��(��&�;�]W�;-�SLf.j����5��O1����B�ɱP��<k��5��,?X<��؍�n���Xx�@/3�M�n �-|�/���d���?(��r��^�r�����S�m��]_�� �×R�.r>���p�S��|JluHRr�����f�9B?/}��7�?�A]i�R�$��(F����𣆢N���3;x��G0/�[�����3�j�Ű��7-?�ү�m�c"�n���*��}������}��/�	f����|��o8{�r�y����2Ҹ?@�*�.�E�@���3��$�	��T(Vy����.��)��L\��b��rN��r��ŉ���z��a[T,�>�v�o�>�ʴ>4�����〢79��ͫ&u��H;	w)@Ϝ!O��(��T
���놾�V_7����
�g��>�~�è�#V�_��c��]�<���L��΁��H�:	���d�
մ�#����BI�p,9��-�:͈8N�=�V>}#�2���Ê_Ӄ$��L��|�E9�L��ڣƔ��#�Bk�?��$�7vƐ�n6ϩmj�o1�N��w]8rmoh������T�p�@�Ao���y��g��Ly���7��;_�-|�f�0�B�+���o���.�?�.3�!���vD�N���RWW#�V�A���{�ߏz5�hs��*Њ)T��ӱ �1�~�U<���P	m�/H7�Hbɽ ���R�����g���7�$"�y��e5p+���R�l�a�	��ޔD��
��$ꌡ	�2�	
0�)0�n:%��*���S��':��`�������0�����ގ7,TU��j^P�ά��G�:�P���sX4*�TO�hpqmH�댥"B��LY?�.T�I�# �뷕���?�Ӏ��re��:,��0)�ġn=�)�ae������9_]����IÓ���by�D�كx03�{�#�����8 �'j��� ׌$�Y�����#���0�yLNW�PcԲ��d�$�R�!S\���ti?\��u�˰i���> g�)M�e7ׅZzP�K�L,R�x��	F��`���B�!�Gv��4	8 �c6�B�)L��3��4\����+B�T��L�Nס�}��M����U2���3=���A���B�c��$���ʚ���N�G��O9 '�o�&&_�spa��o�#���W� ����D���, ��gNN��c�X�t*Wz�9��h�CS����:��}���z�����s!���>z��C��#�V���:G�d���b�٬�~z�'؏m�y��/$��S6gI��<��1qN��{�z7*^.3֤"D�[ŝ�]3��[1a��oJ|4��Z"<��X��b��5
����?�	t����,�u�(�\F��-�\�ɰߚ!�JkIQ��ǜ'�PI�8	��%d�mw���Nz1�O�e�<���. �~:�\�Qa��|�4���s�1�i�k5Nkz�yN
%'�L[U��������#�xv�񯰭*}k���G������7O.������盦�S7�=c���ck��$8�hG���{_`�d�iK*��Y
���W4�zy�>�dT���p
є.�XH
��Ue<ZI���ِ��O�Ë�Tڒz'��M.��� K�3O��7Y|bQ�\�I�ǩ)}�Y$Ǫ��W_���m����?�ՠ�;/�SV�儱���k�޳C+�J�=s�W=��8���k��H�����/G5��x����tl>}�R�y'G��FC�7�u(�q2��e��Z��9�׈K��-�L�)3��4�� 3�Q��gU�̛�S5I�����88x�#d\u�o Ԥ�=s�L�k�� ���1�a\������Ւx�P�a:ՃC�d�w�˝���P f}�oba�>��W��/Cz5'��)�B�E绻g�m>�h�l��`�n
0��J���~��f��B�C#�Y��]F���<����)4 (�Y�����	񙳎�r���<��U�_� #iۿ�o䬦K�._il���ς*��SY��,����|������IDl�`f�I��W��؞��͊�}��g�ɦ����c_���T*D)'ț�\�wR"g��p��p�S�_)Ī�{F0��G�)c���XQrY=zC�7�	j� �<A��.$��M׉Q�/:����V��s�R�sU�J;|�q8ZJ5�	�[���d���/�{�TY\5���	!���4�� ��zh�4��@fˋ�1��zJ��
.G���O{��w�C@FTBE��)79v	�cr�����f�����
=�>f$j*סWf�Z���Pj�U�A�f�4��9������!	��ƿ^�8�s�Y�:}�8F�^���0]�$}]�����ù �5�H�ܴ�k?�h��W�r35���sb8�׎n�k��a�����E��6J��h�@���H�<O����/�ߓ����u|e;���3�x1�l{��ns�ό�ȸ�o6��kp!qZ����K��J�o��t����J��G�{]`N:���=�?ꡘ>���`���>>��߽p�
�0	(,e��Q�X�Y�lEe�U���f���o�$YT+��.�)1�r���?x�l�j�1$�*�H��j��*Ψ�w����zf�zj���5���*@;F~=ngĺ��"Dz#*$�66xW��>�W�688
��y�upף�
� ս:�ɜ�DO��Έ�lh�H]7_�0܉zd�p�0gS������U������r��(���=±tt��;P����+C�vg�q�:��萭xJ|m����[�N��`�O�)�7}{�`�zy�o��p�mY����0B�|Ԩ�C�e��������}oY�J!KZ��'��>�N���c�R��s��p��]��i^$"έ
�0�M#��B(c�]�<����v��A����i�ݸ!l)�����Q*���+IhN�(�T{M�%~ �EQx����$�.���8�^2�Wi�w�͘Vn����(����Dlyq�\��4���ڎL�N��
����ml
0�5E������@��U��k��d�b�ӛQ�#�Q���s�ˋ墾���Z��9���B��s���m�/@�AsqB�����˛�%�n���+��N��'�C��,��Ҍ9Ul��%�V?��>��*|*�	x	�-��Y��2	1N�g���b$��cC2Vmm���ꃶ���VH��>"�B9<S�Pĉ'�
�+�������x��_(�hy}��&)DR��s��V�^8��Pn͟IH��Qw��i&��^�l��5�w$i��C6�XňQdR7��mj�O�ޫ+,�OFa�8z�!���*�~W֦��Ôi��|'��y��ǅdl$��'�a�'򊢯(�F�����S�Ϋk;j�NZ`k`^|ґMk������3�y��_��t�%uݓ�~�G�b>��Ԑ[c�^��+a�<�y�G�>m4����!���=�l�<6�A���0�c�r�UQ�e|�@�K����d@I2D�srm�6�������9>���&���	,�׫�#f&�H+)X�]hG7����BB/������ZMh��E�!���5���C�%E��Ϣp�j#J֐�b��|:�X��)�����EJ>�rz}���c��9{�Jň��]21#vE��5�B������-�Q�Ӡѹ5f��?�\�-*1">�LZdz71ׄd���N�k�!6��:"�b^��K ��α��+�/.S������ņ���Jr.2� X����2jr���QP�<<��h�����mi�-�.�մN�4v��
Я�.��oK[(jj�Ѭ��T[�;����E0.8-���
����c�H����	���l�~��7�U.s��r^�����}/�W#���6�i�2Hz�6�~+P���� (���:�s�&���VǞ0��o�!gs ����spv|�jh�b�<gy�<y�.
'zuػ�i� (V?_?�rH{���<F ��5c���R��mXZuO���g*4���t�l��/<��v�IS8�i�E~X+U���$��� � (�}��6�<���VX��T�Ӆ$\�b`�Ĺ�	���ܻ���$C�4��d�Ă�^�w*�}�aJw�.���~@/�̽�n�8[�˨E'���ܢ��-4���L.�[0s�-i3���B��8����4�Bi�B�D��lĸg�h���`�����Y���ݾ`�,�86���v����V�u��g鲿�!n��K�EW2K�7�=���w�8�Ϥ��[��Q���R����5E�Uj���&�B|m�rx^�I�M�w��4�E[���X��OK�V� b~�jS�KP�v���`�~��	�+sģ;��Z�4��ہ�t_�V�*�-�a�s�c����F��&�ʂ�eZ�]j�pf9S�v z��9Y���9+w͹���5�<�^��t��-��+mo��'k蟻�U���+��_M;����e��/2  8Z~V�`>�%��9I�[�4�>$ȏ-�?+ 6����x�3:�P�J��m�˦�fcEmC��z�����=\#������`ߡt�Q`C�����_�p�D��2=�Y~\[ۀ�[��a��M����|j�vQM���g�{R��ǲ�]�'ܙL���,E�+ �,�Ty�=ۜ�f�!>��rKD��1�C=�W���D,�j��l�2�z��gK��aJ���e�\c��9�ρV��> ]|�k�W��ow����� ����{�,ۃ���\�c�g�~��c���0�+ڄ�������4x�@D���6��;7}�����s�x%��LԳi�Z�F�\42�=Q2O�ب�\�V����M���u�F\�8`�%�cL
��5#��^~�s[���s�Ea��{ܹ=r�Av`� l�-�'�|7 ���k�B9Ed��G�Ce�4��-�
�_�`wl���y�c���QFO4>�l}�.2�Mh3$6�;B��}�WT�6����l�[�<a?q��=%�It���wJ�=?��c��!��a�B������Q����P�����=�}d2��ir��{�D0���\���_�
���Ɨs;��Ϊ���󆻲�~�Ѹ������Ks����u��RRF��[�K���b�L��͑��0�\�Ҋ�V
��Dh�#>�6��C���S����rVpŹ׹)�e����ʉ��� ������ �n��騶O� 9�!x�{uw�
 i�P*B�7�HF��͓��Vm�јBY�U+U6G��
ͷ�f1���|�ތA�x��ʥ�E���mfX^�� �uJ�1��Yݸ�
��-�4���Ȱ::f��`<���vuĕ]���<5T�3��Iq�V r�~9/�t��(�|Jr񠤜r�%?Mh���?���\��]!�&[,R��k�R}҂���7��YA!t���b@�n
�n9���
�q�N��J>6C�<KsuW�/Sw�qR7�][}MOBJ��u��:�>����И>����G�z�e�u=�MqH�$�M��#��3�I��F�;��*>2$�`\�'쭃,We�t�{4&���G��e+�R��[q��N��铚��qޠ�^�ݺq��J1�G�U�x����^��vcjYR��G]9ԥ���g��C+5����;�$��UK� �z����
c�v,��-��W�<��M/G |��v�X�zӷ�,\|��>�߇�t�o�A�R��10v���I-CQk�������T��ut�� ���径ڹٻf�v�`K�'g7ң!|R3v�ʇ�@*�u(��/�Tz��s����Bf`����"S����~���ְ�6W=�`��e�'����{�����XyQ��f�S��a�O�	���k���Q��ŪDM-D��y=p�]�jaP+:��v�hԕ筕�O�R��㜊>�_��_ �Q�P�C�jf��P�(V��8d��ݍ3hX��j��w41L|��d~��.g��Q��?'���A|^!��x��~��G�t��F�eկ^Q'b4��q�����zmi*�P�h�R����K��/J���U}���U4�l�2v��Vқ�� 	Yl��cc��y��Z���P�|�0t�r ��r�e�hklP1Ak��b��p@#��1�A�������CB��{L���\���iB#��L�n����(�zn��?uY��~����Gy��*�N��3�,C%$�-W�J����b�fNX�6ɒR����������]S^�mjmD�dg��خK�g�N�-خ���$L ͇��T�;��yX��v�����*�;jS�������;��l9��������ȩ�״]�� �lM6%��,[�[�J.%ֹ�J������h��-�KFc}����:� 0�<7$�<����&J��8r�d0ߐv�z�
⛉H���.;	��3�L�t��R{�>4����������c�w� ��!2!A�by)L��0�帇C���a3vqMR�p0K).�.e~�|�u�����Ri$r�3�.���rj'��İ�!��@<m�z�r���y���!������.�|	s��QI�0\_�F;f��mA������,V�����e������<_��ʛ#��SC�&Z��$��o�
�y��M��rq0$>EL��6 ��H�������9x�+�m&я�e���즚� 힩�l�
-��vK��3���"ȗ��-{�g`��,RVײg�AS��o)��|۱�Ib�3�9� r	kv���Z�Ve ��.�P"3;�O?돎��!,���ǞT�}9X�dơX�ixzLa`3@[���=��
�3^�<�
�� o+,�ĥ�j�)-���Oj�Wi>���a_�H=�m�{{8]*��ok֛�݈@�̒C�"�[���ٔ�D�9��'�eb������Y��\��&&! ��7я�����c��?(<�S8���P���qt��
��D��4 i��w?u�=������S�)r�����W�H������ݖ��U�yWO��J����6Ȃ��Ik��qn�i��ML�u2u٠���ɿ�j�i��Ѥ��K2M�9�6��zIMz�.�gy��Y���1A��K�&V
%o���X�gA��u\�X=$�e689� WؠƥM���\K�-�J�Qآ	�t��B��2R\c���x�`����f�j�Ϣ�m$�1^BH^;3��3�����t^ r�S@}8��q�.H�U����NB����{v7)�d�Kx as��%�Su:�}���'p�g��ژ�S��ܢӊ��Vk'v�͔�P�ך�IQB�#a��X��3�@`Z�J��vqH"��F@�=�MHA�yo5�ԓ"=��W�[����ch���5�T�:c]Ùs����">�.]��.�+\�,�_�m!2�b�f ��7���u
[�	,�6��B�^�p���E7�>J����)�����mヤ�;�L����갍3��i6�dW�#�[�47�^�މz�+§�#,o�0A�L�XQ�I�-կK�;�����E�� ;���+�K�\(=���
�͓��6��B�	��D#J-�b�{a�@/���$��{�ѵ;#�j��sS<b2z%TH�vql�Hh�������UI�����@��=0�!6e�1�:���fȊ�[�c~�(�vפY�i�g��X3Q���_N$]L�&/��;A�#wt�?|��ُ�vh��^��P N:n.���>�1׽z�ȼ/�j�Η����~����)��q��V�bs�/�˼������_�.�{f���Z��$ar
�=O_��J� Q��ɢ���o�Uy�J` ���3;�4��38��Vص��37X�V��2��!\�u4�Ϸ�☰!~d=��_�����eA���wj��?lj9����-^�
4V�iz}/����I����&�ץ�qT1��i���3g�|�sq���S��j�*HzvD;��RHr���nx�c�s����i L�|��o �w-�Q��,�o1rg����3��Juk�q�L�������Fb�s�����?���Q�
����_�7QH�͋o�Y��H�E��.�d�Q?�g�F���r�y�(�Ke�(=�L��fq��#�:�d����ˉC�����-�h�D>/��YW��h���J ����O+��	D�U�zDLAJ჎��^�_B v=�L�
r���T%pDΝ���c+���e����pCC��^����BZk�fl���߷Dlr8~K��[�8���	[�}��>4�:O�]�#;�Ӌ���YU?�?������n�^"��H����2}0a�3�ge������G�GB��	},xn0�/�)��j�}�ҙ�@>� �������2-D��H!�y��1���@{�(�?i���)�������#z>%U��ٹE��C�k�z�>A�� ;� ��AMS�e����D��Avס"J�+t	���I&�`�@�]C韣]}�;=�	#|����}s$��@@2��>�x�$���3w��h�k���2��T�a&��u����!��yS�:P��v�;H�������Y�``�$B������Il0�Σ�w��4Y�l�t8��tҡ$Iz�$�+t���VhCx����Y�M�0m�&?Xh�h�F|��a��d�������Gw=w���1-�V��e�gq<i�_�=�}*�R�."	w6 �q_��y��K�����7��j��>]�D���XRSc.� �<@�J��>�'��
�1���VД⹪>�����j���λ��p�=��r��W.4������MӮ��[���Y���pknt2�Zǋ/�����%������(��8Ϲ�r�e���$��7����ͬ[x��; *Z���Ą�RO���	{��(�~�Ӈ���H��yb���$�j��-���}G��33}���Ǡ�\�`�|u#W޽����i�Q�eǩ�[����D;Mi�䛔	.$�V|�"z���>P�U�qY~%��	�^�#�X�`̇�9^�.�+����f���DW�u�5Ua��Ǟ�yŦ/R�抂H�.�O;�,-�c�Bѓ�.��^
�e�qӵd�e�!G�1K�z �����F����E�,��|�8t����Vf'qJʹ��F�K��F�(�D���:QLW��c�BŨm�.U��7�˅�ݪ�"����׳��V��vN�V36Ǟ�V#���Dd9��@�9}�ᕘ�]@�1A���������(�i�*��ѳ�eQ��~j���a'��*���� .��$<[�8��
��ϴ�P}��yӗ;�M�/��g���b�3|�M���O$�D"��z�l2�ϣK X/��6�º�S�/QYή6�����o���i��'̈5 @\�N���v�/�}[5X@Z���=���P#��IA������z6�$� ���|{���li�D�-���=۔MP�n�'�ԚG�5��E�uHư�{V�Y���h�̤�#~і5���t�8�a��wӥ]GEЫ��|<%P����H��Vd$���Q�D�?�����&%��j��m��TAn��OU��AǄ����x�z�Vo��%M�,���Z�2�[��Pn�h���b�<�(�Ǽ�l��c�$�{��	����Ѵ�'EI��`�X������[� ZI�	g3��ή��)Q�����@�=�4�����₫�2=0��n��ЫӘ��eE������>���[��8BAƺ�
c�b�����5_�&�<�$8?gN�4M�)?�~zB��c��}z&�~���cq�P�W�Ĭml�3��/�`.�`���?%� լ�],�b��M�2���p�:��
�5����d��/�N#��� �~Fx�^#MMo���8����+ۣԞcd}o��͇"AW<#��6�G��<,K�V��M5����ӹ9m�8���VW�������?Q����������
��赬��m���A�%0�;!����(3�g.�V��,�qx\����mB�#H2�>ɎJ���V��{�&a|	����i�Z�)��-�
�]v*��IƁBhAW��P*F]�57)|�Ȕ�]t3a����%u��O�͎h`?ڂ���v/Gy+ ��	j`0W渆"Pnx�H~�k��o��v#w���b�(�X8?[�_�8l�-�Q�RT�wLgQ�Ӹ��Լ�Q�W��� ��i��a��g�-��h|'��XtBӀC��ؾNK����͌��ԯ�lj��F���2�L��[}�������?�GS>�빔l{�/6�!�1����j=�0�K��C���G=?�G��m�A��Ka��q҉xsݿ?��"�w-�~\����Pr/��~<$��,�ʼ�H�G�?s*�o'�,��h��h�,�<7�;���|2���}~�V%������X�b�,����TH�)9g��D�k�,Y�;��m�`X5�������F�~�\}�)y��୵�D���-z߁��A�`Y~��1���x��eQ��L}tQ8E� (�y��-�h
�T+5fw��h~��f`Vx���� а7�Ԯ�(]La�����s�$T��bk#��fo�1��>>~R��h�N�vW�jρ������5�s�m*��G�>�d��`bE~�?�⊩�u�
�.0U��n;*�p�7�AѺ��9n$��6l�%���:��)�*G,�r��㱞S��΃G��=O��7�Y�W�k���VK�B�R}�Y�S�z�a2;��":�]�K���}�NcY�֫w~o��:�������)[�A��4� ��L�a{�Pߢ�yf�N��p9��`��9_� �h���5d�h)�}��8 �M��$�����K�,�i�D�$�0c�D����a�ǆ�]��A	�ՅdaIU���`mZcT*�ѨQPP"�¿>���3�W�C����ڸ��*��WE1��Ůџ�ɒ�;d��V�X���dr[�7/�4Ҁ]�䍾'v����s�	Z7b'���~0qö