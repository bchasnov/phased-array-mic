��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\����q�?��e�I8�b�Ǽ$��"����ׯ1�V0���g)t,+W���LY.=�(=�SI�}A�S���5��h��P�D�%���Wp{�5+��u�^��:��ƽp{����K�N���h�v][B�of�^�/����Ο4=#bP⯃��{e4�B/�˼V4���#F�G�2�h�lU���fo�(�2�QV8^�D\�c�?b�#�����8��x�"�'�Ŀ�n��G��w�qj�ԢA=Gä���e;ka�#v��:���%)f��M�T�����I+pt5f���_��ؚ5� с��tfO��J�s��`�	�����e6e'�{�[&t��Ā�]�HQ��[ur{oE�r7-sӪ�2nѥ��~g�b�tι-ɲ��j�Y��ܸ�0�T�t{�
4]���_��.�k�m��:SN��,�i��٦s#N��Y����(I�XT�1�gm6��9A�
��IfJ��h�ӭ�k#�zW@ѧD&���P�Ն��X)�]Q��B"f�B�Nq��ˀ1�h����V?ⰿt}�����o��~�:y,Z"ς~|?�(܍���i�M�Gu�w��׸d�V77����?c�M�VmDJM���ѳ:A�eD�X�.9��}�i5eV;ʰ�0N�>�(�9�P�H��0[�A`1Q��6�[`_����S~��x]��0��K��(��]�K��pP�nrc��#�r��Uq�a�U�'��χ����HM)G��w����Gx������]��F]����<�+��`x돍�Q�.y����������%^c���g�i�,��Yl�nH�����!���خ&x)�q���1�t���nZ)�yr���	{�'���}[��q���rO~L<[�6�N��_�<n��&���I�S䈄�������31X *���ƓA���J�X�4���d4�aH�y)���H�Ko|%)�qi��s�I��g[��P�%�لܐ�X� �YP�`�Ε��>/���P�K6�)�+:����w�z��w28E��^�ִ�7�ނ��f�0�S����-��f�V���2�i�U��o! ��H%�~E���5�+� ��X�ݿ�z�,���q���D��� �D��	�{\�ea1�g��*4�>Һ���S��^#ysR�8�+�2B'�*�7�&ÿ�Y�-��Dh�6�a�}os�tR�m��.�W�eb�f���#:�vAd{��!��ciW\ ���X�%6p��;f��_�Q��$h�а�4�~�m���G
.P� S�f�c�C/>^�|�ԁ�������^@�
���՗��k3��Al��!�4�W�E�v�,[9+AJ!� Ӄ�9�Q!'@�G��� :��d-y��r�<�� ,���ҭd,��my��VqJzuU�6AIj> i�xG��1����"�3A$d�ŷ�M%��)��b�*�HS�3���Tƙ����5r���Q!�W��,�~�
R�ٞD~}�V��]J�ȱ��9Y�X���]��9����Q;�ͳ4�����nF��)�a�;���WV_H_�s0:0"n���Ե���n_W������@�#�ɚ�� Fi]��>]������D1pp�^���9�4����e��hGJᡎ��\!�ۢ�ސH����_�	��)�^b�s�d�Y�ކ��_(�-��i�=vqP�����f�=rɒ���=�%�z3cr|�mY���2�_a��w�1_��2����=2���
-CQ
�J%l�=)�G9)����Dh�.�� o��*O�ZN�>�����d��(tY�ǒd�t}����wPX����� ��}76�Y�F� 1��5+����G�+7�K��Щ����϶E���6�hbMg|������ܐ錙��"Cn�+ߨD̟��~�$��\_/�Oǝˣ��h�RE�����|>�����J�N�	�M���;��7��Y2A�ԛ�X5R�1�Z	�U���?W$^��9a�<����g��<
3SEEm�逗�[w�kj�qk����M�_n3(��ۓ����B|�fɶ��G���®x�	�zq����a�6z:gV�u�L�'(���F��%���2~d(��]5��5������J*�u�Nj���� �`��j�0���;h!ז ��r�O��ȳ��x#z�}������ǹ�N4��@���[L��D/K��o��������n?��QG�iȟH@����-Ed�]��_ؐ���^�,G�ؿ���ش�������j���U��+�x�.�����GƍSaW�����K*J�@`�f���ca՞к�^e��.Aɣ!���5��m�2eY\�lD�Ј剑���~���]��ʋ1�DU� ��a�jT@:���'�<����5%�;<=���Ğ I|�S�������O�۰�]?s}kx����벴/w��Vz��2�����F�� ���O�wan�N��EH�nig"�����g�,�@A������!dـt������_����%�� �f�I���[SSG@Ĵx��? &�O:w��vm��UT�MB�Nx1k��Ut#��%��A]�m|�P+Ks�g�� }[�	)��n�������/>L�(��aʄ|u�b�C&^ X8��g����(�6Q'�8AV�0rȏy����9}��l]�6j��撱�8� Li7�7�쮘<��?�
ʔ^YC�>∺�9�6haۦ��>+��[ט�	D)F��O�������z�([�i;!=���HψvH��O�\7u�ը]�@��h��O���c2�YIXrV<{����+�c4�Kz�U	c�Wp-�Cw��RͯO��@�.^�m��s��l;��i(>+�8�����4�*L�RQ~�yLQK��BK2��\�e ��7��i6���V��\Ͽ�z}�3�Ă��6�U�`1�|I*�A����^�.GI���L�H�@"���K�E�LS����A�.���Dp�Vp��
Q��1Iʵ;�'�҉�WDY���a����}
��ūՂ̸F'��X��� 't&?L�c�JT�oG��-S�_p�ۼ!��^=���,��,wu֏����ҿYv�E�
8e�$���?�h��a�f���N 	��T�@����7"�o��蠺�,��qG!�� ���
6ĸ��t7���cm�_?oK���'Re����uI��b4$�Y{���#��Kd��hDJd���OX)>��I�p�17Cn�E�Z�:�^ �o�'�G�Nm�w��-߆q��#�����t�9.z�]����eJ�>Ν���:�+f��!*hҜ�?¸E��<��]l�m�װ+*��'�m�4]r�Lνn&eҴZ�ŀFlz\���3H��ҍ���5IHO�xHNu;�����.�)��*�ɟ���h����A��Q�bmsk�c.��!�=����>��wJ�q�ċe����l�D^x�)'��C��6�0�F3B��$0w�v��a�I�������W �a�� �i��F�$����ɨ�V۪!>���%M���K� ����]k�:�ɉ'��[���?.����Knk�����Y�2r�	4ߌ�ͦ&��/���W��E�k�n��l�3=��VB�0�Z7�h#����B$�4e�A��Բvf>����s�6�tB��d��� 2��K���P��Y�\v�WV�RFÍbe��b�����_��ؘ��c8�:��CL|B���Ȏ�&�S��Vni�<��1~w���&= m[��s�j8�Xٷ�񁞒����e���o)����A��l�8���-��xWƨȷt��"��_��6u40=�^�C��@/����Bp�s�&�mo��*X����]/t�}��r�Y�1	��
��������?�����*K�G5_$DڡW���߈��,��k��T�٤���:sp����nL7����"c�փ��r���3�	���B���
P����aFp�;Nu�B�>P H�e2���zc���hn����=u��	�?��~�-��9kڸ�\�0�ۄ����k$�߫���gLϏ�$ѩ+�t#���u0����O���w�S0��E*홅�MӗT������],b5f,�e�v����d�o�`FMf�d�3�tZ��\�K���+��Zu�Ǟ�_��i����9I0��Snw������G*��92S��(4�^��X<;�������%�V�I^����ڼ#�'���*w�0��eI�{�7W�ô)q�`�w��̡=ZF�e]:O'9O>�<���\D���۪��ku�-X@熧͑T�Ђԍ,��qM�v�
V���E_��C�*�i	��Ӭu3��������!�C�Db}��jv7�C��5Aqq��>�bʥn�i�����F
�j��$y��CG�@�|U�og���V��X�x��PυŰ�n�b���O�y^��(e����b%>��S&��QzT�lad�����]��VSF?��A�Dy4�Q_���ϟ�6x+�5ͪߑ~�������� �V�a��������/3�<�O�9=#������r�S�>�Cy1.T�7��F|/9[	k���-�KJ �U�i�[�f�e��,1�Q!�!�Gؼ�o��}�����ԥz<IZ.��9�F�?�Х}���"�޽4�]f���& �J�^��[�g��p���	2�"��O~�AG�b�jt��v(=���^	���w+����*О&����<z2-k�n���]��~�����qd�[��rɃ��,��w�x5x���v!�.���p�j]Nt	�0���P��*�%�J��B��b�њ
�a�.�&��_�#4f-:�t�0.Y�_.<�G#E*d�!���&Jї��0P�
<t6U3�zjE|�r� 1�t��2֡�и˸Al�t=�1Jv�%?F�}߁���xQ,�8��ӭ���GɦR3۩%�QN������.Q�OoRp\{�P���a�fO�rMx>$�'���I�VH&�Ѕ]H�1���e+�#� 
���I:F������c�@�a!��Ft�������L�;"�>@S/��{AW`���3K�f�� �|^��e��+`���ʅ�,V�����N��
d�Ѻ|���hZ���0�^yX�n�	�#�V��ǵ��8�÷n�H��+���7I�]�P֦nUO��0���Y�nhoi�Z��NQ����LN�}�I�M�\��#�� �z4���/��Z.M�o����X���hZ��m�����|QSqxVk��Ǖ�q��7����������#H�8��F]'� *�E�c��yˬ�k�Xi|�a����dHm��n��rҙ;��>�p8n�h���\��v�Z1���ӝ�6o?@� ɕ�(�W㕷�SŰ���g��O ��A��T���ߪ�!�9���E�w25)�#�7ج���
�.e5\@�O�A>$�:���U&ݵ��+_G�(X��H�6n��!����{t RpYx�_Z���m��`~�Z_KWX�0�L,�c)�sK/�K\3Q(�0�@�k'\(O�&_�:�&,�K�A���؉�$�6$����:~�VD-�Áf$�����ȵ9�7q�[ڽԚ�h�/�)n5�&��.\Z�T���H�[��Ԋ��Y��C���^P���Fl��Y����F��nj�w�a�ҥ�kX�1�7���Ȕ�Ԋ_�%�|�Xw���D��R��V{�'�Ӱ�L�/��~h���#y��5��Oei�F�;����ۗ�%�ڃ����U�hd�����Ků�|X��4�L�C�Qѻ�B�8�s��*]EV߀��d�Q]X�c��_�5��p<{D?����R��oJ�Y�jY�
���n<E(��g[�jH�"���"//�G�vzsI�_��N;�jy9�Td�u����r|�×	�c��b2��Y��P.��Ya~Kc?��q�,�eƢ��!L���~/�l��иL� x�El=ώ�!)��L�_s��a���>,�s��L˲GP����tQ!�+�&��Q���zX����eP�>�j'��A�֋�7�XՃ�Y�w+�B�uy\�~�Us/^v�4��Cg{�����u�#^�V�R;9�m4�9�8c֒�<V��ǯrY��iD֝�w ^dc�Ɠ(�Y�o�p�sbUvSLF���@yףq4'����*��`#�r':���-�|m5f��iuJ���fR'��'䀼��g�W]���y�V�}�e�W��5^g�OK�6�p��Ʒ��*k)#�v��Z�l,^�]�?ZD�>�\�]��V�es3jx�X��PTP�����~.�:}�2v#�q��K8�K��%t�E��z�]��h�10�"��Gr��b/��cn��ď\,�Z�b�Ao7�,y���;[�	���P�9�y`�`s��?�u�G&�9��Q����d�^qu$��	�Z�kT5)�R�2�'���n�;�
���g>E�����I��
zo�dh�e7�"��r�ݑ��*;�M��U��f�5������
�u�����e�q��]>���{2�/�-�G�Ҋ ��'Vq��b�c{�Dwi�g�}H��و���r4����{��l��L�^�&: ���>C���z}���f�s�dsBJ�A��Fz�3�2�Pz��D�-�J>[�9�8%�B�����c�����9e8�gg�4?<���D���ȵ���F�q�pP�d�
�X��Y���axb��Ϩ��M����5��$?��\�t��Lj�if{�P�n1MZ��Z1U
$��@CIi����9N1/]�r�64nI�����
"/ !)Gґr�h��&@�B��������ٵ]@�+�zt�mh�xO'�|v�H�ä�d~A43I�w�ȹ��덠���N3`�`#{ؗ���j!�2����X�M1�%���Y�C�1ɶ�h�eԲG���+�̋_ұc��*�i�96�Ǭ*e���ܒ���L-3uyI{���)�hkQ���Oi�m�o�ƕ�p� J/ʫ�,�*RcedsY���W���]�<t����؇���=̾���h��.��*_�iq7�x@H��7�r�E�-��~g�c7E�֯}U*Z����V�dDؑ}�wB�}��O�aZ��gU_�d�mС0'A�<U�O졭F!�<i���bh����?h E�����9S�Qܥ� �OgJ�p��])���P��d%�P�~�ڦ����oE�-�4�~f�s쏤��/Eׯ��SĞy��7�"3�1"K�E?�̲ޢ_�61��^�j�����)�>ګz���G]�<���pJx{Rr���bd�7ܴ2SU�X&8�M���E��La+�@��r��N�����_�TԸVh���T��=>p�@���E�H�з�MU�ʔ���[3�����U��P8c1�{�L�,*}�3gp-T���h$	��I$��Wy�a3���0^�����e��|�h���3��)��ĵ�뤦b�1JM���3:���t�y53�4�E�n���$}Yj��
i8^	Ɔ�S�s��f[&b�V�6gW�Ke��q!�ׅ�D["��ɪ��b���	�ַOxb
f�7Hว�*�(��K±MRIc������ߍ�s=ǈ~C�V{�jd��"G2��#�Q�ZK��m,�mB�����
_���qH/��Y��B?���c��w0GT��A����9���c�O����x�jE�d�Ӑ#��`Fq��f�k�,�Ͼ���2a�'�Oh_�	y��ׄ����~�:�u�1���Vo���暴�NE���;l�h�4�4Qڬ��H���Y��� �\�Jм��A0�p����qU�Ngu��۳�u|^��z�N����I�YT����Q2�(x/O�g`p*F%�	�?���Zm�j�hzD�\�^�Y�+�]�J�M@H{�D%J�b�9��!qm_Ʉ�{;N�z��p̊����ޢ�e�&����g��؋(P��f/����dߐ؆[������$����ƴ���������%�0oQ[ЏK�ö��JO��Z���{��Fz�e�fS���!o!O�\���z|�޶ً˓�ٖ��Ff.��Uguݏ,��X`X{u�
Yy��Iܡ��Ȳ�iJcOqZ���������DOyY���O}-�t7��6A��JYNE�\�؊-��Ի~7����y��8���w����y�e�/T-�|�5��q��}L@l�G�.�M{�������z?�K�cxѵ�V�:	FU.d(,��v �R����h��>;2U��f�C��/9�Si�DB�}�z�]���ND�H�� -��p�6�F`q���8Z�!B�T�!�&�FG����0�rWȳ'6
�.�Z%��Q��܃��[E�0�9fp8q��e���6F����_�
$�㉞r���؜���匥����G����AhY2ӊB��t,�K*!P��M��^�t�t����)�ydG��o��1��s���[��h;�v��ƫ���vP�flO9:a�y[hmҽ�:�y��|{�vt�,`y<2~p��X`s V5�e�������JU�!�N�u\��XP!�	G�Q5���?#������Bf: (�y�!�5��Xߒ��m�/��ƹž���ך�+2������+���h����!�p��6U0��T��'���|'����-Ĉc�%1�n6d쩘�D2֫U6D��\sO!��:Q�)}�i�F��%��W8�z� �A��K�s���D�}�inY3X�>@�>n�YZ�fu�[�T��5��M#�M�����o�#o�X�kWog���7�M��K������`:C�	���Ǵ�z$!�v�������%._u��x B��d��.�G��$�ݴ�M�k��PYU�8}��w�+"�50�mN�G|O_{P�:�꾞���
��7cg����~�F�؟4�˚Џ�ؔ46 ��#�M#��t���Ny�1ּN���#+�j��������.t)9n�9��@����B��D��b�S���ԙP�\�s���J�[ʰ��y"ʄ�\

y�1f�Ez�p��P� J(m9b'E��N���ԬCb�_��,����>��{�O�WD߇�ςs�U�,\�C�-���<�Ҋ�z[_[�5��2�0�5��p,ZW86[�W?[�AIS��L��a�7�������4]��-�㝈���2=��޸	��ƃpoPu%ɶ�)��ê�;��{J���Y����D�A)�O�^�]��BO�Y}L�l����a&���ш�������_�QÊl1҆Y�Y�l3`V�1x
�3�\���e_�iIB+Ħ������9F�U15b'/򻜛��C/7A7��N�p�dD8w�_!����U�Z�0�$o�	1�S\��l{:&���T�ꋻ7!LK�8��֣x���TSW��@��m�����	��o�R��@A3L�lVz�9O��3c9���0=K�(E���D-D������?�TrJ]�)ߖ��3)�i9J�q3\s�[��G���$��*�y��F�� Dy{V`D�p�Fp�D���z��x���s���|o;&�G�7+X�cZ�:��Cy�u�2X`Z|m�4����Sm��:�%<p��D(��֛���z�"P�d�c��C����<����N���9@+�r@u�,�K�%�a������a�@�T�K�ʂ��nD.w��-d4�ڕK�W'ާ��?�����^��	� X�釞-�@�htW��i������Sz����7&��6���ZgsZ������n=��^����؁����(P;	�����9=�s�6�m������PoZ9cԳ~�����^�m� �k��yQ��d�Le���Bqt����4'?�b�L
��d%*i�7��7��7o�du�Ϋ[k�����&��^��iu[�ɝ�v�̸�D�!7�"��3���,�n&�-Xn�D�X�T� �)׏���]rc!���B���}" *"�xq�X�?e��*̀��=�� ��,3��#��>�x<�k�e�o�:sP��y-c��0�&���.#$�~B�W�z1;��6B�l\aV��R��Q��|.��]$�2si[$;+�	z�s�_1��j3/�!=�Y=��0�ΒAy^	����Ú�Mk��b8#���vV��$�R/�G.��zXr��d�-CE�gaN��Os�h�*�'k��i�a(�W�����Y�A���z�L��>𣲐�����Fx SuZ���+x"VDѮG�U~�G��O6������c���s&uu��gG�CpsX��Hw�f�+��zvs,o; �R�DO6k gj�`�dr�a��q���\p��V]�^y#��~��,hᗧ�OߓNʞ{M�H�c���:�Lpw�5���f���i�d�I5�o+���"���K��l@�qL@T;�t`?�Ky=wN|�'�s)3&v�� @)_��S���fzB�liUtKvH�<UAxV;�DE�qXj��&,�� �,Xt���&�8��O9���Ch�FŹ�;�«�0i�7��A��ڪW�p�nVm��L0�~I}�e+�k�9S��k0u�R�/	bF�����WR�h�7b�AR�SI,�HBOd��K��(�JH�'�b�Fm�����_�+�R:g�٩����dC�4�R (�z7�0�
>s���#����M�Q9_a�4�ܮ�/��_B6�5.r�L��o��qo�f�j��]ע`H��aN�a8���(�?�e��6�$f+!�4�ucXqEN:O��R�����o	j^�2[}z�Ć���q]é� �e������s���$cxӷ�p-)��Z����aRI0N�f~���S��V��4E�GԄ�K&} }��M}*���E���D3[;�o��ʃ��g
Eo&o���ؼ�a�p�±�(��K�a"�׼�۾�:���k�������Rʟ�1N���g�BLkY�eץ��/)��*ޜ������흮qx��,�p��f�_����^Le�a�l
���B����ܳ7UD-.��L��Pfz�)������ u�a͆���|�����Vk@?��O���End�����v*��6��zp�\��$Q�V�Q7bb�g6����=���XwJ������_�bF����Јn͑������ds�gN}��=��z٫he��\^�t��0=����uX�R�Ĳs;"�1=`o�:���/g�m	�h�����
}i�7�y?L��2V\#o͆�(��@�n�v\�	[�	ߏ��k�LpQ���w���%	/6��}�w�8{��V3_ֺNAj�c���|�i�[f0�B	�K4���������/}H����:��I �\�V�ȶ�
o��\�ե{������jt�UB��N{��4A@���3'#_�¿nr	1m��m�_��X�}W^�" �1�7X���a��>��_MeMO7՞��j�6��`�����>�Yq��qn*o.Y��{�H�Tg�ل��yG�}��b��lד��4���!���f$WGEcgy�D�SנT���$/���1MgJ�����M����S��"�e�P�'���SM����wa۔( ��w�8��L�����hǜvPT�A�j�Ò�ߠEa�/�e�ք~̢�7�ts��8gX���ԫ�����;����B�*s7���p�Reb�� �84sm�^�|�<h� ��-��v|�*�A�8�@��Y�q�D�F��J�.Z�>�eg����|_�@���[Ԃ��`�2���}�;�:��⢸O"�Q(�8*q��{���9�[A���m�y�[��q�@ݒ.����4������*�YnuO���׀� W?DR׳X�	�7/�V�������ai�I�r�~���]v ��w����&$s��:�����4ʈlHm�$o�m#���9�/���h���Z�T]W$�L�m�k/77��g�G��u��'���Aj�`�=�y�@���QU ۴�//б[��	2Um ��n��ꑊ�qr_���ZcW�˪NzE�GG�}�T��ɕ����*�����6Od>L�]�w�̄��F��fNuu>i���(hP����"�q-��ͣL�^��ek�����&>Z �=ێO�wtrJ��%����O��u⹈v�ٱ�>-�zlذ�Q�<a���=�-��6�$��_�a�S��ܽ�!�����T�{�i]���łԿ��c�*͋�
j!t
�x�J~Zw|��V����  ��AW��p��y�!�U��65�yuj͡�(ۀ���w�x��ˬG^bS�،>���14^�*�ۀ���df��M���:�����4�fԭ�ţ��v�u�dص�?�>�y>}��R%��to��#L^�[EB�L%�3�����owz�\���&��Ե@�e,'��ښ��%1bK��Q�8oz��CC�e'����!�]���ވ���/$�`�W*N�b�J�u4R-�,�����w��a�6����'3�w�{�͓�«3��9L�x�u���2I�I2���C��5$��Yu�̧�� ,���q���:٦�*�W���70P�K^L[ѧ=��m�n��^����"�����2��4��F���nꥋ�_��^���&����b%;o�^iuHc����%�!d�qz���M�C��#�{Z�y�2��$H��,��q�vI3,��*jȤ�xH�I��"\�O�����K��x*�	^����e�3�D�_Xu2,e���D��R/���7�B�v�����#�Hq|5��^Dg�]i9 v"+]*fm��o2�w�͡�u���^Š�hK����ȇ��ҡ^�\��۬�I�����	ݝ�S�oRE��^I���J�X��7�:�u���@�������:D+?�%Ƃ:�%�*�1����4=rQ	�g�j��f}B"��g�Vt�O�]!B�ƇL���E�x�UO��T��u޽��=�:URԧ&�أq����� \�����;�^?��:d��c�\K�i���u�8�ߠ�9��gm�t"�s��@g�����3��M7�b�XSF���1�	�T.f�6P��	aөY2(&K�I"S�wA��&�� �R̄��YA5f2�N��I�����\g�kQj	�=���;a�4�V����&_9Y_j���j�J#-�Q�K��\��K��a\f?�2�<jr.�>�V4�Zq�P ?Ƽ"O�9�5o�NL����u�����m��y�����Т�G�.~I��&u�����/��f��i���hE��P����"i E[����k����G�8��K>��/���b&��i��Oġuz���nG�6��e]x0,Q�*��v�a��ϑ�a�B^�A���T�\dc�yI|��;u�Ee��)�Pg|}7'�ג���P�s4<���@�y9:`G�4x�?��j�7��������㈔��>���>9G?���>S�`Z�Z-��p}i�kH%�>r��m���:�M�n��1%�@IQ3� ���ou���i}	�:��u��ф�T$J����΍ڤxT&�����ݟ�*3���('��t�'KK��$���Q�Td���zxw0�o4�}�V���5��D]�u����X��q
�ͣ���f1���e$��A�������+����q���ԛ�%�ަa���:&��/��� ԟ������+�W���ë�6�Fgr�tʂ%�����;��lV����
��M�tsv�rh]���&���F�$TpM��7"M�J��\��}�� ���[���n��W�{X|m酨7���V_�A�qV���Qf��M��9��2;�d�����}ϛW7�|�q����v�z�P��'�L�>p���!����^ ��O��!�N��0�4�>cLSgE(Hk��P���A�~Ye�fS�YIJ�Q��󸱠D����:	���1�h��m�mB�:���x�-�)���.��L�
�֖y{Š�d����f�$Ѹ��Y��<0#1�(̇o�Ph�@nuv���8���g\��#ة�Y�����d���]�~���~��Co�kˆ�|iL���J{F_o��rh�rN��I�N��;BA��<���]G�JN�L��K��(e�J�������N�`ݐ���\����p��w�{�*�.��a��tg`�q,Y�=���r�EW����R�����,�����>(�[P���-�<t��f.s���� w��9�K���`�J���Tb��3�n?�����?�̲�L�lj-Q�J�1���:�y
��R�]+��b�%j���hm��-zZ{U]*��*q�e$у�B	-X?��hȴ�[�"W�K	r9���pk۞�k��j"Ϫ��J"���H�� ����A��������ς.�4� @3:�Z�Θ��DqG���v!�ؿ�r}v�����
��������GӅ�P�D�C�e��;��a��� �ȩAj�os���!�`�%:.v���9��u���e�y3���0���@�Z6�/��n�m�SnV���q�'m�,��|���a[��Ӥ�EvP�.N��T���EX�X�:e��b,�wZ���H��&~a%2 �{@;�Ht!�gOM�\2�e��0H\ײ���+�6��hX7${�ϒJ���Jw��$�=��Фuѿ8�*T)A�7��>��jmL��<��� �����y�u Ya{rO4���m8�"��ge���dikg۵��D�@ ��h��/�lp*��*��@0{B�����ejk����{��C���%���`1�o�Ǣy0R���:��j����Q"�4ƌ�:�S �ax�8�C����i���΋%��l7�~����fy�|u�Y�k6����;�t�^���
竎��5E������/@^&>�!ް�u��J���_�f��9,�~WL�9@x������s|�xI���--�ע�>ˬ����R����t������&��lu[��;`*l�"�Uֵ�4���9[@�;)O��t0�Bdb�\�#��Sӄ��6��]4�mEF�=-�;	�{�j����%�ܙ�[��/�u�=o˘n�G�]K6T&���|jq\v	��_|��HM�
!D��\���70�1F�ޮPg���G:�� TZ��zh�:����x�{�r���XR�Pb.��_���q�,|��m�+�n2O�~�z��}d6��Ӧ�-�ѭ^�?�C�Vը�28Ìcl
�3���L}|Ƃ��z�-+S��x�%yf]��}w�Ms�|�N)p���V�3��P���� �@�{�z:�ʲ�[&�R�M��)q_�dx���@��r{>,�\��2����(��'
�"E2�����J,�:)u���"�|/�L�8�wI��]��	��SM��C
9�r�״�T��5��l0�����[|�2ͤ�;�}g�p�Y�&�L�-�8�)~e+��96�>���I��m.�R~��v���� $�%Ic�|�-�u[�0�1z�d@U�nFgl�+�>8�W�w8�U�C��]��h/P��Z�҂�z	Q�d����ԗ�L�������[@D����S��~�!���[Q9�m�-�L��"��3�#���%d��p�b�8o!S��O\�)j7�黂&�\��'�0�*�Ib�0{ښ!"�+���9uPv��j�2DW�7�M�h�2_^e7�	�#�(0�U0G2t|�iZ��=KME�|aM.�w��X	_�V��o�����d�&� �㮂{��J/1�'9�n,��C�����C���2֘�M)��i��9�IӖuܫ�� Ujll��%�;�Eњ�l����MeJ��C�W�>`F�{�g���"�b�H�K<�Lk��t"��VKpge���_
c�"�����7z�a3y�Y�*	���U�w'�<^Ne��!D�]�c��7��e
gF_�CI���:��H���@�7�Ռn!ZD�&��0�S^L�<ډB榽�,�'�4�4�͓���T�=@�V��;���%?.��+;2QW���i%���[��)�<Ŕ�J�����G�_���f���;������4����`ѰY�1ꋑaϯ�Cf�0���P����+D�=��i��:W6�w��-�`)buߋ���|�E���'2���+Z�z�.A�J9`����'s/�4J��R�?�2��{Z:#욫 �� �:Ɨɦ+�"�"I�ӽV	{�!Q<����(MX�CL{�-5�K��@��n��Ѓ��]�J	����v����y�`�[>Y/��EPRy�����_�o�1\ĕF��i�#\㭣�3��r�W��K�#�4��iu�x� ��J�R�HD�l"�2���z"�k�����EU��n��B/^m�l%��.f'P v�T�Ƣ�Y��G�51Ċ.]=����q���Q�����-?�_�Xy�GxB:�w��� �������!5r��etv�5��/���.8�������nC��(��5�&L{�̰�%W�}��A�R}~-@�k=H|�ɧ�>��r�N���M(�)�"�.���\T��a�m� ��C�#���Q㺛�v4�m���l {^9��/U2T��h��ZN��{�C����E���!�A�#U��ݤ)V)�"S�nJc�d�!��$d�����]m+�k�,?�+A�IC{�e����0�2�]h�B�9���ʢ����}<�&W3�Z��HbMG֤��D7�~ڇ���(Ӱ>pdcLRv���b�ěW���s�^0����R���g�c�7�o��cu���n��U��t�)�������+7n�$x;4~��$x���C��֢ط|��6щ�?�7�h|g�h���.���N���Zl�&`%��Z���ɮr4�J�A )I��V���J�V� W�Ԓt%�tE���&o}�E��S�9��U���5C��^u�o��Z�\������߻�p�ݏ��8�3��W�L�w�>�_��Z�6�[���&_[D�-d�͙��Y�4�������35�A�/U�
� '�Ϝ[	�_C�YZ���K}͏� �{�b򼻐��־vNrR8���9�C���Tm	Ӑd#5N�	|�Ry����h @���}�<�L��<�WV$�f�n�zu"?��̻�p-�=E2?�&s�bI$���MC��N��;��"d8^���1?�g��t��w���2����Ñ?bK5��{��ߤ�!�#�FH|��Y>��r���Օ�(9��Xɶ�^��� @,���r��a�l��&�TكL	50���%�fo�Kh�dx0p�;�'{_٣n�E�HLPl�8��a&�� &Zu�(�AL�f'6W���8�X�"`�5�����!����d�]����������Z�	)��F�#�"�i�(�/z����o��-�`[��_S���qs�E8�������#ճM�s1[ʈ2��"���F�c�g����wAòWD�qwy^P�x�@�+-�	��*M��HO z���RpO���0CL0*XW��Mp����W��Θ�es�yI��[(z�q�GyW�x��5�o�M��OQ�s%WP�pS���R�_�YSb�,}�G�4I\��Ͽ���O7&"�q��6��R���g����c=v�B�R�a�u�R��"�9D�+۸T��C�ѽr3hGe���Ͽ}�4F�f� �cuZt�2I���Q�о���A�ol��A��-�k�Ě��Z�O�7]���,A���f�}�F�����;cTj�� y�&I)�D����<��i[�4�nXb��,j:��YS����:�Y<Y/q��| ����E�!I�twP���Q��k2���5�+(�G�au�ӈ��P���
����*�Tz��(�۟F6Tp��S�.�Ӣp�F�ۙ��*4}���|qTl&�*�b)����P��5����ݳ��g�d�.�]T���9��69e[Y�|q�+`6��\F)���}+�\�����,�qJ�ឫ�C8�Jg�h��Ʃ;�tS��+[����r�{6˺Ǆ����щ��&Pހ��[OAk(�jg�Ɵ�����ؾ��ٿ�F��ּ�W�\�r2��Bb�	�cS8Hb���o��
��1���֒�*{� ��������g����;B�|Ը�	�l�=t�U����I�)��{Hl������`�����(��G�Zn�]�%d��������h�pSN�S�,/�m��M�"�Qܘ��3g��� �v@�����W�)�تn��v��_-�
�:��U�z�GZ�L�5�,�Hq�$]�!����q�.��:Y��c�ZN>�fiw�l+~w|aD��+��X���9�ZOu+������g.�&����B���'����h�3���&$�~fvi\r�(�����8;�=Ǧ��H�JD�r���2lp����
�	��v����P�}
^�$%V�8p�J�Kª�.�.ض�?���F�1X�\��I����qh��.�2J���p�s�G#얘x]R^�>4� ��� A�� ���Ry,0�p|j�B"���-�yI^HѨ�ҟ��k���j�J�������`���Jk��g$H��L�Í)4�Fw)1�U�3���^'���-偓�?
��)�1$�p��w����2fL2�����Ȅ������BN�=�׌M5b�Ϭ�=H�^�,�8I7Y6`ct�~5�j��@\k7�=��(�c��ɩ���Ʒ a��pR�m����Z�8��2����h���0��f8+otT�G@�j�&�,�Cщ�(�G��,��6�f�V<Q�����+c��pHļ�]�ʮ�X�~��708�M�-�W�<��U�����c�^���X��:�(��� ��1Ռ-J���mtb��敼t��rOv�*
��S�`�mV��K(�D�����V���bn���R���1cw$Ұ�/&�G�n�^ �[s5�_x��$]�/���s���<e`I�P-��)����#�m,|xؑػI�����j㸗Sl�u�\�
BK${�.��R�P��S�|{�m�EZz=-O���	�!-�q��W& ��#�oL��c&��G_.L��2��ɠ�)?0u]s�֜��dYe���ۖ/�+�^q?;˽���Ѻ���hsŇ,��;.BϠէ���T�VΪ����|�P���2��	ft�'s�\�4FO�ut�0�R�]^^�P��*R0I�v�a�8N�J���j��Md�Ls!���>���J�>�w.m`��-��"�If7�x������+�5m���wq��,����a�����v<y�W�)t�`��+T�1$#WR^����5z�9��g[0�ӟ�.i�`��H�=BP�5�1.
�Q�q#��Kr��(������uB"ƪ��_���=�<t��
�s=���Pϵ����_ܟ��Y(�yD��sm�����O�5�
q1!� ��K_W��&�,�-��"�jOA ^�t�X�#J��X3��* ��8��\���:ndq�:.R�Q�RY0��x��xQ%XO�e��7ǯM�B%Q�֚F1���8Rqy����l[wnP:ЦAzT�v�>..����@��G.�㑬'�"Ekx����tl�A�`�ؘ?���@_��{U�JTj�'	t!�tYT�8�O 0[V��j{����?�U�-�T�wĖ1�ƀ��kq6�$���~i�Z�g��C�Q�$��KyA�b�����M�+E�@�4D`짡�{G��`�O{3��ZU���a�����?y��2+�<!�`�:���'ä�&��3���I�u*�Ka>�YM��T��)<�!2��!���xe��Z�_�K�m���/���j��1�wQ%�� z+�+�&:�r���S�ix�O�㳾�����3���K*��Dg�sqOI�� �Ѷ��Y�Ŧ�LN5#iLi�Py7Ĉ��1$^�P��J!�z��{m��gź��HX��r�H��W/��#�<�S�V��;�A$��l@7��|% ^Cn/��Ď( W��W��Y7}��4�v�e�Zv�N�:��АT��Nf����P�� 5ڵB�E��9:n �����r�|�Е�q@w.ʒ�-w^�a�//�fC�-�� �weu��ӥKvc�mM�	�oҕ�+�6ёГx��arS5�f��vpW!(_�7�f�n؍�n��n���	����,w�OB|����Ǹ�9�L�Suq�Z�'�d��A5��/}Ӌ:\h�羣HI�q�8��,�l���%��F9R�IR�;�� ���х/+*!�����u��Z!l5|G���jU��!��*���r��Z~	x �KK�d�Z��h�fУGa5J��G��̭B�T#C8%Ru�=���ì2:V*�f�� ��kN��gC��n�����:��S�%v�]Ӝv��l%�u�r��h��KE?�P='pFR�T}��~Jgf*ƍH�˙���0A� R�ײ)!v��q�Ͳ�/�^9��>�����F�K��(%"Z�(��S��o��=���f�N���]^	��r�J���k���E��O�Τ�����3#F�,&���w�`�P}��"0��LS%F�,>'8�MC�_r��n�Xp̻�I�.��d��vTi��;��/>�*�X��EX�-k���W��2�.Ut�Vp�N���^�1�a �i�D�ri!�#cg??�����x*��=��'�[7֯I����#�J��Xo�i��q���*=�-�3-��WrXL�`�wBPc�ؗ�j��G>�W��Iv��V���:G�ҥ짣h���ٻZ)玪�p̶��8+[�m���_�橠�Ơh��S���}�>b��T�ZqcB��1-7
M�g��T��i� `�nJ�9��[v ��� }��M�Q�]%�7�� ����A�S���.�c��*��p�1�j
y���L��>-v��=m/�E����ʰ�\�BLr�U�&V(�N
>j_v�5�̜x��|�FC搗_,{�ھ*D�A���w�4�Y���/�������<ۯ`E 0�]H�7���}aֺ�@�Zq�R+ ��;m*�~e�\��{|���I�FN!�	�x��ny�I�����%V;׎����{,�/��=�G�k ۨp;P�|6G.4j�F
0c2�^zɕj��$x�����9��	�;�-��ֽ�JN���?�e��yڡ�W��	�T��9�3��}�&U[��/q��(5����1���F?�lއDA�|	;m_2?��i�!�=��D����#��{�f�[�7C��z�ך�v�h����T)2̿�vG����	�_��ck<]򻵒����N���Zǻ���d%��k�b��� 7�m�Q~�	n朵[�[�ɏѳe"�r�V
���wJ����0h֞"99d ̜��ҝ�7�"���r�f�+�.*#�r:���G�n�)G�rV3s+HB�/`Ç�n)�Έ$�K�|�)n�!c�"ub�V������M�I���~�t��nN��)��s2�Q�d���wM3�V i+uo��ȷ��a��/�?�$���6
[��Uo���}���u5δe'}��ܝ`F�o|]SR\��9�F��`�,x	dn�ۻ�����ٷ�yD0XU	¯K2�i0Sk+� "��[*e�H7f9]�E�1�rX�p���������k�����G�W��0X5u� K��(�Z8�o}�	�'z���3���������� ���M#�9TU6{S7'D1��m�׀�_a�H����ʞi24�ڀB�u��2�@�g��.�?9�H�&|��4��:g}t򯨂�k�!śK����Gq�!6F��.���-ג����p��Q�t�7�����Y�Ȣ��N�c����2�e-='��cP�ca�;�,�]����Q~�IFU6���V5.�O�t4����梴Fu��a���P���kp��g�/�����#��c#q�:��H�V�r�xɝ�0ģ����>�¿��� 7,�XG���_< �������c�}	�'��c+�O��f5��a�@N줻��#W�(���A��� ��ҋY�G�T]1rf��$TO^q�*��E����K��	�� �>�t��6'J��Z���W�Ìm�ǿ�35��G_�8Z�q�����oP�(�b�OnG�^�;�Q�N,��R��2gZ�D[Chd��I^<2a�&�x� ������fŖe�]F<�f��-�:��\��T�
�Y$}��ݽ�O	�TS&���n�"��x� �S� �=w;'���h�R�$sJ	���0x�M;2_�C�.LQ�ԃ��7��'J�=�-�~ kd?���fl艶�?8��<��~;E�@.=��2+Ag�iXI��f���Dn.)���x��C�����j��k��q8��=�{�}�`�ªm�|�#�򍳫�����K�*d�dZ�ZJˁ��3�C!
*�.vx`&l�q���&?�C�KG3L��bX��X��e�2;����S�2�Ah�.��s�Q���M��^)3(��Kn�����t�Q�I�F�|c?��Տ˼ \��W���$>)M߫�O�j��	Pj��u0]$�ۑH~h9��g��m75t�7Z��4��&{�6�6�)Z�[��	��V�?�wy]�¶xY�j����W-���f
�f4ܞ�dwH��@��*�ފXI̻�ߕ�i����9��_�G�ػ\"&�Y�a���+|S�m�P�xd����p͑� ���,�1�|��ABHU��o^�͙l���]��v'�{��́V g�Be�n��,��H
Ew�yX��q�r8�����R�O�hõ��5J�'n�C�!RJ7��X-]v��)��?X5;=��^ʟ��Xa�9�j�Ve�\�y�)��L������X!C���˅`ZJyˆ!��x=�+;�罝O \Y��w;/�Ϥ�<���mpsTP`�g^�S��H�}Ӵ�[s:�|�.���^��gl"tjF�]v�kA����pډ*ð�$�'��V_4χ�6��ځT�.��Q6Jr�>�� h�ɄO��s�:��O�9�r�ػZ{]e'�m>����.��F���|�f:a�dg�f��~cN�Q0�O�Z����X��JL��,� ���Y�.���8�ťM����ŷ}��*���XI��5�2s��^�;B2G���*12�k���C��^����������AڞwFw����>�ڗs�����m5�59*�@Gm&r�f����}���0),����=�f3�k��bŃ�r�ZP�y���V���ǣԚS8���
��b��^E BU� ��(h�#i����G��pDw.��#4+����1�1nr�J/���;��lv-ȫ���b]ň���2����`�讹�\B^�( #����O���cD�7�n�n�=.4�Q�g���{$�S��b�)�:I�����s���F`19����YcȀM�����q5N��ZNV0�K��gd��ff׏�LY	����F��e~E�@��'K��#�ϡ�`���30�HN
I�ג��qw��U.>j0W��Soj��.c�	�`�G_���(�w`�D��̊Dy�Q��i��c�fy����n3��<7��$��d��]�HI����$�LM{�U�y�ac�׏N�u(2��m��A_�`o&A�wOΏ�Hr���1)Z���>�&��">F{����諛����%9L��<��廚�CN\	�**�#=�N�䴼���Ym����n�\" ���L��y�,&	^3�o�����������~[K�������~�eO�r���4�1L�i!RޗGh��+C�;bAt����$}�͢���͏��,��Y�|�sC��;�3��~E1����?��5Q�Tն<��7P�1��X(�\6�Y�EǶ��L0�$&i!t Xtpކa��ܻ�<0]KD����W�����?&\���|�ٕ�|s� ���85X��"�qa�4�ƻ��V�TjK�8
vF��$���Ħ$��l�@��P�i���$-�G{����0{Β�.�N�F�oB��0s*:��/)Q�Q��bL������Z��q��q�:��b�4d�1���j�B���W���5+�4�p&c BS#z���T��9�0C����Ca)[�h$^"\c��%t���)��31�$��������h'�����"'~�੠$���i�%<�%|)�7�b �-J����Z����u�t�gl�+��M�abD>H��"�a�I�Ϊ�L���*��3�pUnox���U[*�j�&�/F�N�ܡ��K��k�zA�v>������
��Y���'1,�)�(����af�^;ޮ�?����B�U�ض��w��*F�l<#��!;j
�ߢw.d�����O6
�R��q#�	Y�/�x:�� �6vF�g���D�D1b�TN�6�{ܔ~���$�T�XG��),��5 ꍶ=�đP.�O@p���C��#�(Ug�^N����:x4b�^���A\Y�/cӗ����:u8ےw�u+���t�_�3#8�RGT��ЄmR������s7�v�-�oț3a��i3�?���G(D��b�
�ޜ<��'x6���c|g1w@$d��5���y�f��0��ř:�Ls�(�,;Y��>,��4= �Z�3,ޏ�_jI25)��]��ä2��d�"��8l��g�?"c�܈y���ҥ��x���
�J��T�̕V�#�-0P_��*IN2����+�y����蜷��1�j�w:��L
�J�!RV�4%�J�Y�c!���	쌕	?4��?E��3'݄�B|���GhM᪋�Um�t�"C�U�p�X��a?�]��٫3F�C�����3	 qǉ����(�c�����AkDM۝R�4����YD�3cWhm� � �
́�P/W�L"��P3��8�2�P�l�M��6��pz�)�]��b���y�x�8�����H���u�9��@�2x�x��)_��	���7ɶJ��H�}���������F]�n�x�m8i[�K�^��l[����tL�-����ڨ嶆��9�2����jf�.���\t����� Lsz�#���������B��m�ƄmU�!�e9��� Mp�#GMO�.w-��xȢ��@��� k\zL������ A�S�f�fP���@�韲KN�Yk��~Px�_ǎy�����ϊ)A���@��2��4.��bc�C�M�UJ���Ee����XH�E�䨕.�~zn+��m^�-�G��4���u����3D�&��3�[YM��`��z��r�J0�XC�.-�Xc�^��6�.Pq Ke�+ʈYJ�`%Y�ڸ��ڥ�;l�Q�!}x4������ɦ��ɚ�U��e�fM�x$	�/y8��pw�����5� .&���@�����!(��V��d�i�o.���d+���){^��|�YM���g�� l��J��!Q��8(XM^䚊=i&���y�26A�˅�H?�����ssN;[GOk�/gk������ͬ�x�H��TG6Ӌn���/4��f��:�FV>��-�^��a�p��(�W��5���~;(�Me�dVY��ಠ׃�#����.h�y�q5'��9�$�_�t����D� h]���ح-���T��vp���<+�dcJDL�q�|+�t���kN68Fg�j� ��(�igQ�Q~'<���� c��(LY
������!_&
xV�_�dW�Ik���'�TK�'���/��{1������_�sX����q�ջ��FnL`VDr_�6�^7ib�7}:�Y+dp-J������� �[�3���4�����1��?��]I��u+�>����H]*ts��Q���@�0�Y5@NMOq��Ӽ�u�[G���a ��v�W<�y1��<��|X3�\1���Ҋ�YvOVY���J�$R[�����ŭ�d<�S�o�/F[������K���.�] ��4����"�[�FD�/G�L���R�I�d�J5ў��'9g_>63C3Ω���6w���?���V|�"�=�i��
|����[�Xb�Vγ&��B��tY0��<ȧc0�L�xh�+N�w�R�&d0�s��ѭ�Ö �(S��9:-¾Fu���<�j�ѷ��fY�Gö�w9M������)cIz�ƿgc�f�L[�>��G�"�����A� ��6v=\���IA����z��	�߭���+�����U!�H���dԦ��~�h�^A���ޅ�^����+��7�K��-EHG�+jm�0�)����7���8Qo9��5Z����1��Kq;3*7xF��u\�LT�""�$q֪ի;�&̌2,5����߂?>�1���{H�kk5w���|
"W*�LB\N�$/M�xF&�eK���#��v��61�yaF!�rH6���Z�ms�J)����.��6TA��X?`=B������|��^K��k�ߴ��/=E����O��.'�.�N����A`_��������^�4��B���ķFvx� 2͋�W�p8�9�<�n�4��Di�X�Д��0瀔P}멀i4uC��]�4�2��?M��W�F����Y�����]����f�O�(�pe�����b$���Y&"@y�m�����7dڥeo&w9��/��=�M����Pn@�-��ւ�v�y
�He �'�t(����2D����IȜ19tq����5G���;���2���ؿ߰�i�5�}J"�bD�-�k�8�_"����a����e�QD�HX�����̠Y~�ù��q+���2;���2{S0Cw�i?7ϧމ&/�a��Q��hL��I>$(���_��6-#<t���+�\�|w��2�i�7I�g�Cǫ㰹+^��)�fx8��PK_�_n<�.9�ޅĮ��TΛ�J�)O\���m7��L�h�/'O�i��Y�D4��.ZC��?��!��5��\t%�I���!k�/	U DE����G����~����w;`�Wcףx4�EaXb"h<h��D�ѫ�T�PH�x��m��Q	�cԽyU�1p��Ʒ�5wg�9SY���%q���)�y��nLƁ��'���	Q��H^��&�J'Ē)rv�56�����br8���6�1g2�Lw���N^�C�:���F7�"!7���5E��F�[�]�<��ά��:O�l^q����N$SQ0;�u_�B��I�3)��X�dݼ78c�v��:�h]uXzx��������`tg4n�g�O[�T����+�/�u���~ ��{�@�/^��Jb������N�l� erK#�*�h�0�e�lN2���*�1�WN��+!-׻3:�K���Z��]��m�t��6۾Շ�B�g�P""J��� Y�t�_�\��M��o�m�{��(�s�ʬ�E��
���R��9��wwiF[�`븐\�����	�Dxs��+������0�R]'��\� G�(}$P�u˿@�_<xp.���W��뷗�f�U�c\�}���V�N�.<5F��\��8Xp��i[�]���<�c��BC�=��jl�tQ� GA-/��e��~^۬���X�5���oٴ&`j�y]��"�9��I>w�������X.+�d��3
V�I��}}�T,+$��^��#j�丌�)LB�!�֬�z26�ڭou�0�f-vE����
�T�]I�x]�y���uk���;��u3�ی�����]�_��<�9��֖q'�	����Q�ҵ8ġ���E�{���ܫ���<�y��1KffV��uVC���v��
�o���%5 5Aq�#e�c�8��`��v!�D^$�H/}<��2# ����
�9 9�!E��+�k
���5y�6g��p����NU�L�Q�#Ms���:hJ��UR�2�2�l#��х _���J�� �v��m�(�Ǐ
T���j>ujk���������he|�y�Q'&.�~�ӈ�+p�b�:!=�!M-�V��bI����F�u�����Ñ��EhM�kV����/����w%���=�"�UP��w+���+o����lЏR�{�q���l�I�l� ��~:�:��MI�g%kg�����'�7j��V�L�8J�&FA5��� \ۋ����:��n���T��a�ui������ㆺ������~�r�J�7y�_J�3�D'��XǸ�����so�w_3H�&GJ��|A��d �sX�|��""��zAd�z싻�?�g�H�&�bv��H v�R�Z=IȟbQ�r�+�}��k�n��(1
ʼ���!����w�~�K��$V�ʝz	��^�U��ђ��Z�,�
�S^Ê�w�Imu�g`��;}2�s艪�ҥ�DMC��'7�,��󙐢 �Z���=ׯ�]@����`y��>yU'%7`qੑ���蓼�Y��k:5�i�<78Ĕ!�B%�/.�g;�yf�z`��2�|#����c�&��pO�U:~S�~��.L'���?Z�{��{tp�~UC>ԟS�`���gM)p#��P[&U>P#�ˑ':S�^�(j�(�脁���"�wm��@�!�K2�h�c���_�%t���Vl&.�q�+/�[��ܞ��QRo�q��*��1��%&N� �ǘ�ZT9�h��i,���8Q��}w�9va��s��v6�p�@nڕ\��I�b����n��Z�]���E5�{(�m�����Oi�)��wP�g'�b�Û+�k�\��W���1�#vgi}��.�{R�X�[j:�QoZim/[Y���&ŉE��e
������ihE5u��Y0���(��ćO��qW��+U��0�� �L��V�s3
����%y�����f,��}n�{7�|���p8�P�3��X�_d��K���O�1�c����IDZ'.O����@d��<���+Ww�Ig�6����a��yᵰ*�#�Tƚ� u[3�'+��Co��Nk��W���]��r��F\;C-��&X ogJ/ټ��H�	@�Mʾ�_}����������?���&g�.�q�"��_^O���������~޹��Ձ����۵�!3���M�A�������$��}t�i �*�_�R�E�U�¯��%'���'}C�Y�E�,��� c��7�97���(0k~,9D�#�x�0�7i��P�]��	�U���j��.�ĨB���*?��+���=�s�	_��^�;|���c�Ma+��<��~ci��L�*>N�}6�5���A��#1�Bv�Ĩ_MAK�r9��ڻ�'3�;��ʓ�K<� �tf�]�~<���ws��UY��x'��>��*3��Y�P]����K��U�Z��t� "�Ws�Հ RO��V�lt&6�řXm��Ʒg�\o}��ҧ�h����:bQd��R�4�~��/C�I�F\FD �UZf���j��<j��SR��'KK�x��M�(�E�=�j�doOyRU=7_�}�BG�0�Żs_�#nvE(�&�����X���4��xx�{����ja}�#������V�ik	?���������� Ҋ�bg�Xy�D���i��s�$;T���Dn��G��%Ѻ���m�v����"Id)� �(�r���LlF��O�xK
�l����u�b0�.z�� ��uTб�:��
����;(�vX���w7��=ef"P5���X��+-t� �˵dA/*]�:���S���z�\��
�>.o��YڍgJ%��)�YR��h�-w�؄9�R��E�hD^%*�;����M�=5�&e�ݑ����o�g�p(��*�����Q=��fy���E�Nh�G,�����[��Wɳ'
��>Cו�.�7P!Yxw��J�����n׆/J���˭v��		�Ry`�`۫󗒐eqv�z*�68���.?�&�ʁ\w�����m�n4o�<�Nyl �g�q���S@��'��l^�/2hrTD�uJ#;_y%J�\�(u�ܭ_r7�PZz��71M�j#���q��J��w�=}eK!Ƶ�ƲUݦ\�O\.�y�J4��A�5�����g�����W�Ƨ<˗m5�f��<���B#7c��*5��C B�̪����y�:J�K�<����o	���:�a��B^}t�J��z���ko��$�i/�
��'�n��Q�-Ϝeׅ�C�l��/�:�@�	������JT�
��D<l����(F��4���*(��7[&��`G�["���J�g� �t���x�ŧ�L;��;"�{�,��}�-W�hH�N%;ܪ�M��5K��`D�~���3��O��աK��
C�8.鱄����a��>b[���2�b��#�P�,P�$\�XV��U�|�� ��R�Q��S���������2m�6ҕ��@�t�a���@�����)o��,�f��Ƕk�&���ʁ΃� W��co���F�A�ES��)���y��s�_�l��?����_e�|>�.N| FL
F���D�u���� ���&^�^��_,S�j�`��O�=�$�Z�4����>�m��o�f�����N��:��us��)�c�t6ro�Ī�����^�;�`�:vf�+98|�����x.ț��){�=�0�	���R�ۏ'�����<q�\n��@H@�ؓ��k�:��&��x�v���uf�!�協,�fI"?��H��M���C��-��6dt�c���Q6PF�W]�����8y�ݦ�,���4h�� )�7[	�;�����b|���q�>Fa({�u>�A=51��%��O[(�<^�0D3`�ͩY�����/YQ��H�����&S WL�*��1f��U�!^�+�:�@Wn͝���1��Q�~b���߇�EYv0?F����j{�!�<�J��j�.1�n�]��Rn_�*yY��I�V���ZU2I�y�1W��C�H|��DS����;|N_d5��_���_����_����"D��ۓ��J�	j?���{��V��p�/�"´���D���Ɛi4�&�_���e�قԃq��"֕Y[�%m=�e}��!E�������j������p�o�<#���{�i�Ǹ�ݢjU��&��\֮�f�J��u�ch���ⷯҝE���Pk�[� **\�]%�8c���/�I���22~I(��F�CZg`1�^5���%|*�AА�#�̦x�N�����s~�
���N���k.��͝���,İ�C�Kí�z��Ά%���I��,�G�uС�(ͷ�r��.�O�(�(��x���盶{%�~��؍�szj|� �$/�2'�(k�vgn�knͧJ��۬��5)�����G�g�������Ъ��Ǿ�*�H>Ǹ�mZ8��!.��=<��"
�(_�Vw��ػ�s�����>�+q:���{�M�9%�X2���g}?J�D��C٥p�F�b���$!�3������Էq>�;K��v�`8ޓB|���lxTVX�Nf�o����{ZF$��Y�K�.�2o��^�f͎&@A� �*�- �f�K��p7��ڦ=`�����L�c�%��I�¹46��sG�՛ӎ��x�@�;|9?e��������7�Xe�կ����0�����$x��iDÊ���%�D�X�(�.ԕ�uEʑ�����ޞ��A���l�.�S�F���.���NB]�P8_D���E]�D���������GKJ�����\�k�:���a���~���u>�W�JA���'����R�>�SM�� 	��~��F\b֎�$h@�K�n�:�`yr""�)�cJEC5��<�|e�ϋ��0������}�ePH3Q�s�J~SQE������Ρ'�:��|���<����+C1I��q[:���ϗE,o�(��v�;m��yH���+�� �lM�qEj�
ǎ8��{&��N�5��Ьt��h.���Z}��}���}�J�q��wm}�3$����g�~w5���f��H�������L���{�g���_S��84�^'?�1+���j��N���ߞ�S�T����C�sU��i1ժ���
=��`Eo*�b�nd�ؓ�|���?i��A��8,�|�}ޝ�a	�б�kU���I6��3=]"������yZ*�G�3������a�b�=k�=��{�����1��������a4r�-F��n��i�L1F�ECA6i�6TS@��|8q�R܇15�E�Tяo��Đ���|]G&x&n�v�i��]��N�Um���xR���*�Ws���=��g�&�W�ܐ=N��^�;��y�ч=�i��J��4�g�3� �9o�Z�� 4r��{���
n���N��IN�H��t!݀��*5u3��d�7M��~l�I����e0^S=ݭ�M*�CO��8ۅ����?��\NƊٕ�L��j*�����*R�!K�zL��k.
�剞���b���}�-��~�2֞���/2*�.�7�-��=sd茵KlZ�Mcy�t��k�ox��m�����,�S&�7gҨN^B`�13s�L��T³ �D�!��d��ɘ,ɕ�$�|�vT؂�YO�ϭ")��B3�'±�X��O�֩]G������Wdci�G�aLo��(��b�̨5S7�"�rw$�� ��8ϭ��@^�*���.r״"��.:�S7C�:WEw`#M���&g��X�ʟWY#��FӺ��-�رn�.2�#^:��`�R�5$�&VWd��Q�}$x��+w��V�|?�����4�w?�����z`����i�C���LA�$��ǯh�p}��x���U�Y�-�lʷ�!2�%�@����Z��Bf�T�ةl4�d�����O�d���%�v�0W����^��eCr����tآ&bw����ޛcm&������5�������J���.�\hcE���LS+ZKbh ��]$[3�.y��D�$� ��j����]�Ea섽Ɵv�e���Q]^G�ZN9����i����G�9��d`�i1�h�}9� >*G�C����|�0��{����$�;.'Q�������~��c�l|B�v�Vο"��6楇Ỏ��B�AvI�͓M_�,'��L/����!�J�KfZ���#]������F��H�J:���$����ZJH/r�ǌi琭��:��f��8��QR^*F{oHOl��M˾�h��tEF�*�i�ju+�Y�CA�>�L��2nv��J��I����ŉ��B#tv5������:�R�7����Q�[���J�����Od��$�s"(����0��*@!�fT�8����q�\>G��� R��9h3ж:��+J�F��� ��,;�5l��N���V-�����5�g���7^�#�k�����E���@��f54E_(�xю5n�1N�&��/]�׎[�,�<��<�"�v�Y\q��:���/�BCgN���ȩ�Sp����7�F�ݖe�hp��n�W�^��d"Q{�����[;�T(`0�gd��1�L��5�D�Ľ�������=839bT���B�t�ِj������6c�������-�a�i{��r�BF۝�!?(�4������b8jB�$(�3Z+�w⡈\���pD�|Y�=�(Jy�Հg�+1�L� �a$��(6C��M-	t���+]ؼ_��ws��v���EB�{x�ч8�(�1��yq�w�X�/�c�� 6	�Mo
��IC=�MMA�/�jG[F���.�_�R�R��]RHE�3�5Sѯ�6q�*zsT����G�I�k��ϡD��+1ڠު��AO�����~Yح����|���3"K/eM�J���N:K�	F(|�i���5p���GĮ1��d�8�=(�w)�+	za`7e���'�q���0Z�F�r����"j�)r�#� �Cq\8Ux�}��i�aW7�`CMZg�+9�^v�aF�6\ᶨ~�F��Mjx�S�Tb���n�rP�5�B�م�z�+�^7�YPy��C���ɯfJ�rP�Np���r6&>����m�qm�@��\*Mp�F��|���/D�Y�+�ߛ�&Fm��ْ���w�)�T=۔�#4_9^]D�,j.��+�>���$��JC��n���@��K)�_�	��������t8���|m��.��rk�q�/���F��<�v�R
t���������Q�]���WǛ�9\G��-�8#�.�[GG�?	��P�ϼ�e��g���|F7=S6�$���$��Ռ����S	��{�ҩ�zA�U�>'o�ڻ��G�P7�����I"�6�ޥ�x�٭0�cꚥ�D���ȝ�r^��EV����fg�����Ax�b�/>���؅	[�E=6ť��[q�ٌ���4ke��!��2�-$�f�fy�Q����zn)u���u�yXۀ�d�/�Q�ɒ�v�P/_#Ս�;�̐�j�D�2���Q̵~�^��o{y\p���7؆�
.S}Z�{k����S�S�φ4�Wa�68<����ɕ�Ը���VfB�Ӫ�mJ'����㙄���G����/�\��N��͟��(�'!~T>�����Ӯ?u�X������]>�fO��

*�.*[�芯ʙh�Ǽ�>���LdV�:� �t��g� �8�]>T�o/G�l��@���`@E�$�B��N�zl<h��÷N8z��/�z�q0ܩ8��/��9/T�J�������-F+�J3Ϻ�SR�lp�T�myScX,G�L�=���LR�֏��vF��F?�ޘ6�%����UhgRe�[Q�/�`Up�1^�L�:>]?���6{z���.�0�X��[�����r��{����LA��C�m�]*�9���χ�y5�^i�Dl�p���a�v�.�ʹ�>��z]�ٴЦ�|'@'JlhP��ˆB(���\Wӣdp��bڌ��7D�٪>���I���dY$��1#a�"�	�"4f'�P��J�)�fO�X@�d����J~i��:��8�.�B�'��qS7(�&����CP�ⲷB屺�>�јhA҃G(����.�Oq����kw?�s�	4!/Y�!��t�z$��_R*��u�~co���x�� ���ֹ�+7o�"�'|�h��7Kg�{cm+بאwM��M�w��32+�F;Se@!|)-��m�~ޖ����&2d�	#a���D�B�?�>�l_�����M�BW��K}ĥ��%]�9�#0W�'<��h��~��L��$ř�%��h[@�#��Ū���g�'�5"pʰ�Xto��co]3:�P㭼�J��)?� bM5Z���D9���F8�q	a�U�!?���t�2�V�(׊Xl�m:`�R]8�����s���ߊeA,m����헲�!�7^l��Z?��B�0Zu!�B[(
\>) �o0$��[��'p�qHxE�6"�_H(=A�9�����7>5��]:�ttU`O���)�أ�/��ǂ��DI	��)+��%��d�R9l^��[(R�S�˥>�h����g��,����4fBK+g�9gw�%���h���@��B���/¿�X�S�Y�����{b3ե&��u�A_�a��[8��e���,s@��k�z�}Dt,Lb2��x�C�v�{v=��L#�JK���>z��$���ȋ�Eً X���۴QQn/N�׺�9m�A}�g"j�I�bv�80�/�-���_	��if:���YC��'(����Ip�!/�ܦKW�֡��S����x#̅������o4�t��rݿӛf��wT���t��Q����3���F�AɹL�5��=�����%�K8�WuJJ|����v��ϰM��_�?���I�Ac�[/_URfU���.�Zp�?��H�F}�E�RB��<�]0)����&%fo7�7pN���V��� Y�w;��}��� ǁ ��kHAԋ�����(�H�%63���~^���ҷ/�G��F��E�la�1��\�π��䵉8��X@�' S��/֜[��=�CpD����9i��R)�۳��N�/��t�'��2���5���|}�����U��g�p(��+�jv�WOL�&�w��Rk����Y3���\b5{nP����:�J�mjk2ɡ@�5����}�T�W�[-�ʲ7ǖ��rb�\�g��2=[5W�n��!W���|)�l'�[�>2������b�7����'��UॲR�+��:�м�1(Q\Z�����K=�AR�=F���;³yֻT���e�v��R�)Cj�\�Ï�a�;T_~�VNz��oi�l*)���j���D����¶��, rP`��!M���:�i|��b�D%1�=�37���5.�٤��X�-�q��-��|+�����Q�E�a��p-@��� ���吝��)����z��H�Fn|e��+k�����/_�x� �Y&|�C���Za\� ��Z񋚛�}�9��hg?F� �� ���قLJ��%�t�Xr7=��$U<"!Ч5 �I����6��V�8ǕA;d�(t&�IA�:�J�����%c# ���=y�A_6���S77�{�=�2�`�\�e���r����!������C��6KUN�̀�K�������hF
�\ԫ����9k5���o9�JVQ�D���bk���E����_�R�m 4.>ֳ��9�>���A��a�B^�hň����t��2�GS�B�gj��b�o�7I�:�1�|\�Jϧ�D���s���H��q�S�V�!>d�	�+W@� ]��yx�����:�����'�I �H�����ש�<�	Y�Z�hd�m[�j��M����Q�Y^��pPL�(�i��.�!>����.��c����&��5��+(ܬ!ڶ��-��{��h}�LI�۬��&l��n��ﺕl�g�=+�cwb����?�J=_�ޯ�/���L �����hׁk^BsX�yGh��E,�NG�c_��1g#���A��|�F�1�4�AX ݇���-ϊ|���Y.y�2�7=���	C�D�c��AY�3VT��J�������{�pt����I��s�D`%�i�bHW6�t���Z^���Nn�4|����;��i��D��vNh<�f;���u�����qR"���%�.y���;�}H;B�V��=]�0N��<)�]�|����+�4��IH�/��(�Ts���t-��q�ӫ���*vn7�� ����/;c�pB��hȡ���|�ƛ���é���H7����D�������K�2��g�7�-��ע��9�C��,d�GF<�w�>Ad�b���g�d��YX��tWv�VvE�(�#5����x$�8��:ƝkWg�5��J�|C�;-ce+d4>?.m]���M[(�m���nU��3>�C���S�M�6������8����(������[��zL'�u���2�b{r��۟���3��$dM=�� �	P��I�ȫE��ۮ��z�$f�n!������s0��*�n��v@y�S�>�{
?mt)��ٗ@6V] ��9� (�W��2t��ʣO0� ���x�Tn8��k�ٲ�B�()7��d�C����q ��/g���<)ɍzt���&L F���=q^�z&��uA�Y�dOl
�&�G���AXQ�E}������m/�5<db�n���v�b�Dt����o~�ܹ�	�&�����A�_�?�mg�>2��A��x`i����~v�Zl��>SD���Fz½2ǁz|���!�Pz��;,�_�����}��i�X9�3@\��tCRpkv7��1Na��|���_��3 j������ҿ��l�&{�����k���f��N�.���{�	�G�j�X�`�dT}�&�r0#2� TS?�&;g0h��h����)� Ⱦ��P8k��Z�tJIw��:+�_�=��y�d �Hm�C�_��47,l������h���� #]{�:���E�lt��J4+�H9�v�g=�x(�Q�4�!^�N�v�vItb0���Y�qS�M~��`5�^�߻:��#Oy�K+�MNi���)�y�������嶟��v�Ld��8JVn�"����qJnI�re�<"Y���^kq��R�|����JV�S��eQ�����R��yd=}b[�:6ҡ�-�ϼ��F�����a�[F��ѩ�H=��!��ڂEZ6*"��\
���R%�4��fÜ<���������������g���R��/��7�@�°F���Z�̙���
.#aiDx�V7��sn�>�A�0[�ٯ\Y��J���'~����=��^'L���\$�H� ��^���;��gy��g����i�*Ƹ%��a��eSD�6��R�9�F/���\���?K�YQ��s��(��)D��rr���C�,�pz�7'&�S-�ރ�F�Ұ���DK�q�{�O.1�w�Xhy�3���|������>�k���Yg������+�,��òE�iۄ�����榟3UW�ķҡ�>9¿K7 ^�\rZJ�;X�ZGِ&��7���̽</=��`ߙR�-��=��m �j��(Ĩ�=b��=���;�.j g��?����6W��j����]��F5��)��G����p@��-D�a�} �����B��@L�HD�SQ�gG�pڤ�px�-А*�O��<��3�A�aT;��>�*B�T���7���m�i8m��'�*Ya�KC�c�\G%y�a��y��e����|*C!�SF�K�ҵx��#���{����"򲶖�C�Lڙ�s'��v�F�R��Y� �>�KZ�v:�#��q$�������k�snM^E��bh>=_��w��H��<m�v6� F�#�|:��0$�D��)��Z�*cIհ�zW���.��$5����n�֌E������Lw��&���?f�*�w��ԝ�}���;��t�N"�O�Tgяt������XV/+�m�,I�]?�6�>�7���X��ּ>�qGK�s2[��c�	�)�{��A(�$[k)���U�]�Q��	���*X۩=��R������K��"\���|N�eS�R�a��mG�H��6�B[�א��GO�l�{#fr��X/[(� *��"~�#'F��\Pq}`�09�֛tA���{U�Hv83�������K�k�;����Ai���0�`3�/i�A���'˷֓��H8O���:��\~������r���(y�Z��w�@�y�P�@`�yLA˅;�̹p4���Tb����BV|Ql��Z����/Y̿]�Su��j�·(r�S�8��<�ȋa���3�?�b�#Fs�*1���&�6NBUP~|!DAf����1)|����C;��14�8}4N2ԕ6::�{�<����]N(T����������*�&�|^�tŞ��	���:}\���3Xϛ�S�:e�I��5�R�1/C��2��&T[����H@X�o92����q��Tv�LL�5ҒV�[i=��wK#��J�ݒ� �}oں���:	u�P����'2"h�Ӵ��ű�� ����>�s�@���k���c��ĥ$ݎ��㚠����Z,������$��%®[�V51�+�#J׻��9�bwDT-�R����+Ao�y(�R�������5�
:���X�x%�K\�ˋ��3w�~��4�M[�!��ת������SԪ���j��#6>1�:��(v��Z>�G �y�.饈k���ۉx��ӕwG�D�WL��,�HL�Cd������V�%�~��2c��HY6��(�QPc�}?�z���L#-�g(\��t��B� �-)�'�pܢG�0+M R;~SJc2�d:j,���h�sn���ڍ���~�T��(��e����4�����T,��p�.&��=M`r��X�d�JD�g�c�SޓIZ�v0��'5_�"���d����	)R����f�-1�����ީ��Ƌ�M'cfZ�ot��VqN�*��󌔈dދ�{�:�,)�������I9�\]�P�dp� �ET�s�]�aomM�)���zc��)��3}�<��¼��#<��i
%\k�S^n�O;��	�v�8g�Yۍ����3��Y�ӝx�|�f�+Ս%V� �͸��ü큭�VU�Pѕ��# ��4��Y��CI��A�^�#}�͘;vQ���ր;A1m�B����zD�ր��rn�)�ԓۇt�~a?�׋�P����w� &���!j�xx�N�l���6�v+�y���ѯ��w͸�r�Q|���Ͽ܏:]�U�K�i�<x���i��kǨ��uTƆ�����w��hY`MIة�h�%�T#-:0Z8��-��Y��^���!رD"�z`�����DJHP^�{�2߻�F��0u���If�Y�˵��@Π	o��Bc�9���P��.P�ge�������d8Kq��ёV�W�")f_4f9Ҝk2'e�f_>g���0H"Wu�=e��i�Ɛ ������o�@
f�=qF$�j��Hv�0�;L���2W��!E=���ʍ,��a@�z'Lil��4����D�^�2�8�?+l"e��	h�0q��2$ �%��k�@o��q�mH�8W8��L��QM����E4EV�D�q���%�GQs�':&o%���G�s��+����W�#=��Ŝ��l�?	z�6΋��	"�f:E�!*d��k[BQ���Z���b������Aa�'��L��('<o5[�ܧ�s�Ƨ�|D��,W	d��iX�y�Щ3�i� �V���'���i�b�����M����+���c4x�]?1 ���G�-A�Й��XԬF�[����rXC��d��)�I���ߥ�x���#oєO}�Il����-��|Lx�E!��'7=o��e�'��_���tdn�6�]qÑ(�!���aׅR�&0���Mj�W��3g�1�`���t���a��Vy�ŵg�|��f��0ia�������#ОŃ=�C_�ѲB75 �Y�/0�}������|�qd�#3���|�(N�1�(׷�c��'*���&�Z�*����s����e���JV�sG����ӡ���oW��aD]��JȌ?\CO��`�sekS�Z��4Q3���z���çd��T��d����g����,:�� ��j P�q6�1	:#��'9�Ԏ$1�$�l5�O#��4|����f�%"t_�:pm�|9��F��7,�O\@�<����h�O	�q`��/���d�~~/��)��"912�V2�4
��s�q���0m�6���CT�����1t�'�]��.�k�G`���.7�1���Y����!$|M\;��ke�*�:��ZH)��-�b�[�:�YqZ#;3�����f�#�<%e�`�B�E{x�����6��n�����Ғ����>�� ǡ�Ꮕ�`��HY�}�!���!H��xve�|̓�#��P�E��7=4Pٹ� �^(�-�A)!x�����}�k	`���1�eg������Ǻ��i�&{p������qr��|,-�t�X�DR��N`"�<-�	��l��6\
0N���w�D����0��%cZ
w3=g������&֦	�"����	w�0�&�9?�i�g�Z;KJpx�T�a\Ǫ=3݋��["@:���oe*���3��4P��(զ�w1E�(���t�u:���|�����������,�p��#�E��D�~}`>��yNC�8"����q�S���ӥ��˵�2��(~��Ǻ��@ ��^X��LmN{Y2�Fa	���vo�k�k�|�0�QN�`�?�c����S����ʋ��g0�#(k�3Ɗ��}.��ٙ�>0�Y�ʣ<������
S�[ᴡ̓�c Q��ߗ��rf�j[j����9�w	���&8=W���uᚪ��w9Hkϒ�R�K����1�s�L&��`F)k�J��q�����7��CWv��K����6'�#�?p����G8Pc�],�VC#���B_=i<�_`����i��"�M�IVOn��\c��2�r�"��=-��S��������ً�&���~�ETJ����#���.L�k�׻��j�}Q�6�m����[2�-���g.\4Ͼ/�	��>�bVX���9� J��F��G�љ�c�
E����a6N}�ux��/yDt��v��K����b+q���\2B-qe]���E�.Ql���z��(j��I�^�u��!��F8�+�$��ӆ���w|O"��a!����%-�$�d��BVs�,�00�ˍ�kϣp�x�h
K�;�h9a�����>�3����ԧ�3h��Ѵ�HT~�e�~��U�dV�__}U�D�-��E[�����F��ԧ�E
/v�/%w���L��Əx�n_O�J8�oRԎ54�� �b�bd'��/0
g�~P��XX`l�^�>v���ghv?�u�`�^�([�X=:�IhYE�)cJ7����z'�טA�l�c��KI^�T@(�}�z���H޾�N1Ӕ� �d�V�`�l�b�O�U�ΣQ7��}h�f���p^����S4c���PI[Q�<�!��^���}�[��6+r��X���G���n(eC@�3�.�u��5�|�����)-�I�$�P�^[~��V9�o��\��rk��x�hz٬̲��$��V~}�Ts��.ϼ�l�I(��6u��4�#F�����F5�Y��X�EZ��@�<�0�lŉ��'���PsÇ
�mx	&E;{C�{i��~��t�}�+ܙ9+�xIɑ������?�XTx�le��h#��7o����?��m#ߢ*U�֣���T���Xt���n�w O
�zG��t@N�1�k#�y�(a��3-$~"$L�yZ���U���tw�K��{Y	�|w���O�A�fXGRT��k�6��`�9��$}�:Qbfۜ�\��8Lja�L?fNV��p\�O�H�VkX�g�:������i3����rJu�\,�WC���[�x��4��!��M]g�o�S��B�@�l�����z��~�
D��Ń��ϗ@4L4�DI�F� *� 2'I�\�T��/���t�#)��A��j� xMOˠV�����l�e�C*�Qc<�X!y�6�Kl�|�m���$��Nz_�SN�
ؓ|����Nf�}��$�%��iWE�+Y��DU]�-�ߐ��wV��(|�Z��"�L8�"o['�r��J��*�@BF����b�g�eey����0�w�g�EME"й��/�Dq��3�Q����J�m�k��j�/��z�.��t�#;a�^ӑSO�D��9�^�� ��:#�H(��̰[�'��64܆�A�I��͢�\l�X�ǀQ�㞄�:�e��W�zg�ɸ�j�ý��no��5�O(��9�_S0BZh����V�X��"�5��.��u�)\|;�'������gɟ6r�n���rcԜ������<Gl�94i�g,�m$b/̣��ؚ�v%7�����+�)Y���n��wV��B|�S�w�0F�O�6)�W�(ܑ[��b��Be:r/��)dX���wi��FV����2��W�
5e���?冺��9̶>W &M����go�\q"��6�x���]IY�2ˠ� �f�[L/��l�}ދU,oN����;� �,!��CfBӭx�����X��h��p��o����>JS�;�fھE56�7b�WG��a�0��P�svWل�0�nA�@`0gE���(B��GN��j�H��@�	��ip��,�!pzÆ��v�G�q�i��<}K�"��<VW Q�e@��e��Pf�!o�V��f�@?���K[tv�R
���)9{ͭ�;�� �gs��t��%��P3�>!	*��o�!��)+8A�,s��w������0�1�*>v����$�ݣ�pg��0��7_t�f��P�mV�Y\����ŗ�y(�.���o��x�?�q���G��I*M�	���Wk�����A�q��`�^'�V� Q	��<�����*��r^�p�P#�6D3�Jg3Z��l#�{#e��z�r~Mp�N��N�R�򿅋�	��~��m!��,ͅ	j!�P���}�A�T�6�\x��FaǞ�#o�/0~;豬���Nٮ!�	�Y�m4;�����	�@ҥl�Um_����/��*'�YV
Q,J��.���a�@��n��-���0B!qA��e�k��_��\�tR&�sr��óҙ��6wM���%�:�Tݜ�ğ5'�Ɩ���K���$�qx����zz������ߊ1��}���7yZ�qd�Y0_��_�TC���.$ U��3����7�7�g J�*V�]���$�[�@nޙu�X;ю;�mp_2�`��bH�|1D��!�<�s�����J���{M�H����y��	�[!u`�ػ�~>Is}���j���q�'?24yQ��n0-�$��3
Ou�:(�q���È��B��褭��vYc.V*$�2��"����>n��]���q�UN+N#�QFLpiȜ�«��Gᵻ�+ť�Ű�A^�M��ᕰ+�b' _�ϖ0Uf�Y�?�ڥNԛ�]�DZ�+���Z�|�a��i����ln��`�6����b�ߦ�/h�����w�P*�:��&\o�
����<�u7�2���>�ajlh����$c4�������O�����#����h��	�%ѝ�Ԕm^��#���gG\ߕl��"&�д�}�uN^�tyۢp���~!'�r���������oc��;��M��#�xj����KX$��Ԛ��:��T�x�\�{� "U�#p��1�y
��N3[I�e8�obބ�F�s�͋�=�)���W�x�a�u�v��T�W�V�4��SAPB���.B��}Isp0݋��n�����=�w��\�«�z�BC1s=�G3���*3b�}��R���ȱ��d�_�zߛ#N�Ab{&� ������.�19D}�x�A�]a��l����8*�W=���6'�p�tt�0�9��S"!tOu��k�9�h�گ����)(�3�ϡ�b3n���熺��ڪ.8C�f��R�;m��3s��NrgVٹ���3������Nt�$�j	��>Rż1�z�>M��0�(0�x�O=a*��ˮC�	=�*����S�Ԫ�P�׳�L�����(`Q%�T{"ߤNv2���2�,�����p_��<��
�!�r��>�~c���k���� �˝X��"�d�
�\������S9@D�V�^7��V��^~�d$]�sr~�Qƫ鎏<�o�T4�
����?^��c�0�����������7����4��� �V�5�tDK�S�F�m �
����x��������u�ՊǇ��T�^����5����o�����c���F�H�!g��|�6�`PC�}
��o
d�KZ�,���G�*z�k�n�����"%?kS��Ζ�j��0��S2ٟ��%��sc���ŹL ��8������~ ���Pd��	^t^�R�o|)h|W��.��2����2���$�>!S/.�dMp�$gGŧ��4��W����*}	hÖ��=��㖚���V�-D��/�ҿ�瓄0�]̞�%0�����M���/�e�X#wO۠�W���⇧�ڋ��5���ҋQ�z��ARL��BBP�����蕤�sk��m�)q�?^-�/��UG�BT��I����c7�d�u�}�S�7w	�Ju�
H}s嘿�ڭ���(��z�����$�PD��ʟ�R.3�������>h+q3����|m�����|��:΁f��el�{b�ɦ]xvU��ɇt��I����*h���Ξ��"�<��ȫ�f�P"!�3��(+��1�Ї��f�7�D��SA�3G@�r�0�z7?����*Iv��=��C�Z��)6q��:����^q��(��-�,(#͔1��ۣ!�n{�UP�V [�Jd9@d;��+i�/-]V��c���>+�#ƸT3��	�<G��˱���A��K/�Ki%j�i�֖y�h��i<�s�`Qq�#N�n��!���B4����f)@�c�0HnK����ʬG��kT���zJ��� �t�w��:���j�����O����:��� Q�;m��� ׫-W�� ���6�����2�}�k��5o76��~9N����~�4%E�x����f��|_9o����+�,!����fs�_��;r}�Ɠ��M�L�ɢ{�vi�Prv�3�+�FYaɢ��%��O�,{d:.�e_�X'�Q�ׇ�=O5=*o"܅ep�K�dA'A�Oz�����<�>�,�r%:7"�h�%���{��p�4�3𡣑��%�ô^~	7�8 ��S�9o�(3rC������W4�$.aۓ�.��5<�iF�
8��i¾�)�k�-��C�@����O ��#A VF�V���
�#�r�Wq�[ ��9���\헣�%�oN��x�ѯy�d�s��Xyr����P��	3Z-�ON!�+t[�4Miz�A�},B��v'�ԕt�Q0eλ�o�oШcF���E�5�:�B��"[���>;�a5���8���8�B��k+!�sj�oi����m�&r(�w+F���܍�}{t~'�+-�;�K�㱴�{�)D�`*�U؊��J�R.&E��)����q���h a=_���WZ����Y����ZtF�[�И�t>)s�lmul�vj��O/d�u���Os���d���T�5~>LE��O'��񯇧��O�ǝ��yS=7��I��!Zh���^|�y�݋ċ�s�q[<a2��8Kp%4�Wu���5�F=�C?3f���F�R�m�������nIw�]Vz�xB� �D�t޷��Pu$�{n���s���΋=rT'�ߒ�"�`[��; /n|��3h��)�PHn<���`�d���O�s��@��ܠ�B@[��̢��K(�r�am��9}�����%H��N&��\�\�[��#���Y�w��M�dhk7J�� Uru��>W^��Ac��<��Dd����)��B���;!5�ßI�+
ğ�����k�آ�l�q�L`f"��� ���n��讏6�FRi��§Q��R�*�����Y�#	��D���n�e�J�ޜQ��rNI��c�-���a�) X�7}�2&�?�9�a��/��`���h	����O�����!H�ƙ)N�W�5��H��3�����av\x�,kh/ҥ�R/#���B��n3�kF��S9���M� v�S؅M�)_��l峠��R�Mu��{�Z�ª"���I�Ϳ�{�p4����u�K�fT	<��o��sB
gW��R[γbח�z�)�8AJj�"��]G�������2�joa~H�r�:[x�y�/��K��F��c�p���Q����@SWWy50��a�qܥ<~E�w�;1*���Ty��a�>`|��nY9�d@aLi����E
��_��ĵz�#��Q1{���%J�z����`��.kDHDOic���f��mB�.���'o�a���qp(8��B��Ľl�Q�r����ۆ %�:{(e?�ˬ��;,�!�9���z�XǢiJ�(���\�7�v���K{�긽���Y@=�ڲ�@��cљ ����A�F1(^s��7;��_.�v���%ER(m1����LA�[l��3'���Mn��X� |Fn�?����G���lo5.��=�9͘ȓn���_�ɽ���V �lb�@�Ukώ<ٲ��m�o$r�J�Iq���ը~�Vnl��K=vv���$�
br�T���&��00�*����~���$y'�kڐ���o{ֺ���`�51��dk0���(���k)
�ƻ$�
^Gj͖�pg�^��b�O(K�"Ā��Dꭑ�,[�-->��~,�����Q��j�i�({]���_���饡$k��_1�QA�L@�V7���ʀj�5B���a|���J,5<J iM�K.M��ק�~MS�Շ�Bhkh��Aܵh��g�e�"�?sb�bːP��sPj�W �]�x!�w�7�:�}y����/����ps�'����o�@�7��AΆ�Nہ]���SM��4־z]�D"�,���j%% ��f?���[P�'-�1'���!�Z��al�!]w��kũ�����(�M�Q$��r�����!X���^�Z���Α�>$B�Ud�F;��2�ѣ3�E1��.+�ukg���K"���PQA�&>�#�e\�wD�lGy��X9�10窸.I!o,�W�q}��|�����>A��f���R�NZ�AT՘́V�P@�çV�Mt��.�
���^�*�0R�;�6�@�#�����E �3wl�� @�4������H���C��+�����E��T�#\�8��Ѵ+�4����k�YJ�$��f���(w!��z2&v��������˲�b�r�^�M%��A���,�G��{������z��0����WI%�Y��K8.p�J��/���f�i�@\��7c��,}� �����&UKc> x�H���f�E=��1�Uh���__nH��0./&�2� �;w�M|�!��+��Gs~fd��=���P׭�R�dN�O��Q�qx���$�ue̽���׈�9aO��zs����6M��t����C��iz)�¥�ʾ�$�4 w�"T�a���wV�!^����o8��"O|�v�hNN��#��Vr�x�3��)��8ݜ��L3
�вX�-D
^b����9HV3	��"�x��$�����D�J�7w��o��+�P�}2�2����V�-L-��ǟ&�G!��p	khV��?��������'q:�E�O���aK���e.?@�8���F�0����D"��1��hw�ˁh�wԡݬk^ ��O�x�ސ30�����7��	y�:�pʱ�.W.Ͷ��߿gPE� �Z�
�ې��~ֺ���7N���;�~.����;��3����@��߾kݶ�Rw�N/�����/�A;��`��<%Jy�^� \�n��8,�jPC��]Iuꯂ����_� �7A��8%��K��>���{>m"!c�/:�Y�/�qT\�[P��=�+�տR|�x��GI���K�:����ڛ%����7"|Hd�H�7�?���R���!Yl�'����*���������������`�悃7�OÖv�z9&/oz ���[h�!Z2��b.��G�xq��=rjT��u/�l���\�e�(��x*���=r����N@i��(3������
���m�/�b��<�N?�����M|C���e�Px��s��Q�꒖����%�PAMZ��>��iu�؄�^�±���'#nz�e����JM�A����s���*B�U ���4�ao��c'��DQ�	IU}ꍂʠ[R�)��V������x��G�)�%#��;��� ITv�~�t��@�6dD��Ls�u�����*��~���E_*�[l�O���A��r�[z�����Oc��ы^��E�3B\M`�%��"Ch�/WG�t���jS�䐸�D�uhd^[}Ao�¶z�hB��ү�D���6��D/E!��Ѻ'[O����e��p.�/���m ��0��:U�1uD��Jm.m���1������7
���-������R΢�Օw'�A,tPT��?���&�H
�O)��9����˾;=U��IeeqA�F�'�M�J�R���ս�4t���qݛw���|�oT���!�OU�N���=��,�]}��#��
��]q%bCa�P�[�L�5���"=������)�1�y���N��h�V-� ��ս�4����$?W����z����T��gmNsI)��$"�����!�~'�����ڥظ��z��
�e���MC5Q`��͏t^��4���lO�| �?��!�	�4�쵻{��
�Nj|����>?]Ы�Ķ�@�Um��qX���,�TΞ, A�By���G]��d0G`��۳G>�G`\R�q���0�F���p&�w�<�Ũ������u��B!,�F|&^��yEo-�̻�]&?Ȋ���G|��׀�'){e�O5�O9�8,���F��:��T����K\V��^���խ6��4ϭ4�ԓ����@	؛I��c'���@�f��#?uƳ���ްx�,����������{���S>cıFF��"�S"9Y%���P��s�=�@���<����n+������
?���;mC��w#������73E'Zf�HB�����������S]�s��f��0�>�J�z R(%���Q���b }��п�R�8l���>SO�.�7ځW���WT��l���˺t�7��\Cg�50]3]��f����԰R9oP��Y,�ű���2���b?YQ_����}H�4��^��k��Dx	m��5̾"5�=ߞ`�nT��g
�}r�B�~��/=�ݨ�Ԋ����L�"�"�h��S�$7��oFK�L �f?���0u}�rt�7���͘w4���ށ{�e��3�ڀ�hg�Q�*��b��6�h��½��nḶ�Z�jތ��Y�Ҥ&�����3��^p|�y��\}0�W��9�*i^PKab�~w��fP:_� ����9�����6
Y�볷g��>�|{oR���Y��֦�׊���F�ϱ�7B����?�� _2�l��dZ��`x�_���	�̔�OR🧺j�
��_��*� 7�}h� �ii$G9��R1�-F�e2G� ��&o�;����Ar'��������с H����=pI� '��h��@$���Cr��{X�F��t�xc��[��.@B�rB�5x ���aLÓ���-o�s�ʨj:o�-�SI&�؝�^�m(�d��<�����=@�Ӯ��#���r�L�cH�!�7x��lS�����r�^S�H�!iyy4Īß��<�E������V�_���&{��'�O$�N2�Y}v��oal�uކ�l��N���p�Q�k�=�d�()�.��c�j�1(7�D���F��0u���}��U_�6!D�!�����(�ppl�y}S��;C3v¸��T/wu�4����_�i�����L����X�^u��II���y�L�E[L����Iv���Eh��Tv��-\�k��پ�7Cp;zx�H�P���n��la/�y|�p�ެ8�墻
��΋�r
Z�r�<*��w��<L���b{
�y��/��E�Ć�V}��\ೋ�=��*���L��/��Z��Ъ�SJHܨ���o��H�+��F*�6���l���4bPYU%ۓ����V����bz0Q����eL&-X-@���bR��*�!��̐�C1�^�+�ӭs�v��gx��Lr�M�c���ܴ�2F�1�5K%�*�`觯ڽ^����S��t�-mj�LrU�x����C�eQb��^�����~���in$��߀����6O��ch��a(�*2�专��No�Qv0n���f���H�^�[���Uuu�ӎ���Tq
y�oslW{
���&y�$~q���h�X�}X�(�[��#��������t�FP!e|��{B�\��L1��g�G���i�t�D��^Z��HD2�s���Dy�f/�?_l�]D��yBnk��<7��:i�όd�֋mBı=̛I��6�h��f��{�Ns����;�*�c���j+h0N�&�f���*!��|M]Po~)���se392_o�PVNqa1צ���0f6)��c+�6�� ]~�[7%�7�>!:��C�0q���+V��9��6�-�N��
�`1;����/S��z�ۆ%��@-�fR���Fڴ'�!�)���iJ�Z�@�P�c�
����,-tG`�m��<x����.�k���(zP)�0����?��v��6����4��!\���U7ڼ�޼aw����d���陁��0����]�w��Hز�Q�A�eM=��5uB�Q��B%溭�7�&�tw����8J���P�`L�3�Tt|xs
�A����i���#94��A�� �>�{��%��B{<rH�Y]�hy��v�mV޺�X��M�Җ�I���Y&�ZrsQ	���I���k�~���m�g�1��΅N`��1�sͅ>��OF�Ov	����Ya�cY��9&�
ʉg!�Ѐ��6_W|�� �#�dDϯ6��Ԓ<(`�B�5os}�$��E�vp������߸�ldeP^I^9II!(�C�`}�,��_|>�� k����7/-4-t�����o�@�{��L�A�A�J'�m�H��Wm�~\.���de�A�G,T�h7�Z
�9HQ^fe���?<��n9��Z�U<x�����@S�߄v�=n���nb��5�%:J�L��c(�rKN�'{�!����YqW�]ڷQ��a�����l�K(���$e8"lz�j�b��/�~����N�.w�ä0e�!)%�[Q��:�`��l�b�`�R$����W�D�KHU1>,�M#�E�=Td'>��7�rL�G�I.�"�*��Bv��n}�V$G� ��(C]�����(d�k�i��ņq[琗����� P+�߿'z'�-%0���jtf��0��
C�XI����6Cƴ\����*�P������p���ep��d�߁�rK9�����3� 1>����ϻK�ZF�jAS�gy�/���z�}�W�z($z�ʢA��_�{�^(��쾑붹������HQc�R&�P���݇2���#5�w��I���:�-<ͱ�4Ե0��n�����t���d�uo#'�Q��A��_g��U+����� C�00[D��T��1=k��j�r5��04�S�Ū$�Dn���A<�M��d�B:N��JL��g�蛌6G��Ȝ\��F���R{�5�[k%�C|�!��Ox���{�㶨����Ǧ\�x��| �铁FɐD?�,�eyZR�1�s)�-��ë�3�6��q�1�BWo���"�T���ď�G�M��w>��4�JcA��/ ������M�\S�y�7�%ܲ���(��'�vTnH��M��q�Z�7��p�Xm}��m�����D����q`�-pO��`�op�b�'3(6{tc@á0H��qf L*:�Z�v7�����,^��\V��,F1�I��V��GD(9_�?�ୗ:�����J8R�?Xd�	��0��3��[ �'��D��7au�M������c
�w�ԡ�����������\Vs�0�@Y ;4X��
�o/#O�a�LPx�w�k�tU8����g�H3�>�M�m�U��E�SA{ĵ#Lr�m��,&���ԓ����$$es�=��'6Eļc�kΓ�< �rMmp�,Y�3�{Wi<��lX]�_��er��l����E�	����_�!Aտ��}f<-N؆-mQ��5��r��z���٣����H���\J�ɜ�&�^�^c3�����b��8�d�F����ĬG�4�wZ�gYb�VX�y�%6f��������j��-EJ%{��8?�#� �;�B�*��`�����-�ߧ]Ǯ�
�&�
_;]��a�F)�Ծ#�_���;�R�ULcw��h�s��M��2�J�B$��u��EuT��NG�C�/0�Mz��[>ZH&����� eeҭڅ��#j������Ӛ����ɻ�&��ְ�����Bq��2��Yu��ȼ���dG�J� 66��V��$�+�d�m6�y�)O�)�*7d_eLZ*���Q<@T���L�B�L�q�S9��lf|+d��A	��,_��I}l�Z\j��5q..�$����i�Zz�� D"�j�m~���+��GQ�_P�RsE?�\n��ѱ�Og�hM)�r�8
|W�9Z�[�y,����gtx�5㌗w�$4\��|��	.!�)��U�~Q"���qU�w�:��ڥDjC�∳�Xέd����]la'�w���LV�������)<N�+aPW7�῰�<�|� s�:
fo��''	�"��AX�I�@�1�u��dyz::]	)�J����F&Ȭ�p.o�_	�8�Ώ���{�@v&C�rRYA��P_�t,�<�DE����$#7
X-s�4�3-���S���[�0�V"h��b�,�G�K�:c�>�����2��N�Q��E5�)PK��ކ�{ 䈨������F҉pr��ɦJ8x������Zo�w{
��ƀLPr��3.t�k|�߮Kߓ�u�Dg��r�]���'3�M�9CC7�p/c�-��^��Ks�Ӽۖ��_Y���/&�l��'��xY��@C�j�#��Pj_HQ����fZ��͍j���.�xl��ɿI�_V���!�.Y��ׁ払\H$�y����Z���f1�"L�H|�1-��/����I�ۺ?�`�1;
���+cv�l��@+*�;Ar](��,4]Oag�p���3E��eR7��$��R�O��(-�wC��7[E|Z�^5D�t8��r�Z�F�"x:��.�-myC��&��&�R�O��|O@�T2O)˧��C�����RA�6f�������]�X�j���k��L�'Lq��WhS41sI��yvGzw� �H��GҰ���!]X��W�̎���6�s>`�!����A�1zӷ��$�BS*(��e�*�f'4��
^������7H�}���q5FuHf�m�E���xǇe��&O*Z�$���A���ڈ�s,���Fזې���[��8;�����P��
$��������F���=����Wu,�̃�x�VȖf�Gh<�0E�=x��}lc(3�������0�.}��#G<N�1%�5�܆��~%]��|�k�� ��Iy["�j�iE{�DP6��Z�(ZK�ب�G���Kl]@D>%��܁�jاyL^�ڹ+XlF9N0�g��F?V%�	辸�����k��t�;�� �p����a��ћ�PB�[;�D�>Q&��%�B0L�A����IQg��fd�	oc:�'�ew�w��ɵ��V��˄%���R�b�O�]�3�E��&\M�)��%H��j�]}����V�PF��i�@�/	n�P�o�sR������S�Ҧ�A��@��G�<���qg0�7�����Oak@n5 �p2t�3�Y����?��k�h i��Nx�&HZVG��<��4?���S�y�a�eU�\	��n���t�O�S�ܷ<!_�XtV�]�C�DX�x50VA�X��_�
��ְ�y�����㯹�ͭ�`k:�r�oi��=H�M���I����l�r�PM���+o�
��рR���3��F���i�B�z*�8�=J��A��W�����������B��d�i�e2�Y.N:�4�w���;���"�v�i�E��`2:(�~V���
�F��"�4������e�����SadY�d��H'OzT�\��1�&�1N�_���E#�犂�t�tbd88�\NE{6���aH#'���|�=����~Nyk/J�3N��[5���=X������eSݺ7z��c���8jr9w�"����}A �2�:�ɾK���s���ԓ�Y�����C�D������o�e䠛��_��1a'����}/���rZg�K�V��n!2P�E�{�Ub ���:2{l��m�c���LZ"���2� ������ݭt����?,���#��E����.bt��w��GM����6g�5�pevq�;|9'�O�?w�� ��g]#8M�����B�=pc�n���k��A�a�F�*
/,���7!%Z�Ő�mc?�O�R�愛��I�/f��g���p�f<&iC�29MB�����n��D���}�|o}܊�Rs+���Ǐqa�����V���wT8l���9�q��ē�zm�>$g��s������Dtx$DK?I1\H�d0��	y7)��s:��~�x[v��uly稫��K��Dbͪ	&T�^� ���4Q�De�T|��Fo�o�z�����u�i�<̪G7����TL6H��3����w&�0�NM�z�b.��~����F�q0�EctT��E^�^i�r V�-�컫�w�:��g?��E�I��/�:Չ�k�ͼW��J��̺ԒF&>����r=��|e�Po5�(PU�Lf~j�>W�Q�&��5�e�A����An��z�S�:��ާ1���9�7ji1�=��ycO?��)\��,�,̤�PMGu>���FVB�==�Yc��t��ܜ�i���)uz((?�y����
��������@�cE�k���c��B���]s��$��,�-s�PE��-N��᛹�?9�S�9%�� ���S74o;3x^h}e"��H������M���h)��Osv�ފ�if3��Z�g6��?� y$`.y����ԓ�3��#&�*[�Wd��u@6�V(�@�����O���_~г�J�$����纠וZ(���k�&Z��+���hR�:��,�o_���˰s�j�J�u� �G��q��)|��6�B����d�%����L&q?�ͬ��ۧ�=��Ҋ�>Ǜ.|�C`c���)��1q�z�s��ˬLQ�7�YH�ޏ%�ƃ� ��>���(�Յ��},�g�n̙�$���|!���~�f��9g��=���`]a��ᬧ�:Ǒ��ع�qu���>!�U�j��'��CGE׿���kec�D�i\����4�&�,Hb��G��#�S��5Fv�%d1���G>�f���ѩ�͟(�m ���8�:փrTTlNm��3���*�S��k�"JC���>���SΟ�?3Q��]�fr�J0�s	2k���	����o�q��:pG���[¿�m���,��t�6�N���,G'���)>��c*!`��������vN�ч�RH�%���h�-,�2Y-!�G�ᖬ
��z���H�>i�6|Z��E}��5����?����-tռ����7��(��(�D��UC<�^��W8H7u����9�\2�Đ�8�z'Y����6"��c$���Q�F�mDz%��t
�`tx{�[��*�����u�* �fE�L Ф:����]7%٢�E��~=�4�V�D6�Ф�85/;�\�Y�9n��Gxm}�g���RS����=ՓG�δ9��8���O�裧�i��	�pXx�I��/1kl�vZۙ���ϵ%��j;���g{^gī-ʊ����A�;��Ep�Ƞ��o�!x�y�4X
6�n��f���a?@��a�xT��{�_34 ���>v�W����i ��rK�0 c$Z�93����w�F��#a+ih��1�/�ϱ�(����\��nB 6ٯ��^^����<1b�C1&\�0�5b�=�U!�W�Il֝] ��>[(�!^�ot�}�8��Wh�HQ`�e;e�R�f&�:�JW��n�4�|P8���*�=v 0'�Y{@$�̾�r�'>w|:E��՚^�>$���IIrԃTt{��;�8r`���8��E��W���x�[��4��xoD1�ѵ�]�^�K4պ��#ؚ'F����eG�TsqZ~��Oq�xw��/���ާ�(^ˡD|��e$������r�<��rT� f�<;1�o�cir!��/�%н1{��"n�D$���ρE^G��lL��%�2T3�fC�cH�:��M��"�]�G4���Z6�RU��Ȝ�jk[���x�~����txK�W�5?ۊ��Hs�֩n7y��uG��۵t��9va�o�R^I���kfb��k�8���-���j'��+~/�X�&�=DK�tu���r�#��*ENm�/+��k�ُ�}��*�b~���o{�:��{��g	m:P߾�_�[�sS}G��m4sN\qV�>C�{m ^�����/�U�I�������X$������!���qM�<z����g�j�����0��4�����Y�OJxj��F��
��E�z�P)	R�q����=\-�(#�u���1T�u��q�|[��#&�@�*���l-Y_������RUNɇ~{O��0�PH�i�Ί^�1�t�&BžUX���M�ɤ���V���s7#'��<��� ���WDdI��#u���2e�8 ��D\�*��M��wN�Í�%pzX���Փ;��5ÒVɼ���/�����+RQ��)�FE����\�e�U���t�Ϸ"׌�^,5��&M"wc�_�7��:����믮�������s������K����ʞj�s�^8�̺Z
�G�P��O�[mcI���EcD@Sr��༌e�2Ɯ�QxVV:媹�=i�N���ni�a��ؕ�!9k����=�uM��I��<&��A�&��V~�U������.��e�o����e����ϲ�esس��k�S�f? ۠u��*#�Z4��}�l^���.��1�+3�z�Y�i��R�i��6�D��ZTu�7��e���VԞE�:�q����+[z:i¬�{}T.�"�_+#��B�69\��Ө��r�%(�:_f�dCi)�^-��ʸ"�lƘq�=>�ϳ<��O(���Ij�TPEo�ϗ�)0k���(����:��-Q1�GA旟)ߟ�Q���?��]����#�r+:m�#Ϧ0�s��#�06^Pb�$�Ś���j���7F},3�_=�0���&9OS�eEH���ȱ�7C�9v
/l �4��m�Yc�)�$2	K�ovM����R��ʟ}�׃��gM��7�Q��4�O��'�@�A{��2,Ƽ*�
?�_G�	��6!�/��!��O�P�����L4��W�@����4�1h��VBBZc���\&��>�IXXsi��Qx<~S3���ӀhV(����#�g`�ԓ��=���ާ5�]:����(���Z�SC���:���b���2ٰJ{M���[�;�bN�_�}����҆�k�Is�!����J�pa�H��Է���0}�Ip���Uq;�w��V��(�lB lqN�� �a�0���vq� m;�S���������'�O���Qlf'0�	_1�eyt�:T�.���ԏ*���>����D��R���~�dS�;[DC��i��<M�� ����OmjVԧG�I�ĩ�
(�z�+y���n-�ϯ��s����U�w����ߊ`�֗t�l=�(;@̈��X�	�$�FwK�v���&Y�'��;�����1G(�\?����W�t�0.�띞P�Z�>��E<��L�0��ǚ������B�AV��p���0���(l	�H/�
���:�0�)��.�#�~:�+�/ه<��Y6VKyX��EH,z��s��@�u�����W/��$:�(E��M�~�!�o�ZA�N��Gʯ��iVWy��ZHEJj$�ň��� �'�h��	ʃ0��;U�N�������d��3.��j(��8TŎ���k�a�Q��'S�} f�3���Q���@g��p��r�HUX�ݐDzo������X�-�k	��_K��m�@����O�)��v�S��BV�Zζ*�}��E~��T�WM�`���=���
��kB�Mr��jӗ1��c�=�U��6z5�}����|w�kn�����L�{�/�q���NVd��=�J �%�����E9!�)[��V|i�|��=<8U�D��p��������qB:�.��M����\�.Pd�/�8�퀅��t^&��,��[h�)�k�b��~���qt��>Y��	��<�y����Kt{L�l}�A���]S��4ʘCr�uLʞ��IK�y�M��fFS�7"�{�ߣ�-�A�'�1�2�2��v}V��/L��:��C�V+�~��Wl���7���,B��͒.�ښ	3/"���C2�"��2;�]�zE��&��btC��Ո��Z����%ң%cq_A)�> N���]�{�c��pW�E�T�l�|����k�-`b
*�G���d�L��I���D .f�n�6|�7a��pM�N:$z��|+5V��%75�t΂��h!�7�`A}G���?"�+��$��S�SL���fK�$�v�&�<x�o'�2�jʹ�
�)���D�`�.W:�e�=1m怂�{j&� Q� s˘��>�`_8�^'
���F8k��Qe4'��mϵ�y�E�wv���+G��"xQ�G�%?��ixS�on��FN��ɒ�����XCS�#�R�|�B��y��~:�A��;��Ũ̅�}��+8�^F�e������l�3�ZC�!�MS�Ӄ��c���C鿎O��;*��G���,IdD��Qg5�s῎��G�ؽ�Б�vK2*���)�թ���S�;�*=d�\�ˀ�SY��xs����eY���@�c���xG3���G\C�]<��s��[4�Ys��(�����z�u��l������}�Ԥ��c�5�+�e�߳sؙ�؞�rYiiC�[��-��`gsIb�Q�H@D��-4Aa�1�GU x90�A�b�"w��\��ސq'���\��biB\�o�/| �B������k�ż��EuHS��h��ouw�L�2��<�d��]�{� ���CͰ������ p��DqifP�D-#�*�/*�sHs�9;V��c�@V���=�G�����ޜ2X� g�1e��ća�`�"VVu�x�2eK:�O���J�P �_����p=������x�	e.�%��rm�V��s߃�#��rN�ň0��0�p#�鐆���U6rhUo>��݋x��"^Nw.����{�r�Yj���p%2.ݵJ��(���0�-_`��rv�y]E��Ҁ�ҩ�J2c�]��=��l�G_MX�W���֋įi�}I#_��뀧��?g#V1���w��o�O:��$�Q>C���V"n�c�-�q������ q�v�U�ca��Ю��Et��&�y���F3��&�I���7k�Cg�\K�Rχ�_�:7N��*i^���o{�@��#����WW�o��Y���֕���� a���q�tٔV׳�~�xK;�ё9Y��p��w�\%[�2Ђ �Q�-�� =����D�s3��%��f�0DH�/����#wN�W���$Z��~�ixL���|*��̚]�h����[��8��` s��x����`��\���,q9�W��''��Of�ؼI�z�2�A��L.6�O3y[A��z6�
�/L�v�o
�ț�n�~t:l�R<�8�N���;���V~R�8;26�l����nS�&��Mj��~��~黁���.��(J���"/���D��s)Ǩmň @�s�nH'�p���[�8���W(8���f�U����ѱi�'r�ty�Yv�Fx�lD2j#�Uly+d4�n�)~�La�&�ˌ�;,���$������N�5�o�a�i��cZ�\?B��A;��\��Abm�m/�Iڥ�����~��!Op����������Pnı�]�a��I	�x8Ön�xGX��oء�5�j���\�.
��+���۷/5�O���nkծ#�SU�BZ��W�X���v�ȁ[2{���"1��3��Bй1�uZ�]�bZ�Uuz)���X�D��v/�ɕ��7��Neb�Aމ��#�Ù���1�y����1��py���ٷJ���&(�2���\�J�f��~�	e���5'A�[S��>�������A�ǲC���{f����`L��nl�Z3���B����[ǩ8��)?�)MoMy�Y��a9D��	��	���`��@S�&��5��}�w|��H
��,����(Re�[�,�Oj%�(j���g�T8s3�Tn�\�͐�)�ұq�z�f�^�U��8-�a��D�Ԙ��EƗ�G��o��坄,l�}`�GM���+E�<[~���42�;�,#�d\�[�\�nO�H�i��ʁTY�-��.'�v�(��ȹ%�4����'t��Ϧ�-A�&��E�ʭ0�;�<b�/�nNA5`��8�ua̺w�����������h�(�UM�Zo���3�Nz2=i�L��G�b�]Q�C�:��Rǖ���C��R��[�;�)�͹6�FS%�Ⱥ0[��0��� ��%j,�y�pw;��]vC�����X���G�8�����`t�C�u��F��fh�w�-3�9B��P,��='N�q :�o^(����o;[�����n<R��M�?��_���HW���n#�քr�&�2�E��e��͸���C?����Rh�j��:j:B�Ց�`���5��lG�YX��A�L/#w��A�x��f�6���)ݩ�RS2nީL��c�ʼ�x�E�P�E�JcHDduT�ى��)��kS�딹��G��m?�=Y����t�An��	V&��Dʵ����P/�#�I�XU��M�-{ר)<��BR)"��Oc��$P֌T�ǰe�hz��RtZ�%�e��X�����*tqm� �O	�Y�����\��x���U��} ���!�u�n�� �� ;��g����&�?��^-0������l���Q�����67��ٸ6��Y���Fǂ�:�f4����_���v��`���=LP,a���{���G|l�� ����|�v���5��b��T�w�
��� S����y�ģQ��#���q��*>|i�����߃�FG���޿,`.�#�5���_������)�r׼t�����P=��$Y]�(uO�tfGeaR"X��l�� �A^�J�V"A��6N	����Y�ϭ�4I�uf_8~�$�}"4��c�=�j��QW���* ��;~U�a�a�߆}����^��A$�ec�t�O�R��0Bz�ŕ�3'�.��?j�2
3�{	�e�ō�P��0S�3lx�}'��tbc�X&l�k�Z􍫑�\��N���L4�	4�1{��)��H虿����s���_M0�A=9�^�9�,�;��Sn�.d ��.&*�����N�<�ݾ�Ac��mŧ2�/w�ev��m��9�z:���2႕�˵bP��֭�JXq�J,�G��SFO��֗��Z=6�{m�y$,ͱ�k�� ڍ��-}V�2�dún���;�Rp21���M����ٞV�ƞO�t��.�}��g
"�)H�A�/�l�2����5y�ޛ� �O2ul|�g�5���4e��2Ie4���d�r�=��X��9ؠ�S�u�s>e��f�>�KԸ�6�*�����P[r*��e��J�}��Y>(�C����t�Z���K��y�3a5i��-������������]��K�t#L.@�4\�_D_d ��^�0\ O}m%v��T�X�m�*�ۥҷ`%�u_}���X����j5����<�ϵ S|Ʒ	1ّ������ǋ��1fIn�h[M��}��bʓ�0���>�/�L�Y}�͡���x��uM@�P�[K�#(}�p0$���ic�j��\n ��&�[_D{_c;JU��~�׿<����l�1'U�)@�'����A�S6��^oջF���j���S�{Q�Ou7n���#V��}����َ}����22�[�z��ovƊ)�^|E+��G�
d��cw���v�,%����7"��W`i� u3�����uG̳�� �m#����$" �;�&<�<[�{�ϩO��K�:�&cm���w;����X�]�~G$��"�@��Z���R�҉*��rT��Vf7����9��m�M|}hl�2��8���62�9z	'c�hl�Z�s�-�\P��=d�	�o����>�� �?mPO|P��Y�����~�%V��M�?�ms�%�\�R#����4{��8D�t��B�&����x��Ok�M.	v�'��`�hc"�|2fə��\�n��lk�I����0�{5���l�A���!g�[R~n@G[qHX��bp��n�G�U��
|QSm�
l���@��O�����ƒ��/�{�$I�}�Rbu�Q����(���4���_�v���Dﱱ���P� R�Uz��c�B4v�y�f�>�b�F��A�N����ҧM�uCW4O�BV�)�VR��V���z�(�HŻH�zz�~C�u�`z?m��j�¾��1\f��Y�=Tr$Ь���~�p,�Gx�.Yi��/2Ű �2�L�dŝ(@�b�G�]��_�-����
�����=�SwY>}�7OU!05��DOZݱ!���Րj-��h�����A����T�T�!�n+�*�q��Ilo�Bk���N��+�БGc��i�
�84�N�<:f^<!rți�5�0Ź��p��?ĸ�!�z�"������}S��3(_ 8E�tddVO���,H���3!Tj�xv�K�e�����esE���v���zR��?˰��Je���GdCK��Ìǅ�>�IM�Bl��ЃLif�u��/�t���t; ��A,�������\۪�#ז�\!`�rS�!��T�m�q���<�f{f����L��m�Oi<�N=��J_��[���T%�^�@�.�Մ5�P���H�P��umJ��c��;��	e_�X����rqw�
�3�)�3�7�;�#$��Pg������`O�ie���٬L ��?�
��R@�7�:�=��PZ�h�`�D+WĠ<aP �	��+	7]��P��V�^�� �w%n&X��ka��c1T<ҕ��,�� �'�Q(B	�J�hI��p��$������(�j�ġ?��)���ʨXM��G��.�.�
oL�?�@Q�GZ�%x��,а�� �h�o�.;�>1 �;fOĠ�,��+6����5uF�g����	�l�l����o,fh<]pMh��7�䮗�ⲿ`�K�%�8V~e�Yo	L�7;N�3�ބ=� L�FӁ����(��2J	w{͍�f�|�R4
�_1�c�q��z���kOw'Iz*mJZ��
��c�<���ϗj��Qk1�q����B����w�dɦ<���l��}�W�,��">�*
;���#�����/*��S�)=�'�����Ip\��dQ+�+����L���R�=�R�Jǽ��"���p�s��1����z��xQoo%��zb���DdU��;���	�,��ن#�_���[&�'��'?��\�D7HPkF{�1��%[�T���1]1,xt\����ޥ��R���KPn�o�E��Ÿ׷��&5�$䯺�~����^��-1"��b�4�7�=j��v�M����0�M��W5�#�����J���Q���-2ث0fίȸ;%����ũ5�U������,N@q��\jb�ʗo�lE�r}2�kP�s*-�ެ��ί�P)�r���>L��x>�i�2qHH&Urbb3���P�P�n\i�u����-�V��#�K{��oӃQ�˥��>��'�m:Dz���q��f�;�$�e�W�#�.�&��I>I��g��-�4���S�������A9WC�7$u7E��H�
����C+����[k��3a:䨛J�o3��L���u�M��W�<�[V�^�H�h�6�\��{1˨�R���$$aՠ<%AS�MZ���{ܪ>�	й2��58Hԉ���0;���u���ʊ���8)��*t��-n�.����m_�$\6q��W�CT�>~��-uOrժ�U�4D�<�y��f�s��qF���b�䉠k; �w��dT՚���U.���S>���G+�mG��鸅�������9�S��ż�,<�9;巴����K� >���������AO�9Ld$J��)Ƹ��o�[b�ݝ
�x�5�M�k�뢩a)wBPhT�Yآ�ĒF��ICy� ����!�T�������̜��!�2�\�׻E�'!f��6�ؖ�.�s�Cr�� ��o#��LO�6OOR��W���sd�&<cA�G)�z����An�=^ M&�^��Bg.4@~8$�ֆs>�kt���4[F��v/SCh�4���� -����cZc��2�yY&+�['@M�X�\]�VU��1�PZm���zlI�V�5��4��ԝ� |�����.|�L���>�ς�.�U�KF�_!��C���'��ث_+�;��0D`�Mi3�U�H���ZI�i�	�M��Fێ��pF�4�VCJ'�{V��O$���T�R�ʂ| �Z��ނ�l��񼴥� m�~9Ast#��"ua},�K���	
:f�e�8��
j63	7)6E�K�_�|Kcؙ��S,����IF�W�Խ:MԒҞ�$�a	tK�0n`]/Z�9H~��J{�5��-($�j:\�4j	 j�A��$J�X̦�Y�a�LVyL�Ef�U� �_`u`lYMǊ����̠���u�"��O]�x*��YO��^�G�e;5��Si���0�̡�K	W�T�^X+��z�ScA�A�f���*���1fd�w1�R��<�gl�gkd�굊�ћ�J		\������j�}4{�X�Α���h0X�ͼ�� �&�W]
@J$����a�m���2QģwܣDߣQA��A�e1`P�h�v��x�#Ş���h��ҸZ��l�e�A8��M�Gr��8d@PGZFA�>���绯�t��"�w�n�$/�]��+F�=�i�t^|ǻ��'��"�P
�e]�L�KﳈZ�6�Fl2��*��f:R��S���0�ߏֺo=������Dx6 ���	�G;$ۓ���1�T�:���DN-V�dF5�&�,�&�+R���}�j:�ro�����RA���N̓���a���L�`����^�T\6�o.����7l%��Y�¤�s�u��-�Ɍ��2--1J߄~c?6D�*?��BC�-�R2ɨ^[��d���-�:�G�d'�%��RK�L��t����F������������"��C�!��>)�� {9L��T��u}��������Gc��_?���P�@��Wk�?:��lǁQu�=���(�idw��e˜�/��~�ƃ�=R�CE1	o��VW�FB^�]�WTϓ��j�:Y�\Y	4DZG��
X��K��x�M���M9��~��tO���O�$�/�29��x}b�9[Z~EՏ$����֠���qe1a�3�����pa)�M��
��,:�HN�JJ��l
�͚���W0�+�v�����Sjۻ��7�~~ePRj�{v���1���'c&�)�N+zv��2<��NI=��ϧf�������c�,&I�˷$�e/�Xm�aKos%Պ~1��3�����l����)0:1��:bb����=�����&����E.��=����[�cu�
��"ot����D��WfP�qg��:�w��alC,JJy$&P^��%�IfR#�˰"]�ZHSK�.�����S�Â�+���g���Uk��W!_e�9�KH_�2H���L���:��Lw�k܉E#�[;���V@Ԥ��p9�'�tN �v�H�;t�6�i���]��?ĝR�A?В��m���EX��V�cU���n��ݨ�n���/M��2�{��`^WeRb�'�p��g��e_�{s�W��������BW�1��ŕ��(?E� w[�~��m���m��c�a����ϣ��z����j螈7szb�eCc]a�q������L�E@Kt?�~�@�]��yҖ	8�VG-
�sW��$��_HL�rZ���	�f��E��t��*ݎ/�W�H�C>����:����%���@2f���!�H�f���i-~�R����>����JeZ�b�yj%�9PZ
��n l)�[v?:��["��@���{pΧ�DK!��y���0&��"<���
��aa9��Ԭ���Q�'�i'�� ��H�1�m�L![��j����ϛd<̩_t���	Ԅ�+o��1�-�.��{H�p���U�+M
´!B�^�����je1����_jh�KrG%p�zƃ�v�����$�nf%�s�6�mG��H�a^u�ޫъL�F���sKN׹nQ�B��8��B��2y��e�v��^ժ�M�Mn,P4�/�A3�hƙL~�ޫ\�RQ�:�{Y�P��f3��(�e���� �w4�++J��b>m]�^�㫖+\{�����X�=4��G>d ��˹�����|�)����-��I)��`����[.q&�g��۫Bd��KJ��'�1*s�F_�r_lSj�h΋T�h�IfZ�I�S�Hn��4���>?�3\>.I��e_U�+ɡ�}H#�
c��[Mxa�L����lZh��"
��2�ox��:B)�8!Du@B��,Mb����F����׷_6bxo5���Ҏ�H֜����6U��؋��)w�q���؋C^�;��Dj��f�|ml"侀N}�u�)��W��%������������TL:g!c���Ďb�t ~�&l)FXw�0�������h�rӂ�Wi*�����T�k�����%ǅ��^�Ճ���)̝D�=D����e��N_��j�R���̔��w�E�����D�2�{Α���� �?��Q[��~ĥk��xؙ�gE��l{��Q؁�>-���u�0XRu1��?�и��*\Y�^/��J)y$��+O��6ρc�򥤑�%�>s`BТ
CR&��{�Го��cB*�V����5�������$:�Lx�Y`e��7]�^�ѮJ����R��i�-���O��4}�V������B�N��<��1ؐiTk�	c�Y�ln�+?�a�I�|"�(�CQ*(�
 &^��%���g�r�m���C���̜�y�%�8vr}�����dRՒ\c-@�����5~� �{	'���4bㆰcR%K��y:,sʳ��R�F����M��DR��H�Ԛ �� Mqh7�~��>
Z1�a6�{�i��2Z�(wm@��e��z�M�U��ڃ�FS�)6�0��1�B��s�a�O�3��-ro*�<�<��5�=���d�*�R�&�(�`ǻ	��t����w��cqBݙa�1�Q_s�~�����ˈ����z��NNF�C����!pP�gShb0�!�r�س���;��e��EX�n2��|�������2Z~�Q�0�pW��2:З|=/%c�����Gל����H�0��~��؀��"�c�y��!ܵ	�\�vp*q�'�A�������S�<�b�Ģc���k���8!55'�n�k<f8��,�|�P'=��%Cv�������������={��nϖ�T�^�F���,���Bi�c�/E� �ȁ���`�	�/w�.��9�w�o@}/zՒ\���>���PM�qZ��~]�@9��%��\�/h��ʁ	�h<z����t�b˝��HD<�:?�g�	vK�@��I=�75Y~,��&5nC��T��^�:����o���؁P�����-|�0��o-��@��o�_�'�h�h!���Qs�Ff!�0U��	�`�f�~��ջQ�@�[� K0���BA�c.�8���FG@+�ٴ�{� �>�H�=�}A>qp�җ�>��aqF���&,�\�P8\o@OˡBE!���x3��iR��C�$�s�2f E�bn�Gm����\#T�t���"�𾄮�~9�"�5�m=C���N�X�&m�֯���	$+��e���6Bf^P�)�kP�	;��8H%+|����v�c���Gس��N���F4�e�C��)�I�},?e~�������_�6�Ӳrd�k�?w �*�Hy�*~]KpU��[�Q��I�V*��0�m���
[��GC�7g'd��6TJ�Ff�g:�q���5.=���1fw�Q�$~��J�^���%�y��N��1|���<��x�#0'�<3bD%C���ʂ�C^z����*)��:d}�µ�%���y=+gr ��oƏ�:���t������꺄���a৾�﷝Ȳ�t0Z�\�'o�]�c���<�V]����HV�%G|������!8>�p�(�%��Y/�yv� �]3�7�Z�þ5����!�{���s�vƞ#r�YH�7�V�`^������$罶W[t�+wo��yJNv�ћ*<}x>П�b�6+#�OV:����c���-�+/#}x��]�9�U�J�\47	��=zk9O���-�k`E���ef�!���Hk��?�βJ��N�sgB|�P��~_��j�КdH�)a�}���!|r���=���Z 4!���j|��t�qR��u��6FE�4
���+ι�QL�k�[㽱�K-�|���!N����+Js)�w�$�H�q��T0�j]�9�u��ҩ*u%A�K:~�T�4�_�{D%�z��e�����X�;z���3����>o�I�U1����"H�R�f���g���n����v=[j��A꧷�����6��ЛijE��jc0�h����~�තP�q
T>�y���9m���X�>l�����a�ܼ�V��O�R��{��'a9�zY@냀Ė1?��G2��Z�쀆�]"�z;P��#{kY�\*:d�F1�I��T���:&�#����qcb�[�rA�ܿ��w�p����-�&����5���6���s��@U������C��7�BE��.�Pur�����i�yCa�,������˾^qQp��MV������G1���J�Bj�m�8_2OtɈ�'w]�*���5���Ud�I�<�j��8�+���n{�J�!F������o��'}9�w�tL������. �����(c�i�
�A��rfu�#}(H�=�w
U7x�b�I���K��%��A�6�jA�AHǧ�z+������U��]c�mU��U�D�b��-=ձ{M��>oT�}��;V�����9��t����3Ng��x{��%7��MA�O��U9�����i��r.c;-�H�р�Oug��10���N{��vw�Ѓ�2��Ӳߥ1�)Ѽ�H4����2��� )�?���b}:������g72mO?:��?���D��#��J��񛙚t ˨�$Txl��3�4��8r���r��h�3�ua�Ǚ�S>�ށ���N�+����� ��7i�
���iHo��W����h��!۩  %9��l<�R�.���T��Y���֒��إш�����?�˾_3�����2�eB�v�q��4�%���i*�(���i���A�~��W"�:	&�Xm����?�X�q�5�eb�1-N
���x��8,���m
^�լg��Ղ��}��v=]���������(j�y�]QR�%�$�ٞ���{�V��A���X+ōr!����ƭaX6� 'ަ^&xgJ��|�oTU�FF�U������p�K���a�P����.�����7]D᳔���'eA�T�(A�S���:e�c(yi�� ��m�ڣ<�cXh���1d��s�����!�Ú���b��BS��ݳ�����$����H|�I��#�Xz���>
QP����>6@E�����փ��y�qn2K�s@�0�yf�b* ��X�)�DK�j��_��i�z+arX��Pb��g�a�tVK�~�����F�3Z4H�l?�rʐ��Ħ�]�d[KJ�]��5����r�B�2�~5fF=7���Xi"B�
;AT|0��������#�7T��	���=L�Ma�E�����Oh�y�6]�o;������F�|�!iF�[��G�J��fM�uXP�G]���Z� QK���H	Dq���]��χZ1Pk|��c������b���0z����u,<?���	]�L��<KQC�
����� ͈��.�p���N�ɐ��:��'�[�?��j�(���d��Z��l��-������5��j]R/����7#M�AT��ʉ �||�s�� ��_Z�,������8�i;�R�.r6��-��|LK��(�=�ywuV{��`�y��o�bӛ�_�J=�m�*���m%g0��K��A�Ur{ys_�Ӯ�%�҅]�v�wYG���s�BH��z����dK��rY:�4Ħ�j�T��G{L��T��]���t_���4�^{@a�!�0}�!!�I	�x0�Y��c��BPx� j�.&��M�K�g'�9�L�^d+(�S��;7�%,���FV�����P,*�d���*��p�EW���g�"�vM\:�Jz�5��Bk��X�����s-xc�7Cؗ��n*~�k��>���{��e<�lN;�)G[��YZ�kW�q���������n�����U��=�e<�]z$�������ﾄa30γ���/Y{�(F�N�[�O��ьD�w=ԓ[�}1�Y?$&2��+%;�+�E�Oh3$Ru��\�U�<y�ȑ�A5K�L���!A檮�	`���ׅ3}�4�m�htCJUy�&��!�y�R�@�D):���E�&���1��[#�W���rV���F�j�����Tm���U�s��f
߱xpcxͿY[��X��9'�^���I�bI�3��6����f_ �nh�N�����KQ�ܝR�R���UZ[b�\��z������Zހ{�����4X�;����`�����[�:��E�y�^���1�J�#�g6}���7�&��T:Ȇ�ԥ�!�ngM�ŀBM���QVm�ǐ�/��I���3YCƐ�9H�Ӈ/����4���k�``'�j���2�W��ٴ}u��L<����|3��� �x�z��O,������%ȇe<ɕ�� ����g����^F��i�hK�泛4SJ���m2>zOw�ƿfk{
�9���h3�-��ٖ����Z^��La{}����ߠ	f͙80:��B�q�����^�Q��
����ܸ�W �Y�ο*��������.	�����z�f1�����դ�X�U���b�ut5��J���`��W��{t %�z�{̨��l�:U��.�����m)�+�#�E�����=G����X�bq�k�ړZ�\�����e#ǣG\�c�*i�f�N�}�3-'��.�9rƶH���J�ɵ"�Dv�Dއ����w^�����l��!�o��3;�B�����"��^=J�V�}��T�3�u�b�pilB�*#���Qi�Xިw#�g3Q3�cȋo�b[P��੔PH_�u�2vM{�{6�ko�8E�'��q��.�����=9&��/�v�H��d��??��N��h"���×(~���M�zQ՗QZ�=��m�P�����÷��@�i&��ƅ?�w����5�c�����_rv_�:�]�-!k�~٨{���Ĩ��T@�	�W���]&��J�A����m���)׃�!��m��E�V������8��C=|Z�
^�@yv�b�L~e�VV�|�P��)�Se��-� >�l��jRW��O@��XO��ݙ������`�Ѥ\��.��8�x �vRx
D�YzM��˱k�L+��BZѵ�I��`������;��==y�ܛ$��u��B�	�0�x��,d���RVþ@I�,d�@�-�v�\@��:�����1I�>���~@rm:Xl�9�8��e.o��Gel�)S�i��}����r�����F).�Yi��?�MR���]���}	�U������G�K�i-d��l�r�= �;M�+��-���Ch��+'[��
��m���5,����) l����7�{�ka`��b��˚�#Bol��J�$�����^�S��l�*�7G�����9�'p�w��nЯ-�N�.�B��,��� �#������������G��?��?�ā����2OCB:#��'KSQŐ�m�J�/��ϴ��4�'.I�3X��#h���2��^x�UF�nG~9�L�qG��` �M}2؛��F%EY���2l���{�L�괰{��� L��\��M�e����Ɣ���GD��x<8�r�\���yyc}U�AT�j\Q7j8�X�5���˶2��_���߁��yf���O�s��z��	�ѫ��ɚ�o�q���f�;�;g[!$�}F�C_
xKZ���Qʢ&[�$=�&b�G��Ix@:���dAZ�ހQ�O�v�����}�Q��F����$���u��-�]w�;>B�}E9�J�oŀ�>��:��>l�X��?�EJ7w=�xjߩtpd�~��׾&z �^RTX��S4dJ8ie(�!�J�MU�@<���Ϲ��jbAh����wg��zt�1���-��;!�[�`H�L���]L�P����kS�7Df�vkhGT���t����L���T�X
6Lo�!3}\W��Z=,�|I��.@m�,P��u�3 #d�hve[�x�~��RK�՘�W�z�g���ܡ��F=#�&��ȗLW���e�0W14���&��@�&�&vSml��j���4ؒ�����=��#�*�2��i2��g�J�����n��p39�aO\3o5F#��X V'�{_&ݱ��Ӿw�I����);�����Y�;H��U�H찐+�IX	��7���*��VN:7(�J�P����Ԋ���ƫ���½3��/�>苟�A�_����
u�.���/}�}��
�%�yEuRh�yX�������-���\�.���g��h_!f��Ops ���A�+��N�L50s���IC8o1���Xg��w���eB��>mxu4��(TY��\z��Y{@,���s����1�]*=���&'�ӕJAk�g[]��`��Nx��.�T[lś��-�'r�|��H��/j��}�� 7�ƚ���D�`#�g_�\
�q�se�C�:�&�	�I��ZmKR�!:�L��3��	�_�a�VK�솧�e���JtO�JX4s�5�cOP��W?�1
��u�#Z�`��i���03X��	A�I��OF�H���"rbƴ �p�0�Pn�勵���ou�4��O���Q*��n�Z����g�@�wK{����'���Y[�Gt+�EK%c&��?[O�A>�B�9X~K��S1�O ���%��O����Ѵ�����6M�����h$eYH}��g�i�8�k��� �g���b�+���!u�1�z�.��Cu�}�o��cnzࡔli��v�r�b�XB�˱,���97b���'��آ}:�uu����		�+��`�o��5����r;1�y~���,��\�b�BSO��!�;�oRSL��3�Z�6�O5K��ݑ�V�es6���6��wKuN Z�{��E7����y=6�������0?�iȪbS㫵��QkjʥG~����؎�\�q����
Y��
Ԥ��O���{.�@����X� C�����/��������P�N⬩�lfg�Z�@��"��ΏH��;9��0���S�|��!'��gh�J��@gU�G��6�L���׉i���	�di��?H��u��nM#?���Lx�i�#��_��f��R��\�Q�7�	6��H���{%Ҳ?�~�y������Va0�R̸.l�Q��'��a�F������Ya�|�ĝ٠�+�Z��#R��Pn�P�^���t(�Y˷��߽�����	��i.#���h�g��?(�q���`L�:����JQ�+�;�Jk��ABc���Xx"0J���U��P�Wa~����{��~�/�ȱ��FY�g7���=��T��0���nV���� +��Ih{�a���(ez����l�c��0n�P����7У@�f�8N�_�t\cڗ�'X*	��]�BDOt�"�g��J}�B�C���ς~A)�;'��iy�H��E�&�T Ǡ���դ��j�}:�-*}[}m��d�k�����5�=P����M�Y]ED� ʼ=v�h4�/�T��ۧ����T����#v�N�Q
d�ch�J�k���JBK$�/�\�7�I�B\aϚD�_���ޑi���
��i�0�׃ T)�̢��M�=����Pբ'���@�L�j+�֩~���ߍ-�Lq�#\
�@	��/ᗞ�ֺ�4�n���R� ��̉#Bb������Z��I��+vC�{Y{��k~I�ЩA+�����K��j<��n��lDC�?��/~&���FT����\��l��e}m�q�����6ӥ5��N�{<�ay�"�䫦�I_������k��J��d%7:}ͥ���C��`s�;�&I0�Pچ�Q<l����3�H�.CnR,Gx�6r��Z������@"T�H����,��`��^tŇ1��
Y�M���*Y%պ���XF��D��J�sW��Fŵ��!ޮ��#xUI�+\��7�p7�>M

���ވ�j�:~A������5�GiR>G+�\�,����a�il)ך��{��(�	��:[�܁��J��茧ɚ�ʀ4������%���j����)�$�^Ɗ�[��x:��c'���Tk����%\��-�eY[\�%���B�k��}�c0�B�ʄ����p]*�J�Z�j�|2��z����\ � �s�<ƪ��8���5Ϙ�$�>ڋ��N�K?�ٓ,�+�:�*Q�m�]P?]��F������A�{�,v�q�:�ȵ����.��~��6�|�.4Z��D>+�"PLoU<"��kQ�^��R��UL@_�[�(g��*i&+�Jr���*lQ�]yr�e��#���	��°��jX�3�;�M�:�i�!��Zx������q�J�e�+��٘Q3\�@�9�7O�k1I��o�]X�l�4rڶ��Ѥ��PWšm��R�~7�]yNnb/�ȹ�L����sN�K༳�{�F�ǉk�Ǎ�8>���>P�h(����t��������_�������Eno3g$J~hHK%%!�����c���@�Q���@"�a��a�p~�1�~2������qI�`�Ni^��F{:���y!7�3~@K�1��	��!rG��ej�%�����%�_�U��q
U~܌��W�G�n�l"�c��P0EIl��� �Q,Vɸ��=���eC�J(�/:,T�
��C��!yg3�h��5��nw�ԟ�
�6uU I�%��Ȗu�%s�枕�A��3���ș�bs`&�e���:�f�^����hґ�eU?)����y��4�v���A�ۻ)��,Y�Nǖ�Qy��391�vZS��&Z�X�͒.B����an@�x_+�@G����4�*��(�>�1�%�Xm蛓i�����b��L�f��f��r	�(��{��іo�ɭ[{�36����8��وt��ހ���~Ey.G�\���M�jw���9q�DhGK�U]�-�w#@�(�<_����ȣ�&�3�q�)β�h'"ү ���ϥ��G�����#Ll{NL�E"*��F���)|���Ӛ3O��~+�!H�FJ���:xf�ӑʧ�ַ���`|1�8�����*�����Xg݇I���de���Guf������U]rb�����Og&*d#�7���F*�@$މ�c��IL:Kƌ��S��$�o�'L�D`��AG*�a�ټ3�7=d���(� ����bъ�̟]���pM.SԳ�oP�0���4�RG@��B/������v���o�]�G�1ț���1���c�a�����Q���H��?�y\\��E��:`F]�-�2��E �ԝ�G|[�+b&����b�����kZ��܏���d.��R�:#��@|��^pxD����c��,$2�⒔�?��lV�}N�M(�e��o�g�#$~�{���+��B8Q�L�J�D�y�_fc��FoJԆ�&�$����9֘�e��6�6mP��L[��8�q�N�aХ襰R�m����C�} �#�+9�߄�''ULM��Ы24G�VY ;�9�/� ��
�xw7W�E������`���2�Xj	޼�}����ݵ� Oƹ�}���	�G������h���rc�:��"'+'iC�4�gZ�`� /Gj�_&QY�W�Z�bqh���|�b�QM�o[o,��c�Ķ��p�7��N�~�l�j������;��o �Ĝj�,%d�jM�N����5�/$�uUn:�Y�_�5��nA�6����:WӦ�[T�Y�w�|j�al��Sn�.� Z}��2CB1(q�I5#�]H�{����(`F4*�����gP���bH��w���y���KF1; ԙ�B��Y�$�F�i�r}9eVn����ù
����`,����MC0_�pwo�����s�xys��੺�o�H/�SB-JBxMW���(5�k�.A}<�>}�>�A�K�S(���/W�mQ�������..C�����@���T��� �7D����kA��R�R����r�!�F�z�&2���*����[�)��`"������b�8����T�Y8
�?��6���t��3}6�`��\ӕ�C�3;`�E�I���u�]����/�^B��(�q��d!�UG���~��?��"i�������s����s%��^<E��9t��C\/�z�T��j� �`�G�fKD��X��j���)J�^^��Ӧ����K����\ ��V�-S�?,�2Wq�I,Sj�tS���q�p0I���I]\�ڮܶ��I����Җa�f{���cp W��0���GL���z�2�o�c8�a��[:*�a��h{[4E%����?u~n�C�� �,�r9��'j-w,"\�<�����Tfg�br �jX�=��ɧ�^�`������Q�2ϣ�9!�f��Bf�;�f���%&kX�O� W�s9�0�I_e���F%����e
l۹c�T6�_�՘�:QF�E�����CQ��Eڙ��
���)ٺ��8�����kiK�}��X.1k_���;:H����q���a�&�ˡ�.N����Z���a1�E�X�?��l�>:���,0�����bn�+��A� D�OނMB�������U7kU[t���工��i�]v�������&�6�G5�F�߁�q���!W'��\D�
�Ӄ%Y�%��͛�а����Y����rv�N~e��gh�Mk�͐l�9��Jyǆ��'~�F�A�������	�Y���hp3e�]�v[N�,}Y��"Ԋ�� ��Q8�r�e�0|��_.�GT�v7󗥶Q�!�n��f�>w����T��`o��L�w��R����ձI�H9�ck�h�ڲ-1�'���� O`
¯W��Y�"����#�)�mV�0�שּׁ:�i)��
�%��#�J\R��d��믊��dc��߲�D�+%\}0�B��4KEe=��*&���3oy>q��}䪯���6�a�D˪-H+�.�Hr�%+�k��"hؿ�����3.7ּ��K��p��v*e�v��&1�3�Qkl!����U.�]�����d���)��R�f嘰���j ��G��"-dxdӔ��J��iK�$�>������WL��h,F`�4�D!Fm������6�~�xح�`�f�+�GhO˲~�Y��=���\O4(�� )�8㩭HN�x�Iы���S�X�l�vv�s���Ο���. �H"ݮa-ch�H*�xd���W�)a,�u#o��?p��I�^�T��	z�MjS�N�K+hd"nzE1���c��~V"��	�tb�7�ig���;�K�l��}�~t��p�Y��E��.���u�2�B�Ӓ���?��/z�o��ĳ���ML���`����x���n�`���oG��vZ�p[��&5["{[�;�}t��Ӻ����2[[�Q��.n��㹥ل(���45�<M��tE�;����B�a��Ƕ�* pi=�"�����#��Y�4�ƁLM��Fv~���?�I��Q�!���A~��5X���\R�)����@��~ej�u�b܁��&!;���p\�?nu�|^�l���
� ��sb�J0G��j������Xi2j���iv�<�1��� �xc�ME`� #R��H�#�`�B��$�� }��zڙ�:I������:^Q=oё�Y^s�J�{vᩄ���j:�LH�]v[�1/��1�<���d�8bw�Rܔog��q\�#���|qm��_pP�&���i`T��W<�A�=�<�{g�����'÷l� 7�QU*T���j��,*AkX���5��}愺<�;�U�B���r��?s��t
=[<�m3��td�iOjZ������� �cVU���z �G���e����[��5�=��7�*��.r0����B���#�U�臨�*����0F�l��nz3���
ha'DA�7+$����NkK1'�3�{���������w�y��%-��w�Ui����e���dA�tr��j`I���zZ,@KoɄ��D�f����h�d>®�78���^�!�@E�}��P2�P-{�D>�������Q��$�؇s�:F�V���B�,6�����2�5�M0=S����cm�4�Y�%1�:s��&W���5d_d���2��*~�X�N1wӮ�pS^�rO�
|�'b��{�Kt m�ko��M�&�r��q�-F���5k�W)k��6-��&�]P�Ƹ=�S���M[Bd"Gj��F�q�zgc��\�
r��ǕB�!<]�w��RQ_��g�dB�݆U����U+m5$�9(� F���[
��G�;
�9<';��/�SS3\���M�%���/���$������" �:�2}�S��(��o��i�V��-`]br����V��?	�LR�t������\L�3���6j�-����8TѮJ��_y�b⁨�E��+��.�>)����LC]���dVP2�0jJ	-���Y��G�xI�אz��X>^�z�H�ľ�#��#~�@�Ш���V<���^$�g!%
VJ���v�
67�\7?>���0�#X�l���i�G�&��g0�OvA<�?�\#��t���hB��h�o�6uL�����_xh�ce�+EU��^2�6��F��������Y��vf��x��e@�)�d�K��D��7�Y.�"�����jvI��f��_坤eAd}�I�afw��>���G"�3�
�����أ�@%f��nUォ�k�7�&��g����U>3���������7�1�����:]�a�
�}�xk��,��LX��t�Q=f���j?��8Q0�D	��i]�^Cxʥ80�r����T��2�_/�T@X���]O\GLj47.z����h�����tA�`\莕�K4>�����r��KH��/�*�S�a��䲳��X�"������KÑ��;���!�6[\������K�R��&��:�jvj���F{Q�㲯8���fF��H�� ��N�{D����N���	���co�;������P��������ٿpb��_Ek�j� �w�.�8о}�)>���-��Y\Y7�<%[J�e�S7���BZJ�m�`E�H��1�P�3��%�3����8�j8;:2�jw�eO�Zz=��QQ��W���(g�p$�+rx���E��"P9����t�١��_�^�O�1���9(97� 	�I�n=-�i�q/��It��-�����L�'�����:�b��׋�C�)
�E�6t�b&(T��ɏ���9,��)�l&��m-,I�^�H�$á'T<�� �_{ hE��x��:+2M�����.z'�
�v��Q�j�;w����[����܂~[
��e�U�C�]��u�A����Ӡ��!2;T���2�	���<��������t��j�ZA�bT+>�H �l�z̑'3K�JCD��������Ԉ�ys1�F��)Z���ܬ �d�w��1� �5(��B>V8@��`�~N��)��-D���!KH}0�k��"�g��g�gSj�gMó�`5�R(�t��n4��p��Ew��~�`����h��0n%��v������_���"F�W�h96t��i��b���p�W�Q�ѧ�[ίĨ����5�-��Y��uY?Y,����a~jk/㪝�/����c9�>E���wh���@f�8O��V7�j�d���3�������p�����ӽ=�짨�Ҫ����E�iv�'�4C����V��f!�Ig�we<Z�3����|1}R�~�	%OH�剳e���?P�=V�׺_�k.�+��c�N?P+��f�^t� `��w��]( a��T��
�>qm�j9�6�d5ʤ����Y	��E*�g�
.�uYg����F�W�K�7�R��;Hذ\��?�A�"����C��a8MD��%�D&�/tDo��)w�<}$����u�+芐�W���;P��S�g.z�{S����ƅ}��M��;�:�i2#}ď��w[��HI�v�-���)��ػ���[���
	&m�/��T��bs�����3��v������]�o6 ��n���%`Rb�V����PB��!��1hm9%'�BIGi�^h�b�>&d���7/�g��-�O��\�9����z�M��5d��];[�!�1)��M�{��-d�L�D�J�f;�م�F��q:�c�M%�4q�X"S���\�%���r+��6 D�(�"̍ZWk��A�Q��O�[<�Zڡd%�Lrh�'ʺBSa¦r�j������-;��%@�9���<��M�N��p�3Z���� 3i&xTzo��ݒ6��$e�0�=q<k�߇�iX�=Fbh��(���'Q%!J?��9U" �5���cuV�B�ȑ��/�|�{��ẁ��2�{(������&;u��l��}&��[kXl��h�d��O7볍�~�~�c(���͓L�Bs���7b�B�ڠ}��`F�(��,Ƽ���\��rM8A�%���J�t��J�ث�x߫�5D<.d s����ACt�B�����嗖��ʬ��Ӂuv�D(t�l�^(y�"Pm��z��d�T��%+������rq$v�Kk)�@�aN�N��G�	*��8U��'ƚ�ܔ����D��L�W��B��~	���]�#��9�d�}4��,S5f�:S�$·��0]���%g3�@�5G@(�;	�d��������-���3����466cz,�
]��3��z�1��B�A�#����/���n*7��m~���`5H��&kp�L��V���=�?����b3i��ka%������@z{S�W�bϱ�}�(j�Y~��3�{�#"F�3�|7`u
��e��J��g��=Hs�0�)ox4ԤA���^�A�P�xwh�m�iQ��:��29���=���3e%��yÿgzf��[ޱ+.��?m_�m�s��{�ړ�p<]q6���Zr���I�� [�%!-�蕢�J=@�a
�W�\0	�M�E��
G*��ŀ]��pPQz�/jK�5U��DTsF���`��'� ����]��~��	��ʸã-���mb+4���Q�e#r�t��K��@�CI�}��NE ��S3t�X>)�]=|���yR�c�a|l4U���I��y��"��P��^={�z���no�~��c���V�)4۲�ms�wB��H	�%2��d��#��r���	lNXȱ��p�2Eگ�mX�m� ��6)�eO��̲��)�>X$3F�' �%9��d�Ў9u�5�r`q�J��+���J��w?k���'Դ���o���j,�K'N{6>91E/��M��̀b�g.���.��I_�u)�dRԇ�s�ɉe5ۓ����j�ӑ�Ri�a���xܶ�X���fHm�w#��5^��
�� �����@�ӥE��\ң��tѐ�-�CHq�9�L�v&v�0���"?�M�wǽ�d~֡ȗh��[�i#>K��u�'�~#����d��`C�H��m^n���
�z���@m,�NtJC zޕ,hΆBB�0C] c��spu�9�^����d7�1V�7����xh����������N>��"Q�6����n� �o������d���R���>���j��������}�g _����ޛ Ƕ��1��b���+�Z�|�m�M�J���TYg�Q�2�����r�Ė��U�3��uf�G�hĠ��[� �Z@:�xPp~��5B����9��$�^AVE�䴳���0H��&�~M�F0t��/]`7�o�2|��z�[�L��m\��da����K�p^Bb&7��'Z61煄������[)I��B9{Qm~j�ݚ�>|���+�op��k���1��
ۧF�-�e<��&�� �H�W ��n.v�~.����Uq���r��oU�����N%Gx�� Yev
��s�����o��Y�� Wg:��ֹ}!�+�K5��a�k�Z2�?a������_����Y �z��b�%m.���i�$��ק�0(�ɲe/�a7����.&O��3��t?Fm/��k �k��@�@�^�op ExX�M}j��F��
�,�0|z��S���b��f޽Ye7D�x5���/-�٬rwKu�������&H����@�rڻ��doO��z���x%��E��^�/�����+��(b�i�un�DQ�ᖉ]$��������d���ٔ��av�JU>_������$�m���Xd9�ʎAOr���~�JC -���u�����'V�!D�\a׏��j%��[��̗�ϓ�N������C�͔�vrM3 h'�)���v��M�~��)����@��S��� ��ķ�k�t�⭀��(�H�j)��T�����_�*��)��} �_�0����o��!K�y��J��.c|*���N����s8?���,X\`'Mw��;uǨ��������-�o�����Nz�Wa*�����e
��M"r	�ҡ^�����$V? �H�NI�lg�a��k�[�������ün8ӧ�n��pn��������(Ϟ6�5�[ek���?MbYN��9@�0�g8*�"��@B�V�ɇ�X��MÇz��s�r��3�`��3y���7��>��C 7���i�{D]�O��^a�0��C��%�[ڄ���䣍�t��g}�hD��-X�?�s�*_'Xh�����9�́�=�)�Al x.��mus�6|,���&��k+�.�E�Zk�G��Ѻ�"�Q�x�n�f��J�+�c��ss5^��p��dOȜ�bQ�㎺&���y��9N�e�N�w�$���w�J���:@`0��2#�\���|F/DU�ǿ�8���N9p��G����z!�ִ7��H�2���i?�z����!�!'�_%Nt���L�'�M��J�'��X��&c�ۧ,e�3�sA�u�\\ߞ>�'}�Va�p�����;n�'о�1����
b�xFB�_jFI�����*]�m���tٛV��I�W����M2h8IM�.�R�`7> ;{��ո���F�c]��t8K։�C���#��	*Y�k=Na��?b+�Vm2Edtb՞�fX�v��w�b$(7T�ⴘ~�	JŘّ�EHz�
A���|T��Z7y�Z�}� �gɹ]+e�ҁ��*���*�A�� �����(_*��5���J����	�İR�-T ��@P��6'q�+{��K��Z��v�B���9X�En:\&��U��/�|�(}�3���=�C$#N��'�R�褫�V�4���Z�tg��1�����7^c=�8�7	ң?��v�w�O�OxX����3.��=�X�M�ې�GFY�A�A�*�(��hMb�������Q��)U�dQ>NÅ�U��Y�ߕa<`Ɂ6��rѤ� �q�l��F�� SxlҶ1��I r4��}*�S$��a����D��g��r((�3X�(�����F��?�tcAPD�����!z~��\��gN�Q ���n�ޮA��Q���k���������q��(�m#��w�b>9/S|�� P��\I#e!�$@d�d]���-6���@	��i�I��D�{ӣq��1�z��ʗ%>�o��<F>r����P�\Ԙ���l�Kx��tv8�D��׀�XZ{'D���A��*H��<X\�)����3��f�u�l;	���Ц*�x�*���O��]��%�"�g*F�E^�b׀U�_�]�)T����4h*h�$y�P§�>­��İ���Ĩ�1�a��2A�ʵ��(΍Lۦk�t&	�)��Z��325OƁ��ȥkk����	�H7�,q�c-�S�ڄ�8݋�J&�����N���s��u�e��oa�lW��RЊ��*�ֺ?w!�7����O���T��M��Չ4�����f�x�B�+3f��,��� �<	�Jy`������6�/�$o��*g7����AD��AHe*�IN����k�QC�w���@>g�9��r��]j���	',�r�9�h�����iS�S�M>š�Ť_�z·�Ri伴�L�X/S��C�h��7������
�'mĄ�+�a��!�m�ա�Ԕ�/^R��"�(�)��L`�I����7��a�~w�^�o�X�K�Gg�_�|�Á�!Ua%KB�y�p����:��uʸ�ގ*�p�?E�'6\�؝�q�/NEa��<���P? 68e;%B����DHE�^���j֮x�i�F#��a��k*�|�=F2�����ڬ�q��vǇ��Z�����)}T�f�����l�_B�6 ��9c��[T����++��k�ى���^�膕7ZJ1@��3�T#hC��~t���A0L���p`"��z��҉�0y��'�~d<<��(s|/���Q�@�Ր6�w�� �Zc���,âM�����4*�_����b;�%"lf��ط��K!�Z�P�b`�_��P%p^���j�)�hpJ�U��4?�o��z�W� Ol��R?����[�6����)��a���PG5�O�X�Y��T+�)���=���9��ot.�\[��q�mY �����*8�u M@��N����}�Z?���2���Կ@�C������� �7�F�G�U	�r�Jo3�������PB��h�v5�������@;�_�>c@UJ�-˺�<�����p}�`�E8��mk��� �9Z���A��K��4A�섲�����N-4�dF%dU��a�z�I�T���G�V����I0�5�۬�F�_�b��D����J�8Ii���4�_B�� \�e�U�[
���.#�<v������~�/��<	Y����<|�ش(E���|Yͫ�V9kw�B��@!�)�B_����&�+���wp��:��}�퉱�ߝ7�ckv/�B0�gH�!���㠲�"����OT?l�4�_S`TثG���am/3U�j��3ҫ�G��b�7Z^��JGC�r�>���ڴnK+r_'��#��B*��RV��J����2-��=�3��O�p�:�$#�<Zo��LIo�+b��4�p�q�����6i��:R�� 2������]c��cM/9� �2���3� ������%�n� ��ůP͘Rȝ^fk �%���ǀ���r��og��A�Yr���cOC�c��_�y��L��jm�q_5�dQ^�O�mYkWs�X�}B�c�]���0�!��t����%��v�n�p�jL��b�����f�s��:T	����*Zs�Ȝ��vSd�*�F�!p�^�˩�s9:}pa
˒08�N���׹����k��C��o}��!}^m˃Y(�]����/,�����L��NR7.�!d�يp���Գ���ZC@C�k�a|�C�����X�ʝj��$|��ћL&�d��`�h k_\=�7�P���(+�l�M}̈́��i��Cԣՠ��n>��P�?e�g-08����j�f'?X�b�7�ڜޓ1��8��(C��?5��� �2�.`�ó�gA��������Z�I�����?f��;�'����6%�Hi�r!B10"iQ�KΝ�MB�i?x���p߷�B�;W|4DjD�;��b�pl2��#Lƥ�����!�>�"���f��g5����F���v��oΫ"��]|hqt����qx�Ř�x�J=a�@���ח^ؤX��>a�&���Ҿ����[��(�l��%B���2�3����P��P�
q�/o�-�x%���Ѩ5쳞{V��� D�;F���8�g^��ݨƸ�b�x��O8�=�k���J��A�T�����w����Y,�^Ք�D�/�
$���-ϯD{��qBׁS���|$���XqOA���]��ani�	gH�j�=�<g���#���Q2�,���N-��׾[:8�x)�𬐗�X�X�fZ��������Q^�:I�>᧔p N�Y`���sn�zZQ��Yg7@�iQ�-����bn�_�0����rpz6�r�X��^,JJ����av���8�l�[uN�g�3X�S�J:22:�:cE� oj��-b��n�<r|/�@L�C^��a���{ptB'��(�cȬp�L=���W���L�xk��ZC��՝�Җ���Q&�ds�T��׊������Z
��,��Z��D&2h��ڻ�����LT�Ao3'�����9L���T�Z�)7���]����+O!ʉ�v��	�N�����[l|SHeʔ+�s!%��^v�9t��vA�pU������XT��pb����?$���r������!�v � s~��(�>����B(��W���<�WI=O��i�E����Z\���鈜�bP&���S�Α��'�*��w�~
I;��n�3�zNS4�ի1s1H��w�b�J��bӝot=H�0,Q6�R�Ϥ�y�q>��Ȕ��w�q��,��F�_����2ݚ`{���<�R���2<��M�uxh5Ơ]f�_�c����u���C:�]U%X��@�SW��e8���2�[}/�ĩk�de��@���ۚ�>jp6��u�%��qZ`�3p�M��Bi��wL�u)�ID�S��j��
_�w4�������pBTfԜ��(t��q�i�����~D+�����5;��'}�o�vhIM���>��&�7E� S�b0�ΈI�Pb���H�����!o�Ώ�_�)�_!�?$9a�-'����O�u�ai�C�4�U_~Ҭ$�*��j��s���tO���d��+��5X��a����EP���U%��
v'Z"�X���zb
�O��aꌷ�n������#Z5	r(���Ev�A;�Pp�~�H�E�����&g��o�$ �U�a�-鴺<yȓ*I��ۻ�)��T�*�t��ڏޗy����|�o)��"����a���lM,��p��G2*��>P�e��9ȓ(��]�]k�׋x������:}��V}č�P����������{�/��� .��p�չW����o��7�[¯Qjwh7E��I ��N�~�H�_Z�V��SL�����s�ᅻVŜ��w�;6��Z��+i��K��]�.;���	G-��UbcEL��(��4㲫�8;��yK�FX�#f�x[�/\8�� �y|U��u�R�ĕ�T(��KD��{��=�r�d��JW/#�+_�^f1U�Z ���c�Z�Ak�-����x{�!~����_ks����o	ak(=��jv]SC0����bصs@��w���<���&���|��B�㞇C�.��(!���=�/��D�>>(����:�7��2֓)mB�F``��m���XA+�G��GV����\�Q���5���#x���q]��߭�6s
+�L��
\��瞷�.<�܈7����C8��H	�iK�9�Ńְ��s�~��l�E��"��ea#�����F1�5�Ee���=�<s��Y�^�m�Vw���X�d��x��d�:�L��������el�`<۵�Y�;�[�1��7D^Rʟ/�
YӢ�Z�)J�!u *	�Sݧ@�U�u�Y�@�k��5��@�B�c����6�^qmv���0a����밋3���҂���MX������5?���.���E�@�=e��U�v�0^?S)�vF�����o��v��c2%��P�U�5nE�@����}ڙoq!�����μ�5�lߏ�<5-�ѽ�$��M�p�|f�C,��+� {��@?�x���>�#�t�����°�o�[�*�Oh��A}8�f]�! v|pM%��<�)��v���<?)�X?(�H:3�K5HS��֗�Ԗ�Fcu�]W3N
�0�G包��*������P9�}�u��3Dc�<^�c�ݥ&{�a�~��c
#`9�q䒫0 ���,Ᵽl����bC�n���HK<'A]�8���w�]��P�uj=�B[n}f�7�Ů2�j���8RK���3��{r�
~���J0ʏ�
��j��p��č��M�A���"o@|�B�t�A
VOЕ;��h���3B�2ZP�D��a�1�tס�A R��gs�W]ꤜA�忪 T/��6.!��b[6̞'��+�f9���K1�-`�W�5�~�O���u�Oa��E������5�X/�r���D��Av�3���N�������Ma�[^-��M
�QN�]�Z(��8�2,�u]���n�	'E9Ŗ6��}Q���1VF�B�ӌȭ`����/��}p��s�J-����
���ü��O��(�`���Tja���w���������w��97�f�oJ[k��U�	�\"-S�����+�4��0��g���l�A8d�
Tܢ��ѵCi�3cs��aX+7�t���眞����4Cd�>xA�T�<��v�K���1p�W#�Xm�6lU�/��m� �z�~�B׋Z���>�[7��	�^o~a��%�kJ"i��>��T�,^�@�R��HqT�gi�⎉汏Ђ���}G����oQ�T1�X�@�k���׀���A�n��l���aņ
�<
��d����X��	cȇ���\v��է�V�=���G����55s�+�@`>?�17 M#{�\���	u'��E���u�
����	���P3*��Ob����c�>c�]
�T�{�( �y�2��aK�;g�I	��3p�fX*d�4�%v�����y+n��4s�̢�u�i���+\�b�E���z�-G��z�h@ �~1�����i��2�t�MI��Jk��N<��C��O���k�D@o��î�٘?�]ٺ�Y^�����L�{Y�\�z�'��������D<� ��>�u��Í�CLa����`Y\��-ex�[�����l�NK�C���ߙ���.�G�kw~��G���S���b���[Q)��IX�ߧ_�JA�!(��w1�\�]�Q��N��C�E�<�\"����>���WUW��Z��#�����l����>�_�VQ+j�&�O�h4�;̠�={ĻY&H���Z>��?�pT�1�5W�&�d�:޷�
�"bm%5�{��n��-�u��45q�lµ�`A-���S�x��ճ�pp�/3���>3���U�y����<��'�4vi�l�91+� Q?}4��{�,��&������n��|�`���C��`d��,c�s�/��b2o�� �����Y��CI�CF��&jx�F�J�H8�JN����(�n��+iW���>����k����fWI�<#�����¨pq>���q�@��ܴ����+��0;V��;��d��6l�&�[TڽΕ_�-�+Eu<F��f�J�9���Sm��X\M���V���`��y���g�e�sQu�X�g@��Qm�ч�!���Z����B���H�y|�O���	�q�1�G}�b�p["+o��PB�p����%��TR ������t�_0�W�e�s�3X���/eK��6�܁�zT��Q�KFE��Q[ �	�!C��!rc�O�)��h�[�=P���i�~�~��2�$@e�Mq��K!�#�g^v�pc���Z��?�?>i-l_��D�J���!;IE*���sc���Gh��!�.�'>��ѡe���%��"���|M���ypF�`�ΞU�ѹ�%���@"}���<wC���
l�I��"�9���n.�/��
�j��Qm�ŭ&u���-���RkK0mWX=Đܾ��\� 3t���\�G~�o#��M���iU���� �5�-a�/A<XV��#G��h0�~E���y��Sao]��p��Q�i��kئ�l`���9*�Սk�9 <;�;09���ɘ��qgqq�Ȇ��S���zդoV�V��B���҃�����%�&��"<�(�$X���o�"�TQ�z�W��1�}=~�U'�ԞJ��r~��/��S�<�ό����Ô��^�|L�;��=�V��@�A�˚koТLw �ϴȆ�����!`���p;��=���"���ga����\lg+ktծԃ!����Chm6\��݊�����6�^ǈz��[[�H�/
�1�$��>8Hg�&S�!+�{�֣5y��M�Ȱ&!��0k���������7Z���t}������%�%���p��G�ط~7c�C7�N@�(��w�U�Қĵ����8CU'�j�U�+ ��L��v8*�[�1@2H�^݅m�`M[�:I�{���#��p�)k��J�n2���ǎQ ��6����fB/@<C������TF���|V������P���s�b]9y?�j��˾>>���5�xS,J�m����*��nw=���K`8�n�)rC�w������}��#;��8���,�Bq�w����74�C@B:���OF6`����l��x���^��:Z��\�Rs�xhZ�Cv��w_���,��A�A`s���hTcE��Ԩ\ aa�p'r�����a�pQ���V\]QY%K!��W��b�u���ƞB��̳?��LRɐ�e>�rx3�Z���!)�A��ȮԤ2';�e��ٵrV�=���a/�˨�S��n�z���|�;ӺN�FMO�c�	��#�;��
3;��`��K�U+�o�)��q��
D����O]sw˾ʹTY���ZH�jp��wgmpob��M�
D�_�rjVUTc.���y�S�2��4-��Qht�ؘ띋~��f�^v Ϡ;�;,�V��$U���Uӻ�3A2e���1�����-�ШG�hX3E�ŹaI�j���"S>����|��8���L������9>Ф,3t���7w�K��T���r� ��9`�,��c�8	�����޾.����j�0A�-I�,�]�0��Ԁ]�G��<
qGq�ƛ�z$v=Nxo]aAuu���Z �lj�������oT^�`_�m���,��㩅�U�������z13��!ŏ֮S������Ε)�S��nAe�q�8��r��������=���[_%C���1�
��w���xŉ��x	�����
�E��.ʠ?�1?�lJp�кn�K�tiFԹtG!=?"P����!�UY�l 5`=�R�t�k�l�G���HYOՓ�}��1©�m�#^2O�&��e�k^�d�zN.��f�}O`��cG+��	Z��/:"
������� ���qB�Z�+i����ʑ��l�>r�h۞|������΄Hq�Ϭ�]d���Ûzm�{�����w��8�K�^�kQN����u�2_���=O�0Sנ1vg��}4����7���� �p�1��
�L�>��<���o$�!��d	�1���1e�'	xi��M�1v�#�>.%1��5 �Yk�!r������#���Ep�3YŜ�QC��U9��%�F���R�#@E7�։��b�`��?]��L�:��]�.e|���d���� �.�`��a�{܉U����d^�rñT��I��Fr��=q��wܴyn_�����6���BĊ�����E��b�vB��Gu���fe/*ӭbaVd�2����Pq���d�������ΡY��3>,�@���D�~���� ������J��,7���,����c2�'�1�U�iv�Gq,�+p1[O��v�"
Ld}MO?H��91�.����.�O=V�x1!7����I��0?G���I������퀷�c��Ժ��@�rd�8SN�ڗJ4���C�62������Ӳ+�5�����W�'�9�s�=A��,������A��S..uz�Y���p��U���<�ł��h@�@�}l��L�-k��"�E��c����T
��s���(�y��a�`��N	FWEuou�xA��ԩܼ��a�����@���J�vx���=�oiyܛҾ�:ȯ����~G�`z�-�2��$ReHqđ:�pH)G
�dQ��3�,Y�����lJ��q�����7ڻ�����Ȍ�)U}��:gO�*4����y�'jJ���5��HC���{V�s��x)���$�?kC�C�r�%v�6�M���T��̵��Ln�@�7H�����DD�S�K��Z4
dA�ٟ�����(��Ҵ�"A�/������ɘ�0/�*=�	gs�k����EI�-�hlZ�:JTI��NydF�$@<��8�h�t3ˊ�g8��јD�X��,����"K�O�n=��Iþ�f�i���_}���ۻ�������{<ؙ�!��Mxd#��0���h}��@�Vlc!v#��2S>r��t�g͜0T~�JNQH������� �(�u�&O������-�X6����R5(��&j��yY��z�.������:k�|�$���x�F��.5�óoa�p���"�k?�5u�0�zbY��1�FŋsAtm�b�����H%+`ÿޤ���JҀ��H��H���L�jq2���`�ˀ���W��:�Y�nl��r�2�(:��p��5�=͟?<��?��_�Sw��P�8�"<~�䕵 $��|�y`QM�,��k��fG�D��o�}��O��%���H�6@�X�� N�DHσ�z"$g�Ʉ��o��y�قy\#�B	�[�W7�9��+���jl��0��x����pמ�9;�� ;�P�p�����->az�R�Rq0�"�3Ԑ��K8?D�)e1���O��L�M(�C�_����FF�L��/1i36Kr�)�ESJp��dLprn���<�]ފBd��O�4��B�{���tg2�h�o�֋YE�%<�z�\n�����	��ܷ��P��'��E�2þ�o1YH(�r��a_RUQ�Pxý�"�m�������&�f�%��_�2��hV�h��Ds�����"R:IfJ=�N����ckmθ�/6}J��j����3�1���<�����֣	s�\7��PW�\�9�Ly
���$]Z�$%8�d�j��\S)��b�h�ֈ]/U��	;WԏW/H��h(iI�x'��f����.C��2�
��C~�uhxY���UH9nC�c����듍�	.��:���w��c�o�}��� ���P����CG�q���u��_ۂX�XBT��A,�✑�[fh�f>Vj��4�n�g�02?�:O��[��l ���:�6RRK����u�
�ۮ�rjz��sR]���UD!�
�5��{f��t����K{N��0�3pI�i�[�����	���Ĥ�O0%����Ψ+}�`���Q�8������F$&~k�7����ܘ�x��FQ�C:�g�_lhV��s��d�� ����3꽧�c��K�:����[y��V��s����J��E�a���L�ڄ
C�g0���|�(�w��]�rua��P��F��.��8�Z�M28܌�����}�"�SAU��.DDHx�9w㓘t�e;��]�N�3g����G�Y�H:��� C�޾P�6�,ۃ���k�B	���ˮeΜ�U��'�`��&]cj�f�k2�)��B����cڣ�G�A��,V}���A�:><\���Pt�i�V��|�� ��gZ/�!���!��՚�b~��@`U���d `�rߓ��?T�O0�s�MZ?����rҘwuK��8�����&�n�>�����6�!�*����dF�4�٠E��O�~�?����+栺g������H
t V��=y��/f�g��<=���\������K��N�q��6
���e�9�ok�FՆ(@'��M����bE�dZ�#���Nsk�әStd��9���ԧ�3�C3��?�$ �Q�!�t:��)����c�P�]	rnr4���{|�KQ�+�N�|���'���j��W����Q�@���B۠6� ��{nF8*����u��nZ-��!�_��#x<��w��c�U���^8���zn!z��s�_�"5��I�H]1RQ����?@���/ ��,�Y�8�#0�/ٜ,܌��:�|�F��ռ�N%l�4��/�"�7+b���rǒ�C���(#���Dw<@fQ���~��
��޵�H���"�]j <tb�X\t*���3�i�7A�(�е�(w�WR�s��-홚��ISQ۴!u؟S��P�N����,Ғ��5�j���ueΧ1<bg֬+�o���Z<AЀ^7�d���4d���~�o�$����B�&�!��mOS��qb��GQ�-�ED��g�<C�������T{�)�
ߞ�E�3��ҿ��@����l!9��ﮯB��q�A]HP�/?�q7�q��Xf�ڍ�*Ttz�!��S�����[&j-M�����Ѷ��r�ez��v���D6�b#5���J��E�Xv�0Hl���� Z��������5<ؑ��iw����V�d��Q"����3N��sa��;���P����+�� ���U�u@�,����,����ui����Ox޲N�o���� �¼/��bi�# �t1��5��W�j@YW�ެ�(�<��Z^j���L���؉�Օ�As�=tR�gXa3�jd94&�i�J�����M�G�jX6���.=��f�P�l�; s_��'� $VnK�l�H_c-���P����b\lK&��o����2w�?�:�me���Ak[�&:SQc(E��ؙ0,����E��!��PR
�f_�z���r� &a9��K��|�y�n��|/;�{`��?�!�R�ioӸ�"���[ؖ�� �,���S�%_��K[�-��#�P�-?��k��o�ӀL���F@��c�$��[F�^T����v���t��^d.�3�^&K8-���H�b� �Y>�sP6K`��^	�P����y�L�Q���Jvju/7�B�┞h4R���KpS�o��2N(K�f�W���ES���(�ʎ=%U;��6�	;��k">o#���:�	���e"[��N�����
pP&T>����K�M� �?ox�&��v�o^W�z�&Vh��{K<���
��ZZ�\r���z���,�p�Y��w��k���f��M�a
�Q9��Z0G7{���t�v)��j��=�,��\�&�'���Q���
o��m;��U�<-�=�@� ��y�7du. ���q9��\%[�Tx��hEX=���h���@�L15��w���+��k�񯉻��l��V�jP.؇��LT���A)�Q�P��5:\�����=�;~|peI�_��X&����H�V�@��/�CCFMS?�Cv|�	"�����Hcc(�#�%�cqHK�WyQ�d��R�-_�Q��[��2?������>_J4�NW�U
Pw�X�М�"�6���3�K׻qI�s�[��T���g ��y��C}�*z���D{[Th,0���rWߧ�X��0�D�s�Q{���l �+!TY��L]����|,�����M
=��%<2�ɸQp���jB�{Z� ��[�
�$�*����B謩N<�\Z��@/���S���^��K;��abh�[Wg�[ZEq�@X�~�R@� ��ʦW ��Ц2uM��	�~l�(�ſ��ռf;޹QA�:��m�b��� ?���uP���'=
��('�l�I.������_~�k0Mhɚ^Btn�z�_�ǻ��^�޻E�������A����o�=d �չ˫K^���m�Tk�	Э�[��K�fjuuK_>�o3pn�DL����"��2]��Rlr�s�nxAa�U�nf���OP�V��Tjo�0�%��%�����$����;�5|�|��/�T���Aq��QD�%0	�j�q��nA���5�a��2e�7�!&n���P6�?�VbU��i*��(~�"�U�(�6�@T� q�tLND\�*p�kZ�c����$m��-i��֨j."�̣l�����ɕ����o�`����1�'ە�l;ڼ���ǔ��^'R�`>�6�{A�����3
�պ*5�I;'p��'ߝ}[%J��~²s��G5Ŭ����L��K�̡fꄝ����$�E2�����B@*ܡ��4��v�]x�0l�Ĕ9j}H;@>|T~�� ���-�e�����]��VN������y1ƠYO�|q�:0�W�ZPuр�]�_�Y_����jn��0j0�A"9��Ueܛ�;'��!���kl�Sn"`1�	��E�����}��6A�\�-!���Vdې�E�IH�Vi�s�0y����e˶��rx�,.�"�e�ْ�+I�[�m
o�ؗX�?�jL��H>m������F<�*�籐�'O�#MRM�2]�ˤQ�
�+r	&�����H|kh�w��>�Uh'|� ��n%#�_0*��3��i~��P:&�&8Y(�YOx@4��1+�6�~p��M�^� 7��lvö��m��>�_[|ۅ��F�+Ywo�����
)��Z�+��LiSu��DP�K��s��2�*=�y���UmaV�բ�>�xd k�0���$�����i���pW2�%+�=�,�oduB\oj�|�����}��x���W�UK�P9SgTl���9�5�oc.���J����e,�_�k
�+^�9m�����f�7��5A�4
���R�wn�5x��b��5��������wm�C/�O�v7ˍ��Ҡ�3�/�K8Fg�T7h�Rc��H�&�q|���Q:�ې��#�3�Z#mc ���f��f�[*�����Q����5�0M�]��ϸ�\k�L4�i��5�Q�K/q>��u�O�?��KT��qIF��o9�B]���C�z��<��)��k�jgi�d�[���: ���T�K63��D&2<�=�'��,�v�r�6a�gLR��
�����t�ER��?p\���|������]����{���v����Y��<#"�F�(�	��o��kd����mE���[�������:W@BE�ꤿ�)���y�];�@&i��U�O��e��J�}L�S�艏�,��[ ����8���/?����⿘O`���19zͱ��n�KFH�����~������m`�Y�蔅H��K�=u�p��NIP�=ݡ6w�1u�������-] 0g��o-�D{�"Ԇ4/4ǐS�W�Lp"��=�)��K��J��O9���~	#8X�K ��鍃	� �	xj@���>b�������%��2t�t��f���;%��2#2g�"H4��;;ߡTC,:6&ιW�Km���l:���p�DgGZ�X�m^��'2�X�/����]��'�$�>s�:��=_I�f�Ҵ��DX�� �_0�� ��!Oo�e�6����K=�e�R��`La�׆���@prJ�����z낥���s����)�h�r�΍�|e�@?wFg���}޷�?��_�ʪ[��Y�8�Z����~�MX��M� �/�Z�cc�g�����++zqW�!2N{�ꔤ$Ii��N��C*�{��[;���Ƥ��/L��#m8}I��П��7���,�V�n:W�آ&��nŔ[��|�4���U:���^	�)#��ɷ�m�>{����F�WU&��+V&��|b��ė�F.�!֋��c�7%�-�]c��z�tZZ�t��F9�4���	v��R ��rtuxfC�?�'���B�er�\�!��k�	ʃ�g5u���˻̴�����ֿ���ȋ�O�oa+�qo6��./����}9w���4P�1{(l��M":�t
�����B	F��շ����L��.�����GG܌`�]'�٭�G���Ӷŋ��f�u�p���e�q^�T��a6�#�^r<c��.��xq:�r�ߘD1�&kS���%����e�>�Y�Z�(s�^�<�DZ����Օ��ylˤ-��-��,�Im6����{���ř�����Sh�9�I��p���3S;G�DT˺P��{BAa`#�I)$�A���Z-s���r\B��-�����~ᾓ����}`�rR�eV�I0���;^T����U��N簑k?�A�.�<w!�7jO3��*��SU�tg@le�᭭��[&(��RXJ�)-�v�h"��r�1E�u[c-��+_�Q��4s9�d������8�q�hM��6�8'�\�@'U�	)��KšU��q����3%�r��{{_j���cƋe��,�k!��Fu�ԗ໅��ܽ��T�v���TI"��#2���()"d�,k@U���R2�{��G^P��t.̞��0s��?=~�@�U2H�C�N�u<D�e��~���F7ӖAR��c��'��U׿l�^Tk
"*����=�<���k)�73�>�W.mQD�VQ�
ҚQd�.��e)9oy���yu���@M�gf4��큣��L�w6j멞�eh��^�tɤ�]$�,�e*-�-��pPBy-�Jy�o4sQ� ��#�͵���A�޴����m�y:,Ea���_�$H, j��8En�wu�2�yR��_|���s���j���9K3�:����Y�B�1 ��?�N����֕Sv���hE��&�J�\�E0���nSѶ��s�7;L� �(.����u$�:��(�nj�B\5��|^:�J@ed޻cBCI���Nj�YT�CO�D7�}ʳ6�K	��Y�/_�j`��6�.:���p�"$MY���x�秱dM�`��o�x��ȷe�����3e�	%���|�͟˭:!�V���w�	iY���%f�z��G�@�a�L$�"6����I���@a*'	����8��݅��@zק�%��m�F�̖k����	M���w�in�����Rh���=���g���Z�a�@��M߱�l�uX)�B���'a."��(��a�-�lN�b '�s���Vx��2��KH����Md�L
�g_|��)1Y�V����K��?��&�������9���7�O�u��#�0�Q�0�u���wѽg�C 6	٩�-;��n�O4H�84�ҍ*d���$b��/Q�Y�Z> &k�T��s~bn���cz&��oǒ�ﰄx���E岣�^sZ')㢓[�9�XƠ��=��mܺ�,K�C�p�P�I�)��D��=��9��nE1tO~R�_JԌ���
��p�
�~Ɓ�{h�'s�z�a�d�:��u�o����+Xưr~�g/��/j��쌙F��;����M�n�_�G� u��n��(���ҹ��[J�}�!M�e��]<�)Vƥ��Q���g�o;��z����?$��AU���Ə�Iá?m�]J���3�C�Z�V `��+V��{�a&Ū��E?U FP�f,%�a.6�I�MB��	Z���8�bm2���I�A��̏���Mg��@z�m[�E^�2t�[#\��8���@��`ѓ`�.F��.i7�g����n{�o|6��j�X���p�.�}���51����l�Mkx�*Io�l!4�Wz/�����>�)��p"Q����� �R[���X7m5�O�V�1$r�΢
��֩ҵ.�C��M����Vۓ��r$p�̥78]kGhE|�;�!�6Ya��	����h�%�Z�<�
�z,���&M�>t@ͭ�%t�F��L}1��n��o�J�a!VI�0����z�	������'O[zɥ�d�l����Y��t�(ā�j R��橪2\����F����R�Z�$hH�����#����5y��~�N�eNwp���7%0�5��E��dCRVSwn>0����6� ���d��j��>�<�Y�+�T$�}W�	@�.�kkz���MhPb�A:���� ��KK��=�n���V�
\� V���c�����"p}@�a��IY����l��bY8/��z܃Cg0q�}�nE�H�J=��4}�P�2Ai�A���	GZ�^�o���\ߞ�W� ]��Zv�r�[�ͅ����]�f�v���e�v����5�0�-=��겥��Uҝ9�p�fhjq3�B�"������p����|���w� �;I*�	�g�DWե�j�]E<	��/k�
DX�����dW�{���p����Q�e�vF���'G
9�τ��}��΃�%Ky�$�h�#a��9Db�7��'d��93
?�s��qR�b/��3����E�3Ǩ�Gl��`�JQ#�V�>^C��1i#QHG疈��Ƨ� �������aNa�NQ��i1t�Syö���K���F��\������8k���YI�6K�U���H�5���KBL�o�<N��9A^�ɒ*4n��w��opC!Wp��`]� ЫV�ٙ��p��iX@H��g*x��&��@������yJ�(���R�g���t�OI�����_t�-^Nì�:�2�Ձ��g֍��:pae�"��O��3<�r����{�b 	�_�3�2��mg�� �+=^	5ᚦ=��|��j�^TۚQ}`]Xy�RD ��T[!�%%����b�V;��h�>ue�:�Fi����7�V�ꙇ�:bQ�G��b��C��;�䣼^�8�G"p�����8w��>a��1�[���<E�Ӷi��C:��@5Zr�c�lB7���J��LD)�!�)�zf
��t�u`&:C�Q@�2����+ןFH�R��;�q�
��bq$I�~3%_dF�WU݃$�u=�f0F]�%C�M��Ō1c���>w���o����t����	��~g+���Z�����	����~�Yf�⭖�2(�H�z���+:΄�]�+م�+�;�sI��W�P[��������؎~�.����m8����Hw���/O���T���=k���N����+˫�	K�r�CQ7�-x��ng؎j`����
�S�I��x�k�Y�/0(,l禲^�@�섅>_����| ܸ�m/)�J&��$.zQ�:WNK6R�P%��g��J";(5[���6�:A�}3�|���(��ۨb#߱�=Sn&+���+Ќ~S�����»�Ι3�����) �J@��@��Ka�����W��[�!��3R]}@��V�9�e[��ݓy0a	v�U��\$ʚ
��>�U�����ҵ��{��Z� u��p|�1��� ��p�����K�����r��C�>�q�B�"w���u�&�S��tJ.kԣQ5�ql��U+cl5?,���E�ʠJ��^�C��yB'&����9�����@=����lf��ƫ�'�D��Q	�g����t�&�o��2ЄlM�s��@8�I�S(k'�ֽ�t`@n��2���g)>\�����{�X���=�ǚ�uֻ�A�}�C*k����,����=l��_BPҭV���Ҥ,�[(QnBf�"2f�>E'��rK�$�g
b�;�gn�
��N��%�4.J��s�`<a{+t����4�M��e,�R}D�{�b�2k7(�x�r٭i*�zD��^��⢩��z�La�t�wY)�������Ź>��~Ͱ�-"���#T��Zdr��z�"���D�� B?��Ej���n���1�m���|f3|D99������[ŏN��6��j�3d�6�8pD6�%1���T��g�T���dd,����Z�7w�gl{~֌b��sv���g�{�~��`Q A 9���_M� ����zQ�N�*���r,�}D�<%��]�U�V`i�*��8�{�b�mL�æ��Y�71������}ۤ5*�h�6�Ҹ�7t�Z���3���6�������hD�@����<��rz����x�~׌��#蜾��f�G�.��F��Ty�r1t���؇Ld���+���6}��zI8w��u�i����<l�<p�'�֜F�e�gB(��7ؽ����_����=bDPy��/$ɖMܶn�����G�}O<�N'K��ܪ ae���K�@�c���v�y��h�mp� ��k���J�/�[r�_
�N��Vj�c�� �������Dy.�{�=���z�|v1z_�U|aW[=-�5
.��q�lrʳլ'M�݁+Sp/8,�ޟ�eմ��:��:��d��8��T^� 7D?���*�ˠ*�cZ>�8Z��rG3�Ӥ@���\M�Y�3�ζ�=#j$>�6�{���U�p�6�E�*G p�)o:��6#�`a4�y���V�c��?-,x�'`�Jz�����؄([�Ze��;-���՞��*�AP�n�hH"�����n�"��>,��E��H�?�L!�[��5�i�ێ�d(7�(�W�q�,����C��f���ӊ苺�iM�(��Ց�^#�0?����;�i��Lr%�G��@�.bm&]�D���;3 �����Ɉ�b��v��@Lo�f kH��~��'O�p==�e���)hO���{�m�����f6d��q�d��`w�_ۖQ�� �q��Ǵb �)Z:)v�����Е����,y
�;��&/����6>�g>�@x:�n6%f5<ȳ �E��&�Idޑ�{�D��=��K����L�߽�wÏ�����g6��g]��[B�(���]������
��PU����lzS�˚=O/�7pągTs3?o~�>}�2l�3��&z��m/R��^�oD��{�Ȅo�+�f\���[�t�'����sV'/T4n�:�_t����� T�c�]eI�@`��Mw�������~�V�
�⣶Xb�b�,|}�9�a�KbX�2�Y��Q��"?����_�h}1f|��2<ܞ��/Q~��Z��7���c�!� �v��ڧu�<E�9!~���ruSw��Ne>Ux��|6Y��m�	�!�u�'�^����-�$�~s��SzͷF�\�緘��-�~��,L�^ �2.�c+��f(g�>�k����?Ch��h��H��\�Z4۝�q���m�͉�h�� D i�M��3��8>���%��`����*��A���<)li��~�����{d����2T��z�gU�iR��h�0#d3������ꊗ���Z���Nl����)f]x5b�9��8*tベe5F�0�����-��(�Fts��0�z�PM��>��/u#�'�0��1�(pVӣ���b��B��L�Pf�;�lөtb��H�Z��H�
�+����m�*�Ԓ�����!f��<�H��y28ъ�� \�{o��5Y���z%ڑ�-���@H�n��F��K򮅔U�
\�o���;��R��`�����`A� sR�Z�8.���O	�P]O���,06��e�]��&T�#���fl�
�H\D��p'� \�\���]I��ѭP��:=�T��fG!
5��5Qo�K��~�����a+��
�or_��5���4��$n절�'W�1J��K�=�q�mf���f�/�8{U�qFpe�a�^!�ˠo��9v���[�{�z��B�ǚO�*��.e�Qӽ�j�ͫ~��I���kiy�ݖY���=�g��Y��pфʉ�u��\vY	J�)q��),�G���.���_ ��O���^��IaPD_�O�sô��z7xB��K��ʭ�s��L:�m�R� ��,�4c^\%�@�'s����x51������m"�7��ǹ�	��q���m�^:߲���ۂ��� Bi�Օ#�t��[.]����J)�w��[]c}��_�M����߾%�s�xTC��r� $���IК��/�Ji� ��+�y�b���-�qY�W���k�J��\I��s�=�e�ȯ>]�0�؃�I3�?��n$�$CV�g���ٰ,).o�@��e�}����:�����#�&��3��vD��ȩ�=�hmW]�'o~��;q4�'|X^���#bed��'���GL��b>��Ш0q56u���{�(�{^�&{T?0u9�:,��<��M3zk)�	��.����uTh�F��jr��=Bl�"V,��E���P���Ϛ��H#�r�Nv�gsU��U������A-{���Q�P;Yv�ebw�c�H���)���9QP=#k�����>���	�SWW}>��(��@��)&4�](�7�N��Py�\r#�kc���;�l����
��G�urɛ@J����)���"Ap
k�����n:X��r���hi�W��!-��e�:����H���ֈxѫK�}�V�V��|�?C�R����r�$P�Z3�M��	F��7(�0[�2��OT�iIx���<ܙ�V����dgɆ �\s=	��?@#�s�" ���QCn���WϚe7��)��ډg�kUv�+Nk��L��C�g$r1R)�߬��o)eh�̅� o��>���Fx�G�2BC��O��nZ�qj&�wL�V Qq2�OǝS��@��o$$�r�ڲP�,���\��^L��]�h@�5��|5"��X#�"��`	ݺb�����sm뼼����R�[��i�x� Di��g�Х����GZQ8sC�s'yQ!P�kU@Pcja�Y�h�8	�|dp�� ��>JW�$��G�B��c�Ι��i2��Lfй�5Q�Å���b�U��s������0�t�{z���Aˋ����$`��݇�v�\��5� ���G$-������X=��P�b���6uVo��H��@K��kJE.���s����
W����ʕ������j�W1��oY���w���q����*U1=(c��fZ�F�~��B 4E�ť{��i�<�����C"U��tMOg@*��8<h��e&��`=Ć-p+Z]pU�|H��G�������2�Z�M�*Q���+�\(���/�/:�����H�ÿ���J�BFqE� -��`���Z��z�p�%Jj���5i��4}Rz��F��wU�̸���΀�͈�h�$�'��΁N������/�ޑ%���M��vv�	[�Kel�@���M��t�o��{�#�]�����'K{)P�Y��m*kk �K�=_oۓ�w��>�x�#v(�#i'ir|�abVL��lFt��V���=�T���i�FU��Us�'Z�=�2��g��?Y��a�7e��Og��X����ܾ����)g_�;��˳7 �9�nQ�Pق�C���*&;�H/b�r�g^~Z��9�5�-�hv����_*"+p�4�[����t�x�oYw�1	.�QA�q�(�1��NV4��ꡫ���5x�(�[FK0��0�Sh��g!1V.�1uz���Op�Q��f]����S=?Y�I�~g�d��y'I�;(����PJ,Q*�(�������̐jq�6��Jm���}�2���>��ۻ�Xhf)�
�Sm-'��O|�d��%���k!����\7q���d�����}v�\�p��| ޖ���:�|V.e�N�� \��f>�߿���s����B�w*����N�|����:�'�����S�dߜ�G�kv�LdZ�Y��-N���(�WX�ma&���f��`�QP��8���};�@�#Mg"�o�+AP�H~]ߞ���vd�"GY�| +�����|�B��}���Y5p�b�}ׁo�<+��l���q}ΐ�OJ��ڬ(���|��/��fs_y���	���h�"y���F���v(�%;�*�3�  �t6񬵚a�;����ꅊo1�|�6���