��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ��nͳ�R[�ظ�_����Qq���G�]~��\�^�W.Z��ke��X�?�I\�zA@���Y"���a`MBl��$���X���/~%�cg��OU#,��;o�w�F�~�wy�0�Sa��qC�$�_됲��ݗ� ���D��.����v��C��k���<�$J��3��I
����<[�P�}&ʁ_m3�P{�
A���-X'�H4Eml�}-���i���[�f�c�:p�D�Vp�[�4��-�UHM��G�j���2Fsaб?�ﻗ}V����g��2*3a ű�ҋ��>��	�SR�B�}����MT���E�nY[r�%D�rN����&wst����L�
$�S�����M:���m����4�Ƽvߣ�4��l�K������7�U�!ʼ�Ӝm�s�߈ 4(J8?��/B<�?[�7� }�һ]ٍ�Ć@�� ���S�g"U;���	�GZ�-/y�g@%�$PX�l�5��2=O��	�����^���g��y�dg\�v�4)9s?�"Zy˼�P7��!�=A+U�0����u
�^�J��^�y6����(:;䑆u�O��cIx�y����p(�OJ9��00�όխQGY5ą�'�(M��W5r�W&����ν��m��*��Wf�h8s��7�����-���W�x���稟?�R���:�tl�Ȗ^�%eu��hC�J��m�y{�i�Io�����x����(|4���Ъ�s~����w����b\�w�!�L[3��Ԩ3Ɩ��y#�p��V�����+��D��9����,�'R+��κ�/���&C�]�(��� �\Ȼ~��_�@������4� �]@��H��Ё�k�yv}y������v�����qvRdx`����B%�̊5zn��D�XW�-�e�V���ݰ +���U�Z�G���4tkI?���;0�ۨ��_���tV��okԯ����9c%����ʄ�P�B-eH���3� ?N5$6=>�1�j۽���@�!_�~3�$R��Q�c ��C�y@���k!�#!t2<��2clgrۚI4t*�o�o3��2p�v��>�o�\�&U� Y	e)e�7��"+�9/�V�W	�nkf
����G������F������l��/��wY��eCRucR�����z,��,. y:.�Fm�2��4j)����|�8wN���8P���,EAx���(�"j�ˊ����~_�R����b"3v4T+v��G�/n[�so�!��"1�		U��:�O������J�p�����>�iH�3�c�ϣ�b$�������/S`��W�x��g���ǵ3�vk�Ad&�8�������a�V� 6p���37�7�B	*xĘ���ݿ�`s!���N��)SG��1"�*U}@�S����Exv1`5�-��������~���L��y�Z�zF��f����&u^��&�-Bg��f/�jlm��Tʒ_4)_2��dU�Ε�y�N�ȋCu����&B|�߷)�}���5p]��c<�ϖ?�W�]e��%���ե�la�~
��Y�����ݹ���W�0Ҭ�?��KjDĳ�[6(J��\(� G�.�l�߿�j�� �EՍ���B���SBG�/M
�o�o��|Nx���w]oF��4�;&��ˡ쁏�������I��r��"�r��ڜ =4}���-OiL���z�H'���v�-���X?�K��>�M�@�S�/�*f�f�F�}Lu��'T��`q(q3z*�X ����V6=m�ޓF�ک e#��=Čت��9�k�5b\��](��V����F!�D�'q�֟U�l99Q����iR��ע:㿷$���&�۳�^`�]Xk�C�F��ƺ1چ�;�w�<>�Mkԕ�J����N��6�	8���� ����Ǡ���$�����A��[9{�O/<�;`!��؜����Z���r����� ʵ	���z���=�j��%�C̜~��1�1� o���
\�#��p����J~�٦?G������L�}��fbj$��3>8�sLy�ӄ��{�C��)H�Y;*�����1:�"?v�'-
b�^x�A�H���\`nd���
6���D�{�T��Κ�E���`��9���r��w,5�s�_4ҳ5x��}�#�`��Ѣ?Bx�;�
.�?bݦ���5xPPC�2,���.l&���H����zeG-���y�����5�T��| {z��Ϣ+�d7��M����(�ѫI%r�`T ����`��w�fՊ�K�RJ�;� R���w�5o�·��[É̜�z]aH'� /�l��KGmu���ڹ�k���AZ.����u�8�!dR��2�����Ԣ���Ʃnɶ��#�c\�Y:�#�pa��i: ��.L�L�b��D.(wj����2��Ixc/l@�����E1�N�1�0������m*�C�7���?�=M�*]k�� �$m
���0��N�5m��]��_��o�At����^�:a���q�P��& +\���Ǜ}�A��7��G7��X�$!ow(y�q���D?�HX���Ɉ�����1R��ks7�u��-�6$���v0I#k��w��bqh>�8���(b���u��i�y@�E��Ԕ���<��� �$�x�1�V �ߠg�Ĳ�:��Vua��U��[�[�F�˳mcj�n}�,Ʋplf*�iY���P�a�_o��Z�G.�����%�A�A*��u]�x ��G�)5�������2!�{�u�DP9�YIC��Fȴ?h+���K��Ep�)?P�q���/�_�	`�MVwļϕ*`�?��&���*��l�<�f�[ ��7	�s��h[�1�6;#l�~a�#��P6Zc7xc-��T�&Yc�s�]t�o�ݮ�rU�K���J�s�x�Q!��wX��r�+Q[?�g#؀Y�ԍ�1�e�ގ:0�xK߅XM��_^g�����K��oG]}�d���R>��Gȑ,Lz�{Z�|v�?a��?~���]�^b��]��XT���=�.��Ċ\?�$���W%N��A0�j�����&˴�������-�e�;���u�m��3>��x�c�����_�� ����;
�C ����H�m���k����d����1��␹0����^��l�}�(�N �JhM�O~N���j��Z�$�|Mw#���u���p�C6�O^��yKP��b�z����7�,�j��i/g�����%�bt�UO���8}w{)eg$������Y���p*P����!��Q�%���B��:��{�=�b��tj��%���Q����Nz�A�>8�4�@B��Zk�yL�7s̺�8����z�C�q9J���F��K#�O��e�M�*�լ�U-� U��%A�xvO�#��` ���
[ޞ�>�P�A\����u
�Җu$���z��}^K����Ѻ�rџ�;���vracy%�=ֹ�,�k��w�9H�����6���Vj��G�L��c?8�9�NƜ'R�w�Ñ�T��V��C�p�j�r�g�a�����'��/V�6,���Zܶ�T�0bн{~\��8�p��#�fkMzo��5�33=��>�2��oM�N��x7�#������&"��~�T�ۙ���`�b>'�p<�De����Vu�B�X���ŽBHG-#w���$&)��.�	��	$`�Q=1p�BJL@�0#Ni)L�<c ց#G������#4�`$��|��Gs�.��?O���wU~L��x��ª��4 晴O�I,x��$2-�N�{ĩJΆ��nl7&}l��^���r)�Q�Ӓ�����T=� �D.�~�� ޭ�3$x���ŚI���Y�	��6�l�|3 �.Y��.��>$���X�MO�9�����Y��bL�+�U_�9tyj~���9���ƞ� YSዋh�Z�ጹ��y�i�ޅР�vYX1�(F�IůiH�^?����X\��'�K����}\� ]�5��gY��W�2��rf�&�`v�Ƣ��`��[��3E�1�hq�@�(cJ�;	y�G)�uW��gd��_m���>ӎ��
ۛ0}�T>���	�e��P�Bx��W��,��h��Y��ZMi��|���f���3�Lbe R�P���p�?O�.˕C���5�:0	�{��s�N%���5"N@�%p�j.hc�[ �R?��#�`�4d�Ϧ�ݛ9X����r�F