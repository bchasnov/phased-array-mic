��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,G��U�	�oJZ�@�z�����>�� �F9!�/_g�T@_hm/a3^��(#z�dZ�E�����v�h��|���-�>����w,.��N����9Z�S�p�ւr�p^������[�G�C-�Dʩ/�Pm��[m<��#���/5��X��i�|��ߖ>���p�y������CP��� [�FcC2�YJ����H��d�4��!��_^h8IP�/���e�4Y6��Ơ���:����ԚM!
χ��À��]�v�xw����@>��p���,k� ׉{E~YnG�Ǣ����ik�1:�)����Д��C%\�����kC��p�w��=�$���E�2� ����;����UX��Tύs�R��8�7��)�`F,'�� [��D�K�uT4����)v6�b��(�߱� Ox�U����Op�9�W�����H�Z�읖H�{T��hh��R��p;�$C~ }�ܾ���!�o
��ӈuE���
Q�緪M��ʌ�?ݎ��
:Q�В�:z�`Hur�FҪa�۪,�[q�k��t�9-�
&���ZlP���0�'�B��w �J�N�w��m�ŋ-8+����)��|&0q����9ݑ���T�r#�K��_>������Dq�wdy���o����'���8�p/|�wK<�����-#�s-�	jL�:��M2P'��8$��ː�lo$HB���L���v��W�@i�$HG=Ã�A��{�C�u�̱)iuSI��x��G:p��(�`��.	�nf�]x�A����h��1��L�+A���_�YAs����<��R�3�O�z�C���ž���KʬƁ��xP.�����^D�{�f�Jnb{/����8�t����ɦ,N�V�9h��I��������L�7i�8e9���{"od,�W_ƅȹh��hiZ��]-�d{e)?s��h�hBK�Hs��љ��.n�s\�fk�JԆ-�1��$<]�#�/���]9{�K�:�(�2�]��8���K:҂�W[\|U���W+&�~]��Ssc:��=����?
�)���hTm����p�h�}�2a���oz�/�+�N���'�!t�i�=�18��v�7��;
�?������tDpM�(�3�6�g�Q�����f�2z� 菊�
2�βl�Y�r)7�@}�+*���)/E���u��r ����Pj�� r�)���3��O���=���7G[qJ��r�6�{	ެ�[�X\q��	\�j� �ܸ��{6�4��:�V�:P$p�"�����i�YX�W,,m���n�v,�i)��j�K�N�v7���va��P��`{�V4V[r#�����'R���I��_)�[�0���߲�2���G�du߉R؆u�-���������~#S���"���u��Ҡ	p��2����L���D]��w�����5�>�!����K@��7�J� ��8#������<9܆�`���V���Z���7�z
C�[L�������>�}�'���]eC������a��%!<`������h���l���ԀIc[�u�ni
O+�:��� �r���
��|={�;���Q*�"�$���s���+�sV����v_��ȍ���$����?[!���u���3����ĚI���5�f}f��En����Oy�K�w��/�0+md`���̑m9U�s�ǥ����2��8o��ebd�g���������a���A���p�_$�vGl:eK��V%_&�,$ń�m$NX��pS�mu*�ѡ����?�CJl+�-�چ�X��Y2���Yz�]����)�}� ��9�U�zL�%Ƥ�o�� �5��o�l���h�|�o߫�Lo/�	��2�*2:�U5n���~���ll%��R-|�C��Α�yE`@
�E%,?�G�|�Ь�qK��^�
u�˰<�#��Qo�e��?�/t�sz*]+-�O_�[&�Ņ�V�9x N��r���w�ܫ�Ұ��+k� �/�پo���AX[
�1;/��&�����v�!G��mL 2g���C8�5�D�7�>���z�Z�{\R�XE{;IP����ř\h��k>)i�A�b�h+Nd�s&i��>�|�g��23sY�F��`�RĖs��h��r��,�xl�1/�"�W^��?�& ���V뫊��Π�~�!����<�L(< w�QW�}����;w�F�BQ�щ>�h�y9�H9��EFsC#ZE#E��W	��q��p"�X�����钥5JMY�K�3�Qj��pg�!�_�{§�m�L=�ُ/v���"lU�`zE��RM�F*��s$��6�[9A�1�D����G$��-N.(q���G��۽CF�a�V*��s�g�2=�ިY��K�]����\D��D��)<b$�5��>c˚q��B~N��q����'��$�~@	cG2�<�NP�YՍq��rX9�th�b�x1A\�����S�K\��6|U�S�m-���R���_�.����{��#;$m�x�Q�pė��fL�kX�,��]iW+��q��`��6ن�4W�+Q���r�ڵ[W &�O6E<J��1 O6	$�@1��~���zy,��&R���K^���N�h3�0"�#�6�n���)�"�~���k�ť@�d�te��E�9�Q�!_˱�x�ϧo��Szv�
F���r��A���tI���,I�Ԣ�O�Âi�<Ui��e��hݑQ.�l���:9��s��s��Vi'��"(��|d��<KTt�
�$iHOǿ�|�,��`KN�O���=��NxZ�f� ?�����_���'����m�@�|eoO����1�r'�Q�ۑ=(C��ML�Yx �;��#?�_s�cHiL��)o�U�l��į:����~�����Gc!10pQ�n�~���e˻�ײ,@c��a�]�Ĕ��I��Svʿ�%D�mfu��G�� �(��	��V��q��f	&�E,|�ż��j-Q` ��Q�h���}L`��.��"
W�L�c,v�5�����:��v���E���p��h�܃�R�;�k���f(عH�hk ���X%���d�
�n�Q8�C7%�DhFY�L���m��/���q���l]g��H�If��w�L��X���4�G�2��d��"�N�z&.�IAӢ�������� iv}gQ�z������i&������v(��02�T�4.~� �.����e�K[���[�k]P��7~��'l��c

#����� U&}�5R�ݴ��z��A���˷�2	{5��v]T������y)�O������܄��� ��u�-�#��Hʼ{W�Fu�fW*��<'���FS�Bt�)^ݬ䃿��v���^#�;RL�~�_}E�Gj�)rJ+�|���P�3�Bd���~��� ����G�y.)t%+Ӝ�Λ� Ȃ�yK�r*J�8!�@6�(����������?��f}a���l�u��е��j�r��B�\@�bH�5I'��7O)������)o�:a웧a8��T�C?�	-C�%D�����㤋�d��S�Z�J��8�gfT�������Ǖ�V@�ʒ�Q_O<��`���&;
h~D�Q؉̼轉�V��"S����;��}K��wv��ho�0>����%�O\����|��a��u��B��#��(��T:�pA͍�P�a�И��d�B�+�"B�:-ۂ�5��V��M�v��0	�}fP�o�T-F9a�����݈n����.����͝�Je��a��}3.��ǰ�Qy&،���b��AlN0�/�4}Bi�,)m��+(���mZڛ]�9�>AWc "wrz�{�ei��Mɿ�,@�Rۋ���h��6<��ƼJœi�ʜiX�Ҳ���F����,�L���� [��Kp��G"r���1 M����Bh��'����Է���v��2�#m�7�^PX�:ގޖ6���tr��9��3�ܴ���}zS������Hj:��	&���PM�8j�.�:���� �RĹS9A����v�$:"5�<� ��F0[�\�~��]�]�����6��U�ΚV�2 zc�����ƴ:j;D���=BaF�l��΅y����B� GRR�/��9�047�.-�������͢�s ��9Ð~����n��j$���d~{׫D�/�2g��$�ű6_U�k<����i�'��CH7L���#����du�ȸ��v�����Rv������������w�7Ԓn�����/ո}���X��/#��0@V�-��9 ܔ���v9�ٚd