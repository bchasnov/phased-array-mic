��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1���e}ʲ��cg�t�ϙ�a�:�KR�%���ݧw���ȼ"~m���7��6Ц�~��e4��+LN�u�ʧG��$�h�lK��![J��q){�~�H�@FY�=;#�͙��&5�h~� i�pnt�Dv_�Lʛ��E5Ҭ7eR�%�E�mo���G�[��/6"1��Q�T9]6{�%J�@��h�ȕ7"���L�JQs&q��.�K�=I�|����q�q���n���.�{{�E�\by�x[�|���n�AP������{*�b��M����T΂�g�ڀ{B����c.���:��3R�91d<ǟ:�|�ϛ����U#��.w�������+�P�o��G
���S@U�$,	��l������y�k�������k;)r6�Q˔� ����*+_��a(S�DV^���lԧ�.]�T���U�I��n��/?�5��*��<�$Qp��$�y�
�O������E;����00�M[E�*<�-s9.mA�m��zW���9%[*)&��x��<�D��_i|�Y�P�n��C����(��e�7U�{R�ϥD~�5K�����QK}�5�&��dP
��(S
[s�P��Pn$����3/: :��q�e��ԺL�؋U0�=��F���d]�8�g�A�5RJ�����6k_�#p�v�@�T�-�g��v,��B�^7p.,C��+)�wǦ�/���.<� �
�"Ԫ0c�^[=�  �8���*��h��ƄK��a�b�sM8�K�ߖر��x.8�����Z�eX�(r�!t,w���Y�su�6:! 0��en�A<����o��~u8�UÕ(r����Q�J����q���%��	K�-)����������&6�t�05�����l�!ѭ��GoY7�#�d��;���i#����I��t>�M�Z�_ά���7���1tk&�g�s6����-��Qty�d��Ϸ��7&z�C�p�C�zE��_!D���V�=^�	`�����nH�������D0��+��A=�F���K<&a�6�@N�jL��"p�;��? 6zt�4�9|h.��f"fZ�'�}�!�O�Gm��~dO2i;L+��+1�MvUQC���O��99_���w�LD�eU>����
�t-��`^% T?Pb�H�_�j>1p~�/9㘳P�k�.R�r�����M�~Jonc[��	�M�/�s��B�.(8?�+6�~��IZv����H�(.}�'*�"�݆�B�����4��i�=���c����L���-(�E�[��5�+�`������Oj�$��P>� ��\��k���?��Vt{�ۮᆂ,�c���F���g�`�,�͸��jd��<�����ˮ�4�57P;��
�����P%�­����4CM�dz��������2�]��5i8��Z�hv����pP݌�'`<4l�-��"�`�W���Zi�����GSّ�`\a�?d�ht9�m�vuL\������|I�鉺��� m8�v-N���w	��T���V���Ww������%6�精�lTu���Ӱ�o����*�� ��S����y��*5Д����,<L1��ˣtw!�&�EM����:D�[P�6�����D}f	S;��t��v��"�F ^��u<yPw��~��6j:��6\�E;���z��=;�Y�B����3�n�*М�OA]�o×�s�����%�KNR�^)��_Od���2y$M�
��d����4V9��$�$-�>��j�Ħ)6,�P��K�� �<A:L!�F�;�n��~A��	�h����}L��楶
��)`l�*c���X�
tJ�h�����t��S���b�;���!�	�^A0������Ԫ��#S������*����-X�C��߷�E����I�+��<�1wy竐�ϐŋ%��8/�Dŀu��a9���~�Y�/�vHX%�� ���^%�F��4����eo ����G|] yRLu��VSb��'J_��:2���_��1KM�b^L�޶��e��m�K��Z����$*	2e�|

�Av��4yܦ#��$�o��Q�I�M���ێ�6�?�Ϛ����`���NBL�T}uV���p\ɖ�0%s�15����dS�L���Q��~fG;k�`p��@Qʚ'�M�+[+$� �XGw��}O��nTL��Z�ue���o������D�Ѫ#9�Y3�I��д��Pѐ`}���}�T�0����9�Ð�1�G�	Dq:
X!F��
{5��d�����$�kE�w;�F�.�!�JoD�mP�� ځ�\����pɵ�[F_p�j�s|�jVOD
-8)�⼉�����?�Bs���%"��Pi �`�-�u۫D{H��T�lH�qoH����L�����j���ٲ�L�2\3Ot�t�8�Բi2��Q�[��]o�L�Q��}C� Ls�K�l��8�S�?,��wwџ?�2 FL�,O��U&mF\����l�D\��w����z�ô�%	ަ|g��Q��&��f]J�e��0��[J�hXzIݻ��"E����X �����M�vK��?���N!��9b�  ��w�����&<�BO��߆W���UW�v�Zz��;�G�cC��A���aϷ�)��{���Y@&���g�}\��C�U�� �SL|�?��q���� tn����[�ck벢�am뾍N�i����^�X��UtWk*�9�L��vx���x����C�eT����Bs|�u�1���H��RXK�O�<9n��y����kl(f�i���T&a�j����h~�y�0f�T�.WGy[t���^q�93��ES�A�N�<���c��,1R��������UUa�kD�,��囝��'m(��m�ȿC��k]i��L��zˤ�W+"��P[?�2��O:�`�W��6�D+�l^'#[�1���Z��`�����;'��yZ/A4n�������;�6*]RH8���x�`n���f�^w��>��9O�E��tf怄�\����(��	`1Ա��i.���Tt7w�,Ò�'�Nb����>̍=�xl2|�s�H��+0R{$kM��	��}�O=���R�^H��ʑƕ�햻0�˔��Pz��4�a*g�2�L�
b*(Z`�Y�u'�v�'C�WY�v����G� �=�9��ۉ�$edb+���Pk���ɀ$�����oZ�v�6�O����2���KH;½��L�#����[�������LD~�}yX?_�����Auo󼖼�qj�ŰЉ{�6*]��BW��ݥ�F|�7�M� %�F���pӕ��N �I�܉��Ƥ�&�� g�&n.-�ab�μ�����?%�T�&(~BB�����H��9�����R��i����-��Δ��cO�|8�)�N������u��	���>�Q���pH7vq_����hD��fU��5#A��Q;C[f��j�t��	_0ā��̿�&���&v[��e.h�!~d����*T�B���E���t��tܘ����F�]?�������c�~i�^#��轃X��Tkq78zlw�>�G߽'��n�j*<NE�.��?b���_�y�����4Fy	]��v�j2��5cl%F�ݠ���.-��o��*ԻȔ�����J�	cJ�#P�
����"�n[��@1�~��&����F��9�nDS�̾.�K-�T`)>|�����@7i�8о��"Y�Y~)Z.���F�W��郫�FE��b�����,N�Y=��HYh|YWA5'�P웞]�S��U�ٺ,�%��V(����?ȡU�5�'r듺)�����%��ˇ��0����?l�;i{.���^���!���a���7��t�{TW�x�]�������!�����������q9tBK�Qes����2�y
�m�3� �C��'��С��Hr� f�����7��䂵����
��yX��\l�}�6��\�+��2N����J�[�z?�h#���ˣ)L��83�jk�j�_[	[`�tu"�8'O�?�Jgi#Y��D����h",؆a��re�V�+Z��p5�uN�+h|���E��昪�����
�A�R�}�"����<:31�i��~!�ù����;��a>��B��[Iን�j]tv��He���҄u�Z{m}ڦ��ͻ^�s�m�6Y��SLuB�Q�i��u�W9]��]��</��HTп�/����Ӭ�EC�Xca�k2��R=	��H�E\��K�9��7w��,_��1�I���v������>έ���7xb�aeð�'��=QdN��cM�����)aQ��2XN��Ų�����(j�u��h�3e��]�$^��rXlͮY4T���.^	O� �̜c�o�a��$���S�1�����{E��˲��Lfp��uU�����"�0|�B,�����YmU�2W�A:�vfl2D��w#�>`��fӈ�.��~�&#J��7e�����D�>'�Z�A��@�h\��i6ui�YTvc�`�8��u���:�'�%�$�W1�T��cD�1���.!�  �Ȏf*�Ԡ�&Qx�Dk��!-���-�]R����]0���b��$�������АYS�/�gԆݒ�Z�~�3����V�|o�KlCϴ>
��#"����ݽ�] ���GӐ��C��X���K+gS��_����`yc���q8M����=���r���qJX>���:
���AT�U+�y�(��s�s[���x�N�q[w0s;r��"�/�!���\��^St A3��-6'SAؒN����"7�Ż�赈�k��M�ź�Ѿg�2k��JR��9�6F'壜�,�1��[�Ck�fN���x�Y��w�+�^z"���u���R�{ähH2�m��#y߈�U��6)cF)$i����Ɠ�EMJ�����:3�B�u����!���7�X�A�f�)���jū8��}Hٕ��ιo�Ό���Z��kc��3��#������B��VwR�a9��*L"����[�!�%���c��ޅ�6�8ze�:��-u�?x<�Ѧ7�7S�}�r}�`�IQo�����(m�g��Q_]!ǈ�#"/��t�0y�9�w�����E��٫��5!"(U��<��,R�g�D��$�#�P��&5�@>�ȫU� ��z���~�xknB��f�.���/�<�< �҆�}u���K�(����v��(��j��P�G	����u����=�}8Zmu�3�����2�X�h�Ł�(�!Ҝ9�/�`e���G[$k��V���ә�M���e{�~*�4���&���Q6��`���ߋP|��}:]X�DfK��8�a�yo��
�����������{��f�Q@H*���zym�/1��bϫ�k7k<J���G��2�k�j[L(���%e�ʩ5t��V��ԩVi���'�F�EE�Ҽ�X^���h^pLM��M�,���#�fs���G2Tr��37!s��iK�_]���Z/������q[����޶����тT���|���E�~�}�%D�B<#H�A�XB���PW����SC����E�t~0��l�6�r,�?�4S�~�&Z�#�����_^۱����٫=�\��JK�:^U g�H�.Q��Z���q���Q�f]���X�Ŝa�1���
%�� �Eoȋ�i�i�T׽M\�ZGe� �y�JG@�,�Ǌ�+��i�q�:l�9�f�mED6�a&I�z�
���u^�lJ.�GmP�SE)��o����MH��(u5ݸЫ�,	����es���uE��L��rɶ����O�`!��|�ѩN��������ɤv�tC�F�:B�EՒ���Ja�F���j�*��x&O���IMR�����<B	��{�ll�J<�MD�h.g\
��C�|����[`J�Yfp��E�H�.b�-�q+�����U�	�`�('��{y��4Q3�Y#oK]|�[����g��/YHgoK�w�J�[���j��~��=5��Z�Ʃc�n�ڃ�s_��s��O2�	�y�Rx{��~(��!�D��'�iQ��q�|,*�_�=��c>*��A+��;ٷ�{Z�������*�@㓽7��.�`Y��a:3:z�p��7|�������6n�4�JGV8ܼ2�Ǐ7"����l7u,Z�tn_~U4)���<;*g��	8����{���P<�=u?G���Ή��Y�t~'t�=��jzUd�oh6Υ���ۓ�7��^q�=�^C�\�4Q�e%k������=�b�2��r�^�����`H���g7dO;�L|���U�z�ys~�yDc�:ߋ�t7�z��,��2�lna����!�J,sk�)z��Y��O��k��&�#�\c�4��1|�J�M�z��d^~�[&��z��*�75�F9.P�y�%�g��h��薠*)��R3$�]���A���h ����F�˻WL�L�~�)��d��W��^"#�V)�u��3a,<�v��=)}�[}8�lR��#M��?��]��c]d9���x]�謮�2!LJ�Țm����R&�92�y��=f��h�3��y���y�Q�U�ڭ./�~�\9�6��q6��#N�`��<�fr�����VwwH�zHv��/��� �OL��a�����+�K�}7r>:HJX�<%�h;����ܻ<��ɩ�� ��#�H�Ī|�����H�?N��͎�r�an�s�Ar5��PA���35]C��k�W��G���k��Ă#@|�%��rbz�N��\�u!�>��INy�6���]�M�ח��81jժ����Ĵv%~�2Z��aE
���)K;���nƂ�ذ+�1{�&��{��H�4�����L�O���Z.�NwSinM�B�Ǥ��2�����-�� ��D8�B�o�D�:��cf����9u��'(u��G����~'�p.��Zc�7��:C�}����Pw#`Ӷ)NG��g�C%�%9#WF��ȴ@�(t;D[?F��m*��qkU.�aw#J�y��������1�^x�t.�h4�BM/k�'0�)��^�"���Jh
 {6��a�t��tB��{�+���a$9=�I  }u}"�N�69��{�2��r�%���-Yr6����>�a�2x}t"6 �-zV}s/��<������)�`�3��(�c��D3N~u��r'V��a�P�n�����������wG�v�+�Lnͤs{+Lg��`��/�Ғ���._���ɨ��$B�