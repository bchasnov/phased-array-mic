��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\����q�?��e�I8�b�Ǽ$��"����ׯ1�V0����a�ڡ��ˤ5tׄ�`A�/�%�4�ڇ�}XR�b�����tiޡ��[���1�\i5
��c�ӜFFi��"V�;Ȋ,�w2S���_�N�'�B�e�hS�V3zn� yY#�x�����Վ��' Ƴ*��~�wI�ᐒaʵ	�:R���2�^���v���xr]�e��l�Y���A` ?{n=��U2�G`�#��uI�/���3QJt	�-������D�m���"һ�4�9�Z�m�e�� ����S���x/�D�<��s� �G�����~!���{(�=�����EB�#>[�;�J����)��?u�j]e��o����ځ�d͞�0�������p���F����X����#�3��e���{FI_z�B h����4�����ţ�0�"J��4�⭤I|! ���g}S����R0��3��C���:�8na�*����>�-�>�Y��^PK	\��E��#f%������XK7`��z��).���V�^q�,�M4[����Z\�.y���׼s��8�a����G^#����4�PՇ$����4��Ǽ}6Ra|���>�c��{A9G)�����"zl\���Z����*��ںґǘ1�E�,��H���+�VRd���%J�������`?C�����b�_���i�ϻ~&�d�ۘ�*0��N�m�k(��J'�`������f/�yV���QB��VC�2���r�d]�F��2&�Ftc�x��;��������R�����Z>b�:� O���q`.���Bܥ��S�̥����`�K 5�@��|-ɸh�zO�M��U2 �S��
��5����O
�h�}K7�
$�����v���Ac��l���#���~���f�F�E�U������V��0�ա�>0_�w���B"�-� "3Lͽ�o.��tw�sw� �k��/�ʍf�e�&%���-i�� .5Imd����9ς+��%�H�����/jςO���ڞ߉�u�hǜ�Z�UO�ׇ�0]�G�k��K�l܉t�؆|_�x�?���^�jꀗD0J�c	�K��9fp�ū��B�5� ����^�~2q�0bZw�R�Dh
<��n��i�ҊW���z\�u�:<^/.E,Η�s�Ь�@Q�����Pt�D䭞%����m��������0�2^o�bu�� ��^m�@�5XT�=�l�REc ��.۹O�c:%�[�L[�X	x|!��MPgJ�ȬSW����A�O|���ņ��9�����	�1kt.i��kPdG_m*�)"�~�Lx�ڭ��'?@����c3H#U�ǧlhX���Ұ�<8�6%2�X���J�Zۨ`o�;<Zv�^��S�q�r�(B�� \��p�}��A����
�:���������M`w1���yT����𕐐ٌ���0.*�F��r���b�S}��}�ʝ��nE���A�����bƢ%f�^�u'Õ����� ��-��gvn	$��o�VSY>g�9��3x�:LV�	�WK�9�|�s I�����B��^L�cE�F ���W�T�q�dѾ>
2=�v�xi|�;�b�i��e�S����nf_�p;��&�����,0ϖ�9�ѴW����Id4��脬���t��c&G.L5�$�9	vC��C��7`�������Y�\7�,ʆR�	��C֊ɬ6�*;��rY�H�WC]�F7Z�|�U�H�(5Z����|�}�� ��ԉz���Xɑ+k���!�g�:�*]g��r&�l����Gy�������`�M�+�,�g��Rq���"q
I�y;!R%Y��H���+W#��B�o�r�k��9�ؙ'�!�fT��2�E�d�<1!h{nƜ{ǀL���iXFb��[����G�z�|��"`�(���Z�9w���bs��Y0����@�)esM!iB%V��_lϛ���B��]�����!G>"节�;?@[��Uњ_�7��le]F˜���^DL̭�,���^>Ⴙ�Oa�����<\�����t��h�D��a��w��0����V�ש?�`���O\�n׎��긼?�P���ʻgߚ#�嗕���� ԺDf���ZC�,bq&�.WY�yko�(� ���)���T׍�9gg���H\#�8�/�z��v�
�Z����3��O2���ޠ�V�!%��|;��a$��Y�%��k�O��	_5%�=�w���D��`|iV|�;�f{D�-��_���d���2gQ�+9-"$:g��/��J;ԯ�	�R@ �R-��+c"�,6�]@͊�z�7#�zyM9כګ��RJΏh�vF�Dȹ2SA�xc(� 
Y����
�+X�������m�+[0:��Rd�{���(c�y�i�lň����J4�b���O�NJ��$7a���]� ���� ��VRǸ��5Bh�a�
��6`2i�֮�u`���V�:�D�r���8��2�Z�TϹ2����-�*$1HrIf;N6b�4�����y����s�D�\��.��$|Ԟp�j7t�(K������Z7��N3��JD��y�B�Ь�& ���*O��I�/���L�&��R�$�d�<&~lo���$fGE��,p�������ϕ�1l=9-MMUfc�[��6up �g�Dp5��+L�x��$3�_�"�v�����|H�����E���jx%I��.����"I�P�����`��0h?VZ۩�R8�mq�W;p@�d�#��GZZ\�H���`�N(C4�9�g&�
U���[r��\��\Gr�����i_�1&��Cf}۬��NWzƗ����p�
-��x�[�r��.j�}yV �.xǪ5H�e�t����{��7}K+�f�}��?��-�����kz��z��o�]N�5`�$���o4=]1?�VoMW�Lz��(�	A��ztg׬�P����e������AMI$�Tf�2'�[WZ�G�C�����} }�����"k7�'�$�� ���!�l5X��"[$'qڈ���|�҈A�E����+� �����c^�p�iA\}��SR�y,�k �]�<9��b݀$�����ｄ� ������j?�<O�%��12�w����Ϳ����Ɨ���C
ۓ=��'���R-�	�ȧ��/v��Œ(�Bh1[�?xm;X��f�]P׭
+�9?íuC`ɕ�]�����/����7z�;��@�D|Z��&�PDV��~49�٤JHqo��7)h�	F��H�39U�f4��sx����_��Rn��p�n|�]��loz1U�0���2�0\s(�ȓY �����Q�ˏ�"j��W͸7 A�ep �ږ�񇽎^h?J���[��na��X�U�I�2��е�����Nq�3�����ڐVŶFe�YȄ.A}�CQy����S�����R�#�P����Ԗ�/���+�|��<��y��fk�T%E� ��8B5I��QT?���,l��Q��vw�Wj\��vN6{p%)��(E�k�a>?��W�u�8��khY9�Z���/��klD�_�,ee���y��&uX�$XD�SU�Z�^C�aO�C��۳Q� �y�J���&Lq��,�Hp��j�gv�ȉm�}�7��J����a��U=oA$�p3�UM��PiF6���=WeKF�R-b��g�������C����/n�Av��&��&�Z��NQ7��\���Y��@/(ՅG�*x媖���O��z���a���h�˺Qx���G͒��@�	p�;Q沦{}��g/M������iL[Qp�s3 �bI�����X���:���q����@|�1�wk{����;���W~H.�8 �C�?>K,����4J6��S�^��}��\\����7uh�+|���/��ڑ���&8�s">8|���~f��j���A*�-�c~|�v�+*8��^�%�o����ڄJ���b��.���}�,�Y�T`p�]_8FZ���6ZP>��q���)��1H: M�f��Q�,��&�/X��<7�m;�(��n/WR�.�40�[���_j���'1b�*E�b��*��wJl�<���p���9�YS˂݇��LJ�IKZ
v��\�K>6��=
r�:�j]�<Yd��H�{��R�����(ZV���RE����W�Y�b�Z�6w� o�<m�0�:�S[e���b�S�n  � �%�Y�" &�����$�Rc;Nf+u�������v5^x�p}�F�%�u��g��q��tۊ�j�gY=��k��/e��{ڊ3�^���-*�����y�ٞ���S��]c�k����۬�R|h�m����L�QC^K��m7nm�$�@�b��O�w\�m-�Ě�ξ�!M���gj`-V$�?_1gy��i��#�e�K�jNv�w���w[ ��鐳�ҍ�������*��V�,�m �x�K�>�PEVC��Y�(Z��k>�����v��n�B�n��^]A�z�����-�_��p�'��|��L~h"����oH��M��l��|4�,]i�����n�UA�L:��.K׊d[�⨜��t���)�0�^#vAt�+͑�t/�ɼ�5�1oy�9�l�{'��c�Օ�%-F"�%�����I-_��L��~�6���k��F�n�qW~-�D1�vݟ�7dZ�b��>���O?tUiBpq �q���}5���ŻЅ��9�:ݾ�q��������Y�E"�H�8�A[�I�ʫ�����2�
s�卜��E�\��O�2�����c���8g����-Cr��/>0��R�旕תe� �^��Q�|�7L��x���wo��%��!�%��i�e�vg�*��KX��a�;�������昆l ����+Hr%�,1K�ɜ��'��ބ<��1��*�R�`�ġ4#<��-9�уL�+C����3�x���@[ �%�H")�h�[�B�4��ښ}�Y�xq��
|�΄/��U ��3�E��J��J㵲��h��uB ���|2#�?�0�! V��g���s�ɭ�SQ����5�/��#؂��ߠ�w(�P��S|��q�Ԝd0�c:�%6v��� ؏��񛱝z'����>/�p,�r(8k�9����{�d� }:L���o��o�$�]w��Kr�#M�8���%�2^�7���D� ���vr���@�^��O"ʹ�{�NSM��3�ā������&Y�vp�����\��S\I� �5X���F�S���ێ���mS�q��q�C;��8~�nB�1�'�����JT���,�M���L#��4N�5��4��Ԭ��vB�nI�"����|�5��3�I��0#��	��/&��!�*����3-�|����D8�h��>����B�{>ك��)�?�-�hK|^�i��U�k>���a��f�xf�v���~O`�m�4��Hм��A��3�;�2����}c��6��2#>�$���!��6>i x����I�*�J�2������$�hb1�{l?{3�yZ����檚�!�7�A�����ss8�oAH���1������!ӂ�l����(f.��:��;����9ia�]�h'˓j�FiO	-�*��t�Ӟ �
���<�~m��B�8��}��(��0� ��}sC	�Qeg����4s�V�����drz�a��M�٫vL/���;q ��DMJ��R���EL	��59�h[�Jnt��4���G@V+ʆ�p5"�6p1�n���*�k�d�V^򡇢
ч��Xk� �8s��.p�(�^O�+N�ZA�J��n�	�6������5�8A���LIm�}�j�ǜH�wJ��F�h���d���+�`�}��B�z�AYo4T}}�v�il����X)�e�J"g�b�<>�\?��?�4���i�	QX54�w�w�8�I�����@d"�Gc�DA�D�F���� \�c�;E�+�C��۰���G%z�y�j�*��"+�<ud<��z��յ�\L�ңi�%���X��m����]1I�nƣ�9��!���M�����L����E�ri
`C�|�*YV�e	p'62ёr	��� ���_\(59r�x�5��L0@ ���;��!,���;���?��E�~�m���e�!X�
8/kjv鷦�Tp����SJ�Ā@*��t��t������_���V�2))���܂%!�����<�f/-Y��
�qhUC?&�������
���oR�02pD{CK�q�����%�ÅRt�-����8���Y�DGf��n:v��%�9��ɂvַ/���i�貸����]�A+,��������;G(1 ��0:br�V�ɥ�\y�k k�����E֐�)~��_��ᒸ*��҉:�e��6]8��f\���^t��To���	���Z�
PV��]�j������ظ(=��|�B#{:�P�Q��}�Ul�q����/��et��hST^��x�գ�:C^Hp5΢|	�P��Ye��?�ډ{��(�d�~0:k�
H	[o�e�^$�m,*�Q���>���R�Qj�N=����I�uZxǈ����.j��B2�|�\�3��z#��4*�]{�4���˥�#@�]����;�[.�%�%�օ�F�{�W~�M�A�������P �

C��>�iH���V�*'CO%���g�ȑ���;�?Hr�ˆs-��?�^Y�$a�i�K�p�nq�����gc��v���������e�����ԭ!�Òt9j��>���־ZZ|���淙ԧ�x�NJ����0���3�d���Nj�����7�1k����}�c�
(A_@d�W"]3ثuH.��p�V�@�A��n�������]rOx�����5��m2��ߐ�:_�/��d��f/Y
�����(�FH멏x<��v*g��\x����d�sU���~L-����$�a�;�6ⲥ���f/�m8I�i��Ϩ���G�%l,��	c�C��E��L�L+S�i��_���H�����P�;�n7SH�7k�r��V�~;Q�r�R�1���?j�[�mr�	|�;?� �Р�{^ׄ�x/j��Q(,|��PF-*&`_$�^%�y$�J�c]4l�@��~ݻ
�Z'����0s2n�Z�����Мl�yA�Z�wf0��������Y�-@lm���$SL����8d8��)�Sx7��B�o!5����w���&��M���X��8U:
�a&��2�p@c�O��5��{aN�@0�`�,.SI�Ny�"�7���]���sK���څ)�8���]U���|�*_`k��,��R��5��!�Ӿ��j �!��7��
��
���mJ�Є�7���)p���!��>�"W���u�J�!^(��)����[�1�����Q]�;7�醰��׎�E�����xܶ����x��d]�V05����5� �cn�|8KM3y��(�����eNp�l2;���`��T�vTdoz�a���s��I܅6��RD��:\���.t��D����ؕ�<�\]
��V��9�j�������u�|��
��9���-+ m����j����)W�d�_o�}Ql�fBԼlR#U��ED�U{���5�(��^T�Z���hw<O@���fQb5�nE��i���o�H�
Ӱ"Z���u��[������<_h�UA�����	�S_�E��%��Y�#�q��z"��&]'2TOq��3���6P}�IbCYU9���ҡ&�Y��=҇ްI1O���i+�/��=��Jl�M�ؑunh��'c�"���\����\�9�p<\��Dc�����.˹Dz�0��!�Ԇ��l�}d8e��3|G`޸~,���0o�g�|N���\��QN�#�n�Y���s`�7�|����{�EV�=#^�~(�?��3�Ѿ��O�O��:�)�m�6���_��ͬ�u CK�x��I��q��"ҍ�Ŗ�H�bK׻ Y+����I�bZbY�w�x�5��,!�����T3�/�!��UՇ��/5h��f��Xh#��J|ſ�n(�˪d}Isg�pF���Io.�ɞ['�gX�d��9����n���Y;�Tv�������ن�&���p mVB7v�� �%�֠�O�4r6�ʼ���i���aO�Z���[��AqsJ�A@�DQ�7�7�����N��D_���1`՛��a��;�}���+����2A׷�zc\/�W>��h���4�w*�wE��^6����o0�n�)��Ih�{p�qRD�
Dd�a��=�  �OM�E^pC���+z��	|ӱ���U���2����Um�3h�9��-���-7��kJ[PH�;0E�+S�X؅���Jr;D�k�dx�w�ۖǤ�Mm�h5$gte��1�7"�w	��e� �91./�����"&�/���hІ'����?�E/2�.��%�R�$F�]�d�M�Qu�|8	�~цzD������9\:|j;`� S�M�E񎿞�y�_�U�2��q�y�}Yd�&�{��A\SЅ�l!k{�3R�3@�V���sq����/��'L���+kR���Z�k_"c.K���L����#M��S(7��%�R���?��W���=��7)^g% �jx�뱻,mH��
�*��({��n��u���t��@�����E�!]�>��O��q๿)!�8S�?�),-��4*�m����s������D}\���*��ɓ�jhmв�}�O�2�a7���byO�a+���	3H?�)y<������$4�yKɋ���L]ۤ�o��D^�q���#��嶯d�pɻ��j�E0�?nH���M�F��d�iwX�4$6p"�O�ը�Y�J��:��	��H�0�V����~�-s�6�Lf�����N3�M�ѦL�\ϰł��:��v@wH�a]غp� O��{*k-Og�zq��Vr�G� ��t{}#>kj�.�F�l���fŷ�s7��,�C5{�\ĥ(�9���} B=�CEmʫ�h���ƕwI]�ma�W	�R8�2�q��d�J|���+^-ܶoKDQ���%	N8q�I��e�����	�����e��z��͇�C �Xϥ����y8�Q9�@n�VW÷��u}�97d����෡T6nG�%�HW�"�$�Η���d��J"�x�N��X��_:�����g�w?�2ʎ����i4˜�}4�ðeR6��xs�ȝh�?ˣ}e��nL�?�X��6;�f�^��O/��pLA�����[���߾�=�j��f�_a[<R�pZ��Yt�Ÿ����:D-�d|��r��q���K�soǢ��YC��U6�Mݜ�ނt�97�O�NP�hV��D�(�!Oeq,�b�j�hv9�L��F�|D('kd��)�K�{�� I��9���z�&��������q���7^7UA-&�㦃н\h�$&`������3��4��5dPG\���C�u��N�=E�̨���à��8�rI̍�ݕ�9�>�^Z�&������/��jT�Uk=�F�R����`�:�� �ٍtج�^�T��%���N�4h���?p�d,x���^t|D�l��A��{J8����Q�憁�hV���7�䚴>�T�5c�HQc�'��_��A �@����|���AJ�Y��I�2ilq�2�jF(��b��E�),7o̿v���;�Q�d� `)u��`��hT9��/u� �x暍A��NI�1�9�[��x��%��,�%��mЋ�B��[���>3W�I�I�x_q��h�5p�(��kP*��jY�U�v�x�>����R�u���o�V\ī&{˗��g���(��S��g�9fo�w��<:���.Z��M�	r�E���Η�뜦��n���A����ЇP�!t��%����'P[T��Pn��V8 ���ұ��lV��G�SN^m��x���1��/W9gI����2Fo�S����wv���ۛn���L��ꤥG�(��0������GZ�M�I�ÍHe������=h�a�� �i�Q�H�s�� �E�m@�r��6(i�@�s�lt5Pȃ�
�o;@<yl�p(���V�Ŷ���y�Ǔ��G{�B>v\<�B
**z����_P���ױȼCMVk��+bL�c�VI�������\�Qb݇�4����da�&��8�c(+|���s�v���$�X�ֳ[=�M�
���p������v�����-�'��A��E�K
�&�O�RB��_>T�^��t@\�21@p�rĆ�����\�;�
�6��J	�)c?��D�.��y�l�m�R1Q�q ��J�Kk����;���?�"w�/�V�\���A�5�e]��{Td�l<Z��b�5)��G:���� B�)z��r�*�|-�V������W���Tsy��TZCȾ� 0O��P�X}��i�NAd���h��`c��u�!�����}a�