��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\����q�?��e�I8�b�Ǽ$��"����ׯ1�V0���m�a�I/�$к�Agۺj�L�$y�m'�&�,|�\û�m~b�HaDZWm6�J�}��eᙈvGJ�6i�w����A*�cדz@�����N���{iK��/�jܼ�JU��b��n��U�#�9o�v�:pF䡩��,g�"�{��~H(��M f3 ;~/Y�Hعf���f��h�ݪY�����h)�u@�UÂ���(���24a0vʑdB;�8*[C�%�W2|�����Vr<� ^�ˮ�����n��\�"ދXf�N���̛�6Nt����S<9ĥ(ޝ#@�b&��֩������AQܮA��/�dn5��ͱ�t���f�[X�m�ׅ9E��ތ�ѿ���d�G�peC�7��~'L<����)swJ��d��G��4O{H_�Zf�
���* ���榇{��H��[ޏ�')��Z��e�+�n��S�ɨ޼aE��;��)�[����;�-=!_����RV�������m���N��ܙc3�׶��	w��)��'�(��|a���3X3�>�ɃN嬷T�@�QL̀���$�Y�S�N��P@s���)�D�MgY1�:ކ�8}o�ak��|��aĹx2dD���[��)�~�(v���� ����ѻ����
�j}��,vUG�W�~�F�_��Q��J� >f,�䯯(���|C�gZ�5T��Q쀾�]�1�{,�aH���j���6�7�7��`������q��"�l�5f߻�w4�|�i�=�T{`cF����De~@	t����R�f�����9�7����t�/X�M��z��b�.i��Œt+Jle]OK�،�JKn` Kي�Ҏ���Ag��o���T�0Y}�kE!9xI��x�����`L7�4���Fmtb��{�C��4��4c�_��-k�9�j�>������V�ӰDM���xK�"�_?�H�����|*F$d"d��#��&;_Y�6~-y�/6u,*���,���՚a��c>F}�y<�=o�7��b�[��AA�E���޳'�p��B:#1��uۖi���b:��:�Մ�7F�#,K`WH����+`B�g��ӷ��Z�.��Mق���˺�=��X���\�]����
ێ�we5�ap���MA����~?�������"a|#��@���>�lE|�ӓW�	����`�� �gӹV,�:?t^|n��$�VW<"���do�M��*�cA4̹ $�;�`0"�1�Z���ö�SsNb)�l���s�%��5 �r{4�}��.��4S7'��DMiN捑^%����Ub��dp�ނԂ�������Bi�B��~_��J�Ч|�΅z&��&�g���W�p<��*�����p�'�h�k�#�hh��t��ջ�%a�L߬���o�ü�Pffr�j�]8τС��#�/[�Ge:�hl�|N ~�Tr�BHR�����W��X��ew�r��b��o�l��W���+O�ːohU�P�u�/q3�iZCƛ����7={ ��UVTq2�䂍�Q���0�Qf����񝨮ڣɹU�I���z��O�ne+�͂�}e���C�Lk�>sG�J����eL��z�x{���?1?g�؂��c* �^�UK��TZܜz���	�n�lg.��V�|$�]�	_��fӡ$b!h�<_2�F���N��7�Y���~7����Ѭ����b�[�OV��{l�Q����y�����dc�K��4���H�ݲ�F2P4}�該|r����#{��Ѝ��C�qgC����!�V��ت�]Q�-*��D�<)k�!J�yL{Ҹ8�O�Q�v������	����u��`��d]�,���ґ���c\
���RS��z�^�9���x����G^�	}-���hZS�٪�'�g��3�y��y	~��0f��;gH�*/�qq^��	�=�);|.$+�2�As�����"KAV�m'���Lz,$/�/�\!�#�[(��lBo����kj;��~bQ᥅Z1�������wų<#_�����2��SW�Ve=4L-��_)g�!����u�@أU����ʡ@nF���H�ߢ�/�*����7��p�	c����f�� 9�Q݊�[�E���4��s��UzWa#R���hd^��<ʯ���Cpc}��̨��S�	2�I�ˊ�Q��C	��T����Q��f������(��������<Q���홞8]06n�O�:����|g�:�I}�dKҽ�?�w혊���l�OC�%�ϣ.-{8���P�3�����},���b� f#�������n��J�JZ�����g<4�a�o�.L����eS��ܨk�7�-Z!���� ;��&	{�ל�=����7	�8!N�$v�z�
�/�� �3�B�H�Z'�:`CN�87��jޡc���A�*�����+�/~n=��7�g(��j��*���ܨ;��JUt�
�G;�]����$�s.έ��$ZXU ���R��k�Z%�!Y����w����k����_����xNL�lЂ�v�C�Č4r�A�3^q��k��`W|n�E�F�[��ʲM׼ɺ}��_/"[��7���k>l��c7�4���V\�4G��^5�g�0u�69�����]?ß@%}�˓X:%�؜�0ɘ����D��#�~��=O<t��<J����I��S��ftT��!.�{���M˳x�ط���b�|�~&�$$��A�E�܋>a\0����8��L�c�-f��6���qO>�'�0{�v��ԋ~�
Ͻ�=�-�NĴc� ��ΐGӴ���6��ӵ�:W`�CN&	bfR���A�?���,�zL�?��r��ؑ�����&�ǡ��0D������Jl�>��
k��؄m%�L����z�Xa�|���?�F�&����LgZ]%�_�Y��~�?�L�Y�-�GH�;g��`z<�i�~LD��_Y!U9��W-�]���^���|�����(6P� |��K
�'[I��܀R[L�q�O�`������غ~�j���έ���[\��w�_�0�����~X���\�ؖ����p��y�2��.�,�<sb�-�����j�1w\^��c�"'j]U���Z[~C��A��hs�:��9�ʤF!<���#�S����?�#�$�l5	<���2���ysc�-Q;�g�u�ܻ%h��`�����*w�q�ޒ�'�o�"M�,`p�z}��儕8�/i���m�	|��C��XPPN�h�@�d��b�,�B�x�7DAm�h�G:
?']:L{ �:�g��� ���r]?���0�Òl$������Sl��Ж��O�c���H��B)�o��t�)�"ŁPub�����PԳ���'F�e;Z=�{ȔX��c+\�2ϴZ�u�G����C��ȵ��W�~q3���R�H�J�if H�adC�h��� նW�w �b�Lc��IED�?�F���7�		���w����T|9�oΛfq`��o��U[?S�ۭ$������8=˞~
��3���h����;���D�۪��t�IrME�^�P�l\��g�E�*���:�_�����&��nh\�a|[[�WƆ���ε	�u(oHGkw��&�����䶰�(�JQ�}U����'~�$&(����Y��9�>:�GВx$�!ܘ�_^��-Y�y�ݔB R����ݹc'��x+!��d12(0Ie9�����c4@ʰŮ%��>�_|����]a���G}t+(���X��˒�� �S$R4�lf
��V��ݸ����EG��>��]�����򥈚x�����7/
d�\E�0Cd׶�:�2��WW�����\ĵ�ru%aG'b� ��{P���+i�b>(�o�ӎ¡���X�h��^�{��_�ϩ:ҋX ԱM���>E�(=�&	����j���]A �bLg�{����Y@�;@����m��l��|W������E�)�8[~b����t	�E��El�P���N�,l�^	�����d��RV����y6�~��s\?Y�a�+G�ag�n�(��۱�\�4ob�hy(SQ���,混�22�ce_�8��VU�R�S���Ș<Q��lZ�r_�l���+ĸ���$���3ժ�@�H7�z��z"��uj�n]�g�_�"��fU/��T�9����������8���p9��z}pn+	M4�������j��Q8TOV��_���� ��)Ş�r����`��xב1�_Г�uye���4��s?O�4�#�K��`Wq����UU�r����S��5�Q)䕣��]�nʈ^u乔J¢w�X����!n��O���.F��4��K����;p+{3bS"'.���'(��+�rÖ����ft���Oĳ��R�Mq�����X�v�>o�(���#�-�yA66
`��	�14��kh����a��kK�9Wnn��S%_��C�KE�K���������n�ڴ�S��тlWC�V��S�Hћx�'�_�H�+�i3�ȃ�A�9�#�Ri�����HľMo9��QY�#{�<�B�]���`k�}������eooP�H6�L� ����@�]�L��-��!x�ڗ����+&-��q=��ρLj��z�B�,.D�ml����
�KQ>��[������W�Y���'�C���=�.���1A���9~ oa8@��i&�.�B�Ze��p�g��9��qz�q�"F�2��H��.pk�hu=n� ?��|Q����G��8!�&k��L�o	_�E���<�n�����aSx*��R�.��sO;l��u6��X1��K���� ��W���oa��8"�m=v3�V�E�c�FM���"^�` ���D�[tX�Y��R[;&�5$�N	/�֟�ڨ"
b�G���^�ʕЇ����h� ����WA՚��:�C��	ހ_e��vZ%L!���e���E�)T������-�)��ꛯ�ͳ�R�&Ye������e�.;^��i����I���;p֋�{G����߭���φ�ik1�ql��mG��9dS�P;-�p�-�ԑpͷ��7���'^nDPK��ЬI:>R�/W~L��|�_�������Eɟ����N+'8��}��k�P�S���yi4T��bu�V�i� ���fm��C�Z��5����u�����&��ӏ��Kk�K@E���P�o�t���`!x�����L��;E��-Ñ�+{u����ɥ-���'�:�@��������&$���j�,�-ᕶ�t�"kRksO� ����&��6u���ڜ�.��w�?A�TO=~G����\E|�'��Do�<�����l���uڗ���K#�6;`2C�I$E-eN��p_�2=rE	�1D�uo����K����e{�є5�������]Zd��ᶃ9���bKJ/�d�:�N8-L�("��S���c}<����?�֥�*G���V���%�-�hrtd��"�������V8~Y��yhk�����oZ�.(���E,���H�`��60�^�{n� V.�B T����`���� O7����f�Eqa�E�d.�r\1�_D6|��Rm�&�5O��N�ű=��P��v��D�u��wx�VoK�26�$�[�<�LPxe����� )=<��o��pS=8'Q�����������چfx��x�<ռ�HQ�Ǘp_���>%,o�_SD�r���[�����*�p\!h���H�p"PN�~���3\��u� r�&���� Jį��f�l����)����P�_'��+Ct/��B���M������q��*8���~¥rE,*QS�Vd͎M?�г>'ĩ�RO��$���*e�(2aG�r>w��y)E7���a�`8�c�a�mJB�����7�ll��{������7T�?-$��-�v�0��+�����W�Ƥ���ߧg$K�5 �j7CŰp��|�#AI-!����|A~E$_�@"�_e1�t�U4�M[���|�Q��Oރ/d�/O�p]��c��ߘ\DY|M�L?hn$�	y�~�r�{y0k�Y��4�.uz1��_\Op�'�o��>;��ȥ��γ/3�Sc��ޔ�]����K�����!@*$:�"r$��Ncek�-������i���tI3u�N����ݜ����5��h���ڻ&� ����:F�(ݚm�o|�p��ܨ�l�ƳҒ[~0�u�w�!&9�L){��-::R�g���%+t���1������Og���LJUgY[ǮL M���,��H��b�%ĭR��Z�
�BeHp���'��L���K|Y�u�8��|�;Y����'�����]'�n��pƅQ�am� �f0���i�}��x����Y�?(���?�>,������CVM��=���D����lV@�s�b`��g.u`X@��щnDNWC��{�} �n���"�Z	�F����<�4;�r�����0��	��J+߲�B�'�տ�ڝw��c�vy�d]N6y�`�[�V�:ơh��B�w��%)̀ز��[P&�¯L�*/�jÛ՚PL�f�	����+ko�4,�u�0�a�x��sa�˔!dkS�,u����Ԧ�:R	,�iٓ�:�N��2�	+߈�ك�Qd��^�I51����i7W�e��ɍ��}�0��M�+3�CْhU?�[�N*z�y����:	���.�O������:wP+?��u�W)�er��� {��o���=K�ߊ ��U
���ek`�J��q^q�S"�{�k �0X_Ѩ�܈,@��f�fhV�>�{y1G
�W�n���W��?��(�n�%�X��&��c��{c�hp�0���awu3eI2�}*}ڣ�[9�3K�b���XmR1��h+@�IT�
��-�)����l����U�M�:eͨUK�xjim=CE����]�B ���!�0Ձ0�������W�>������7�lQq��5�5JnE�����+W�[�*{�b7�/��g`��P>F��0������6N�s��:~���cM�v��E{h�٬8�߳`��M�[�Cj֐B ��t�>7m���bm\��tj� �C6�)3p�e�{����#��E���5=�ӯ�_���$�������(�v}�e����ݵ�Κ�G�h����NA!�H￶K<��}^�������;H�Y4�4�dZ1���ǭ��}��A=�e����D�_�����3E�YefW�tb�3��$3Z��k��jBo׺!�6�9f�S�Vr���đc�,W,��0%!�%�;�����}��$s)FW����A�����զ��NA�k� ��ʑ6���AY��T�_��"W�(�y6x���WЃ�X���B�(v�a��΅�y E賹)eu�5tUSuP)�6UIkB���s�"7�c>�U�nx��J��E��R�!%�149�;Ecu"kۢm�DJ� ��Nֱƍ��(�*��Iw;8�Z _�l��S]Cv���j�5D'� ��0I�Y)�G��Z5��K���TV34HP��<�Y��<�i�1<����H��/�`$�����~l��EFB�� ��|������+�9�|�љ�K��_3��BY�%��#�lF
eqy+���[s��7�i��5�Wc��<���<����jN��E���n��|&�m���+�l��1X"e����p���*���ϾU�Jo� �v](n{*y��3M
��>��G�
��)O�t�K/��P�1�/�Ӻy�hG P��*��5v���#�]�����>�ow��ݕrr�b+�卺 ���IZ�ұ)���~/����L������I����ܥ�uro-��5Kl��z���%T����M��+�p�*!���-���_�n-Ѳ Yg/p�ӝKOh��S8���s��J٣�<�����ƛ�w�KM�m���b�kZc˕�l�^�՗��1oV#���-��wzRg�%�3��OdªF
�����Ä) ��wWն�:5�d�_�s��}����G|~OM�	n=�K/�_�*���Ud��HH ��9r\]�A��D��R�s��J��1ު]$<ËΉP��2I��P?� �G0l���$�������j��Q&���2	!��Fww�<��6 ���X���VJ��t;����[� �?�n ��Qۧ/�b%��g�S�|73�����ոsr�(0Ӂ��#�k3�}q�7 A �7�7k�_Hr-h�D�C��tڊTO��m���&흚��1!��?�ϡ́����|��WA8l�cĤ�f �����ߚ�7�]�'H����ͪF`�����)��ᐪ�հx�f\����滩/Kž��A�7$�ٝ��Z8��I=k�Aܵ��x��$HrL	��>��r�|��{�L���#�ð���a̾�j��߄8����:�L��]���&y�7��F��x�m^Y{�Y���(c��+�D����9��2^�^��!�_Z��E��?��\����!$K)B��䯾�B��|��Q8+ƕŵ��~H��o-�$Ag�5�����i'Cx
�%+��V���$�f�����>=�̿W� �n��1�¹r1	�:����y&����ƊL:���K 4T9���w�n`�����tU�<��d^�t�3J��<�u~��zL	���R�u~��T�+x�b�z�c�^
��h����#��&Ѐ(I)�����4�N�
ү�H�Ԃ�뒗i-���S��)HU� ���
?�%���-� ɏ���)��4Kw0�k��C6$�m�T}o�b�������yQŐz���x�'i�L�`��W�c;Ea�t�>�
�����_ڛ�ǧ�'�^����0>��F%A0&i���UӲs1�P�Ļ��쇤��780��X*0_9��U��\���+���w���Z�YAa
�ۊ��kz�x�kO~L> q���MD����K������<Y}s$�!�M_�rF�{!�4X�|�bH�To}�����^V@�~����-垬P�Ϫ&#��_�=7D��v�J�8�Ć`���t�ӆ�?�d
�y�2�T��	�<9`�:�X^�E�ך�ۆ��,(�"��o"aڗ���pb��/�C��ܜ^�|*�[�:*[2r����[�@�!��8v��ތ�/���=�#�AI��[�rH�m'.�S)1�T��g�;D0�K��,M��E��{'m�O����|Ԕt�+��*,�!\�)�۽#�[d�Xہ��
�����l�W��7��T�w$�w��R*_��A��*��aW�n���\uK���7*���Z�'���-��xdv��P���{�g�ZK�A Pu"�67��j���!��������O���
ާ�k�6�)ۣ�K�C����C$ж��|J����f�S���I8X���������b]�Rw�{g����0��HV�-]!�^���:�1�"�m��vOe�c~�}0S>J�ũ�!���qړ��x<��JA9`EMK[`��Z��NF �4��Y���a��@R��|����<y�&��,�6F��k�:��CSRR{��JfXg�y`�>(u�'�<�Ӌi�>
UD��in��C�`�y!�$�%���{A�Y1CH�ʳ���XO�m��+����8.
	r~�Z�W� �����ߔ"��dvC�=���'�v��������"k�B��w���;�J�)�@jʷ��@��B�U$;vܞ;vYKZ��ǹ ��:��IZQ >����)�F��q^�`=����V��R�\2�4ӟ�]���3:�A��Bb�W���ǦW��g�c�H��^?��+�e5��ڀ����#L���Ʀ�H|8���������,�L���iWW�7�"���(lzZ�Q�/�������W�R�qz��R�3�0Ob�4����̐VRq�:���@�g�E�'#ǒ���H6�x��a�����*H�P'�=��W���Kp+��സ?�H!>	,�O�@���<�7f�s/�!GT?�K��-�)�9J���+���5����jwx	"��ޗ�TQ���B�TQ}8��
=��:&�K)\�^��L�[��t8`��{/w<1ʔm�}��r�%�$}J
5�Ო�y�=Ǎݡ`
�JObf寯�ܼm1B����b��e4�x��ƶ��봈�� �J�:o
Է��*���sPYZ� �}�)H�?=�����oܑ�L[��z�A��S��2S�}J}����P	זň��_���4e��w.)�%�1�u�����'{��h�����dk�n��z�A�A�N�S?���!貟��;�N�4�a���Pr**�{Р�!�Ω����|b���u�'�|���� �Q���0R컻c��8�r% <�z��=R�b#VH8�:���u�y��6A�_�� ��#E�>��zQq"�&���d�+���	@P��)0K�g�x�
���z䅰��3@���v5�}�O�ؿ�����1|�U��H��}�R�A{�5�t�(�4Nb�>��6��Z��~ŞAh��:Q�4䨫H�p��F6$�KM��Ƒ|�Jyb4�<��2�攵nxp#f�Ҏ���FvT�œ��s.�ohN_9Ѡp�}w�Z��Xm�wE���ߺ'�t���+U<P������q��c��n}�j�u3��c����]�8��L�r��z�c�Ċ���D	]��[�Rp7~:HE��%���qf����T]�whO����>��=7.\&��$1 ��F���z&�L_ǉ������(=&�8I���/0�M?�a���u����n��p=��K�O��]�Z|�.�S4��2� �A9���l�Q�0o�A]g�t%=vG6E�v��,����"�ؿ'�=ɹ&�A�G��HZ����3�J��@C�p:l�jYm��)�1M����G�!�f�KBo�@r�E��E_�x���V���̕�D�Σ ,�-���{T7#�3M��j�ל9��n�QN��<T���m�Q�{�mU��ttx�t���?���7�/�l,A1���5}���y�G��_{;�*0=���b���TC���|���
�P�
������0M��v�B|#���a'��;%]v\a�U�ѓ���a/���#�o${aW>s��SU*t����PP?�XjL�z_J�{% �����d�0,Lxk*�rú�#�8�k�e��%ХY  ��Sd_	����y=���
����8&e�"iR� �T�E���X��+�R:��G��0�8���?��j0�ʠw�x4�N
Bq-ㆆ�����Gj�*����.�@�Qs�lH��z�j�]9a{%�6��E6c�%^M�nc�%�I�5r����LV�7"	��I�;�i/�I�	��眦�=��i�غ1�%�E���6:���4���L�(J<��5��F��%�{Qd�@o�������l�f}�"1�r�� ��i0mO�gdN�R�҈w̻�yݼ�}��v��e��k���<Bz�b���1��I\�Rq��_VR?ё��j
K˙�
E�`�Q3��
^?@��D=�[�kao�'	�� ��c�[`)��o�ꁙ>���K�!hJ�5��)�����I��P�@������_B���C$��9�|���i�2A�ek�_��t�[�*)tOGE��(-�q�Uy���c@X�_(�1���m��7O#0�%�\�����k��A\
�a;�"�S0
�±f7��G?=��O�G�!��?��,Ra"������wvۑ��X/B�d�<sY�
H������XX(�L%7��p�=_�T��D���d#K;���C���KT ��
s)�0���'S��sհ�i`�����kv�Ӯ14�s5(�t�,�"{�|�Y��3����`��O��@��M���s��C�+��:�2c<*�ޙ��w�BR显�rt��P�A�\�yW*,3�W�$��STI�`2t���J��+�������]CS6@�5�[�Z��<7���{�k2�ZMz����\Ǿ��#�C�����짣�]=�'��ԅ%���gr��%��֠_J��=�{��ͩt ~u��O>d�[�\mq'-���Uv�dq*���)�D	�Ӥ�CO�����S=���2�vn\p�8�����鑫z:�!hC����9A�x8�Xl���kۺ9����X� ��Ћؗm�s�KۭwY�;Mԓǚ�&�n��%YF��u�C��� ��Z'(�� AV���^L+q �'�ϧ6ש|h%���l�,����������8��,]j�4�㙿����<�h���wH�b��}}�ƛUs�N]H�:��Xw<��P�X����Đ+�7��N[!�(f
yP~��^��m_n�$��]$�6gw��G��`���KLs�4WjX�.fv|��F����~�6e䚲�*�GX��=��9� G�uSn���?��;>ֆ�x�O��c���Pc�} }^��L�u�>9�~����F��͂����n�?~�>o>1NU�n𔟻���p�1�����sp��^�x��7:�Ax��t��j�S����yZ'4A�Te��"�a���I���z\;F��^��qJ���Cz����Xag�@R�N��i���������ې?dUp����B%!�i��5+�w�7~h��[�Y	HP��ipJ�ĥ�p+x	��04ẫw{/.�+�'�c�᪸wg�#�h�����Q����=<�뇰kN(������<' �������'�����'���CFod�dK����/��G�.�7+�]��sSUJ7���ً۩AB[$�h���N�)V����Oٖńp���)�jjpҨ)w�s<��)8sp�l;�{��t�5������>�� �9{��7j�%�u6���������)���t�W�Ҭ�j�K���ζ�ZI7`��f�N�o�n�&�l���b�LO�/�SK�+<JX#(o��<U?o�k��
��s��&*͌�x��8T�L(�Tc��	:�J�����4�����
��&�L�&��<�|"���3�j@�0�b�˳/'�K8�+���)�S1�H>���E~ϢX��p�f�w���o�QԌ�E���Tܔ���|>wG�[��Ƈ����z;e��-o�������7�q��
x�i���bq����-ƹ2��H�ö��<W�(��la촻5A��f�'��vSね7/��%[�_�8q�櫡O)�O���ѐr*}����sTa�hoi�L�FW9!4ld�2ph��i�/dm��;}̶\aؗ�}�)�]I�ŷ�+uȽ:��c��T;���k�z[Ar"���n�G6�J���!c2a���e9ѻQ�;�����;d
�@�_�ާC��"�p��0l>��4����.���	*_uѢ=)w0,~�����3�,_w9)�v,.X|Lu���ǌo���Y���v<$���Lp�exoy���c0x��Fǈ��fB��� ����gHyw��d/ܽ^�1��#��d ��X>A}�>3x}^n-�����+n0�����4���+`�%#�ɵ�IH�i�N��QP�ܪ�	�#QZoV�n6�g��VJNZ�+�RE����5��XZ��O'����0O���(-PבI�O��9������ �@%�6��O&˽w�y�׹ڱrB��G$j���6L��lK�ɾbhL��3��O�!'墨\D�Az0�I$r}�*:�m�;����|x�gf^ɪJ�a4{�S�����b�ķ��t����&�u���fסo7�]��P.�z9��O��������o]�Jg�1G�t|�����|.��n�����-U�ζտo���.����%�(0�Gg��FC&q%6rR�@p��*<|J	ڀ�����o[X�u���i�����<�({.v=���|���1�N�"~���V:�>1eu�CpE�S�T�ZO�;�'�t�.����U�@6�!�����w	�ꂨ��I:6����$��4���U�C@�~�?� �Mg Қ�%��n"�G�_�5`�}�4�L��I��:���O�Q�RF��u�ǿ�g*=� s f���s�M �H�Q7���,L�֑f�b�|�`��b%dA��ܯq���p"�Z���^gIw���H�� �O�tkA�P@��G�B�.���[�
�?�`���Ơ��ش�������)nv��~܎_�>�Yb�Ŷr�-��.;h��[ŎU���}��~�u����J�h�@n�w��s���ܮ��~)���u����J�0��7��ߋc~�[���2��#�,�q�[vb�[�f���")��M�6��Qei��31�c��>��3��ِ�������e�=����v�$4]vٯy���4̲���1���Y��X�>pUo���A�bFՕj�I/C�a��=>��K��T/�FݛUčQ eA�G�,�n�B���*U�2�I;�=�_<g����=��꽔B��j��fK�?�+H���v?�1���cЊ&̥F>��C�uV�(��C�X��T�#��V� � .2���w}ng��z_���&�������ɬ�� c�T�B�w��5�v9���hFt��%Zi!�����]#�Т��X(�TQ8g��e;ܲ�:\r�Y�I�6ME�l�Enl@���՛���Nu�C��]Pw�]BC�e4���TQ�D�C��Cd��I�Z���J�w0򲶫�#��Zl��:m�X�������C�h]Zj��f�T/6�ˁ�{(�=�7�3����?�o�^s��'�H����i����SeR�xH���b��m�����)N'�h�]�q��`�����u/�񥮣�?�!a�&jg˼�d�E�;U����(p]'t9��&ww���{����>n�XG�kP���x������J@ �z'��,��Z"�Ќ�}�RH��%��� ��t6��.65vڄm��-���������p�@�t!�~(蒽�q��HG?+��V�e�� #gt8tm%��˗zO����%ꪔD�%�R��hE��H��)*�ztg&6[uQ��w��W�lgp�}�P�G�c��{G�D�v^9H{�8�9I�T{�����ޑ(<mRܷ�� eOp��Я�P4�0U�@�(4�W���4�d4�?���OGKH������`�+m]�8�?�
R�W!�B�ð3�D��c5��ބ�
v��Y@�����8tXB�&f���*�s]��69������Z�}I���Gd������)1%V�Q�q/�#J�:rG@���!����,n��z�&�B������J�PtI�D� m�Y���6�A\�9`Zgwt��%�/ �5�n����c��Eer���qˢ��$��w�!���k��[�竫ۙ&���.o��k��ޑ����^��''W��G(�3�)q�&�zQ/���#SeC19M�ѯ���l?���we��c7��A�L�����s������/h-�L~������1 ���Rx4 }��0�)Q�pӠ(��(�ji���Wk�������11F~��A��*�6���Lʄ���a���_�zKLT f2��Lx]fOx5 �N f���t �I�,�D�)�%v'ҋ��A�Cě�I�W	}6y��~`�ă�������n2>����s����A~ouU`�au6/��uy@�P�ŷg��I3���Q$�uЋ V�'�3�K8/� ��ku����rKi��1cdC�������K0	6�{\'bFsz��v��^!}�ǭ�c�"�'%E]\��e���47xn�SQ��,ڛ\�g�}�Y��9��R(^G��Bo.bZ�D�gH� ՀX�p�"���3����uŵ���D`�k���|����쬍d�(�����!Z�M	߶�����~qGt�(����{�6�VG�KA�v��*;��x
p���K�g������W[���j��\Ȳ���: ���������l�}�Y\B10x5�K��^k��X��<v�o5�S���J��eb]0WT9�{Ѳ�.S��>/#5��G-�������rr��=�u�X+<�N!�+my�Z�ezB�鋯����N��Y�~ ��)�Ö���'����q�S�m��:�/�]X}�RdYfA ai�&�O����"hS]���*�X�81�q2����)��7�ub�FBmJ�7M�����$S��CYJXf���bK">I��	j@E�k�K[���G� f���
^�Ix�2W	��Ԅ�<�3�]�����W�%9���ւ��E;���eCo��a�ix�h�>����<\�ֶ9��S�"��9r�^�s.�����P"�L�^2���Z.��\4B�H���3���|H��_�M�L=�S)��y �B%L�-��6��YW�Ŧ�V�}��#��[Cz���K��V`/�3���.AFa����/u�o�0�\�nJ��n����q
a�ao� �Y6o{�4x�E��S�IY������8���v���m5��r�f��� ��������e�U_و�w�jHL	�}��3����Ƥ�ϝB}��9��⩔T0Kz�1�]��@�ߑ��֏�D�_�m\1�݂a���U�u@�w0�Q#������f�B���z�5�f����Kr�f!���G@z����p��&�g�-r�-Zԅ ����Uѕ#&aoegA2��cПf��o@M$�6a�%��̶�*�V�O&J��n��q���h��%a]w5�������3���9G/�4I2�h7�ez��:c� иއ��Y���s)��d[؎���ZX��!J���[�|`�3Q����w-29�pA�,93pM�TѱsB���+��uSb5�{�����f��Lx���;��	qՄ�Y�^�}�������a�rg�(y��C&$�B�R#$g��Eu�Qa��W��Z2,�/lV����K���E���4l';�=��K	��?��I�Uܛn��S"هg)�(��@��mK<���m8y~:��e$���h��ΐYe��m.�ˆ�ln$5��,��y�c�e�[u��>7,���x�0\`��3�]w��#��Z��\�C^����J'W�3!�]�.���Q��]� 0xMx�V���/[=�#W�j���j�DsN�2��Ԃ^��yr�s���<"�p���vR��0~63�W�X#��[���Ц�
�Ml��� ���#oh��p��u{��&8Ѹɴ�zW�ә���� H�m���FbW��@���Bq�/�K�'NXI]�"�i7��h$�~����ڍuu�3uld^�ol���K%��Q�~��H�l#�WV/ƀ�~(];�Q��Z�3��j.�_����oK�Q��Q�Ch�|���#���\_F����ү�c\�B�W�͇3.}���D�ɈE]ə�8���.r�p�w�j�y�${C����yȤ��G��Ю����ֆ�4���y2t�n	�ϖݩ[��%1��8p�?�pr)�~�����y��Ii�+�A��0(x�j����B�\P��LZq��`c;p�e0�<�;���EM~��ͅ$>�gߋ�g�B��>�rS*i6
�7�B�+�>�Y�55M�����I�Q�%h��:�u_�\��BL�m���O�kZ�2`� 0�W�s�X�����r�N��Ŭϫ�g��s��!0�4�ȝo/9.Ѡ���I��2��<f)�.�c?�6��"�P1���N��"��=�L���k�|�����d�En�Y�W��d���R"�������,A]���Me��D���ϕN�߫��T٧�,�:A˲�W�Wg?�\����3����$��?4T�䝶���y��g@۝��	o��E�A˸]]�����>�?�ή3�l�����_�4���+��Ѕ?��'t�NJ)P*N�JJӀ�t�L���j�_Xy_#zfd �<�Z��e�,�/��ӓl�e7��@ }�oR{���]6l�&�CѴ ���>�r���F���Fj��$����Zɧ�Jm���*/����A����_���פ|N��y�S���t����9`4������z�ޝ��]n�����
�Q3�h@%j�$埝1�o��=\�q�����%Oad�Sﴜ��KhHp(YRL�SvS���d� ,w+q'�<G<o�2=k�휚�Y�h�w�� �K�E�z��Q��&R�`g�/���0$��7��iq��M�7�
�F�"d1݊o���|խ���LH`Q�4W�j���^4I�L�����Y.�� ��$�ä1"m;]�X��ڝ�t�z�5��9�q"��6�D�_jp�D�;1_=��@���:��}��2S�b.B�ۆ�]�~��\���l�[b�G��f�7)��)t�/"'�*q��[��3A�Z�J�'qjA+WI�������t�q�уw6v� JV�
�>t���|����0x�tgvUw��(x�ŰY��s
6C���[o�E�r
�m�|2���lHV0�/D�yX�^|�25��n-�?�k�b�孡5�MK�5�W���[J��R,�G�IN�9_ҁ�W2�KJ���� 5��/�_C�vA~�J���y�8[#�ն�œt+X8~�b&L��7'h�rQI�&~��l�g�;Q��MTq�/L���O�^��!|��Żn�]�$~) ���b�
�� �_ʡfa�V8/����`F��z��L
�=:n���<�=����� ɥ�Ϧ6���˒�I�IY�ΐ\��M3�}�~�6=�A��=�䓴&��=ې���o�F,�v%�}��Q�>�Q�.y	�.��ҟ�P�/�$ˎ �k~uy�I�v�2}��Q���=ar�@��E�Ts�N��J��.�2`%Jw�tA-Vcn8z�~��3�y)�|���7p����0�ZH�f�4G�aV8:��Mb��<q�)�n�㵠�hi�ye�����X"���n~���}��e���S�~9Tל��ړ�o�ކ�+"(��t��}
e��a�h�\�����s+�XJ�_W��وď.�4��f�����_��}m5�.~Ԍg���*��N�lX�l��p����Uǵ�MP�st��+D@�@SF����?�����!��bj^����H�p�.╞-c �H��,����6d*M�gr�aG��|���DKER�m_��N�⢻�&ո\�G��?��	��T���q��:���赖�r*	}�;ayA�E�=z��(�!��D��\��=����锑��P�ĭ�|ZKךW,����&S�������k���&��U�O�⹲�����ཝ4Q{���,g�J� w���bʘ[�'^��䜞j��(̅�Ѳ݋�nF-Uw�}�{���xe@�kP��x��t��f�h���Q�G�:+-��  E4Jׅ���$�fQI���+�7��d����{��(�����ȫw'�е��@�*W93���-�.u�o�T�:���	s���'gOJM	1��U��v�"��mT򢎍l�3�90s��%|#؁EǪ������M�� v;B�� h�/�-jCZ$���i��	�j�]��ͺ(�X�@x7,%�\� ��t���bb�j]����jB�R�k� 6�fTpr��%sS�Յ=�Ӈ?��
��¿Q������KQ�_Ѹ}�d�t�x���ֳ=�A�41��:��|G�1����NI�z?�DцE��x s�`� �`<dG��[j���o����b���䚀
��'5�߼dU_��ƞ)\;��t��H�M��8D�
"M�d}��{E��v0i/z��;0]��(vG���jy�#��p�N�!�d4�M�&x�w���k���?U�|D��$U���	"��T(�a�6L�Ri 63��DA="Q��;�?�؀��ls_y�,I���7(����X�߳p�D���c�K�?.�A��e-����!JKә�Y���gV]Ì5C>~��G��'G-��c��7P)�yT���7*,����k�V�U�E&Wg�ۼ6�r��G"�j� ���3�{�P��olz�ॼTF���d��@X��QS]��Ü>��E��D�.C>���V\��R��@�0!�e*�#�G��XFK;���M[�0�@y�6Ϛ/�;�;�GM{�I%���V�FWV��:��Icfʄ\:�h٤l�&��^H�x��&��M�`�����/�tH:���r5¿s�&���WE��)~_���/-��n�S���{n5�w����l 0�~3�����6�M�{6YO���~ۚ��/�XE:k��so�`�ҍ;�y�Z��1ͫ�(2����ߘ5���Si�h��Q^����^L�A�����U^�Q�zT\�H��@���k�BZ�+���)xhd_������F������g��;7R���gldg0����pR��-U	��H^"�A$���C-Y6�ڏ����� I/i���Ej(o-Ng���&/J�,ϧ��I �s7a��0��f�����H�� Ħ����p�p�>����Eݺ��jLC���z(F^���j<^�&�V�ΣU���L���B�Q�y�jH�Ԧ�N�ؿ>d�A��3�ѯ	�%HW��5Φ�k���dvm��"�����_4 �4q�
~y�&�0KUJ�9��BOOp���z:���H_� ����wb�"���ڬE��|�i,傟�VF�����2"��`�wS4��ׂ��c>�sc�yN��(x�z)�|�����mo�
���B�-A�Ź��rSKԝHvn� ���
�ڌ��߸����N�v�%)	^��݀�h���а�L_��;�pEY��%�(@0�����J�bW�������""�c�>�`M��}���8>xynN��J�y���vIB��g�@�lV��Wd����L�|�e��R ���~ϐs�x�e���a���ė(�ϒ��6�=��mj��� �a+L�L������pĖ�W\�8@�dY8Z�}�u�j����I�Tb+��Q��uc[�!�Qm U�ӟLҍ�N�ꯁ�srB��+m.�Yh"S��� U��0��M�Ĳ/�A5A��&����-G[����7}.nf�d�m*�97a����0� o.�m�fA}B��Q}��N�`G�m�����a��)�2�z���G��+<lD�����D
:�O�EhR�y��@E��E���2�3�]}e'L緛�$�ɱȴ1�JU�t���<V'"bk�"d.�C�[�D3���Y�?��mT���|�*���OY�"996�B'��/��ޏ�\qp�KKj�[8���V��w�����H�F���+�'��".�4�Sc"8g�Q)�K�k�̊���T�i�r���oW�1���0��!�)lu���+�4��i����(�Y���	!]z���[H��t��;�x1��zbv�h��5ֽ�w��âI�U�nk������:�[���A���0�|n�B���L�4m$���DLå@�+�;� �9��H���� K���G�	���跦��T,��Fb�e4��O��e����<f��D2�R�5�LԄ;4�(בtK�3z���1��"�X��AFQ	.��|j�'͛Ab3b7�f��B"7.yt���1
yW/���������ߋTv�?T� Bx��j[_�t`��[���V)�i�h-VM�C�*�������fu��U�` �C��+��>��5E�M�&�e,5����#lB3�H֍��ϑ+H�����x� y�F��]	}��7�9��nV��[HX;
O����B������Tۼl�2ΐ�#/��aE�*&tɒX��<�R��k>+s����0x��Y2���ۚ�^� ����\������xc�y��A{������0f$95��8��>vE����f���$Ո�)�r�b���xj܅�����~�a4a�uw�̍����dU���-f���9I'/�@��S$�Vi�b$/�.��&��0Cp�nb��{��]WA�.����;���L�#Z�WT��3xfa���G���V�X���h��v[Ҭ���>Nr��g\u��>*�N�L�Q�����l��a�7)���/��Y�{���&��G}f�A9#����f��P/'�*��_ )T�%3d��29�og� )p\�@-ɴV�$��#Xێ��h��¥ �]
�޿;2V���"aoc9]�w��7s]q*���Ǝ��5�Q8��rB1d�|Q�ɤ���.J�صt���u ]�ͨ���h����c¦s��B����O̡��S��Ao���[C��Š��C�g��������3}���ߋO������C"J�(��(�"l�`�G�-���x:ՔU��D�.���b6b���&Q�.�вZ�R��3����z2�}����"aX��O��XkW]P�T�tA2B��-}>��2L���Q�7:����)�sW� [��F���_]�ve���#��BvZ��d<��on��&x��t��Z*B��EӎdW�L�	�^���qեTP��sJ�6����τ�!�@��Yk/+�F����2+��7�!psR��;>�C���3���kW`�(�9�~G���4�㉬&H���?��~R�^u���w���u[-�*O]�&�?H���N-�	�r@O�����i��/�|�ӹ�|�#��wWrtN�W�>���]��goD�z�0�FU5�L�ߡ�_���4���$h;V�1�=b%LKY=��E��c}� v$�f�;�������f������M����r��m��A���\�zY�l�U݋�I���4B�K:@��<�*�A��O���*1�	���F�	<)`����ļQav���������R���!m�6���s�%�@�:�9�Q����Jgx��s��g�"��cp�A�A�Ne��#F }c:r_�i��(����xS3��͕;��{��᱑H�\D'g(]�8>	Hm*G�@g}hP�C�Z4zp��:�'�U#M}8:�~���IuA��OLW�R��=?��!&@���ĽU���]@'�tu�	Q����4q
��/t�w`':���ճ���ł�7c�ۊ��E}]�Z��y�	hqď9�;�W�[��t	(����T�-F��;�sD�4�	^q��!<Æ�cAɒ�u��������7���B�A7R�>(�d�	*��~���U{=r�jl�D�N���~Pj�6z*�ھ���Z�F͸^�IN(u��-���~��X:�~SX�;�4P��5*]�]�h��9���}ܼ@ϟ��\k	6L���77~�W��c|@��5�i�$f\ҵ<���Q}�GK|��U� 74MH����݇oT>-����3�c�����:���"D����cr�ʾl���*	V�Tϓ��x�M����U1VM�(�ٔ����0Y��u�����P���?��?�J��b~+05�/}�>�و+}�jL��\&[0�~] KH��k�H��@s�Xc��l���1�=�Y�16)�T#1��0b������\��%=�Cx��H�9��ժ�~��;��.K���:���]9s���s3UY#*!���ȍADH�ܸ�L:�%��Yh��b+��T�!�y/.������%L=-+x�+2KN��T�ꢪ"J��F�8eQ�:�]]ux��>�$��RrZ����`��)jR	��",�R��qa@�N+�8ȫ�)�9߫2-�x٩�kR4�i� ��0@z�ZS��*��)_;ǚv6�����op�G���z]�| k��1i��F��,���	9�rUS�S/\M������Y!��=�JcT�c�P.�cg(��/~��l�:��[ۍr�#���13�"�����Ku�K����D�no6\�~n�e�L5�~�B�1�$bn�fS�0�෨��M�9��`]����r�㲇�� ������-����敾���bYXZɄ�����g�`  #�!y �|5�<��m+�IuE�uy�	~�`�� +��ւ)(�QZ_p��I�Q�KQ�9ݟе�n��T�Gc�Vvc��<������ڻ�A�as����]d^-R�@C��̿@w[Y�{z5��#z6��Ȍq؇��w���3��Mx[i�;�4ɑ�P�Θ�Rp���M�����i�<�q^mŖÓ�g}��zi��t5�h�
V��k �����5=��h"98�y-S���&̚�1�_�������Q�Z٭W����wݿ��|~�[n��l�(�~5 �	S$݌D�Z�_�ʑP�V������+p���;gz���h�E3p�U�%\�n��u�"�n��\���ӯ�����Tq����JM:���e�o�E�*D@Q�MHz�C��s�T�om���E��]r���^�BĔ`�9�|��X�
c	řz�Y����2�Ϫ�h�Ū�Ho�IW�4� �_Dd�'��7|�+�jF�	 �o]v�p�2���q��q��Z�V����$h���S��"s�P(��B��\{}�	�������V=�vIG�b�B&Ӹ��"���,�)6���啘9j��u�H����R�޼_��,fn�A+�T���znkR�_�~؄�b4���V���Q�l��c-�y���|��:����qd��Q��o�+A�v�0�x�:�@� !��������@Rt%�4�3�&.���r����O :^c��\�4^�`!�rS;�'�v�(����!d��H
8��iuw
q>�^��\/���2Y������]�= ��?V.IIT^�d�W���su���^�6t����׃��p)L�Q�.M����^��\vj��M(,�c��������"��o�Z�s���bZ�g�j"���/ !61^Ӣ�1KX�I��p�0W{�?[��3���p���6�E֠�ʧ^_���˃nǞ�q!����GB1��A�mJ�a�L:H���R�od��������T�K����n�zt�}��3�2���wo���۠l����~�2�PB<5SH�d�f�,���ZB��&����ι��M�M�H-��/�;�m�``������ޣNh��T6�5�h��ڎ'c�ZL�@&�9d���1̻Y�����]ZeK�!!�\����c�[���,k7���;|/�I���A�H2Kǹ8�U#H4����L�c��k��Ӌ�iN�?�%l�A4�����}'��|�8�'�~)vѽw7�^��0E��B"e K�+��U�� ��2�ub��"���Vj�U��cw$�������Ca����O'7�w���#jJ5£z����|6f��j?�W�����U��1]�[�m�l,Z]�MKAՂ�I�2��V�-���H U]�.'p�L��-'9����?rz\ʋ��8��vT��q���A��t�[�(� �PĦ=��l�Nb��M�W��Ǒ�j/_kT� M��9��j���8�
W����iw �	�҅����-N�_3j� ��*b����v��-��e�~�㲡_JI���B'd�7�&?����D(]�q;BȐ�E�.�pU�����u��ጜ7��NBBD�l�/ K@�4R=P��Z�� ೧]Fk3dVl�M�\���@���z�L���W���Q�K-��a�L����݊OH����S�����v����tg� ~�]�����g9�F���n(o�[`W$i�V����΃&�o�x!~���0E�AS�V�B"���m��#Yw�����I��9�g@=������ySG[d��h@q�6��G��|k���s��D��Ё���e��B���jU�\�u69P�՝p����1\G,Y�*�iN�Xp�ۢ&,���iʒV����翤��uC}����#�b04��<8%5�D`0<�Q6�x4,���W4H/�uϳ�O��R٦��k�y{t��9�c���]%m+����j�h^;�Z�{��G7c%�t1N�H[kLB��G�c4a��9��� +�0;!r�i���Sh�M�W��F`MBJ�A��i**oJ0HEi�����@�L�k8��z�mUݚmKf	 �sR�
EԦ���J�!<ERe�9*�=�Y6�}������6�z�D��˙�}��52|�L>��q`&!e�� ����Y�^>p'��j�Ry�A�x|2��/엿ʮ���{�Ҝ�}��>�;�� ��r�m
B{i,7l5���:���cn`�c�<1�R��y����Ʊ�<�P��{�?l����sj��C��2�n�:֣��;_>m�0Z��C@��WO�������
_3��j�t@�|��J���v"�%:�:$���#�]�Cr��z҄��O���3�@<����C��9�}�X�`�N�����[~��[$�I[��W�r�&,&q�Hɼ#�k@wOQS�X�.��tc�@�Rt�O�(�2���-��J�x�y��q�����
�-^Z�4c��ßC�/n�
}YS5�L���9�B��1o5Ck-��B�%�|�Sd@�l�l
r��Zo�hd��s�ٯ��L�?>�h�>��?���Q����*נ�+׎�\M4����'�����&���+���f���µd�P[ts�!��&�S�Ő�w�|��|��K<�s�){�&;�M�ۂՈWQ�0Zy�M� 1��(n�5�#�?�4QQu�hl�9�J���	�!4{��9W�
��lӦ"�D���,c������ ��B�OeF����r����ii�2ǿв5*����K�-����;�sP�}ע���4�xf��W�z!Z��'�愃%�Y�{vɣ�Y���	B�c�Q�mv!&EjNi� ��]e����+��*MX��'ϼ��]��*�9�b�F�N;k��A}	�J璐*\�k}��?F�+I*m��k���j3�紁�gQ��,OK��)�0z��<�0�Յ��q>8��K�_��<�f�X�0���'�_�rSY�`��^��grK�Q� �b��x���rC���(���t� �d�tS80�O��MĻ"Õ�����b��lCWG�"\Qb�eE��5g�r�����1_⊮$g���&��"�`ו���F�l3\R�
�|�� �w:�~�c8���f��U��(tTP�K�mJl����P����f��܌�!�L+ؘ��|���<�	��"��iپHn�Q+Еؗ��qNN�)����5��3��7���,�.�h�}��>?:��*)�O9.��Pb]��Bih%\8�ֵ�#^�m?��N�{	;Z��n��Ҧ��:���q��*0�m���	�e��)M����� ��m ����EGXi!GF_0�ҵ��{�qKY���&X�a������o���XSc�J����,X�K/�mj�?��8��o�!�����F�+j@�w=_g«#�ma�G�q��r+��be>�경~�-xL�_���e�Z|w8e�\�{aw�97u�%�:�$d{qi������I�D���h�A�ɡ���6���͘vhr��A���˟|��5h�}��)xn�w��XƱ�M�lyņ��.�(Ї��e�����7�4Y����h�.��* x�瑒dP��y�����(��/_וmI`�+`k��9[����#s%�@Q<*����1�1th��G��_曊9�^�:�c5��B(<$r++)�>�3kF�i~_�kK��È_".��;���[�H0[Ş+6ի�)�����Xi�$�,�#]X�����|���Pu[݂�$�:��y\b��5Ծ8�kP�w��K�SO�Ha�Q������cH�$�DXѽ
�~�~3έ��]�������6�գ��Ϊq���sly|��Bq�E�g\��R�et3���lqi7�~���@�ӭ*��!��Pwo��g���|i�Zm�|��RBR�<�&E��8�~̣a�c�w�8W	fNtl����y���74z���<p�H�m�%{`�������ɫ��b�����Y ��o��jgv`��yR'�;�w�u�+�$l$�(��T��7uFf�m�4OW�7ߖ��lu>>��/u�ÉE`��z�{+ˆ�x���,uT-d���%qD���Գو�-޾����P�(�e�2x�9$�K�'�#�pV��O�li\�w3��Ud��X�RzV���o�j0�y7�g�H͛hD���*AZQza4[��#��)��8��J�b
�T�-c���34��F��.	$7;���a\�pN_龷���ӊB"��E@�Xgq7��g��Q��
�y���Z�ʎ8���z�jb|�IP>�DF0�Sl7���J7AyN��6�~���·�Ă�M���cȤ 񉜄���y�l7�YNZ�����zI�(ܙ:�3�%�8&�C���)��96sAc;�\]J��jx�s��0�j�LL���:�;)2��h���<an.W�H��hV$��REI��Ux�ԟ.\dU���[�=�z�6��0ҧQ7S��f�'��:�������M�s�6��z4���ru0Z=M�N�7C�����u�D��)�6��H,���ڄI/+��U�U�J֏7�A�t` +��AϔE�ex:��������]�~Gc�e�Tֹr�K~Al` �P�O-NDuq)������[�e)��z%ٕ�>�'̱shRR�b����`q�\|h���1+g��qE���T/H�1dيU�Z~{!џ������į�S#��Y��Pǘ��@{̱t���:9��d/yM�AGd��E����h抨���ұ�z��u��]�ԁ+��z΍ "��聺T>0�c0lT]q�U�4�y�S=8��� W@Z1���d�I�|������u�m���𬁌��.���x-f��C����;��Z��_�|.h1Q*�`/�Q�}�d��)�+f2�K�;�*���@{�V�ϛz�P-?ծ����|�}4F��9���x���O���8s�s3Y���b�9���-⿭�PX�[�Z�(5)w���;������-B~�Qx���� ~���/��u#��z��݈���s'/G��	�`瘌;�*0A_֡э����j����Nzh�-Od��۸5۵����Y�-?)M��g"Ý��$f���2x�&���wջ?�����<�����;��Ȥi�!�p&�\��y��ЫW]���������A�@;6-���2���Ǻ@���k��3����b$��q�V�q�����8M�T���F<��":ܙ���[��Ak��AwL@�L���T�oP�\G����>C�H2CF	�q�k-�'�'�[���9����!S0�9��E.��4�:y#3�Q���%�{��<{��}��w�=�Ώ}�]d��۸�`�g�t�P���JG���r@��f�\�ΰ���C��5���B�C��͎I����r(éw��"앎0(�w&G�Ҥ�4�H��������e5/�9K����_Q�ٝ� �:/���_E�-M�����XI�,"t�&>�����e=��	ҵ�: M���?���6\]+�A6ouY�O��
>�*�X�Zv�^- ��Eܦ2��b�r�����[��_D�8#��tX�#&��K0@�7�OȦ���lR�[�}u' � � s�*ˬ�i�j
im���O��(×����01D@�R�F�I4/�秄՗:���T�����?���`�ʚ��gغxHH��u��q�Q�;ZLv�k�U������t��V����_�E�8]&
�.O1�i�?1��f�q�D�{K*��rN��^�Tw�H4O59���4 p�&sP��N��� Yb������ǜ�� ��0V��z�76��WSZ;(J�v;�_��V��X�����y���RU����o�T�Lf~��)�UW2TB�.�p�����-!��
�O��%1D�E�B��z�|����@�LUV#e�Y�n{��KC.�6<�z��L4���l�4_��إ��%f���Ӭ=Lh�Y���S.z��eV�}?Z|S�l�G�,���S�r(�L5�\ʗX����u�X
s)�юQ��3V-�c�8�V��)6R�KSq��^�rXR�jDS'w�n��%�i�yQ���q{��ߪy����cHp��F������K~N��"�⛏�aq��]<a�˛�P�v���x�X�����	|�.Ix��2oz�/B�?��u�3CE���79� N��Q<1��A� 7W�C��W�3�8��ᬇ��z�ԗlb+-�㈣G�7W�)�*JB�&� e[��H�A��g�{fIQ��@����\qJq����ֱq��@�a������1X?�]�ʯ�U�������>�R ��5Y����w]�~��\I��4B��b����$M�� ]d_��;��_R{�=��y�}u$yQ
���U����Jqp�W=��AeȤG��<����_��F"���w�� 4r6�[EW�ϟ��ο��:O����*�� Tf�݇�.���|s��ے����"
�q �0�dP�Ǯ�u�I�͂35	���!ͫc��p��Kӹ�dx�J�"C���l]N�`�i�>��b���5ph��N���s��ZEb��J�c�b������F	�&�"���(����؝���SF�	�r����b��{�E����
ԣ���D�X���p��ii��x`���D(�W��v��w��.�2�8��V�� ��T��jw�U!�5ף��7�d˓�b�R2>zD�+��$�b�t��r`Vk֛��9�-Muι�g`b,�;g���~��z��;D�W�1	NeN����S��)n)�9M3�8��������dCb����w��%aYht⦵Q}��ϝ0+���G| ��h���Ṓ<B�clwS}�ہ��?v�(���G�_0`���Oǆ����N�����E	?�U�HKю��k�
6���'����@��+��^+`��Q�^�Y&�V���Tbq�8���,8+������}����W�H�R?%÷�~H��~߸��EJ-*����z���`�Y8g�)SFaf�O���r�$�([�ٴ���[�T�6�����I�Կ���'^�ӧ��cR��ȗ�Z�'9c˿����2FI��El��Fu��3�|�}����7+K�o�
i��Zeg!�;@3�| �0uU�!> ���MA�b��R�aX�+��.?\�r�<�E��˂j�0w�PG�/~b���1/�"٪�)�̿�R��B����T5f#��È_�Nq<���L�4lg3��y���E�A"4��hl*�h;�Rũ:y��z�kP�a���x���N@�D�id>W~c�f��J��'j��Q�$�#�����Gp*/Y�E-V`�٩6'V96R�E�n�У�e�9�m��߱\���_5�@��c W������쐋ac�L��l�J�����!��JM��;:��_7�/�����
95�
���T���,��A���F7����%=�y6_����O6J�����A=�6o�:u�0�vm܀9��Y����4=�~M�c;b�mqKoA>���=����f�y��~>�������`ջ�B<��.[l��h|��`6u&89(T�ԅ�UM�_����*�h�R�\�Q�B�FS_a�߁�A�0l*°*<����+W�����g�pc�iρ�B��UFa��$�o��C�\H+'�%U��}M�ʮ"I��.����;U�cN�D���I.Ï������pu�^1i�F��X+l08F�Ǎ�s!R�>���P;~bɵ%V���:��[|��b�wM{v,F��O�l��dh-�r�璞���]ʷOF��=44�5ӷ1Q�ה8Ĳ�g���#^��c���,�a��9K�/�M����ѥ��F|+���'��&i`$V�f&�'_�9���}�Ry�ca���Rח�`B���iN����Ѫ~ձO��9U'���j{T5�Bb��g�*(��?B����ȉ����_� ��TQ#�k�0DT��
�Ny�|��R}ϝ��B��r��t�/���:+Iw��_�;�@mއ��YRP9��ę�CQ�.X�H�R�_�$�X��5'	�ۇ��O��3��'�̭Ő�USS�[�R�B���ٴ&��l�y�	D,��&��Q ���V�vZ�a���db���i/_1l�	-A!��#K��z��1�
��q �+����w�s�N^�)��J�?�Z۴�δ���w'���j1P���g�����lpjW�����E�q�YL�r9P��Ѯ�o�f�U�$%�z[��f6�\R�As����9�%��\�3d��x�1,CT{u�_����� ������ę;l2Wt�g4W��H�w�Sq}������}���`�fں���Ϭ����;*��
�W3�̖�$��d��CЄ��&�7q��勑67�%Fa!R�VO�)sT�9Ev�1<�1;0���^�A�䭑�.&Ub�
]s�i ��w��O��Y ASGxl��4�se�.,|�u����x�GaeX_ ����u�0xf�,!gTo21{�7�i;W�8�U�YA��$Ha�-l)��vfPޒ��JUȃUԖ��"["ے����^g��[ƩsuKl(�����tz�h%6�p���3����ۧT��Y(Ȟ(�tj�O�6��V�0���V�#�Q��\�Y�'�|��Y��"z���M8��x�-y�H����
��P%`�6��뗐e�x3���}p��݌F�+
���Փt-|�~�M�#?N����u��E�g�x����q��4�>V����<-�xt�%@E	�۠�
�ޡ�M~�����;ñ�
R��f��b �_6�O?�W6��Q�Z����|j����K8��w6�j���	�݆�����fLn0�	�uk�jo�� v��؟2��������֎5�Iq��5eyt������H�V�J?���!�eEh�~WK%_�:�x�M���bise\�8�H�-��31O���M_{L�3l�&�q�^A<b�Cf�<�b)������ӑ�%��Dg�ji�w�i�o�Ff<M+b��jt)CGV7a���>0��(��xV�����:�Q�*�I�g��{��M"��E�I�&��*A^�S�ܴ]D��$�MH��cF4W�Z^���{��[Г�uI�����-v�|��n~����5��:P}�He���~Z�ã�����O��D�ڛ5��#���e�qG/n�J�˔��j�NXG �t�+U�E"��������/����n��<x���1�KI�����SB�z3擀+�!�yU���k��V��@LYJ_���2���2�o,�����y+᜹�}cJ����ay:*ϳ����+2�T@�q��#�z����T˿��.���ͳgQJ��E4Ew������ٸ�gD��S1����*��\�@�$�2�L����1T�I��a��:�]]�1�o��9ȠÍ�:�	BÑ�J̳a��O�4�h��~m��h�5��N&咩���C��ˠ���]ǈ*�R`���eH�D,��6]��߄'oSj�X�:���	;�* � P#W
F!���O�Nl���O��B����z/��֊��>V2��3���s����	Q�7�9�*+�HJ��gçQ�yK��z ��m��Re}Q�C.��-�O|K }&�>h�M��J�p�h˭ �P�1�A��Jn?^Dҙ�N�kk^���h!Y�JY�AC��J^���Oa�	p:�sBNF/wD��{�ϴ��NcR��/��	�`{6�P��aP�&X���)B���HQ7��>`W�H|mPJ��4X�3�T��f1d?���r�C؛���a�K�*�1�K_<��̓����n#��I�2�tG}3�+�]Oz4r�s� a�J���$;m|5� 2`�n!�EO�7��_�䣩Wg�5�h'2����A�_`��Q��)��W��S]�O��xx��� (aY��b��߃�m�Fg��qp�U��S�3�l�K�)�iS����E�`��ׂ�_kb]!I�J|�[�xCZ3 �g'�K��ɳܿ�����'Ӈ}&�n2�w�ʦ�x�7�ܤ�B��yUU�%�:]/� 5jHc�%�*y����÷d���/[���_�ӝc��-�N0噟^��s
��2�̚�c�����)8T$u9��]����|y�Էg�s��Gv;=��%}#�05�e�\�;�mC��޾O} �IZ�����~���400Q��Xx�����I(i2`˱����h�̖W���]zKmz��]%yZ	>$�����%��>�ݝ"���x%%����[��g�7�w�����i����c�x4�GԸ.�V7y|��s54C(��X�լ9���U�U�Ǌ4[��ž0&>=������`���[�	#+�CNH)�#�6�O����NG`��x�#����`M�Q�緷E�gG�� �&�%L���yW>ܣ�����*JPL!���PRH�������UF����Xv=��#e�5X�vD]a�߬p}����?t�}C�8��ܙ�W&Iu�,�ѝ�؛�Se���wۦ�x���sl���>�2�� ���N�XA�c���|�h2>JX_hJE?�*����3c���]�J����]�u0�O��hqӌ��;���ƨ��[s�0�fV�S�"��q0�����
gt����A��l��g]��(�Wg�o}�a+��S�P[�9�%���N����5��ֳ���^�����w�+h���3rm�d�[�k�빋e�m\����_u�nÆ�̩�8I�	mE9,{XD�U�>��꠻~}ќI�ݑ�YЏc��V?zm[�-�׊����d&��P'����^^��`�n�-����`��2M֜��G��K&���{�,0�#p���/�t?�6�e3m�
)<WBh;h05E��Z����5���N��2�����	�	Ke�]�x�7�HC��27��ܚ��6��N�6R)�=��(�o��{,����UZT|:�M����> A���8L��Q;l���q��c�`J!�r��r*gPw/�[bY�4Q��bF�F�}��S+����fC~3�|�����2L eh����*�תA��i8��1���{�B���6U*�:�_ U\��ׁ|�JBv~;�n���-��gD�+X>�b�E���x6X���Kqc��v�Q�쳇�fY:\J���u�ʿ�g�������(Y�T���.�Pw0�X2�ɰ��T������poDbj�" (+O�`�nCN�ߚ(��!������@M|��#
�j�e����?�c���<������ F�rw0����85J�fi��� ܁[�SauZE�j�G���f�'�E<@0 �(���6PY�Kԇ���m���K-�����;72d���ލ��.��%�����ME��]��p<i��2��Z�UޒYj�0ys/q�-�CE�\�Jr�S ��m�_Sn�=��n���G-Q�ͱ>��(���ß������M�lVU�^��ޖ�2�f7yt��?it���v��ޱN9g�	 %H�aš&���]�6eZo-6?C�]��|�d�}%�4B�YS]���`O�W��ͪ��9.J�=�������x^�@�ꖹ5���BT�:��a�(R�Og�z9b�&,�.��.`�XX��b��_��VS����K��&����-�t..��;`lP�c�|^"Mk䋚�������睋H|��Y��>^�j�xm!2�&�Z�lN0b�R>l`pG%OO�m�u��^�=��J�m�ɆB��{w���
a��~�r��(��u�5�y-�d�r����-~z	�U��H�BZ��g���Wp�]�#�5�U:�TM�(���Nk]\a��}�VE���`_���]����a������p���
ZYٺB�x	� I����{B�[�\kpݶ�F��I]%���� ?���§_���Z�?�d�D�'����R-�b@S��dW";#���sJ ��/�j{�F��=?6g/���4[~¥ALg�2�R�S���'�X8��˹W;E�������{ЌW��P����VFI�ȸ�^�/z��3N� �g�.�F�ҕ��j�X�����c��K�rt��B��mv��b/T���%*qoCQ!����{�i�f���YU4؄o�ʬ�x\�$71�#�h+J�f���6�߳��:,F�~�
5�d�m�J�ݭ92�$V���q��:�dU-�X���G�cJڟN��WCc�}ҏ$W�N� 0�SƁ�K��6'}�3�K<��fP�6�iU{�;�uc�(�
F�F��0�s	U��&!C��1t��
�N��<�*��`CWl���A� �I�VlX��0�V���7P(|N����ӕ	�CS�aA�h���5�a�&�������P-{<g_�'"T�p����[hp�+7N��!��0�O�iY���ъ�R�{����;���b+C�A�+h����k��嘨�D�|}U��~�����c���W��+B�<�QIM��{��S����E�k)R�w���<ܵs�.�7`�c���2YO����W�*3���h,�"F8.���f���qT�4��=bׂꃂm��{�͑� �ȓN��i�I*
����������0�K��R/=�"��8F@�I��=���W�Dͭ��$ ��#&5�F�[{����&����\E�6���]o�O��~����D���f�ZA���|�U	oV�MW��@���\mfW�5;��]C�Ti�ǚF��5���u q�^��:#�����R�GU�5�a���q|v_rӓ����3����1-���H\�Q�����"��P��C؁���~��5O�S�&���s �n]�KS�"�'B�?c<�eն|��B��BSM��B�C�ö%^g�u}m�eb��{�ۧ�?��Ozm>,�z2��M*��	��С�H?��Ɗ���+�*
 �o����.�|��n0��G5�!�/��B��g+�O
��>�,�c:ᠸ����E�[D�-y�
�S6a_ثvT�j&Oh �ym�*g�_���c�����	���U����e����!��"	��/֟��敌Z��0P�q���M�>���#�j�-R�ɩ0�Voձ*�	���11Jo9jd�-0����(^}� �ǥ�J���@?�k=kRpM��YQ�����ӷ�o(�;.7OǙ�:z�{����a�h�i���mwe��V�W�n�H����_i�4]1�a�H;�\�j��5.ʟ�t_跶�4��)�"0=�������@��0m�m�� i���n�!]�X�n�T�͓w��-���"�`�00�8k_+ˏ~d�I�m�a�+�6�?�+�XԱ�I�� ��B���dVؾ7�BG�	-c|]��9(��-	�1����c���VG8���HäӋm�gIV����PLm1�F½�%�,5W��hr��3�'-H�le��"HB��� oL��p[�KFA�a��q���򅠦X%��X/�s!��}��}�,��md��� �0��]A&,OH/=���P��h<'����pn�}���P�H�m�?2�. �eKu s�