��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\����q�?��e�I8�b�Ǽ$��"����ׯ1�V0�����A0����S��<]�x:7v�%֐����ƶu�̸��� �u������Q����k�k.CY� �F^�7���eIb=�B�tA�F(_�ИC����Ô�������{��*���P���������f���Y�k�2KI�o>h���EX�|V	-8W��;��� 6L#N%{�^Q�u$�1���DoA !I��R��?�cЅrp��+=��u�����I��6l���ֶxh�&��E���>лM2���p�j����+��y�BY�w�sw��E��|,���l���Xr��'�c���v^���ۗus����_/��R2'*��t��q_�[�|�xO�8M=H#N�s���@��T�RH�͋�f%���-3�9fC��R
(�Dr~@����*"��X�&�΍��hd��+j�L7 Y0ke�ZFg	�8���r��S<Y��Z�a�B�MQsݜ<�,_=���dGb�C�"�7�e�:��T��W���9m����g_��Q|Y�|
/��ȿ�B��<��xsD-�e�Ԣ�f�9�_�$�V��'�P;�@x��uU��h�z�W�(�0�U��Q�06��m���t{�md��K��#����b'�4�F����b��}q)�ۨ
��,S/���A��������̮(Z�~slt���J�s��90v>���܅���v�d�).d!j�T��6�Y��)� Q�DE_���/Z*�r�a6��A�Sî���e��G�{��֊���]�L�1�JiUkA�X��Ucl������� �r�O�F��ƿ)u�	MZ�������Q=s��t,�}�s��ciRM��WO��.�##�Ɣ2ʇly�1:yo����O�yGWeX9�1�>ǇR!`��iu���5A�;�
O���6��F��6*/M:�S���@��X-EaG��8�Ɓ��ކ͑�	ysc�s׭��ws�,{���gu;�F���Jƞ]`�istmG*�mLt��v��UW`I�O�o`JN��eރ-u�.��6i�\�2޽� �%��K�2�2$f��ޜRk�G"��!��n�;�f�|��Mg=�jr�?���*j��������-�B�R��m�KrY��C�)Ƕ��-�f��2 A
�cS��tZ��43嚈	c�D
��A�J&�����R���>�#5�wϠ���5�5��
��q%��+^�"�bL�!s���r}P:��ݔ���.uG{)��*������/Y�.ζ�'�b�B߻0[��1�2�:���VXSA$��I����iZ�����%r� ��s݆���C���<�iN��.`