��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\����q�?��e�I8�b�Ǽ$��"����ׯ1�V0���@�Zr9����!��`w\M?���*u%�Sz�$����p:���u��l���#g�R�b.� _�U"���2��l� �
� �c����,�B����4н�_�w�mF��B�\�SҞ����VH4f�Ш���d)M��������X��ż���Й��9#�v:k0%FN%A2Z��r��?<���Z��� ��`&9�3͑�Z�b�gF3<��E��M���� �p�t�'
��*�p�ӽ'�^�4h4��f�L���W=l ɎV��� �p��$8���xR��tt�޴��D�����e%ϛ��m���D^�N������m������D!�.�s?G��ٱ?w\F�~G�o�I�C�r��Q�G����F6F�$.��~�ӡz	��Qr/5I�PR%]��B���8CJ6ٱb��9����Ŭ��uI#���t��	1�M$v��9@y��>�
�=THo��ɱ���5|'^@�2��.2D�YK����ψI�. 3?9KT�C�2V`�� [PJߑ��IX3;QeoS�; V�l�)��7U�;�,j�b��艰�R�$��
oՔۺ���H�wAA٩S	��秦����[;e3�Ӛ7ɪ�xW�E�skN���������F ��ebM���k!U�~	 �x��F�-GX���-
I$������� 1:ʄ�4�����E�H�����a��!�ʮ��C���Ɯ�X
��c�'�g����J��TBX�ZF�mQ�̄t_�'	`�!���������v�(g�@]`�v	��P긽��Ξ^{NZ�����M(Ŗ�!��yL�[��'��^p��*�x����˦_���*ɔ�	��n�&a���c�U���8�����.Q���[�/&�� �h���~�k[4I١3���t��s�ڨ��*~(U� ��/ ���M��=E���?6Բ+� `���?u�u�dr�9�L���*��hլ��AՃ=s)�:��v�j�S�݆{B���Z�9z1���O+���I͍{\�LC:V����}C{�R�@�ܻ�aPac�\���9�2�s�:�,!@be'��<���V��a����4o�4���-N_��Q�����W�>�,��[د�}召xw�dSӫsq8�>ⱳ�;;���ىd�Q֗}]xAK(��=w��*vw�& ��,
.��G�0��j2`S�j��k�#��\ե��Q[#�-诈LS�������6{�p��dW�!u�s^�F�EH@=���[α')�|�t�uOZ8NSdFf�h1w��	\z�[�ڵ����w����6"ʨ����*���)m�->>\��^�(v.5l_p�B$�g�T(��Z~B#`bY�Vk��^E	�>b�%��p(�;�l����9����t#�L�w:OF�u�æ�ؗ�	�����4�<�k7��UMc�۶h������y�e_�E!]�ϥ\���k�yS�W�qg��H�u���4�fۺ��~�ͽYM(j�M�SݿQ�*���W��McBc�~�o�]�״h��:�X�:�GN�\7���\U�ݔ�rn��h���@\%�qs�޻���ה���
 K�M����W �*�MC�8rsl�YX}Έ(B�V'�*���i"f���e��^��Wv�q}����R5���J�͢��EX�'n��9G��ś�k��"���;�}+:�f��"��;9&�����@i_�7�P�H��՗�	���.���:ɅA�_��&p�'��2����Z�+7���=��`ݓ�ZM��צ#il���R����:w��%&��T�5>���L��r�O�E]��,Ee���-���Q�&�B�_:��K��yc)�Ȣ�<�2��﷛������i���Ӛ��Z�.����v���p�6��I֚�*!��/(E��(Vc�X
�����[?�o����J�@��<���}���7�*hrVf���=����>�[3���>G����w�l8s�r���s��#}���d[�-��s�z�U�/�"�]onx�m�ԩL?��a,sބ�l�b��Y D�����qv��_GR �l@1ǐT�����ǺVˀ��hp�r[d�a:�>ׄC�������&ekm\y���l�~ŝ�'�G�Y��f�s@�wL8W(�wܬ��yw�F��۔��PZ�˙��1:���e໅�����G~d'�(hf�~z�#A�`���l卖up����YsM
"��/��[���s`-׾�^Y	��c��x�Ԛ�*��0�|I���X���3(n�2�J�IG����
GI���^� S����g�1��Lc�U���u��*	>��:�"6�*^�黛�����n[)^n�&u:���,�qT3����8�/3$�1�/��Fu���T8�V���b�N�x��Q��:F�zV�ӉNM5R{�,i xP!�V���-�)ަ��k�������32�#��i�iİP؂��Xu�s>�2��1���U�p��/+�K���a���H�(aס�z��́z��G����Uh���]�Hl�oD��tP��1Y����f�;�?ַ��Ka4�eq��C�5L�D����6�0r9�,�Q"�l��8kb ��鱟��I$D$>(Erʃ��@Z�wH�^k�0��&֥ia�N�k}j��F�4(�\���P`?v����C0Q-������En9T#��N����zmO��m�nu�ƅ9��Gu�<�+�ib���!D�*�d4.2�'e������MтOn�W�#�]��;�$�ʽKe��ӓ_+"�p�}�K �nN��%���$��A~�}����"po2&������m�[y:�a-W�;��Y�l���'������+?v�ܢÕ�@�2��f�@}8��)�n�n�.��6K��j\���\�v���;-���(�%�R&�;i�dwinB@tԁ��ۈ'�
�gJ�x?|����D���S�6&�!��[u�uY�fn�
X>g�q�9+ݤ��f[�3֓���-�����
��@��*�0\+3�GN|H�{c���2a�D� pF\�T�~☩�p����n!�^�o�����BPrD;4���<��U�*���t'r����"q&��a7��~��;U{��H���)��5�76��D:���ސ��ǉ�u��HxmY�B��\9�c�"(��lI6�8$�ჼFb���@[3�P�"�����M��e4�ā%���H�A��{��ZY.- g�7
��;;�N��	�5�����,�y7��%���=i&��|�1l�1f�N�"�G-+ͫ�2�6�~�,^F��Us�e��y/3�
���436F�pe�΅�Y�e�{��� �t
��ۊn�6"lnάdg��D�����lU���q�x����Ea�"U�F~�������֣���+��.��p����v×E\C�;)�$)�lcx}S�����R�޶f�8�*I�3�0�{�&��?+'Eu�qU��1��)r޶j��5�0���5�v��1쇯��GM����~����DB:4�Z��j�cꮾ��伧�)��uD�to���M��~ē�7�2�O9���_%��L)D��6�� �7�nsD�N5���n��A|)��SFp���ݿ��M({d�,˯����Ysvae�Vv��v�xB'TJ��qFK{W�Sߴ~�~�J��^��'cwM�pT�#��a��'��ȇL�>B�u$X(ͺ $ܧ�|�M�d���@u.���J>�U�^:Z��K�C`z��i*�uÎ�}����q��la�U���À�d��-��=��}R����Y�ʵ�N� TڛhS(0�/GL������ܟE�lם0���A��+�G��[���L#R�5'��8)�����'���
�!�ƍ	�ݹ���&�S���[�䞡I��r[0��pw$�;�_]����z�-�i�R�W�jv[j�"=tf�r�A���^�ڟ�$���
����8Q��n�g�s�W����¢ܐ��J�sq�cE���{ڰݎcrp�c�=Ȑf|ɕ`J)g������J�ٞM��f^�A�w�=��H� ~���S�g8h�����v���3�2p$���T�]�Z{C�ԝJLQE�B ��r,Q\�̠_+��S��8N��TD�n��N|g+��7��h �Uv
�l��F�>Y�U�,x��zs���V<��$$��t�16e(]u��ˁ3EA:w�\���0%osԹ�F��w���[�?#�f(��t���J�{0O'
Ĺ�����c��ŷ��tz�?\`�8�Z4�Q-�S>t�,͡�d�Ր])`�3��������3��u��H@�껹BVb{��ٔQ!E?�"�)��u�bvm�uI~�MN��>�ҵ�fa�v������T݈AAr�˄c��TԬ��1����]�#����۝��w����>+�:�I�W�fn��#��0�kP<(�[�Q�	d��Ӏ�I2�AzBܚ�����#by%tK�^Eꦃ(�4!I;3�Ɇ��@U�HWD�WS�m���'���{_�2viu���ˤIF%(�%o tX�碐^w�U��j��$�j|��Fz!m[�������@��60~�-�ٍ�j������Ӎ�_z�}��|{�wǢ��4�	w�%�B!�qٯQ�<Ke��L
��cQ8cD�CO��+<�lWpRp��u��֓s�w�B�k�+`���X=��8��4ҩ���|E"��ju�L|a�S4:�8��zE��9F��r�H)�~����˓�˷C!x=�<V�t~j,�����BE+��,i�>�j?��x��3�*
H�뫘ɼp�i�_saF
�BM���F�M�>(Cj��&������8qJ�t�q ��J��^�]��S.Xq^g��?q����k֫A�i;�����zL���m�F��	�Mz_H�n��^�i�l<�q�h��m�g��{�E7O�쵔�����k2b>b-��C]�yN��F`�\�P���@�W>~u!�r�f%jb��g	�A҂�aN��~�g�ho���xCi?�֋*r�~�=�¶5@��K�{��mѴ�Y}T��cٚ0ֲ(u
�p?t͆�ٱ�v���^c�ЈT��w?a�@��H�q��,��٘��y��r�h��Ɲ8�q�Uˁ�lW��u�(6Z�:ldBOBE�g1[�y��<vý�q(w�{6;r U��f�{H>�	��׽k��Nc�@`�����ے^�zi�j��z4�gص���_�e��JЂ�A�b��s
�,� &��\g�򈲇׻~�FV&:�A������'�m��춵�2�������I����l+��I�2/�˄ ��=P���cs�SX��.���4!Ǖ�z>~�4Έ��$�'I��LmY3�%2=�9�c��XB:���c��,�қnѿ��ا��x\Y���<	~&�a[�oC�z��C�ㅃ0�-��܄"6k/՗{�c���m�r� O�Rj'K�)b�I�L��s$��U�����,h>�i��R���~�l_���8gً":�I��jyG�<��7��,Sxs��l]�To'ۣ����|�_/�a� �Lhk�@�lg4M8ϯ�����]��^'
�Zc8��ŋ�o^�ip�|V7�Y"Z�����U.��-�8��6Ԋ8�
�*z���
&AkH�Iv՝��Fj�̷w0]�cth�C�|��XA��Ħr�D��*�z���H��tg.�/�V+Am�Phj��J|5TH����XZ�LJ��g�8�-�۝w!߫m#�AX��$��C�����Z�ߍf�;Loh�mpx�ضSWpev�.���$m�ϴ��2iSf<��rE�Վ�:���&��1�3q�>I:=�H�\V�G��#�k��޾G�S(u=�Sk�ׯ(�C����na���Z�X)L����}#���x� "<�M�+X#�zK��Ir�%Mŋ<Wl�uA� s��}2q}�P�v((8v�K��/��Դm\'�����}�t޸A��>�#�$:q׵}8�Z��D����g�[�-�����ĹKd@r���A�{�B
�l��aSL��k�L��s	�VM��\}��x�?ܣ���&�ŞJ�ī L
��+.���L��
<�3�U@�}z�W�-JI��Uc'5?T=I����^�]8�*�P:Bu	J"p�Y�;��"MZ\��e�;����uۭ��k�-@��y�F���}��R�7l�?g�qEL�)Q�S0+�'[��^#q6��à�@{%4�`�oz ��z��j!}�0�����Ed��=?��]�1�Ϣ�#)'����~d"y��E�i�m ��JU�̣����+���>Q�=Ng"���$NĜTI��5��⒇ݥ�K� �o�[�D�a�QY!]��ĕ2pح�~�UPT�-��][���Mv�q'H��U��j��F����4~�m�����R�(M�b	7��	�^>����0:a{�)�q��Dz�:+D񁎚�� }N>7i����)X��`���G_`�H�̡�GRz��M�����"� �6$9�ZG���1j�;�6|Γ�Iy�Zd�դ�@M�����.%�����=��@�������Ev����\?��f\o ���{u;!��|kɁ;���i�u{��\�H�Z\�^	�=�=u��T��cn-��5+O�Sv4zV���'I��(g+��)HT���'����b��(
sD+ˑu�wcPm�g��.&l��i�^�͟�V
�H�,�u,!ɐ�X�ȳ 9�HBw�(W�} ����Z��H%pz�"0n� s�v}zȢ��Ո�Z�X�㬁�F�=ܑ80��pV��Ei�������-w|��P�,�R�7��u���y!Vsa�Q^������F���WOjA��(�z��	��c&)������u&�+`�3/BO�P�J�-�p����ʹ��ev�d[&6$�H�������k�����	��昅����*rS��C:Z��[y�1kL_��4����m��&�z*��;}D���E2e6�4�7�������V6��i�!��{�` #p\�#�8�>F�*�|%�����P��v�_���[�s%(1'���:��c�����vCW92_j�%y||�`.ˬ㔅�(Ms��S��C�.HE����ǛH[3�NPЂd�[��zf��q��G]��ז #����/�"�Er���9����F�e퓽0��Q�u= �4�d�H�4�Iߝ֘�Ql%���7
s�v%o��H��O Hl�O�+��ܑ`�JSsE�\�,��<C��`��m�Kj��B��z'	�.�a�/�PP� ������N�ݯ����{]�p����W�iL�/
�;�E	OdT�]"Ts��5�3ޗG2�9mKN�%������7w��ie������t.�+Z��`�\�(y|�|���e����N��Z#c�pM ���D��6T��kR��3­=�J��ar����f��u@Ƞ���rJa�q}�A!v�	�!}b��6���bp^�!�i ��̊=c=p꬈2xb��V��r �|�Z��W�&��w�!|z���ph������T�ԝ3��?)j�WZ�}����9y�ȹi�PV�C0)7�Tb4ڭ��r��wQ�:����ڻ~��l8�h���/q`De�;��^�,����{����HluxmU&�-PS���O��i)-nau�+�c�<Ҋ��^���[���{�c�pw0_L��떣�'��y�i�o����,�i�����e#���X���t:�r&xV�lq�@s�4Z�����5�x�V��c�]k���2��{���I��d� uYl�y�2����	:
_�l����J����^;ڝR5����tFMW4��8Z�y
�ڻ��E%���A�`_�$)���H���ÑUԁ�`��P���@���Ӗ��S�Owjkc,��:[q���R��;Butb�0�Ɯ�NL2�Y�\z��J!:0���p�i�bTә)�~���Rq�Ɉ-������+_agztg-��{[���h����iW�G0bl>=H�����ʦ9�������_�� ���mÛ�Q�d��CA*jl_K��?�k=�5���y-�V���μ��ț�Uj��>��[+â�R�<�圥�j�[&c���&k�.�9�!M�0��s��Im�N��ʵU�DWV��o��LA�܆�S�;2=�G�q��36�_)m*�N�Q�a�lE&�9�I���5�>'��By����k+�if&�AuE&aN^�U�dTe�i�������	�Z�#y7�VԼ�{�ɇh?�+���� 1�Ң�����c�o6�ƠՎJ�,k���um7u�1��g�H�D�W��Y��L��!����B��Ż�G����3��DxP$��l2�>Kn�W�����q��Z�mq�`�B
���2^�E<�I��Z������@R�=�9�>�,�o�����_B�� ���zo� m�%��9���T����vp����w���S6PJX�8b���7������م���H��]Zk2/�0K��I)f��/[�k� I��"W���R�w�r�T��o�����s����1*5'_���sS�/���̿~K�۸����T�sJ�zF9?/ϡx��qj�8���,?Ұ��}��&� �v݇�d7cx{�]wqb8YN4)�x��_#��'@AXj�lR������j_�â��x>4s'c$V	�Hx��>�b�-,��d�G�"��3��ū�����������֌�����A�q���~��<w�}=��zũ3 "�r�n�Ҥ{Hؿe��·4���d�В�.�n