��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\����q�?��e�I8�b�Ǽ$��"����ׯ1�V0���Ս|0(����vN�,x�^����EMhV�������4��X� t�c�ރ��H
�Ϧ �|�P��~7�X#�&��DYPA��S�A*��j�>�f�˚j�D�KQ�za��4�n�^��>�^>h��<���Z�y��-�����g.�vʱa�7�e�L��
�I;N=���q�#�e*����Tq���۾��a�b���b�V���`k�����NgUI��Ej,]=�Pw+y�2Z����z��Fqi�欪��q�щ�С��o����� s�iz�El�p�M,�y�$8ې����۟�Z�!�5���y7�vN�ѻS:�&z5����.����ߋ�uFPX��+��	���$�D�����:��6��z��I��]��-�YTAQ&��?�-����DI�(-2P �Cq�2�:H[83�Oi]#%�)i��fx�n0���s�:sX#��.��'lM�����-Hަ�2y�]ü����?g/fU�;��rK�<�Sb �֕{��]:!I���]���3��1��;��>���#�v���Ml!T�R��P�n�:��؆��N�{��l\��Oz5$[!��S�fЁP��c�������v����a�f�i���R�7�q�p{[ԃ"�ˢm��R��W�K�"*�_��?�N�����q���."*�m�c��Ss���r�tԐ]<q3M��Ь�W�=������ʹ	G��A~lÁ��YN;V!���s~�O|��c���G`[�Y��x��w8���N�զr�x��U>k���Lf�O^�)tr�����.gY.� -���Sz�jkж~ə�p1;;�d�B�d�q��T�<�N�"X�hx�|�W
����HE�
�T�@>b������"��0��(i��N��g�W'`��ۖM�
����S��܉���WG�_�����J�$mCU�p�Vdউ��;��Б� k��;�~컍�Ç��TXуD�l-}�B
-�1O[���'�u���Vhö�����`9��J��f��A=�x#z:�=�Qx�qd����ۊ���ʝ0�Z PI�A��yc�ˌ�%�IЀoT����k��l�:��ʉ'��gUs,:�_�B�_CO�*�f��'KI�S�%�I�v�����*���0F��LQ/Ռ6�ݖ�����=�-z�ԝq��]Y��t-7l��-�����[&4F���|��(�U� ֑]�m���mż��뇘k@�&G9+��֙T>��x������ߢ���z��,��m1������:Ǎf�����׉#�
U�<�JEܛ(~�?n!xj8	�#�1йg���PK��&�v@�ʍ���ӽ{J��� ,/�W�r粬����]0k�@��R��&�r^��=�����3|��u�'�-��pcXf�Gu��ol�!	��e���O��s-1}���������A+9f:t�͸�������N�#R�ކ�o�;u/�����{���jP2��(�O�D���MB�@�D3�`m��Y�O���o[6>���E��M=#��_������R��zC?B�)R�$��L�o
Y��E���̙:� �Ʒ�����vj��%��te1��6���5�L*O�w��K���C��S(@cE4D:C����ϲ����I����3�t�M�-\��tl��O+*9�����<�\I��	!Y��!��RϔD��%���h�c�f�y9�x(*�S�I���H퉅ϲ��<K��ߩ���vg� 6�4LY�����ln&�-�
�;�;��b8�$��.�|�v3�AA��NS�Ƈ��ٝ�U���t���ip��H備D�R���t/{�����ħ�B�G�-+]<�a��6��{�xR�V�"�3@?��f�nы({��f�
� ��ޟ�>Eu���PGރ���+2��ǒ��l�#�L(���W��wh�	k��E����+����g�2��ľ�5�nc$~�穗<�k�0#��i��8�?��'=@��!��MI{�ț�x	�^�L�nK��q	 ֚�v����9�ՃU�ו��۴*�L�D56̝�E�yߍ�X��i�<#.���n�b�&�au��rH@�T�Rv�c���$�;���*6=	�e�r/�$�j��H�οP0X�Ej�C�_�C�&�m���脚�J�����Ø_\��~>�F��v���F��&6�7Rm�{����:��֊�hx����g�F_�'�T�~3�4`���%-8����¤��|}-��Mԧ~������̅�K�D9I>��&Y=oL�X,�a�e�L�i���8�\�|/ �s?�}σ�񊋋MG��
95�q��E�6{P��5�/�U|]�<oS:N`m �:�S0�h%p5�ׇ點�\��6=�{2����� �F�&�ב�["�$�+ąsv��Q$�t�9�kd������4B\A����Ʈ6r�F�tqw3މ�Y�k�C��d��Ya҇�P�qM3�_w���~`�%��E������dd���kqg �ɼ���;���G�n��+��I�*b]/��\X4]���>�jjC�bFA����-��ND���`�c����/�-G�����{rRZ�8]Ԭ%�2X�O�f,T��K"t4<�i�qf��؊�����X��f��Y�Ylz�/l���xU�5�@d�zuڼ�=�����F�05Y�Bg�� �ga���mޅ�5G�9f�G�hhM΅�����H�Z�#Q��e$B�*���m��L�4e�b�d*�>�@�c��$"�"�K$�Y>��B�"��/[��,���a0���'���Y'U���0������;�۲����t���[b$���x�$lr�� u����m����tF��`qB�:�ۅ�+XG��{|f�g��gRK��M7+��.���w��^<�w��
��:����o��m�B�N.�6*0��a�kR)�O&[����MG��5��`�E��-[�玱Ɓ!�n���HƟ��3��D�����9����y��A@̶H1�2�+hvLd�W���)��l�=���o�f��냣�޳b6-���f�^�]�G.V3�-E@�	VA�������X�udW�>�Ē�Ϟ�(vh>mͺ�F�)I����]:��E�D
�V�˸A�x�z-�^7�?�dN�f@H��`'%C,� � ����Z��<��Y*�qzV1q/=t�����^?�?{�4�,��mm��A>��04<�Ł�Z�v��z��W�E�	�|�5t�+�P�׹��:��Eϑ��_a�=��YٮF�џ_zt�iObkK` {��D�2݊�!'x�q綸\ң�A°)�˖-�Am!�Kv�wl*J,�E���qY��d���1���!�W	9X	h��E��0t��+�m��B�]���|1ߩ'�q#��r�@�e!1U&�z\��Ct�*����wY5�V���������kF,E8�1h`}�mC��y��h���'�>��VbPP��lGl�y'�����apL*&�z���aش]*��#6R�J���T�C&�73��ĸ��+�bW�ՙH۵88+��6�e�h��p�i:��#{A��o=$�|����_Hǂs����6ZH��3��a ��К���Z�CcV��n�iu��b������4��7��Q7 l3�S6H�Ӆ��B�@�1��W,v�g�".[�ʭ��#�0u#$�pXn�=KXB!0%K�00���;�u�NBb ���	r�ٸ�̲��.o0���X42������䦔1�$ڀ ҕ��L`8(I*Sy�
�˅�v/Z�B����{Q�lZ�$�F#����1��x��#~��}`���e�͎z�[4i���&�(1?��x��,�J�<u.��/��=V�[�M9�w޷V����g�t�?�F�)_�7~�c<1�ֲ��Y��%D���y��y�6/f��Փ:QA�Iv|8�4g�H��"��q�-(�R/�J�u��M����1��B�b|X��*��]�����1��!�� lw+*�Q��x�E?=)?�}�[��S�0��y`#�'P���J���a\a�E:��i5�m�4����s]�(�+�p�%%Rp���h�����R�궅j�.��%���#T�������_��n����քq��ד �����A��A�pI  f�s����7��?qV�#竝��*�D]�� �k,avP�^}6���o7�"�*մ�yѹ�\_b�9�?�f�:����04>��"����\�w�5�E����5Ϧ�7Z=�Cn俆.p��*��1�ء8x�a���,T�°�T��Y�p�_<x��T>iz���_���7e��W6��"�jH�䱃X�$���].�$�/��rT5��-Tf���9�n�v�y�>��$d�80�y����g=��R������^`�������������D�����dP#\��bMQ	~8���v�)|ᝧk��\.o���zU�ɓ8�<�z��'ό0�pG��"Dq{}������9�ɞ�T�8��dн���O)����X\X�~m&|����>'g��`Mp�\���C;�Η�8ʔ��s܄����E�����"Nr	�p��R�CHc�n�"0���Tt6� ���>����)Һ�.1fs
gy���)��Un+�y@�i.c#�v�A@�����S�*���uqa�x��tH��<��д�]w��QU�g�9���d��ɘq+%�7��O�<V�'��]�fי���OD���w��Y��o�^������[9W�k���xk+��h$�,1���Ә}~�~�Kv��gzŻ�w���D7���p��J���h��EY
��<�{`�Nt(�x�q�30 4J�E��;*��]g���,���QI��?A���FW�G�ϐ����,1R���ƬaW|w��jd�gх0K!!e`U����1�V`��{�-6�	�TsՊ�T�10����ɪ�-�xu摷4-:.+{�"�^?|U�|�����>}���:���rm�;y7�̜x4A�Ub������W��1��MPA�����6�0�ev��y�6-���c^\��R�0���x%V�3~
��-�u5���\!@J�Ue; ��CS9ݯi5��l�d��Ȣ�t��^��_���V���C|� ���I�����P�?�T���Y>�d,\GB�����f1���?�<ˬ�"�Z�x�`���d��+���wx
�^ �J7�	�i�:������Q��0�g�BsD_
ś/�	�����ҵ����t6��y���T��ے�F��0H�Jp-^���bsS)�v$h#M���pz�׮Ч��ue	mF��f�`��1��ú
�r�t�#�ez�[6]Pif�h��9�����\���u�q��r�X�ɾND��1kJi���/����pN1�Q[AW9/�&��-A��v��E��&p�b��mؐ�P��0�G�"��/ X�WK��{
Q=��TP�G��MdHN���L���%� ��=]���S�6�3�@��
y:o&�n=�^�v;��q21� ������(�Y��A8�a{��n�"��<����D3���}�9Is?��L�/u�Ԇf����}$o�,��F�^@آ�Oc����p�gGJ��j">v_	{�=���gb{7/�J}�
�װ|-��Z��*���~ܺ�γ���إ��J��C<כ�J$G���ߠ�6(.��}ȕv���B`�7�(�N��庹�������[����p`C����[��F��V��u"�ȴ�nڜ��,'/�iZ)�{4��Z���Ċ1h�A��Y�*6K�=�,�;��y�5x_=�%�,A�o
�Ӧ��.�<)1�vB�H��H���AW*3K�hj�(�0^��C���&�� ���[�n��Æ�"�!����x[I��E|�ɤ��5,�cA���8��"�;�}�B�Zw�Vf�G�Z��)���3p��`�����9|/�`i��N����͡���'�X/G�kP�.]��g��B� wj�r����~�\4�M�z�w�LI�_>9X?}��m����}���}�D3w�Cj���py��܉T�fO��m�sT�v0=�ƾ�Q����`y��*�z���������L������b`��yc�Rvq7R�H+$� G�C�b�:>7�8��х�	#�Ny�m��i������*�u
epc #1�P[����^6hC#f�H��%�&�Bx4(�~.���-�}Q�%�� ϥz�����iO�S�؂(t*?9����
���w9(y�;F�Q��?�;�Z�O dˋ$ʛ"|�i���!6÷��;H�ƪoփ��2�ӹ��%�]v?f�]!A��6�{����'2����Ww��:}nTā�ć��퇿p��	�J�X�fz\u��\{'�4g��-�r�|a����� �.yj�Ȣ�m�7��NĪ��A�?	����@�n�\13�>P�ӧ!���y��<}��v���>`(~7F��v+f�%�>�(w�2���c�k�Oy�.���Nʮ�h��Ϟ����7(%K8!+���$�c9�|��4M\%�z��xHk�c�2XOf����]��\S��w5��o6�X���N�a,� 5[9���n�4rT���eߙ��u��M^U��"��Yc$�؊q	�# �>�����{$���<�H]�( �m/��ӹ�X% ���	���'
�&(��o}���议A��,+�Hhy�YV�˚�w�9p�J�`�J,�A��S�^��o�X/�R��'���n�K.���)󟬗���&
�i����d�� ^���)C�Z�ַ��Fp�E5;z��5�9E=�	S��8�{�< ��9�T��"���d/���E��fs<4�{��!�O�+C�����6h�B��N�J�Ӷ?�Ůa�C����ʷ~�={��k�6է��lc*��}�gp��!��o ;�2"��}���W�>�ʰO�
-�:��V�q���|��6�lz��g�����UR�,E�y�1U�֙�wK^u�!,pA��9n|C�]�(O��yG�-u��HJ �Ag��3o�я��pQx%D�߷�~A����,)�2�'3�:���z����ᙣpP�����?7:H/�oz�~}������{���m�����ڈ��=H"#��h'Di4ޮ64�[���#�u#KK��0�eC��땆"$�3�S����"��Oך �7�	��g�e�淚<�l@7�,*���v�<��-Z@�������ɌJ(�2����;�ŗ�Uy/]�<���:�)��PQ�~�	+7�lc)Xqssn��B!�����`�ߛ��o�Zr1\9O�
;�����Ҡײ��3����,8q���?�2�v������kE�L���+L|� �J�df�)�oP�Q�2�c�/�s45'g/�r�GE�s�@�P|�z���l_g(��cE~�b�(Pa��ȟ��_�4���9�.�Ǯ����+<,9�}�_�EFi \oQ{y����)��(�' � _q&����Ny�j���Bm#vlpEC)v�N��� �%���ҹ'$�lk��w>HZj?�jy���9yZ����'�n^f��5��Xi�F��V};��Oܤ��M�GO��w�����fs�����p(�<�r6c� ˇvi��[ʙ���-�8���T�M��MJoۘ�o
q,��nKr���s7Zڸ@�������U}����?WhX��!ɥ�^�f*'�ev=�����I�y����p���pe΢�Ӫ	�7�2��CU�Ҫ�Y���+M�s̾c�h�8�ԝFJx �K��#Ǹ���~��B#Y�xb�n�<�W�<0N2��<�lCG+�_�r7�u���A�U*k������w�� ��|[vU��