��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ��nͳ�R[�ظ�_����Qq���G�]~��\�^�W.Z��ke��X�?�I\�zA@���Y"���a`MBl��$���X���/~%�cg��OU#,��;o�w�F�~�wy�0�Sa��qC�$�_됲��ݗ� ���D��.����v��C��k���<�$J��3��I
����<[�P�}&ʁ_m3�P{�
A���-X'�H4Eml�}-���i���[�f�c�:Z��� �B�X�p�v�ww-����9�9�=��܊����\j[F'���\��ӝ(�c0e�Ɂ�4aP,d��-��C=�#�룐���n�zRJo��%���f�yI����y:�+�og|�����}�0M=�\�&���F�>Oj@{39"�3�l�[�c*9�Ac��-�ŧ�s��Tpf�h1�Td�'�d�4�j�_���%ȇR=��>�5�z
��n\Ty�������9o�[V�;�sy���t(�g4�'		'LݒCL`����	��T���Y�����[���
_f���:#�@ ����qmV��Z\,�n�-Bs���QKVD*&�� W/�?�ݶ���܃4������P6~rg�����O\��2�?fS�H�=Lq�Q�t$�}�p����Z�tuX9,l�F-�m\���2���L6�F[��_�0#�Y�;�G��ͼW���5�HP˓t�(��r�i�x�M7q��Qe.��?!܀հɨ�>��nVFԎ�Tn��4��1�ʧ8ӻ�X��-���P�o{���u���q�B�'b���G��V����!���:��s���0�&��&W��&6���+N�W>72�~4�H�v~y�-�瀳8;�ىC;�Z+��#sX���2t�Jzǩ��f��8�W��nR���&���^�[bIZ~�����tOxң��Od��SG�+��_]?�R?�����!�����iY �#���!a�7G�\���� �L9�ɪWH7��s����_I*�XY=w��͢��6ɠ�9����ƃ�8'��ר����?�-�m
�%�ݯv|�J@l�N�r�9h	9#,��	��Y��:��F�1+s1�����B���]���0���diƹs�qZv��3���\�p���J��(1J���ZYUpl�����)��j>&p�vn�GjHZ�	�Z�Ye�@��O�!��cg�/+i�)��w���٫�
�'C��F�|q�b5�|�Iss&i�(\Q�2�)k�T��d�e-�Bc�O���H�9��{G{_fZ?����l�I���k}���xP��w����|�d��TE������Rt����B�X?���q,K�a�MTF��K�~�֋�<�94�X�ʩ���0W�:{��Ϳ:��
H��z���Nh�JZ'3��d�U���d ���BZY��oSq�mHE�5����&���q���ږ�vR}�O��w��/���bˆ菘�[J'y�%VOF8�d�#���m��B�o�	��A>���'�kO+��C�
�hp�P~Q�����E��I����Hb�/4&��rC����2��1��,tF'����x<���;�!��6��q՝^ǅ��Ӊ0d�5o��l�N��f���cA7<�c<{���R�c%X���m	lKA]���Y=L��*C��e���*��A���gxU�������E�����Dx��i(⿦1m(�'��Vz^𩶛X���3r��"s؂�iߏ*��h��Q�%��MI�����b��z��ZW<5g�d�8�p���3ځ�k�XOS"����#g�0Q+yЖ�"�i_Ej'�F�dӸ���\2J��}=ݧ���CB�؛Q4���P���f3>�����3U;���[0ɩ�la~��G�-��;v	d0����rҟ�)>D��BubXT��+��_�,2�e�IɅA ��d�rYMIRJ9�ʧ��-�s?�JBU��.�������tt�q��#���h؉���Vl@?���erU�?B��6�֓�6�G%��W?i��4:ڤi���sT0�Z]���Uݨo����BԷ�ܵ��I��G��0���tC�[Pm(Z�+��J�d�ŋ���!�O�`jz��r�V�>yF_�RQ�Ѝ��2�µ�	��bZE��Ɓf7���oVAZ���y�0%(��3�R׃ν���Nf2�K+r	Fr**M+�?��{�Ƞit���m�H�#W�ېJ�%D�:��u��u��W�!�g��h=���HK��P�h'pBgR��Wg�$�o��?MR�;3p�?5'I�2�(�h�M8R�*Zw��Q����HS�5�%T�tY�~.y�"UA~~�׌�X�����%������;�����W�u
;PvRo"�ĸ�#��С�Q$�%/��v>���\4Fُ�T�CDS�f�dC�a��YM�e:�@(�r�M��H���1�#�[#���+Xs;J���x�SC����q�b-�d;gq%������in�1��:���w�6�
�c�k[�n�/�csV<�7%���d�g�e��1�|PDyC�Y3�K$���qtG}� �y>&T�z�!�}�p��G��UKd�.\a�=T����){��|P�,C�m�X�Ѐ6g�DK����vl�m]�.J�[����4�Oq�J�S$Y�RZ�K�WB7W��A�)ʙ�P�+�<�U�w���a���t��ΰ�5>����|V'�@�ih����~:���p���	�fG?�~=�Հt��P@z��ݧ��WW��(^�j��f#�0�:�_�ݷ����M�[���B��Tk���`��L	����� �CC���"����N{V���p��/�=�z��4�h�s~�Azw��:�J��o>���F���ޜ�����*^e���'����GY�2�0�K�0n�(1#�N3pu�f��c}�Ӵۣ�hq���u�����;����*��v���=?V"����q����D��t`
��Ը<]ǚ��`�P�%�,E��w�\y ���od��
Ow�ش��oe�צ�&G`��+^h=%�' �ؘ���c]4/y�`�RU��;�m wɝ�M�BH��R�t��:;K
�b��&)~�!�Z���-))�eG��yv"�>I^7�d���r&t�~xȟ~�����MS��
{o��������_W+��;�R��-p�-���[�&�>nJs��X��2�����
+�ડ�����C��m�|,_�>s��.��h�'B�m����[F�g\,�'D���]�u�%}Ĺ�o�*��>���"-�?h��>�V�;	�j\�([���L��tv��?f&��1�a����e#2U������>�N��� Ѿޯ�������"^�~J��D��j����Aǎ��"��un8ZR���K����{�&�=r=d+�W+(������1��RnR��+�\�O�Q�o��ZX}����g0�����Ϭ��-`��bq���,Esy�t������E��x���r���[�߹�Z�ğ��	����&`6�y�$A��[�9̖T��T�uR��њ��x��J�/IyZC�Z�趇6�$�3҆��cQYxȴs����\��mQ��]�`鷠Q,�^��� 8�V�û}�-:'�4AỀ
kڃ�Zop�2��|�˗���$��:��6�F ݗ�X��ۗyǛ�����n�Դ����ck,[�$�v~K_�N��[+�%q��K������йY�!�9e���@���/�<4�1B7�S�u	i�����Xs�sUhlmXi�X���n���c)�NJ1�N��P=����")�S�U�������Q�y6H�B�3E/�7\���t�C��[k���ԩf�u�:��C�q�	�r��2G4D�c�%]ޔl���ɀqL�A��@q���F�&�ws	&x�@�c��8�ʹ�����n��\�.U�u����N�z��l�, ��ݯ_"��~.S?Z203��KH'�Π�G��(`y��MꥬM4*,MF���~�a���3q���ԗ`�����>A�����N�"������~�m�~?C��,��;�TK�5[k�TԼ=-\�]47tisV"�U��29SB�6� W�<���ua�	��̎^�GwCi	�l����+��9����O�	��֦��p~{l��,��בTZ
�X�y�L[�$k���PX}fg=G�bj��cg..ɪA�t<��JPO�_��v�I'�ZWp��z�{6Ȝ6���=�є b�	����A�2v�q(b���#Bg]��z#n�