��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� f
���O�Q��Y.#�d'���J�"����4���d�"�Ŝ9͜����
�~�a�rN�����o]y����1���nJ�]s 3L!��,���zَaw�{,���{�b�[;ҙ�u�\��������.7���}����H��ΰ�&���ے9��y��y����͍2��ё(��7q|U9��1���i��$>�[�G���^#fU����S�"_a[7B��7~ez�#�5��-������>[{Љ�v��G]��Ew4��5`�|x}��4�y�z�f�|#�դ�e��5p���1��L��d=�㺔��y���h����V���Q���t�̿�rբ��6�j�mcP�iT
���c�j��5�j�KL��tlV��d��x�Z��"ks�kCK�|�i(�;�����6��12�XTeP��[��'�0u ����r/X�<��/�]Gȥ���%N��]84����Uwp)
���un(c�Åf��J��f`9Fqv]���+�<�w �N��fѧ�h ˞�C;4��#�i��T6n�Q�T�����ڸ}�rS3�*�x�٨�j���y�~E�s�~+s�G��'��%`+�w+.}��(Jľ�$SL�2-�M�M�W5~���/%��t%���0;��3��G�rq�Ħ@];
!}ˬ � C_3ZjT5�ъ���29L��>ԡ��I�#iDn=*oB'R�؍����v��< 2<���oc�M Yx�R5��ܡ�����2=ړU��oLW9oq��4S�um줂f�X+��t)�a��� R��M�Ć8��,=���LIQ_�Mi��A�C�qW�����&��f����J�ӷ�&��u�6m�����Mjs���<�R\�Qs��wm]�	��$�a��DMW�0 ��=~��SipW� 
3��5��B�T�������O�fb�`�����67v���ǹ}茾$�Đ��z�=«+��u.>W��v����'-"���=����#�d�N�c,!8u�@������F:�ø-�l̶�sDe��_$�B�6�ҕa�ygϢ�AXPY�q5�[1�HNEj�[ ��a�t��CT��Bu�����c-| R8��@|M�:�d�{��Ͱu�s��is�V�V�����g���!j��@�y�2G���:�՗�!X���H���Hl	��g�:6S�M��~E�kw?����sV	 (u��~����ʠKML�(g+�:�o�K�cw�Gc�~�C�BϞ������v'^�x��|H���<=��b�ŝ�O���L'�5ޛ�E/f��	P6ĒbYȠ��>�ٽ��宰	���RL��W��Pݐ�ę(LR��2z�q�hK�KP�8$c]�ttG���[;Joz����ľG�h�Qv[���R
��	#�EnV᤯6��}q�Bv�y΍�����
���E�]�J��瀯�)#�@�_�⸆��bB�?�����9�e��߽����e0,��+���ֶW+EI�E�dN_6׭��RpW@�{��G8�0�x[S�A��8^F�f	�Yǅ��e1��toMa��U�9��3�%��� �ƍ\�hj,��7�|B��E���� ���^�Ua0B�Цծ_�X^�@����,��3��g2��������e3r]O!2wh� �Cj�7�s���_/�=j|��22�z.Ė��8�{#e��F`h5zڡf�Fj�&�d�8�>��c3�	
�M��A׵oDU���Ʉ�J��H���) <|���b�� +9|[����������@�8� /����J��
9��K��z�����;h�Pp1�w=g z̏K��P�q)0߬�O|��.LX��E4�3�Lz�C�8wd�8l�e�rǹ��D�����P�n��7�*���?�'��^QW�?`�%�Q�0���0�ӯ�@��"77SZ_}��o?2�,���+m�t���p�K佳qa�j�y�[}���R��&G,*���!r�}���s[��iw5gr�F���)�S�g&�Q�7��S�ڃQ�9��Է�;�7�.MB_�+��	�V���l�GO�iT���ԉO{��^�`1
����LP�/[��m���׹U�d#��nCpn�[[PO�!�̐�&�������.2��X�6!��ܻ�Pn���#��ЯljNP���L5>�W�V��n FJ�V&�,��gLˊ\�������VߘJ$���f�Z���{�㾤���vG07�������H�fLa���4�����uaDI5��0�HۃZ�G݋:����/f��:^�*?ъI��(e��
�m�)�]��9�<"��Tk�d=ȦaS����"�B}@/�w�f����.�l��FKm�X�6��T�Z��.T�2��u��}a'����Xϊ����@4H�ܙ���[1�5�[��rke�ְo�L?�Dm�a�c�BM�l��Kb��8]���ӫ�;	ʂ�"|���������W�^��.H����p���D���]Aj��-�P���:�)H�2$:;�1s�Z_�T߮��2�/� ����ر|�����,�Ł�K�J��(+�s�Ym�(X�sP�e���8�7��0�
_��P.��ȟ=m#θ���?W!�("�b!�^�}"����X�O�]d�-��cU̍l_��z�a䌛T�x�
��0G��LY�e�O���:9D����l�������OaXvu���₠o`����u*׊4�;(��9�`�b�X� �̱�D0���lIk��}P�%�Ȭ�(6�S��� �y��-������>��!�n�l�J���� �vgfs
V����c�s�YY�&.���¬Ǥ`e��M;_gN���<e�M��.X&C�L�3�LM���,O�g�*���<�3��p��^O"~���ds��LGA>�t���� �ˈdjb@0������h�B]����c����UU
H/�U�g�D�iє!�.�4�I������l��`�<��6m��>!�W,޳-4и�]F��[��V����ꑟrn&���1}�
>b��U��������@�s���COyֆ�"�f��X�;�v�[�ц�J�����3��PQ����	�
��~���D��ugKV�A�