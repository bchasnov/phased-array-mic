��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|̪��q[�dZ�db����v/u�iw$o7n��/��>e���t;��5<Le,=7�<��l�p���'����35��P�����-��0q�򲘬��8��$��s�Ҕ����l��`E���so��^�h<���R�ն������]��b�A��}�U6w�iQ�����"����/l���H��ɰN,0�N}�TÛ�b:=]�;�fE�� �hϪ+�9S�Q#n��tf�ȸ��^�@��N�U8�Н�id�RL��:[���m��X��a¡7_� \R�喢�˞�L(�򀬖�ʈNe�;( [�sp�~h�� ��
���'�k���&!{� �+� 7t�;���1�Z3���_�1>�"�CU��\ޗu한/c��'t�� � �2N:q��?�Nv�>>7|����@�Kd�w���A����J��d��J�Dq�i��N�؝G��5d!�ɐ�	�R�KL,Avv!��J��膎�����7(^��Tw�4��/���,� ��H���B�U`B���e��&�ͼ-ܙa��w���K'T71

��'�L�����z���'����D�Wϲ�'��?���Ŝ�*Vl��3@aYNn�����G��NW�ܱO�����_{3Jd2�"���(����y���*����߮*��� `��~��JSM�ؙ�j`zA^�vy���a�%�'�+mx���)
�{��PIJ��Z���J���6��#4�_�sZ�56["���\���>�݃�;}�®UAoT5O�.-�{��è�NJ�  K���Q�9�L��b��DS��������֓TZI��=Z�wca.�0J쎷ʅ�ګusJ�n~u�Q�!Mη-�(���ܗ�����fH���F�k��2u�\t���#7`�
�����"�bV�N�i4XRl)�'�q�D�IR�7��)'�4rN�K�z��J����ueK n�������e#�J�!�"���Nx��Ƚ�>�Ȫ�TpQ� ��b37�"J6aM���/�^T����2��C���Ù bQU�Xvy���H�>5���y�Mbg'3D��/8��V>�`���mf�m�x�s�.����
�Ml�UƠj��>��l;�=�?�IT2��_��F�E���H1��Ȑ����_v�(E[8��=�)�w־UF$�����DZ�YH���g�)���UU��S�W�������e�^���������?!�#�×��N�9��g��w-�z7G%4��w��@-q-�J9��	�q��x@���9HJ���bM�Vg���8�֎|������$婉�T�:��r����]�]L�@�b8����!�$��f�_̺�^�8s��?}��xC�W�A0������b(̅������� L�լf�:�7���8���-�;����u���<#���$��:��M�z���kf{<Q{�������Ɔ);�ɗ8 �v"�+ba-RT�3���Xg�dZ����Eɮ��~�Q��A���X,�שk7��oK�(��K�y>���x����3���Y�F�͞Sa�7��n�l�P;d��X�������#&�����kb׉J�:Z��zX1#%���8�����
%2㩝-�6�
���b��}�#��67"����A��,!u�ٴ��CH�2,-@�^���<���i��mA�`�ػ�� NĎ|c���(������c�КXJ4W���(����V:E�����1_#;���>���xVa[d�N�?��zP"6t��n�+����ȍ��z>�̖���oh�XƖ�=����,o�Q��s��u^n+��bOJ���܈�~lIi�|7�r:#��ux2|���p׍������>K"����2����P�S�j�t�7����5��F���o'��I����u�Ah��At@ӄmJ��!���ْ&�̽��"Җ8��j�=�U��j|	����yn�`�IhM�2wY��3����I(�	"�~�v%?\c��;fUy�5�\���W��ӄ��K�J���wB;�+��U���{�ʍ��>0�+�['�@�"����:f}�9D��U��\����᥇b��=�=����Wz(ʴ����O*}
/5{9����X Q*=�b"��E��?�G�I�ˮ�u#͋4"ώ@� e�ض�"_T�y��'����r�G�|��
����X��b_�A=^a��!m��>��g�!��^�Ƿ��X����@O���+�쟱tr{{0��7R�nę�[d=9�d1�/�3���n6P'��w�}���|���bŋ�mL��T�������
�)��3AB�tC��l�د^�B\�g��|�a@73e4Q��v��[��*&�yC�������@Jf���\\FVMJ��_u��|u*c�ָ�����R������B��c��~h4hP�i�����;�v�?���l�<�2�}� �pk�f��6��c�u�;ze2���,��Г�C0��'���v�ї@Tu��6$C��F�_��B|���(��w[���g����`M��\��y��1b2�anO=�n.S���]����r��f�	G�H��l��Q���Ap1��V��z>�1n-�MYM?�=Y<���Q���K4�8C�f���?�}�Ymn�d�Aƈ��C��0�'��^(0 ,�-�'���zН_a'�cC0�.\��O�E���+~�<S���꣯;�ru��z���Ϟ�c�t�&e�s.� Q�.�V��9��ӫ�/=�w��CD�X����òZ�D׋�V���zǎT�<��ʿ�E�dTD;��\�F���+�̳��Eտ��'�2C�A���T���1��1es2��1��gr��>�.%>���v���``ԅ�~H0���PG����R���*`��A�%s=ߌ-d5?K�H�vY�#S�%�j�Mk&Fu黛�b��M�T�ƽ �Ni4��T~҉G��藈	gZf� TV��y�E�O�p�׉��
񩋐X�g �R��ӧSE�����/0�>�D�J����?6��� zܕ.�х�?V��uE�b���|�Ė7�c����i��-}��S�a���8'����C�΀��ڪ��V�\���[�w�i��VS�ߤR϶@��?ҽ,ˏ;*�-<���ʖ�t� �I�����d��b��$���#��?��`w6V����/AL�BX熄&i��Yi���0/?[P�|�����*�w�)����I�=#��'�EIh
J�Ȫm�����6����6�M����q ���Ac�� 1�ߑ�Csk��/�*��\�hÄ��rY!;�n�O�X��n&��Ǣ����R,�A!ec�6��:����} ;���K8���sM�6%'��^\��h���-��& �b���I�h�K⿪��I&�/=�-CL�SM�`]���h�;����Ysmۦ�d�H��V�O�=z��j�͟���Fj������K���~��RY%���U9��$����"Ac$'�P��^2���/��`�b(�3�v L�Fi>R!�	w���q�i�3ϫ���~̲EÝwar�4#�~%���"�M�_�x@>�T�|%��=T�~5� ZE/^����f;�&bVVK���t�Z�3�Gѱ�{iD*s�z̰���������A�o��9*��ͩI��ª���9��n{w�����s� �)�z�J�g�bDj(�ՑB{�%G�����^9��*����$苟�8��a-�^��k�ZIe3`{�i�WWa��4#H��/����[8��M��A�K�{���׹�:�� �/��0�n�vH����:���I[�x�R����DҊ��֪��d#p�ȁSg�T�.�y�������UN����j��R]��1�cU�ꙟ�$rt+�:�=>����&�nK1J'��`�D�6�r�@Sh�[�b��#G3�c��|/�&� �[[�XНB��P��J�{Y���w�M�/���{�1C6��9�;�F$��yF��^4��t%��+Tiϖ?wp��	�b���^�?�Kѧ��e��msͤZ�p�4)%���&�{��[�o$`oʦ����Z��̼/�S�ȵl��1�"��s@O?2�Fr�ݣs9*]�́"5�6l�7����B�hY�&���I�}[6J5!3�
�Df��@��@[���t��> �ظA+��~�n���)����
�cē�F[��+F���R�Ҷ��g��ɗ�Ŋli�<m@t��@M{����t���>�q�pO�S9EɲT.w��\�;=�o��p���~����: �����cl֋N�� �Of��"���c5��p���ڪ.i5���J`�t�g���$���@'�4�!Z���H�L��U�`z|1��Y�U���I��$>9ɧ�u�e���\A��	z� q��a��k$�=; ؉ov�d��r!��{�m{X,�����l�<!��^Ci��F��Io!��~�����m�&�o�~]��g�ڨ ��\�%���<arMbVrT��߁��0VH��(ܳ�p�g9^!P��������_�q�Z��L���0����Rb'&
�]>���NTM�Ri�o!^ V{��GA����������&�r��3q#
�	���?�,���jE��g:�vۜ�1��<v�Uw՟b��x���AD�I 8d�F�,z���0D�'�2^}8b��pq����,�N�?,v���Mý����~r��,���p���r�vhF)�(���>��EL�_y���|�OO4H.I�%bM��#�.�p��T��Ni�s�>�N��]�g�6�hY��M�&a�t��?��c���2�{�oa9���Z
��^h�A3X��$�MmT`�PǸ~z}�V�A��v�ꥏJ����U]�8zq�Ey�ʢ�Ŷ��H�<B	�U{���P�11�h
��=�y��p[�#�Uz͸qkb!���-�]��qO��Ӻ�a����
�m���뒘�6�kL]�!��)��qo�檧p�mg&�	�,7I��j�J7 �Q��)~Z�� eue��+�Srf%��8�y��5&�!|�p��d@�������*�\�dT�J~�U���?��v��ȬU-%ct�N��R��ll�6����jX�0̋H�� M]� �'��:
�|��Rr�[2F1\����Ww��Ɇ����GD: 2ђ�z�
�,�p��p>���� ���^�` �M�\dB�V��IW��Bn�H�V������_�8B��o[��*��:<x&(��K���1mН ��%�"���.���b�8c�D��a�=ʥ���OrE��|�!5H^ �_�|k��b��+�UjzH�VP:����O