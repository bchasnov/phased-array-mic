��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|��We������ƌ=�_�F9�p�Y2����c����K�9�SNl�@\�\A���!��=3�������+f֝�Q�h�z���ݡ;��
`�V�u���#c����B�[��Q��Y��:�3yy�z^��ks<�`K\2��$(�B.��7��n�{=��$�OgU���T<�<��5��y��R��j/��JU� ��T�V�Ard·ڞ��]��4gO�X��Ml4���ab�	t���<{[���"�/UW���p��&B�<qV�ݺ�&�r��v(z���t�>\��� ����C�4�
$����oo�;g�\���V�g���Ԟ���(��9���G޴�:�#�����@�{�8�è���9�_�x?���G�L�Re*�)ꥨ"�bYm�da̘�/Ф�8�CI�����玽���Q�ٙE��2��X��,�}�o����S��þ<��(+��K͖.d�}=�p�<���ê�\'�r�WXS�Yw����r�d����~�e�o��p�U���!���0�l�(����C�6R�Ѯ��u�n��)Y�{�������d���'�[}`Z�I��\��6c��c���r���9U��#�Ə*[���k�cC��$L���x�29�l�͆ HTغ!�aa�����+?�o5[��M�j�B�8�@����c|sӥ3�����ݓpf�U�.�u
ks�([�U�B��¡ڧ_�1Ƕa�={���g���mI��\�����K������#�MCk�%�#�A.D���,�8�/�t�
�A�{��Q�̸�6|�6׳.�i�N6���r*����H�RALY�[:����ו�񴺩�����/{��y���uu��[��s{j�rw�'MΚRAj�O��?�[�l������CV@K:����Y��]~ā�E��+r�9���r̋�Kڅc�ֵu�~�l����N��#>����<���|E�}�m�:���������E���	�j*2�tR�Ӆ;�*�S�W���#{|b<��􈠟̣4��R��>�}N�~���"!�%Ĭ�-g�P7�
��U���?n� �Ѩ��ѩ���	�!�+��|�FTp�AգLF-���^p[��I}?��-�VL�[�X�������Re�mJi_��E������d*�E��'���>@�����iH3V��>9+�F)�"Ȅ�l-��3�3��I*ܲ��+_0a$o;Q��i�Psn������e�b��(pR��$v�a�dN�-�o��e����ބ!$��á_V�YCT�`*��~B
{e�K�|SZg����k�bt�u�j�5.v�p��ʗ��q�@,�'��� [i��ou<�쮓��μ��]
���́���<3�Ii�H���)z���݋[j����t7�Y�0�݉E��
��9`�s�,Ӏ�trOtR�{];5M2cQ!�P��^���+�ƽ���O�s��}���٠or6�H����JJ�w�KT��VՖx�n_>SA)���[���l�*bw��ț�A���]OMH���/̕
8��+���ZG�R��j�ik�J�!�kn� ���5��]��e���"g�}����=֍~�]��qY�U����r��jg��wZ�|�[��P���fpCI����+� �����T���.�J��K��Jc�E�=��g��I�N� �"b�h��XR���E
Z�Dyv`d�>:M1e�9X2���S��[�:��pl�fZ�$qm����l�����ѿG���w�77��m�U"�yC�{���"�.�"���Cb�䉷 v�`�?�k�C�X�3V��`�0�\5lB�����k�(�XB��pjq�̌za�'���~�A�Gu�y���c/����jy�&^q	���������U�}B-�h���K�k9[�����}�A);�vF�ͭ�&��Ѥ�a�m:�ۥ�QKl�Y���K�kw"N�,�ka��.�|i�l��L5c�����p�kaQߎ��.%�C�JG
DpJ��>rO�+-���AD�JNF} z`g�[-�����4�/u�U��5�N�^�H���-���Q��BDGM[}��uϤ-�P*e�u����d֥�1�""�\�AC��c^�;oɴ��He�q�!�w�JmEVc�s$����G��Qg^#����w0ڠL�eIݢ"/���e��4s��핖�}��c�%W�y���(�@�_m�����K)�vں坘�n��68�#A*A*��nv��ҵ�|�G�F�¿[]d>k���ީri!���7��'�����e�~��G!���=������B~�h��3w$�zq9�ѪH��m���$Ĺ����l4��ﭕfu�'���Ĭ���X�fAAQ<�ݒK+���cv�� yI~�G�s�u�f�<��'���ѓx6#p����Cb颒��/�п��LWlr�^a�D[( ;"I��yz^�@jV�Tk۞?�< Ӑ8��Y��`�|�qu(����%�W`�E�NB�����#�I��3 �w  FZځ�3Y�,$���⡌wD�sm�mY�vu�9&#��dD��S�	���qz������ȥ��~_�xc$�N�of\�\r�߬e*B�Ȯ���IZ���ƭ󅐥�}:����t�p%j���pwhx�1ʴ�ڰVPk*9��9��I�e�w}��l�:30zϟq�37��h�(�1~QW�릹�]�c¿��/h�w�L�b���4�f��[HzUp��<W�牷 qbS��y�ۗ�t�ϝ��ݓ��ֱ�P��0����&���w�_�#kK �+]�%�+��u;lп�+������S��,�@5���faGmqOA�SQ���?�vzh�?4g��lc�%���@)�g��qړ+���_��'�!c�=�18̻�Ȱ�.�zqq��/0Eόmi�]��@�v���&�c�~�O�ُ��,��-P�'x�U��u�h�5��_��;(��)�Q5����O�����v2���C@*��2w����O\HeC��=��f�bpΠV�KPV'hg��0gN���U��g�~V%E�p+��><�K��f2�l��ߵ.��G4�s�C̃5�O�Q�w�@�����2DG�����H�W L��B��߾�f��P�j�|�},�}1<ٽ5�j��\:�N+�G�)]{n_�[�������Πg���D�=zHݱ�AB�9�?�z�=�-���L�}��g�/>��=#�O�YP5��Nm��U���F^��*�������\�8j�:L�y�$��eWπ{PY����a-����Ť��/�P]�+x��(�p�--jY)�����s�\哚G��uw���4U�=sפ���q�v�� n��|�1������Waƞ�=޲�3��[�CКG/Ʀ��ӟT&H��'��}ӭ����ko�����K�m�w�K`��:�������0�+���E�Aa��1Њ�z���7e������8x��������I�/『̍�ϰ�mr��Yi���A)G���g8滸;��'#�Ӕ��ֽO#Ԭ�à/Dj,�ĥ]2[�������lǫ���Y/g��Y�/�MWAC�D�z�ƅ����o���w�B�_�$��c��.�0Ѭ�f���ec�W��Q`He����@h�!�B�|G��)��g7�p��@�5��x{�t��&;�RCs�eM���V�"Ȁ�jq��JLR�z�ųj��K|* ��L�3k�ם���D��ʓ%�@й�h[gd�G}�_�Zٻ�x�=C&0�N����l��ڃ���@��PD=�d�Ɨ�s'#z�b7߃����zaA��#�(����T#^6!#���s)+n4Jw���xy����e���i��:��������*�Q;�'	����LP��L!=�3I���/�EXfq�5���e��+�A��~�1��c��,^�і�X�w�K��:W��TQ93�m�p!~�:�˝_�L���@jRo�pQ�H��g��P�} g�5�ӕ�T�2�f��P�b#��V��A˴�)�y�K���1c���+-|�84�g)�ϭ�:{��n����g[W4��*e"XL���(�-�hu��|�,wW�;�6�Mv��C�H�:�:�X��5�XIau�1���:{|�����+??'��N�I�����v��>���\E��D%�o�
&�E̴~�z���'�ԟ��Y��Qd}^�0�k�A�����W��Z�9_�����̛t(�X�a
���4M4���
9]�[ǳ�h���W��f�Đ��"ɧRm����8h(=>��P�b����mK����ZF����Nf+�]�W6}w9�9����՜A�En�
�z�bV���\�,��-�L~2����Z6��c؞%��B͹�Q��XV���<�Gw��wQ
�kfJ�?�^���n���x�<����uYV`L�L���脆�x�3�_�e��w}��.�=Ӳ�[����?�.V��$+�p;�ȴP�,ӗф�p �E��b�~F��4ꉍ~��G�Q1��_�J�w=N�Z��M�{b4��D�����Q��P�[������ű��#�Rf���C��'��]���TC��!�[D�V5)�������+_p�
�S�u���;kC���%q���� ֿKHw6��� ��4m���+ ���ZCAl_���B=�_v&����R&��*�Ƈ�����|MY��݀�o�k%���A�9f�QQ�¶�9����e�����k�Jlb$
xԎ0��Y�E����������!�V`hDtݺm���?i�2RmD:3-�����0Sb7�(	
W�9z�0槂$����ފ!�AESh�V�Зz����t����lI�;��p�|	�J0m�s���������� ���FK�$����h�te�G� Yw�.X�����rgvP{��?�:@��b�;p����WeW��� ��I�,�����hA�*���LE��T-���
�A�aգ�Z x��q�E��l͇EjS)��߮�dL<iF��ͥr)��\�A��a��苵��;i�:���Cѳx���
C�!ʄF�V���?��A����8���3�O禵`�9ф"<�����7Z��n���h�v���`(ۡwLE����l*���	��1�֕cl�^DZ�Ǧh�t�7YZ%�BZ5��@�l����#=#Ba�|�>Jm��oԲ��x����mːkcX�/媎�s�FÎ�xÓVDr�ܩ�б����8kr[�a(��-!~^����o��>��.�|�m�:�Q_@y�[9�BrgX�G�� ����y8��{*m��3�v�ve7���m"#�x�/A�{��%%ԅG����������Ei��S5"����6#�(%=�KFMљ<��EF� ��2�	�g�j�j��O�װ1s�^�iΝl�mbfv'���H��^u��.c��(��鿵�^���l]Hv~�P�	��C����d%����g��j}]��R���D�U�>��Z[̡k#�0�t��g����	 ��4��b��b�qZ��� _dÎj^C�R�omd��q�!y�wl����K�u�TY��u8.S�n�H]��͕H��}~%9��7`���B��Oy,R3�I�A�믳jQ��p���aȰ2�a�Z�;	5��d���|�:Ó�����,���6�'W0P�����}��Dd�ޛ3� ����X���'���,ʸ��?ψ�Ì3�iZy�|��O[�e,d�+����
2�*ۢ����	�m�.bnNI1�RC��r���&RҚ{�-��*\/�wB�h>�<�R�fx��p5�����͓ܷO��k�ߠ]R�l'���V��-�:~�6�=��4?V:�]9L�@ޥ�I8o]���?s+e-�=��๯m�S΂�ԧ�SF�4��R��~�Ug���7�L����y�7L�\n�l��p��l&]�cQGD˔��}'�I�P��P�$%	���5'���"ۂ{�T��#|Ƙ���0sk.�L%���n�����6�*���1���ږ�|}N��=$����Sȸ��[h6��^�S����"�;9	�r˰�nU1�C�������r�w<ډ15�c�W�.w��NyR�L\�;�!�+��-��u��x!�䧙���Ӿ�׀
��7=.���fVJ;�w ���Ұ���9�G<QGj�=e��#ï�?����^���`d���XSv��D�C˞����R[tZ-���Q�j��-̓�w��i����)��&�d�
;���{���JH�ۯ�f�.�s���)�~Y��S������Q%�:^�8�6��c ��:���U��(&�L�2�wP��1ཪG|�
ͧ$Ie��[�DZ�Tb��~?�ǘ�GQ��zoP����D�Sbg冽V!'�Vs��4ɠ��4�U���WJ�Ly
Z��\��I��g~J����cw�C�xrI�Av�DE�Q,e\�6\`�6K������Q$�X�b�6��[��k�~i���o�c�w1WH߄D�)��;������T/9��Λuvf��GX�ȡ���C*}]��JV�+Z�5�G�I�G=�@�L�-U��x����fO6]}��ǅPm��@F����xS���T>�97>�*���ȝ����d�ټр1�����C+�B�$�F�g����cժ�*͕z�V�)q?��Kj�<��Se�s��=n�'$����ŕ0�BRG�yMݭfH�2��B�ήos�g�����-����QY������{�S4zH[& �cH'�0�52)�]Q`���j����G�;���W��Z{�W�!�|�r��J}�.y:���$��T�\�o=KP��ʒGjL�`��R�К�~k��1������r�k�ۯu��5xW�k`41���o�_�:��or�+O��a����9��2�U�B=��l�1��yЏ�!�L��'_W�j����P<�_��)�2�k���F��A�ڰ����ו�G�ݧ���ݜ�X�Yu8�:H1Qw4�@C����Ys�xoj1����x�����ŋ�'��\v�\��L�)@YC)2;eDН�w<nV��"ݣ�Z����jU�\�<�~M��:ʹEXi��9���>apK;O���;����z���S6�4č�׬���8���H�yM��^h�e�}aBL̛�
l;2R����Ue&8&pa��D@��F��z�X]rE���nS \�������0�׹��Ia��4�f&zߋjm��\c3�iQ��'#*9����!<~��K����C�Վ����E&�����
|u�tW��g�੥�&.�-��T\�����!�X�U��§?�3�Z���Xl��1,e��z���)�q��3/^��uط魫P��Sy�=�V_�ܲ ��@X��)�� 5�9����V+nV��p@J��1@��
��/8��y��Ik,��K�9�{plx�S�*%;��xG4�	VM��د&��X=`ӛnVh�M��$��Ge�?^��s�4��V�|QjY>��Ԡ�)߇���Y��y����f�[�}��"b��9���#�n*YG\��i��r;~���������o��|��ʡѨ��9����J& �.n۲\v8샩>���rQ��v��CX~�Ī D��>�9+��QXE��i�����)v����"��*�p&cnÛ�}~�\ԃӊ#����pF��8�z��������_�P��A�u���4g=�:���A)=)���j,ww������ڨ4i�����bh�_%iz���2?�u�?���9 � S��|�΋=�`)��|�rN������v�Z��!1�	�����lY��KS�F��� YKK #4��3�3?�������_��>^��m"هmsu�i��BY�'���像!\���(G��P��	7J�^�����O�dZy�&Z��%t�/uh�s��W��شֽx�B�8e���t�hX�Y1w��ԝ���9�`�OH1Mɟ�ٲ|r��tM����+�}����Ƕ���֔,��k����$mܬ�?�Ov��/�KX�L��g3ڬ'U1�<İm�d MX�xXAk����q��߫�ۃ����7�mʧ��p�N{+�r��Ue���MD+n/wh�h!��U��U5/��fJ{��J<�f*��ь���C��8�	��	˄c����v3!G��4G\t+hv���f�����[w�J]�
�EI��ʌ�P�C���?+�x��!A���ưl�!:��,]��������kt[iりQ�:Z��C�N;�_�T���-�s~�Rtnx�%�b?�[`����y믦wu����F�1L��lu���!ԂYs����O_��i&��$]|�e�TQUX��{K��4�찘����0��C�0S�� �l�ݹ��h&�O��t"Y���D�n̘���Pi]�!Q�-nK-%~����f[�.i�=9f���B��q�Xa|9��I��i�8h�0|5!1~��s��[��YQ��[���a������X�@6����?�k�E;X�P؊D��J��i��0 s�˟.��U������R�sv���>��L_m�y�ԅ���� �� 9u��`���%$�\P��7g;g���������T�]W@+{n�&����݅Lu1��|�O��<��u*>W���}�E]]7^C�7�%�Q���.O�9��u��8���R
x���s��V�2�����e �:�.t�I t����2?�M��fY�煂�@ޱ�&��w�2�� <[P	�x>%�;L�����s��o�
�:�Q�����
������J<p�S��y3Ӥ�ଉ�0�N�@�HR=�p"��J��-Um�}��]�Y5���)_���� M/ql�
���oC��_#_v�9�%�%8�������/6�{�*SH��>�d��	.B�Ked�!�ʀ��n�ָw꤃�>јZe%������_J�V�F8�Mv1���.M������c ��Q^G���(������;���)8t�ח�۩Ѹe�,��G��0j�&o�P.Zi�O�D�]۾�{ ��T�O3��`j؃��{�B)x�{�����	J��#���E���	Q�a#O�N�ݱC��$1�L�,)��i��<��w��;d�oU���iVH/5��:[������G�T�SV�m1x�ڋ&�N/�u*�Xڸ�X
7�[���>0�?/簏:�)zg� �r����j��4#D��6/�*��jn�5�f��H�k�Xd�^	���O-�X?Q����Q�Gp��J�mV��rUe ����AӚ:E%b��%g(A,�<�|�y�W�W���Mw_`�~Mm��4B5��Ut9���t��S�/�X*����j��[rNV L��Z4�xJ�T˕KJ�Ӭ's0��8A\��x�����f���.��"v�[��Fx�J235$�r;���[��d!u<.�̡�q��7���?=PA̿��Mx�3�n[�r!��J?<&2�!nb��\��"�"����l��aYhP%��7��_J(f�y`Pq�a��oR!��K� ~V)���y�q`�]ҝa��	�y�F�N��@�Ԩ4���O��T}t�ң��ѥ<�\�S���Ur���y�{��%9̼V��Y��C����p�&m��Rn!��oHM�3��E��8֟On	H6_)L��l կ�m?9�t���ݲ;-㿎D�|�Ӻ5^_�¢�6�o.���g`�❗�4��a堄����P�&���K-i/^��f�':�GO
���3n}L�@�#MS"�H�Ǳ�^�E���4�|�#��On��y9UP67{R�T2���v���&t�R����/��UTa�~�����`���iǤ`��֧�%���_Z&l3�|G6��^3�gV512'�cJ-��9�蟓��J)G��%Wbq����[�+MB����yu������W���.�������a��4�T��zW@�S�M�Lmf8���y�N���e~�R�V0�@f�f������D��_�=�(���3�#^NAGw8#`��)+Ϣ��v�.��N	�à�x�RӢC,�c�����h��8�+�g f�G��C���t� ��z<�KdB}�z�I�慗��7��L%�Ԍ7�ǳ�<�FyH�zà[&5\���,[�D�\��j��2��p&�[���T&����l�4iEmC��G�&�KCyA��{Y���(�l�ѽbY�Ѐ �W������#(ge6�!� j����ba��l�	��}8�����kA�g9��n��b�s^Fd4ą�uF͏`z4��A�g���
~4�+jj��,Ď��LSȻ�[�_{�"�u�.����X�x_O���Ǳ����l��*�C�e�|��X�c+���Ee��rB@nD�1������H\q���Y97Eu;ڵ�;˅6~�X�e�w;͵z�(b�\_�9�Ւ��`�r�:-�=��LK5�,%����i<�G>���1/4�P��ߖn9W�i�@w����������3�p�e����$��mqý��3"V8�*��9�סLn��|��&�\oٚ�[��}W~0A�m���A���?|DaxU���ˮ$��x!�ߧ����V�X���kE��]=��I���L��YJ�3z��^Lm����:�'��(�_[�\W��pJG�_`#H�jW��ޔ׻[ԥ��D�u1E�ɋ������E�̵��sC�T��~��C���<����S�^��Z���[��Y��!��O��Wu��+���|a�=��i��-��ϬR����ܐ��.��z��ؠ�jC��A~,��r�v|�+F����Z���K�{s�����0=�'*PT���p�,%�9��5!�SZӠg�����uT��C��4�fgaħT��k����im<΋\�������F>��.g�����x�ޔ�W, 0���V�%������Aդx�e���@f�ۭ.a`y㸊A��Ҵ]�����̲9K[:��Y'�8%�A�(E�>���`9�	��S��2�.���gE�'�_*��>� ��1["�g���gN�pA�r;d���v���G��Z�?�,���S.!4���