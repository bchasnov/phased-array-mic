��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\����q�?��e�I8�b�Ǽ$��"����ׯ1�V0���'�#����#G��n�3`���wx;�#���:�@��^��큸$yL�r�I��Þ��П�v�����9�`� ���x�����JTp���'�IaUq9��<1d�.��g�܎��1��H�I����'�wD`��}���8m�ه������Fw����	y�TǮ���	CObv�KU$s#P�QU�{�����e�
���+.Ӟ��4�w|��'������{u��z�����+r0�ԯy�	��AXejKw<���@T�h�>����gՑ�̘�Έ�9:�#� �o�� (1:���pQ��(��)�C���qM+Ds8�n�*#,�v�	��~�)CQ`���f�bxg������N<gQ_N�*I��M@<~;���Ba����:@�>���k�n�Zs=���jG��s�0U8�
�K�n)��,�7�[Jt��B��7��m˥ kՇ�pe~�"�2��K"ic���<A�1�Y�n|�Bl���i��D�E� ~��b[�� �G@'�i����\��קe�t�rNE���q�pǮ_����������6��z���M�1���$�ƿ%�e=dU��m�-�Y����~�	���is�\�pg.Q����P�����}5bR�N?�	F8ܯ�;�m��/l�����\b�f��F� q���F�������5�f)i;u����p=;�!�*gh�h�&>��������߷���Sp� �����`/�Q
��4\cN-)O^���~��е�D��>!S)n�9��#�'X��d�$�i:!�w�c��u*YV��D�ᡆ�T	��ye�����`�_��HH\�=�ʦ���;p=�)��!C�>���wjRWIH���5�z4�/Y�Jo;pE�u�Ȭ�A�{��X1�QWV|����s���!�9�� �%����&O�,���ؒu4乛��#���	5�sH�1�V3�"Z��d��1��z��T�YQ�_"-??�%��ԧK<�}��$I���&%8+)��;3{.��a��]9;rr.#��l�W��ͽg?�W���]`�W��	'�*D8E�W�l��ʨ^���$씆Q-&>��~Y'7�f���
f��s����\ᷯQSCB���|�&O��\�i�_R�ڦa�:a�Z#�1V��`�����Ol������R|�o������(#E ������&���FO4�;����F�E�Qe����b��|>U���:��:}0�̉`0rM��c.��k�/w��J���%r�Ճ6��k�'���컥#�y�)�_�ܐvS�������Z�།j4�5g�����t$����o>|��4$a�!V��{멲Ǎ�w�~B]t���!��Cj5f|}� }q�͉�Yx	���A��p�����6n����RG�"���x�N}��e	"�4� �֠�B��?l�$���M[���b�#����GW�@Ym��9$�)�o��O�@�h��pۭڏ.�����ӱ�������C�g�6]4��s���as��
`)�ROfg�(?�g}���w�䳐;��ir)�Ø_Z"b��_�e��My/�r!#|�l�ƽ������;ٗ ��H���@2<��3C���mH�� ��zP��E4�.�A��ۼ%u������/���x�������!��L)�2�A���{Ht꧳��rHm�1'�9�L��6���N�횇%�tV��;�0zZ�GK^bXF6�_i���o�T`�.� �"�������~�\�b��/��)^�I�0��J��O{�y�l"�4�0�k�-����dh�����$-��f����xH����'��%".:�:��+�n8�ѷZV�~�)��;��_8��(Q��O	��2�j<p�Ae�`����%�$?�#i}��B't�b[�;�:���k`�`ӓog�!�]�C�Xn3a��ǳU��i��P��EEhzfQ� Y���G�;>��i|�xB�fB��P�*�s$z�����d�@늚�`I�K�1N�^.�U�R�����d���	UB��ЅV곲�x���Q<� '�Ժ��$�l��޻8��D]��Nx�o�,M��O��"�g8����oZ�Z�2i���)��8��$Wb���}<l�h��1���V���d(���^�@l�	/��eTކ�}@��֬�w[W��Aa�><p6\��9�7�r=&&q=!z�#	�^F�ԏ e!��?y�5I�J��S���Ŵ���2��~UT�\�X��M=ն�j�R��t��1��N e��T�
�ԃ*���X�+��6����z�:d)[:'=�n�;+�H�#pR��z�e?v�A	-��W�N(ݲ������Zy�^�" 'L_��u��N�1�AM���CzY��@.Y��Qel�dÎӸ%{�9R�x�����[^�.�h�8,�� �A$��s���,B�q�GOS��/�)l�>]�FOj���Dn�p��ѼP@��W��3_���?��*�3�?���^z˚�S3h��fW�c�A�����ۈ��ӛ)�3��1­ל)��w!tm��/�8���ի#��t�G����ZȭW�d��N�����|�<����կ����l�Ĕ�ģ��U�#��-�Ӿ�q�6�'Z���B�!�g��5�|�|IA.rl:Ƭ8ǎ�ڮ����F����͝���+�}ե}�̢iz7��:���N۳�^b����>�����fTĘ�>V���h.r�s���q��\J�x.W�+\�r��������^���^�;���bn�1�T�t�:��/ӱ����H��<�j��
���ogH�hcb���|{��C��31��� b���Dx+�2�¦gem94�ͬ �S~�&��?�L{8lN��y��ZE���TP�q�f[|a�K����9����5�Y*��
͟a?UC�hV�K?e�oR)��33��- ��xRǃ��Z��⓯�mW��{x�?��<H��C�uT��I��~5��T�w�XX��@yzZ�;)LI���4�k���7�Z� �G�c�Ϊ�����Bwٗ��4Y�(�����89�+�z�`^�V��ǧ68	?w�;鈍-�/�c���4lqt�t-n�zq�Ɓ�D�ؗ�/ɤ�}G��� ��I����y�^�T�Ωc�<j�:�}�k�7���y��7�$Q�x�@e�V�V����؞/��"�Z*k��`�P�M�Đ��sM�@j߶&�o��{����,&�h+���P`�<ؓ���Uӈ�u��h ]��Q\���#WO��R�p��P$ڹ��<Ai�@͎&�s]��U�m�ַ��0e='�G5��Ԗ2Y��i��~�z�=0��B�-Å�����]Υ�L|�5
4P�I� �rDo%����D��Q����#qI�|+9���i�����V�.b��9e�3-��Qn�a�~�(N?�9�Q�	��7�n�x��c��\;���lE�t�зneF�`d��'i��k�������]�v���K�>�^3.����w&KD��ܝ9S���޶�����矔+���Lo8���f�ڳ��`�l��k[���vH�W����O�/�`�P�.U��d�q���P��i�[���e���ú�H������e^I,͛�7f�� ���?5�i��~���*�Y�b�[:��B����%�i�|��e����r�4Β=�:���J*��E�c@�h�_w`9��ss}��u䉿ew�YW7��5刕�VE�AН�T�i�fƤ�ӽ���|8�u�}�u"Tdgb(��%��M�U��pp�27+L�������g8p����f�)@�u��w���i?�1M��fx�Z�%k��-�E�]�:��.�I���5�*�����%P��!x�ń�/�z
�"��'5���7��2��08�I�M�Wz���	mJ��$e�[�'�_na�B��]03����'�h�΄�B�NxV�O�N:��١Ƃ����^F�1f�j������`���5Y�`5�D	ðFEW��!�]��H/�6�l��C��P�>�p��j�rb�䍁g5ב�����kM��{ϐ������н�B����:I0��H�)?$"�ıL6�8s�6�NUxe� u��L��z������=�5E|(�_�������j|��HŽ��;(�C�b���0����q���A�%���ͅcI�4����_0"���\�*r/�6ZiKʶAb�������N,.��*pSxk�(�4�twnY-`����o�;�L�ȉHy����H	R��j��T�d枓S��~���؆���M�ç���l�z�,̱�q��*����r���Z���q/�a+nԍ����X�x׎���@�i�D֦��"��j��N2��{���3׵�k��z��{��{Et1����W��v+�J`\����2�0�Z�|�E���?C��d3��h|a�����ͻ璙���u�| ԇfq§�h�M-ڝ�|[���P���,�+�<�옠�c	 MVL?��I4��z�,{��luV�ȭ�}�Z��&�Y��A�ֹ_P"v^�0����Ek���S����_ȟ�!��p�_�)u��d�J������n�[kSDE���2�4D6i�@����$�|>�m�		)��P'X����O��g��y>_b�e�_��;�EPܔ�S�W�<�L@�*����i-b��r����S,*�p����q��	���/�h��_�G��pi�ݰ��j���`��[��ժ�t�Rґ\�����Ql}v]��� ߽���/����1ç�4����1��E���	G��� Y�^�i�]����ҹ�"�2��=@��<�R ���Y��$�cE�R���R�^h��)����D�lZ��@�	X�#Y�7_3�ح��X�I��v�yk��X.�,�4?(եiR�!��6����ezX�d�c�y��$��8�������NI�=jR�ГM�����8�[Jy��j
�c���*[œ���C���,���B�>駼(� ���pM�^��͑L��7��9���n(����эpӖ�2�:^��QY�@@|�ݩ}�UN�e�D'9�����Nq�c�AGvybko�D'0ֳ��G���­.F� Q=�ѡK� �b4A���=�M� ��'BL��Z���?FvQ�����