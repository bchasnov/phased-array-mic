��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�P�;�{��3�OT����n/\�@���V�F�	G�V��]� z�`t���y[q����a2�QG����c<iU���z:fj?�?��	1פ��s���$ɍ&�oD8-��\����6 *�+�I���LYx��"qJQ #��\}�; ?8m�)����7`���#��'���9��O�y�bs}���횞��bwk���D�|����l�8?����He�Z|���jo�㒝��� B��HO��bE��۔�=���)�k��BW�Nij������%&< 5y�Y��	����τf��K�V�R��}1�L��W�S�ʠ�̰=�UqUc���x�H��{\�ӂ�|������@��~��z5 C�H>
/��-o�G�V]-�K]A"���|�k9�k��Q-�Ǭ����SQ
ݓv&�<
Q��uee���<�+j�۷,,�
+P�:6�	rr��o��k�F�^��\>�gX��Ѓs�Z�c����|�'�</�q�������^�t�����.$6U踙�t�N�րS��l�����q�d�@�����D��|�ɇw���
,W7f�k�@��g�)f��������?cad��| x���mlރ���Z����,�߾���@˔G �pK���^#�0T0|�|�����UlXr�\�����&�@�Gjz<�"��\npб�;i�oʱ���C�y�LA��8�%��?[��t�� ׈]d8߅ŋ���:���Y��u�bԂGS��,z/�T'�#��bx��S0vm�q}vV��x�S��?�Ӗ�N��9�a��a��X��i�j@�k��>vMAe�զ�v�PZcc�p�����tH�Zs��D��K>�U�O���}�+��9C�;���c�I��b�Y+�w�%u��F��Z*�;&J�}�f����{�Y�EZǦx��49�I����+à��Q;��qG���v8;d���p�$��@`f���%�)�یL� ���^�U���5: N$�q�����H?q��Iq݄�k:+<v���n��*$3���b3u  1�z����,{z��D�~:���b�."5E��w �$Eȋr|`ȇ�BbV���Á�q�����'����aI� �e���;�U�%3ʤ\3���:�FN���n˫-��c�&�^$�ƅ��3J.|f�Hl��}:]�*�X3��@=K�����n��6=�|uԍ�G:k� 3J⿣�r�C��W�g�6�� �_�;H��HF+M�5���R@�dh�#<@����B���o����6�����0V��Y'JU��H���l%}����@��xΤ�S7 �#�E�!����P�ޫ�f��Ğ�����P��0�d�3�51{Y#����E{^��S�Ej��wIj҇�6��)�ڄ�p�#�HF�8ә
�5�.���M�}���9�z��Z����b�U��i��+1�C�K�i�����&��p��p�8,-1���M�b\�Z�1�R���I�6�W��A-����wM(o�&#,c�G�k+�z��b"�H�@��&������؃z�N
7��I�(�-��1e���n�6�~�!��!P"�w��N�� $CH�a�� ���zK�Kʩ�����rve2��:M��ݼ�%����bWu�uN�ك�]K����:�Mu�킪$����F5�$7�a�81�g���H�c����(����q�qgM,#�do�>�ٱ�
УW�R\cڨ ��Mo�=�Na�}3��V�8�NaJ>>7z[����^+[,oUj��W�E���Ş���]�5��C��J�=j�FO.&�L9�'�ϴ���g\�sކ���C��-Z�������6��ɒM�{�å�ݱ�^�4[��n,s����̸���1�NVܕ�wn�,�_nɤ�(2, ��dp�<� �9���C.j���]�q_���zAgć�k�5�L��m��6��+�Q��*{Y�v���}4d�($���d��G����tJNX�W������oW4�����Z�maA�v��όs���d��m��:�Ư1���h���x�+k��g���
Ƴ�=�q;�_�/��I{�7���{�n7��
��4�c��."�M����hWC�����<OFԫL��Wl�`oa���h�hؼ�w�gGS���H��0^S�9 ����Ċ�~\t]¿���Y<
�]%-�G��i���4[����c��R�a�4h-1�=;Y�@�ܝ$���s���aB��?A� ݽ~�t潸GA�<خ������cs�T�l����h7���$`'��%��kx7p�&�����y�2c�-��`������(y��=e�X�x�P)
j
�Cu i���~�:^�Z���Ä;�a�P��|���_C`2#��|Éi:+�BKP&#��G_��F�����BV�u.	�>r����"jk���UHg�Y�8S��v벶MS�4�Zqfѽ~��S�Ӕ�Z���ZT������$ X}A)4c����"OY�����������|�"������3��j���[0o��32�5.���'�79nq��i��}�dzVA��f�H��F����u���s�g���˴�s������4bڏێ���A���ܟ�;�&U�ZapZ���hnC���c�	��6.��3�����R�J"D���ʔ{���@._�|�<��r�-�=YK:�2��K�k���A=�oy/�j�_���h�8�|`�Y[�\����%O�FN�}���߁�<��j���/���=�1��A�W@<�����#���������^�e�g��ԙ�08��F�4�����\�`��>�۩�����(DvA_�r�!L湫�N�����B7�d���	{r�i\~��ܛ���"m�t�Q�!���v�LǮ� ����U��+�K��7���?���ߍC�uE���l�^�ŷ"�A��{a�\dAûZI�L�b9*���j�$���ȹ�m�sч�R0���33m��/8�6<P�Π&th��M�3�ᄴ��Ie%C��HD	 ^C�����-��n7��#�4�I����˹������`��?!V�����������f4�1b��*}ZZ�>�������t�P08�	�%������f�ή���ti���qm��x��r+*�tS�W��G�ow�Չ�3c�K�[�+�ο�N�`$3�X����ݳ6T}#Ͼl>�e��ӳi��6�S8��}� �p��!Y�)O�v�9��.�.��CY$��j"-�<���KW5	Y˔<���}3������ޛ��7�����Xlr�e�D��eo2Ҝc�2*����+����ߡϼ�#��T��opPβx긣2R���G��h�]@�&�s���I%�`��h:E�����=��5qFTF,�[��V����lea:}xg;�?�@�'ٖ��Ǝ�5J!0��+���8����R��g�]��P���g��ڗ ο��rJ�AF?��<�^��}|8��^��#�.`�lZ2�U'��E4#$�P&�4_l�9�J�m�X�4h��Z�ak�a4c/�R7����۔�����ذJ!i ��|v��uu:b�!޵"�¢C���Vs��U��L�HF�g��a8�W��^y̚������{wtP�i���//�T���cApWhL�L}۶�T�g<�\ �k�f�-�s� �iZ�kKiMB��@������*����5%?�~<,o�ӓ#.-�����Ў_��.>@�ͨV�?�Qm	��m`J��sڥH�%o_3�QAE���#��]4�
�0���oy��e�L����m걭cS�b w�
X�[�}�H�){š֔���s�-}�.j ���u,L�E�A����ջ�\��Nby�F"�o\�<�dd��R�4���E���f�`]1'N��BVm�65�I��>���}��)C?�>�l����h��A �3�����.�����Ӏ׳�f��)��+Ð4
����N�)O%��<am���9�5� �:�!+sOZr�Nq���>8D�fx#4�Z)�kK#7�ޢy�4� ���}��7p��OkG�3�Ҫ��v�r��1�ј��h��4���P��;ݑmӤLC��8�_�~��r��!6!(+aK�Oҙ"ͳ�l�t��� gs�pbZ�䮞
j~׷��Jv��|}���HO>����T�^#���r�\whq��PF/ �������9���-�Qo׈�_���_Dx4����?�g���Wgʝ2r�թ��,>����	S�F�X>����2����e}W����U��q�)�����Z����*�Q����b^8��dw�W����a~� )���hf�2h7m�biH�t�礈�A%�e���>�bsZ��Ȥ4�ft�3����A�J�&jL48��[��ʚ����k>��2J�q�e$�������˹�G�D&�Tׂ�/G�#Kh)\���b��E���eS(c�I�t�~׼��Q�jS�)8�=]��,7��7yl%�fv���S�[-����J��Ⳙ�s�_ȅ�H���)�1��
f����j����U�)�F����V�E9���35)�����FL����7N�|v1�@�8�5�dM���_u�/�=R,5S�E�\�<��?�P�-�0
�]{:y�o)s�PM�T%�@r�G��ەt{�Ϝ�O���Q�n{�GX�˿�,��N�~HO��	���9����i�M���H�U��hF��S��ƩC���\�U�ʒW��=������[����F�TI���j*����7y��B|(*Y2<NL��"|dr�%��s��)���!u)����<��&�'�E��uN\�{E��Cº-���D�H��P�K�������A~��W7���,�p�����7m���y+�"�<�Q����d4[��	��#ۦΑ�{�ī�:[1x�Aa���M(o����ad�C} 
�?w#Q�{���W^���\Z4J��{>���Ό2�c���4M�$��7����	Z���d�<���7H�}5]�v�h6�Cx�Uә�2.�M�Yp�@��Gnn�����]�J˶\\G���oF~l�����/��-�LF�)C�+w(P .<s\>�ݨϵ��ͫ��Ԟn��b%�����i�2��FB:�$4��(X����*>���t���P�2%5ĉ��7�(pdF��'Ё�	=zңVT;=��<u�ۥW����'T���L�#�a�.MC��|s�aֹ��A����vQ��ډ�]��R@���Guen��_a�˶꣘��}��a�H%�~�g����z���3���s������72��2�e��Ç�zp|\]1��E+*��7��Yq o�jIÏFou0l ����Sﴭ ���fEw�Ki������
�w/�px�q?飃��Ì�o�h�����C�fN.�U�+���Z�j��`���&��	�O�ga/O�ߡ�Рwܮ�NΝ�|��>}d�f%�ر��o�K�wD&��|ƫpԠ3��ݒ�����J������i��6:{����g�� �(��Ć�a��p�L4c@��2����	���kB�ac�V8:k���Fs/
�X��"pK:���˷	ޔ7�,)@'�a�K5� ���9	�+.#��2�:��׭�zy��G�KXL���ީE9h�T���|��B,�AJ;iu|��J��#�����Wy�ڣ�d��Q�t�\��#Z����q=�A�90�i6��^���Ԏ�$��3�Oj�밽}���xyR���)�)}]�;}~�n���ܼ�\i���'��V<�Q�%��>���^#e=m�ʋ�W=G�����DEy �%/o����˲po�}�Q(�#�:FUxh���5/%H���dd&M�kL��S�JW��M�<9��6N�۔��/����JY�m�_�y`�`�X�<%Y
j�:��o����m�^nX
���q�W��ۧ�҃��m���n��\�$�d���d�X9���p�F�y���1A�Jx���1���ӯ4�ѩiݺ��e�Y��@Y��M���]x m��ӓ�g�u'L�
׏�nLYt^
���0f�ڍ�
!�u��_U�Z]!��Ґ_���Cڜ�G3�L�5v�АCY@���p�S�jW���*�-ᄖ
���cݨ�>;�^�|����[[y����w�$G�0��n>��ԘL�#� �ϫ��@�X�ױ��1܂!a	�7'�ȕh���9IA�������i�`/�&�DQ�e��W��H��䮁Zlњl�����b�2��hL�.�&��
�>�m����҄-p�}���vzMؑf$$d˯[MY���/�03!՜�����Y��O�"M���(��#�������-, ��R��c/�x�a�#�j �Q�2�{��6�� ע�x�N�%9�2�H�DAΛ�F�w��:x%cA��mtm2NU2��Ҋ���ݪ�&}�5�bqd�c	�Yx�is AA	�ՋI��oi�w�
q�X-��?ݗ$g"�5E�#ɶ�P���v��t�J�BE�pI��[�<��$�e��&_: �t�4x%hDFѴ�����N���̡��(�m��7  Wq>�����p	���4 u������]��\���A/�q�j���#!�+�Ix�)G ��K]�v�h����|����i��}ѱm��O�1K�I(v���_wyNO?et<�Oat���F��X������^�FMt�se"�mi��fK+�ǝ�N/�	��ٴ���	1�y������4jc&��s951�Lu�Kѩ +�J�a��jV�?�;<��K�A�1�4!+ɏ!�.!��f�,Ƨ�{�����)����B��~&�<�����M�0��. ��T��1���ڞ�4�Jβ�9�Yy�c@�r�'_���Ӿ�Zf���z5[]���;�n�my`g JN�lΑ����f�
bKK��N�D0z�7.gW�m�)#Q�>�ܦ�`���ҩ� �����<R<o Y2x�f��3q��g9�s↽�F�	 �u�!0�oϊ�V�ю�����}/>���( �:�}]�`4��`��e��_���7�hk�����o�hT2SB-��#O�j��e�Q$}n�j��h ��Z�͋����$�v���vRUf��Z������g���1�rq�ӱ9�}�v.w�$�J$��K�ի�9r�h]�B{3���xnI%�iXŕ��Z���s��
��9��Uy��-Ie!ь�.�_n!�,{��
����G)r�-���J�D�fX*_�.�/��}S�oϯĊ��t�Q���"���TiN&7H��w~g��o	�D
����i�z@�����;r�a�^��5�b���p�]c�+Y� �pU��J�1Q�z(k��U��A��"(�:�S�J�o\��,�.�a��K,��@�Bt���䋡R�����c�~?~�sϬ�Y%��c`�#D/�,'��o7�	�W�2��e��HU��B{'B<U��'�� X<WN��&��U=�6�5;��I[.��O�b���"D�~����"�c[0���B$�Wv	T�� �RqŪa�܊���Le�Z�6��C4�8�t
�fj��t�{wk�M-T �H��j�(l#l�A�ƗK|$>_������'c��������	J-�z+�1lE[
�pfH+
�AR�2VFb�D� N���><��ۮX�4���(l��^�HǦ(Ê�+��'L�̦�掌�n��$n��f�E"P� s�:�5T��_[#|OE���(O��>�g�e�,���V��RU)�tGmL��7g���O0#9x-"���fw[�<T�?�P������%��9�t��=��:�X̲6,h=�#y+*7V>8|BlB"u��O���_;�$�iGA2h�e1���2�0�d�J�c�q�8�JtK),z��v��0��%l-�:v4Y���id����؃�X������
�hd�Бu�˱E�`O��wj���\o�0lnuu,7,V�Fma�+6��0�uA4D���!FH�g�{����%�(�nf��������:鯮�4
!�/D(�
K���w	���[�!�xK�>�_*����PxGf�ɔQ�8�YQOi1B(�γ��6�8�M���Z�5E|S$�c� �
��Np�cյ��#:�*SN�7��J	��<MZ>�n�!�y��H�J�7.��(�W��%�E�8�$n5WÕ��Mx��Ma��i�v�M�ls�
�쟢[���P��)k�W\y�һ��֏!X���Պn�$�cmu�)�E	
�ȝaÆlɲ�V=+��,�<������J���nܝ��?��<"
bbJQ���dW��c������4Tako��BoG,tĉ6`"�w���ƅ�=]Ί�Ȫ����Mĝ�Y����[��ϊz�W6%4I�
1��ZE2X[�<�%����aaD��񪫭{KB)���^y8��}>�f��s��E
| C��R#$j�'m��N_:tox��ƕ@
��AصZ�N�}�����[�P�n���^��m����N���0K��[�9�L�)�͈�F�U�3�D�#�o�-�I^�o����1�ђ{��Ǔ�ߕ����kv�8-ך�>��Quq��M��lb����K�I�AUHh;s,������"#�@%�:.�N�����X�7�yS=�2�.��˓���p!����ҙx�y�g!	�3Pj;�Q)��I������ Y�p<�}{暆A��oś���<����z��P�07�����5	�(���jm����q� O�:(�|��0\d�w3:�z���a>��˻Y�ێ;;:��v9�c���&��Pǽl�:��T�k���ձ���`�	�ܬ��P������{�$z1���͗(�7g��i uՎ�o]�����rW�s1�ѼW�u��=�$
��)�]��Ң��wx���k�C3�v*������$����}�h�:�KJn�qh�±��m�/����Re��K�]�/�*�����Π��02���Q����e�ę�b��V�#�}ctTU�c*0�"�Ӎ"�+���T-Ua�r�e#���5Z��פP�	�[��c����$��iQ�����|@[ ~���5��w��L�]�����# ��Î0G�>Fe����sRl-<8`����zM�=hHq�!T�k]N��^+�-�����4���_>s��}�=f��z������n����K8Jd}"
�aN@��ӧksn�p^��x��&���RS�C^\j���4�W��,x�q�ˏ/�fӪ��T�R����_z�$�4I����j&Z�|���	Skoq).��M@���U� D�5r���t(v ��͘���|Ɓ�����B�>$!�� �qR�tO�$�g�C@���B���O�mT%U�ԧM���O@�wc.&U�ÿ�k�D}�A��m����̖����9roA��!~��%r�]��jJ;�����(^n��$`��ߓ)�0�_�17�'_����uߎ�?/#�w�;ϘE���)�x�'�>g>7�����ex���Oz�NS`�Tp�x��J �݁�@���^p�f[���u�ri�Z�����{.v����!9+|�|-�7#Ӷ�?*Q�|��k���Fش`�;���S��v=�������M/��Tbg,�a�(�K�V���������L	i�Y>$+v��X
���q�3�����Z�yze'�\Iaٱ�/�s=�Y�j�YTm����:�TG���ϫL	�x�n��@wp����)��ǲ����{t�}ua|Uk��W1���b�2ڣ�=�$*WC�"=+u������:��쐱��А?��py3���0۞�9g�����Xa����S'TL��V���g�.�{�����Li�U�����e�u/'�4�M9��R�)�\ԭR�?��-K4��Ta�s~��i��#j`Z2S��j�a�A6��q	��]M�kc��CP�����S�TA^{���~�G�=��ز��$6ْ��٫�^���0�&51B ������ǚunT�_h+�.�fҞ�@Z��ȅ6֙�޼J���rV����^�˝�#%
bc4>2?4w�ؙ�I~ˢ ���|�8<��C���N�)m�`� ћ�=Ga|Q�bkry0��p�7�b��-��Z��;���H�����xФ�A�Y�f����|v�P�J�a�����>Q�^�I$��o��bhr�������1yQa�P��>�k�������^@�u	��DI�=�P�L� ��K"��}�x���8�/l;��ҳVh��d�{�{��	z�.o�5���MrƉ�\Z�3qZ�=|�n��E�����h��JƐ�gQKr�ŧ��ӛ���1+Ƥ�H��.��uWsb�Z&9���Х>���e*gq�=?���+�Es<���x�e�u���M��*����&]jP�4��T��2i�Γ�RA�C��E�(�	�����#Z�%�)�5�������FB��?�w$�3=l�p�s�$<���<Ҽ*":R��|�d_?1c�����jB
q�ګ��9���	�O�^`��1+��[���s ��Z暠ܦ2����2<a�y�Q������f��Lm���eyt� 3�'���X/��2ޜ�7� �93�`�U�!��.\��� nm^H�� D�ؤ`&�����ۧy7O��;Ɔ΂�/�s�7~�sm���9����b�|�p�E�t����?u������J��Dc�+"�6%�g�|;K���LF��.dvE�8�wk���uP^�t���+��9��/;(Bt��9l&I�� o|X~?goO��V	��S|\����������/?�Lɪ�R����_�T��%�}>�X"G�U(ݬvY�6�{���u�P>BD>�mh�C7#��s>�W�(�� ����<��0������'��^D,��x���,GX�tK��xAH_X7����ٮ�l�N��Ir�c��������;��eEZW�bq|Ͳ�kΦɱP��H�2���Q��ϕ��<!=U(���m�=�#�GD�!gA�m�)	�"O�E�UpIG�X��9�r�,N��(˟�������MW�l�zPu���ȩ�uL*n�ʴ��9��\��N���Z���X��n674��~[�5��#����
��b�F�{$�Q0����z�1�Y��X���c�j�0:d��c�܏&fpw�P,	�8�Zi׃�ܛK'-8IGۨA=>ab@z��T�h(���&@Xk�B
���݃�2Tb���|@�;i��D jH;�[A��p��h{l��G0��������ovLA>��J����{�%k��>g��r �<_pl5�T0�)��.�~|}�bڶ�o���Ƃ�0xj�8 Sݔx�t��CGj�m%ea��i����pu+=-`FC$.�g��}!��l	"rպVm��V�Y\�����ҍ���$�
�n�D��z�(��HA��u��E�8�=���T�i�Q�5m^����L	wj-���h�m����)�5�H�I6	��sг���m����}��?�Ǩ���{�9��s}+���j��%C�
�ҠHe+�z7���A9�Dò�):Z�0��
Qw��U\sc G�l�}Ym�آ��mpD�uC�Y��ý�`�v����N���W�b��o��}Ed:ϫ�	�R!4�v�	)����PÆ�_��Pj��H6����t�+�,7���#�\��2(�~�mV}�}���I��F�{7��>��^o~�ɛ�D�Jp24w�f����"D���h��rX���*�[�P����L;H&{^�Qi��,<e�>�APJ�$B��Y�6r�e�(��i��a �1�Pe��x���=p��M˿��

Чd�
������wa��k��bAv�R��;���������;�;���?'ͻjE��ѱ�?b�K�� �MhJ��mQ�׬_��;�����6d�YA�^�;�q���$Ŵ��� �DmЎ�7nx����D���ܰ<gk�skc����� ���U�E;�~��,�o��~����{up�&�`gY���tqQ� �s�ȝg#�$u-F�y?�)}�klVi��	��=��Q]�&)���W��d��Ԇ@;"T��At���|V5�WUd�ǲ�I	�%�0�q!}�+LXZ5�@�Ew�:�3حU	c|�ʫX5�J�[�lz\�m'#Gs*�*|ϱV~��1{dI@�'�Xʅf(��橖��ˏ*cn�A�#fn����,�S��:z8�ĉj�-��L�~3AS��rx��s�W󋨩�胟��&��{%�!��Ƥ����B�\�|����Y:�J� ���/1*���4Fͳ,<8�9*U?F�W$=�̉�[�|�'�Q��]����j�m�����m+F,�P��R券�1�����0{J����>� Tq�Y�z��k蕈��@�![g�K��fkƛʂ3����>���?{��{�
2l��i�������Q1
�O��wԓ[�JoЮ%#Y�8���f�2p?]��)�n+d�Ε9�>��l���_`����L�o��0O�u�g�& �gI���p����I�� �Jq�_�	`8�qO�00��n��^�"��\x0��7 麩�|�����e�
���Xa��$����Q����@�C�9n�َ2���X�踈�	�v��ӽ۱��5ʑ�ҋ�;���b�6C]2bud�F��	g�0p8>ha%�3=�ȏE�g�&���8��.���,�K���0%���)|8Vlp-D� ]l|�����L���6�m�Hҥ6�׹�	�%{����b���"࠾��'�����Qs�?'�@c�E�!��������R�P�ce*��X��6�l,��2Yn��j $b���'eDE��-?M�~�ԧz��2��	.X4пu	كD;YF$�*�sM M*-3��
��)8���{��*P��N.��q־ |�@h��Y�;asQ�R��nCObcG��mA+
d[6G�H�f�Fo�|�`uE7�����خ8�0I2��C7"sD|Uof�nx#`J)A��:�y��<S��'>��
1�0�B0K��N��_G�Mφ�i=�r��� A�sA*�����hD�o����!��I�Y٩�X���֮"��~!���Lh]�ӷ>\���p����uAˉ�9�}��dq��cr"��V�y�ݮ�
�W�$�(R��s�.�K���	�@��G�p����E`�Jx�I��C�����i^F,ښO䯱m_AP��9\���ZLqH�b�����t�T���_Mɰ��_Ty�)�NS� �9G�3���h ��}�ǆ%��bN��b XA�/d��^��ɹ��������Ñպ���lʛ���k���B
u,�#Wٝ��D�al� �!���iPW�%�!���i�����2McgF�'B�&l_��~f,���2�}R�^"���z�U���1k�$�3"K��_H�]S�4<i�;ɐ�s�)�=�����)U%(�!��/�&�k@5�'�][&	�b@{XfU^�f�.Aj���&�#Òl ��w��;�W���*�L�	n���ۆw�r�,B�F�G�n��d�K3�.x��>��檴	ø+,](���ɔP	-�4m<�t�W�����H�|���I�c��t�c�Su,�L���(��mc�ѹ'����ꘝ�~F��рn���TO��0Y��v�ʷ�z�CaY����f#�Ia51lM�mY���@i���i��c{��,g䖡~��%Ξ�|�^3�U����!��?�N����G�^z�>`��2'�/�M3l�X���-�����;P7�3��_5� Q��T�>ކ�U���Y5IY���s��H������	���OU]��8Va6���LL��0��$���bHp��
���HV�t�J5��P��o<�[~%2	��"�LM���v4������*olQXݖU�ᤥ�4JE@�� @9���]�I�ǝ6�%�	��/8�v�	ZW���7Ed��0���b{؏y�Y!��)4��U�8�ڴ��	i�����Ǔ�:����j2<$�h��F�ny�Ѥ)�(���'��9��cܴ�1��7��V��n���p��D�KT�tn	/x�;5��7Ȁ>�_��r���K��۱���������B4��k�A/���7����rY���˞�}��ۏa�(�L�a�C/����5KV�N�E�$h!�	�L,L�����ap����&����C��>��139�X$}�ȳ��M�s��D�5j���b�?����oJ�~7.�N���|X����Q|j(']�hL��	�Z����&�q����s�`z�g(�0�y���
�Mz������*goNC˺�2u����>,7و�=���'U�f�$ �q '	HE����J.ѳ���Q���4��z����H�����dF����&ӵ�����z;$�
����op��0�p���jkt\A螲�"�9S+H�r�t�<��p�"���k? ��x�Q^ `���C�*(�u�/-�n�e�掿ɫmR�5�O��mn2@ӛ���w���~�,�JLv] a�߮�a�{ys�6k!f��2&�>��sh�����/;^��������X����!�Zd��v�k�c���d:q.u���]��=.�����^��(��*Dg����K�biǕ��A�1,6�p�l��;w�b�cy,�ZQ8����ʏ�V� � Y������h:ŗ����L^Ro�E�o�E�V�T�8S��oXu��V��p�\��Ę��JW��ڧ���9�:j�L1�@�
��Ţ���lI\^�9ҥ�\�V�N�O0����:H.R�m�����{_="t���@��t�c�)c��V��
S�h.kd����pC4�^�G�����5q$�M��k�U ����ҝ#��"���S�s���^�ᅸ� gg��վ:p��&�/Μ������<�?YБ��Vt�NN�e*p�"˩�x��_َ���r�̉;���+��]s���Hk�����n�%g���S)�ܿ6.�6���|��5�Ŝ�� ���-x�}�߃��Fr)������V�YWT�Xv"��qO#�!��r�M�Y��\����4Ǘ�&���"��3���%��6�A#{��AAֹV��|�Mi0f���(��u#[߮qzr�m\Dw�{S�)�Y���gW�m.��1o7� �t��P���b=��R���;Yb�!ԡem�)k���� �bf��+QT�	̟:��&�o�0:�Oބ@Ҁ��Rx���a�8��m�¹79�)C)S9PJ4�Z�&�ථGzCԾ�k�����,����3m�Q%+���OZ�p����"��(�����<��d	�S2���QY3�\D_���[�C��FU� ��E����M'�l:��X�i
�;��FZ�^f��Z���yw�le���T�	��d6�r	��=`~����)��wN�!|�]�=L��2M��	w&:��C|�����p&RBU����2V�d����~��8֩y�ت�1f����=a��TV���X��f���Wg�m���$y�O����l�J�BL���h=�Cm�gLN6�*b��Y�?VB�^͡�("��O[1f�X裕��V�B���MWhY�'1��bJ�V�V���s��-^��BPЏ\�����,�*�����ٲ�e�A��@�Dؓ���囕PW��"����w��EJ�I�^�5 BOc#&��,Wn�s�Ģ`|����d�)J(�%ίӬ��R���C)���&ڡ��{�s(��� D,(֞�5_�6D��'�e�j��;��S6ͩ�w�]b�@�'�dJ31�̢x�o_�<�Cm�\-ǔNWo�_U�Qn�Z�Q�����x](�t�ː�⯳0����Z��e��V�����v�N����N�ܓ^GC����%2R�x�IG�7	�)�\ ��9����N_���%ޮz1[/1��J�A�?�Y���wm(���.��Ϛ�i�0a��s�p�M\���#MH뚽�X����{'�����"���O�2���9Z���z*_��cҚ@�Q��n���2��$��M��Eq��!`NZ�sFU����%J��&P����V�Ż��nh聀"�8#N.ʮ�8�H�-����b� <�%�qM���-�k��LQ��e�����^!U�N�F�g�,p�[��^=��%�L�N�uK )L�XV�y��>7�X/h�i��
=	tŖa
���3��K��*�7u<�j�E�ūf�/Y��R���,g��r�a�$9:b�Fm�5�؛©��aC��|�i��VF�'Rp�L&�@5��4y����9��EA���!Ģ�I/��>�F2X�Vg�OE|Z�HA��5�8:.�Ł�pm6e|\������.�R�I��������p;�\Vw�m��?]���a~�7[3<S祻v�GG������{��0:,�f��-m8Xob6B��P�39����C������v)o9�f��Ast�Wљ; ��h��(kyU��X �egX!p:�r��[�O2����;щ~��zX��W1M�� �y�/�2M\4�@�8 ��~m�-�����57+i�����Hs2�!�0����CH�	�}W���h|��`P��L�� F�!���k�8;VE���o�=Y�VpܘI_REW������B��a2�%+��(x��u���6K�U�GI6�G-m���6��\��^9���̗��®d�ش��ao��e!�n34��}�U
��-��2�ܝ٤u�H�nܳJX�+��[�+��B|O(��(�|s3��#�w����\]*;d�<E��>'
m�������hP�P߆9o��ܲ�5h ���7�Iԗ��(�z�/�+�ޥH��Ny�_ԯ�[Ho��Dk�!�f�>�_��4Y���=�.�]�qg�0��0??�����[� -1,������WS3���.�$a����:��i%�sL��MKw���ںk�7���p`]Ѣ�qj�6�G!˛�1:s��YQU�/2�h�G�5��/����n���ǜ�nd��ޚ`���*�\����Q�<�[��&��٨�eƸ���PZ��?߶����G�LC�p�E�9�s�����o�Lhr�61!��E�]���B;-M��iO���g��>L��� �g�*�ԯI��Mm�d�l	D��O�f�=�����*!BъEt�F�����������\r�/�CW׺��QL'K*��"��I��p[��HcA��������I����|��	�`��.2�jL���d��H�Y]��Ӽ I���_p�^�c3Q�z��%��L�����?|�bX�g�`s4f
))#���EQ%�$�BM9|a���Po>��1&�z�`��	앓)�rgl���6֮�����0+�IE
�㕻L�zB`�^|��s�n�����s_��4�1Zu����Qp�z����$���ĩ ��M���k|��A�0\�V�-�c�o8�������qY�:&e1��M�$	G	$���$�k-�h���/r�����@�<A�Օ�)��	+#؉���<m�2�H`���5睬1�w)��{�L�"JB`�ڏ��Kz2&D�̽��47�4��_s�Cx�/�S9#�V1gk�Ћh�9���Z��6��ceGp�jP��ZD�Wr�zv|l�'��$yF�YTβ��{�\��Y��N׼��m�W�K�A}��o[Z��X�Ϭj)%p�~��y`�uzZ�q� ���hz�2���}��+̶�0iŅz;0S�p�u�n�����S��xQ*|��n.�^���̣~O@���{ ��/�1*��E^+�Z��!s`�o2e�W}���YD��ˤ��J%�z�^�C2y�8ٺ����[<����ն֣ͮ�W�Ԓ�"o�^�B�?��	S+}t����X.��^xjE����,l�쿨���+�x�IW�޾5L���>ɣb�U�b��bF�w,��U��or�� �
�m����n�y����%��UΞ���a�\^T���@&�X��dx�i�8�VX�2���\��ѫ��c��uC�׾M���,�j�6��h������6"�M��R2�S\C�R���\�4gӰ��%��FY�N�(ɸ�&&s�B�{�U\#">�Z¶vc�$,? 3�����ĨߒKy�
�'�f+��A
�� (ڨ��Ȣ�9Ɇ�"�C���t-�G�,V"�_�=�\pSbM�/�V�2'��)_neoq�Q�V����u�3"C=���y��z��BA:E}�Ώh�w���������x���7�I�� �w��,R7��p����
�����Tk�Q�0c5>�,�%?��I%r�j�Q������};�GW�t��"3
m�*�轷_Dv(�ؚ�v߽<�@��NR��������5JN9�#��A���pNA�PU9%ؤ��@~�����4AZ�b��^�as���u�	��j 8Y��Ǧ�g��j7�H���J�DL��3���������L�|k�)��(���L�d4,��(�<�_Ф�B��"��`1.Hrze����$P��&-c����|u������=�9uJ�� AL[���2ceɁ@f5����v�hFs�����UM W��%�ף�Y_y3���m�ڡ0?n`TDO��⸌*���1V�QG����چm��Gײ�`��������s���u��[�i��I���Ox�/�G �����~s�Is�QHݴ=�*5�����y�`��zO� ��(�����ݒ��a��{0J4@�@E���ƨF�ʘ�}�B^���`O?��a��2�:��PmP�4[�i��f��:�	��5�ٷ�=tAp�m/`_1�;�n�l���0Q��8�*�F�?JƁhJ+Bpeq�+O��<ӗr��6�K��>����`B���K4?��#N�>�PKu^���ݸK��ɉz� �Y�n�y9���=t�=.z���Q��S�E��P�Y&���.��b�Z`��j�Յ�7wq�A������*�F�?kp�/2_���.g����R��7~��No�w��2�?�tuU��A>5����v���T�ݴ����Ӷ.�!���և��7��N�Cyk	��ծ�W��&�� ���`� @ie��0;��9&�w�(E>�e�DC�t}��bɵ��b����$� {�&R��^:\'� q{�D��'>61a�ojUh���b�k�g����ԟ^[lѳ�#���H�7��"����x?/����Z��Œm��Y��)�0t�}� zD^@���"|�����_$��������Ѣ�G!��cw�z���Z)aǆ"�q�|�}v	�$�D�:7�X�h��ʒ�ɮ����|3�wD.a;���57�^$H��G�(�I����ת��X�X�]](�?���Y�ؒ�<1.:Ww^�RM˫%_퉊f?�P�M齉��f�/�hgk;*��m�I_���#s��m!�2��-�p��i�)�vX��hf�R���<�G2"�:�79���;�h#3�A��yBm2u�qߍw}���T���d.X-����11�1��pm/� ����M�'2�2�f��|D{
EUd��Rڃ�6��nk���!��Ҳ����P�w_���bU1�G���vu�/���91�mհ2K2@�/A�A�|:A�D��n *�U}A��Fb�m��Ri�
�R��v��_�s&(�`�f���M�:\��~��Gj�&�z\�
����a*��H�8:ӈd�6 8Ʀ��
���[�OW{