��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1���e}ʲ��cg�t�ϙ�a�:�KR�%���ݧw���ȼ�cD�|d�4W�@�1 к�?��L/,��7�/�Eh������##?^�����QKA�f��Mʖ��3fK��ْ7��P�\�����،F���v�w!�#V�mXM���*��S�6gW�I���Ȍ��Wr�*�I�m5��iR ѡ76��K5߲D�x�'��^�:�Qo�o~G�]//�a(YZ[��V4<K������"(��p�s����cX��IT��>}1��Q&4!ʁei�.��7$}�# x�Pb!��u�0nΨ�ΚJv���q��T�_����ȀQ��޼��ќX��j+ǟ�3�eo�[xj�t֧e��y2��-Rߝ��g��T4Q���s�AT��x�A���4�5�3�F"���R���k��J��cS��B�S�_�Q�����~��Ɍ��D��j�C�$�{��v��m��څ�ب���O�i2�6�l� �P��|9��|��Z��b䆒��n'�!��+�Q�����+<����MBG��Z�x�{͒��a6�Z�P��	R����Y�}w�^�D���N^�K���=��f��gF�uĒ}���ұ�J
%���Tqs\b��X�`��X�O�S�޹�*#	���G�ڑf�8����wV=-��52|��Y�~T�|2I�iߠg��Џ�MA�{��I��MW�o�.m�e�`fP��5'��W�x`��k|�@����6��Z���MXVS@��j�����x��s��S���'�
cCĭ]���>�n`�b�����1�p�a��<��`ź�)�� ,�2����z�j݁]��Ǫ�̽�A��*���x��T����(G]mV�*qm��iL�����~7a�1�̞L�-f4<͠^޾��k�˓<,\�kH1�����O1�j-�$�.������-'2�K�|��IY!Sj����<R'0�~�Ηg�@g_�V?��T0���x$������^�!aO���� ����pa�R,��.�,��0��M!�#���tp��Y�b4�f�t[$	���ir� ��c�`��w���H����}#�>�I���}���Y"�鲖����ص,�w�.y�C��Cg�
�'���&���D�:2��5@��{��ǀ�*!�E��T�������@.��_��a�e?�{P�G4��Ν_�%�n�ևc!N*����na��M��C����he�������W���/��xi[i�V �?�'L:��uu�� &��8��#�s	�`*<�R�n�H���=$�i4K,*$�״H������P��E��n<�q:����' �������z�-$.�p���/I��?�K�Jn]me�Eg��
F�u����T�~%����>Z�Q�������x�w���at�E8u�R-{���h	��O���2Zgy0�˓ޟ�x�A*�M���R�g$���KpgD�^�6O��-��>h"XO-j`)(����6�ET��i�^p��[�aT�.�'K��z�ʒ�8K����6��i�A��;L� [�B�~N2tT��#����H>P�uMF��e�%|/��nfqҌjZ�[[h�/m((_fڋ��!$���֠�s
��y��R.������ ��W~�0h�sZ��{�0ˋuA�e`�"����y��F8��D�a�;�)-�a 1�%�t6��:��o+6P�����n�9��B
��4O��Ay��[�������2ק��X���X\��K�!�P��8���;�Ǳ_eD�󀍋�5ѦW�0`�J5�<O:R��4�ޭ���3v�tk�U@^>�h�\�~�@�%g��<2��"t�vJm�����(���-P��/�f5�Gf���op��l}jA'����|�t�@!Ї��E�.!����Sw��|�`���0Ċ�\Y�뀄�xx
-�8�)0^��\�xq���a��Euh~��"ʗ
�Q?���ũо�]=��wԑ�v���޴S��~˩4/4�[�M�L��k����s���glD�X�ۙG`a�.̑�@&ҴrQZ��h��g��.},����"�&e�k�\��zJ��5�����P<�Kr``�C3@�9�%I�>�4��~kP�R=S�:��v�д{$��Ll2lŮ�=�J� ��_�dk�+�(�!L�<�R��J=H�h(��������_9ej��T[�
qMyL�`k��a6F��J�sg	t��'�y#\�U�)��&�P���4'��PQ$�t�:R[�A�H���GF��*�֦n{$�j��l�Ncר��:�vIAEK�#��B��f��cF��o�{��䷲l������z?�K��g|����4���
I�y\S�U�q�HX.�Z
����"G�O�+eQ[�U�i�b<���~��Z�I(�V�)��՝�]r�~�a�Z���\����e!k�!�ͯ��|�d���V#�k����}s��z�����trc���8s��nI�=?����*�[����w�!X�>\S�P�S!ތCp�p�j�����o�b,_?S�j��m��?�ʇ�JP���=I�ܒD�ֵJZ���32`4���� ��vF@�Y�#�e���f�~l�B�[��Yf<^�[?%:�#�������C`�Q���XL]���l�f8ȀT�2Ӽh
�O_?gW�]VT�x�<@���̛aL��;���Z��x��JR*�K��l]sЮ��-3@�HFz�5��Wό��&J����$�%�i�j��G0?}��O�2��BAT�T��0��6W\�R^ �s2Њ�uR���� �u����:�d/(O�@,Ь���K�[ܟ~vs:��'-Z瑙�#�~�����֑�����@D�\n�J�L��Q��h�u��G�(J�QK��lQ_�$�b���ҿ���C�JF�����%⺰e����^7H��� ������e�Wa�Z" �.�!�������1"�,l��R������^]���(T9���v�c1�-v��5*FKJ9�s�	�s��v�}��)]_ =��h�[s)��ɑJc�%�bu~��$�Sn��o"9Y��v (�����S�X(�*<{�^V��
�n�)�xת�y�K�D�Ɗ&2 6�J
��Ĩ��4���P<~MX|�HՎn�J�+#ϫz��L�|��WJ·̲��n��y4�<�,R�
�kTd�a0 ��m�R��@�/iq�rr�:��D�Jظ�I���j��'`��l��y5 ��~�Y�?�.���R�"�)z&'�=�e�J|P��B�3sb�	v��#~$���o�֊��1���3��!��&�������$��[0��o���4�u.�p�DU�79���U;r�Z��
�����4����{R�r�Es��8���ʠ�ʓX������I����S�dYj�"ݬ��~7���)%�t� Tv�h[`EF	v��w��l�����]�s�("9�^-o�8���vC�4K:z.�V/wh&S��s��>6w�x��)��&�ė��#k�����jv�[�:�= �	[g��%eA�]����N/�+���h�a��*�u��j��)�0�U`�Ů}���mmm����ê�f�<8�Q���ܬ9԰nO��g�R�rR3�o�l]g�}�w~��G�u�ȹ���H���>�B�F����߅�5��. 2�Б���bI��{���ڣ��m����mPX\ɯ�������0�5znD�ߋ�yv�>�V��`��P�IJV��_��������}oMB�}������*�1��;�ǚ{����n6��gph��2p�(d�z�C �36��`��~hm~��ۃP'��'��
!x���wz���9O���%Zr���kɠ1a5Q�����{��0�z����PCe�Qk�kό�^�Dd��.�\�g���2��U�$���`��ˈ|���I\a��������W��FrO�;Њ�W��=4�7U�J��Dm�z!=a��f�@�S��ТjN����m�<+�?�Wp�E狆M���_*�W�
�u�$���tI���r�������Q\��ɹ���[�|�3��d��OT������Q^���F�=}l���l�T��ӥc�.|���|3]�*�G�O@9g.��K�ʟ�X���Ym(�������̠�	��_vA�:�Cr(u��E�yK7�;N����q�w��X0��D�>{��iwc��tq
����8Q��g{d�VJ�e���#�������-P_k8?V[�:.�!��?�B���d��.�%K� �T��h��E0 k�O��Y]BwD�1�a��Q�6�c���&>�7��*`�{2J�̃����;_^yT��fY����0�^OW2�F+>�F$g��4�5����kK�`-��p��c��Y��X��Q�*���O͘���.NCAVeA�w�Pa7�F��<�d�P�y�@��\h=N�D�(�N�z�it<�T2����u�>Qբ�YM-M��>����_�9�U!�����9]����iW҇�r�6����٤�O���l���k�����	 b�o���]�%Ѽqf�j�I�Tt*�y�,S�=_�A[D���A}�zAz9��)MSp�w��=��v*ȥdR����K��x���%t��oK��Z:��6�3k0��J�)�B��đ� �����l.�x�67�o�V�P����NMXO͈����ܒ Fa�MTY�X���UT�$��X�TWg:�xV��J"��C���L�#j}���I�?!��s=٪@ÿH1.~���@QG?Co���?k��49���F_���M�������7�����2X�U
�'���u�+�=��R�n�?]�s�!���*�����|m���Alge�����n����������|q��I},(i��äLu��hЋ6��y��e����<	|5g݃ŃO�J��"L�U{": �W\��c�Ј����J͈�>ŬT����H�n�ۦ�[���:&Rz/)�]&�G
���ϭ�M��D-����f��8���BƉ?��C�m��&Y��:Z��\�k��b�c%�����کP�[����� ��TY}1Q���;~��#���,���;�`�s]R��(!wx�?���B���
kw�:c:�A�$�ؘ�������ձ��5����1D9D�#�+�|b|e%�m���/�j�Po:Y�렌��,hM<g�|m5�g��]�Rj'{҆X���uX��Jircϑ��{&�&c�x�9���.���=��n�B*Qh��2��,g�����.94���� &F��aŜ�N<fN���>oY[L�y����zCh�WKq1ɻ��G�o��%ҥ-d��G�ف6��{泊6�t���K24��NK�� �s3}Y5��U�>d�6nNl̥�B�w�A �V��)p�
��]u9ox������9\3&f�Όu��aIE����	8Ĝ��	?�"ѯ�'��It����vͻbP��R�
z���/�$��o^�Pf������9���eәmSfI�9����+:�:�����1%;�m�%Ѯ��8�F~�G�3{��h:��F��4�"����1���.Q�Sw"�I���:�|T(^�Q�4�F=n}��S��Ⱔ(��xW��t��L�Z2�]�U:N��,S^�%6��o#S��@n�,����)�^d{q[-��1ɜb��=>���]]�<ؚR��E�{��=�5�,�XA�?=�[ր�4Xl;CJ�Y����նy�p�+'��sY�.�W��Aiw�AO^���X H�<7d9������1Hr�ϭH�]�g�_ˈf�)-7�������L����0�Hy[D�{U_Ű��wqB构����[)�'w'wɥ7�����v����aK�o���p���|�Q�C�	���g�����e�����\>����K�H�\�w0��Ê�(��N�-�A:�Ҕ�x�����JÑ:ɦ� >�@c*�n8t��ϰM|j�B�fT"1�Ql:Zۨ�k�*���k������W��6"R�� �h�s�Lq��k񥊉19�p�	R&���>\Jz��8@;Å+m�'�o���PJ����hp��[y�n����`h�y�/�鉖�8#h��ޑ��@�3�� ������uW��z��;
��8�J�#��� �k�9�paC��(3���>VMV�_�e����#A��F��+���I�=�Nh��*r;r����版�qؒ�0��?Զ�R"�'���˪��9�J,�c�tm"�������࿑}�1hS���\��Mт۳	���Z�e�O�� ��}���v������%���f�Z�X��s���
&6�GOƐ^�/5�Q � ����}�.����4��ɈClW�P�7w�7�)�:���(�d�&��nc��mK�I)f�T���-�@�I�TO���kHv�÷v���sJ|o��D,٭���?dX�?G��<���j֐��:��\�#�#�D|�g/���皞�KlL��S5���f)k�BÖ��#�Tw�%oT���`���2RrY�Gi��V�԰��{����P�IqQ|�Ĩ)ca�/0���hfm�� +˶C����:��]#��3 �s�ë�)��đ�X-S�c���~�#���m��9.��چ�>��XF���h�k[�8��6G@S�E;a�h)袧�濾&:�z���/\��zæP��������I�k1O �p�l��\�u*���a;x�d4����]c(3�b���־�$ؚn����/�&thθJ�Mu�v,�Yv�u͘12��&V:�
�/(CCw��<�����
6��Y��CI[,�E�����Rr��O��|�u�#η�s����	}}$�c=�.�����cE��5���?@~��&��d�����Vs?? ����Z���I8d��w�F4.���v��I��<���O��f�k����-���k�.Vծ�="�?�+�ˮ�9�W!��T�R�R�r�9nP_m��x����1��qj��$��Pf��t�_,����SeZ?�g2�2���W^��[7�g�׫��_��&�9�r�yyr�2��*���
"^��Uo�:�+۠[���O�R~`-���M)җ]�����'�� ��b���H���bX������_%)���\ghmu�;��<(����E,�����#����͸7������V����O3��ȷ!gf���E�7Ŀ�����@v�<��M.�����Y޳I��LNBC�,�뉘�ߑ;�)�u/�UZw�+�!t���� ���+�/�P^�]	�h\�Q�8���/^f�"��*�o������ٺ<�_ܹ��̏�Byjo���XZAdX��\��x����5����z�n��G��MBi'�ln�U;�s���v�5���ќ��x� k0yvʿ2D�/(�uˣ�	&ͯ,���N=�.�N�1w����Wy@�#��}8�>wjy�n����1���1iŬ�B��^^\&�e6k� �"�~+8N�;C���� S:kN�[��O����W�b��r.i�bɋ���q�V�B���P�JF��r���z��F=���v�������-u\s�\ @(�,�L�#;~>�D�����7lx�t?�<�SR���ݿ�з�ڛ�s�E(���-�,�q�X�_v��,�2ˣ��>�(��v�Z�<��k��@+4P��"�ZO�F�I��$�V鰋^�$cd�Q�X&񪓑t���+��[�aO��,&o߉���؟�{�e�p�r��#���4^�/o����9IlMl	|��.n��'��*ʙPޔ��0n%��уf`�a
��)H��7MKt1Mi���l���h��k�M��`s*�����/�|$&���ȟ�����E��`[��V����a+��Rw���S ��*4ן&�I�%��d����I_����.�����Y�ɶ2mi�+�ÆA�i	i���� �g��[&�l��,�r��IM�JY/���
8�TpK���_Q�������ɸ�G�z,��yD�.J6o*�4�HL��4��p;��Y>�������Lw?{۰���eE��'���H�s���i�QO�3�Ad&�-ۈ��/��{�[��8p	Q�
/(5KhX�n��X��ð2� �3��;�]/bj���W=G	b�E��>�5��+��Z��#�(���&�W����}����Kr�\�@�,t��LX��+��s3�@8�r��TS�3S���&�<�w;F��8���%��З��ym�Pq6\��i�'+��;�+C]xJ����]Jx�7�*�$5��h��/&�����9H�a�?�����@3�(U��aQ�9{#���y�{]��Y�\��U1�����&�jy���?�n��HAj؟���rYU��ѣ�O�����l��@l�d�q
��:��g����*=98�L@��Ey͑>Ub���x}�|��AX��{x�Z�BI� ��r�?�:���s�������iGq���4;�]��M���Z�_i7�p��Ti�h%� ?��t:�N��,
�%�j��w{�=*,��/��e%��?�GV��-~�9�߽�L(O _��g�ca�`Ϊ�>i�K��/7���U����~s��0�;f�HF���J�t�t��"���p3��\�����a$B��b��z��GS#vm�1�N�T���LN��L���Vb�MA���'c�T�=tKL���pi"���0���y�n��}���g%4�*��V���l��� �u��1yP��H�o���NgN\J`$�D��)j�>�Q�
���_�QNW�2ПJ�}��H&Mi���R$�:8�0W(#�m �+���]��D�~zX�&�F��_�0��%�_�^]�R���q�������F���V�lzA����&A�Ĩ�'�o���y����EO�,�[�x�*ʠ�%	%̗������E����	Òj�RF4 �������	H؇��Y�!=�O� %&�an�I�c��Aq�11q�:)�V4~��W]p�:�}]K��5����&c:�g�?<�B�����`�41S!%ْ��h?��uZe�T�QN���B�v��A�'#U�����߬�(1~�]F n�&0/�U��� <�g�_!i� D*��Xy~WF����fu���.�ë\EH��%8�A�4W�1�`
�j�)�c�}�	Ї�m	�2�����GYk�y�O�J�:Q��[&��C5>��%�qY�+"�l��0�?d�FTrjV��Kl��V3����mo��D�,����@�o�x�Q�7�R&[z���k�GL�3�����@��d�R̪U��p��,�Eς�6��M���'�|�o{9�y��5����D�����Fv��_F���H~�
ow�����_��鍀DJPGs8������Iϻh8��5'��U���������Nb:�3K;�ٌ$���5/A��s�n�<4�¦ʓ�r�-j��mI����Cp�ʅ$�����&LR�F��#o[|��tc+��Ft_��~ �^���PFS����'E'�a�^�	w�x��e��|��ob��P��i~	m�Nv��NS_g5�/]��+V��6^��������=|���M�B����a|:����w��ル��q�у=<A9��&���}��l���8��̞z>}�v݂2Y���Nb&Ř1�;6Æ~��G��*�>Mg�I3q�Ci��*�E��[�VL�_8DT��׈7P�9g�u{��9.�K��%'`���pH�j)q�e<�"E���C�[%�k�	G��	���$�aRL�/�eUF+ö���p��;e2K>���~zc2��GM�d�[Ԇ�YXI������2���z��,$��Z,�`=����E��Av�&��Q2��R���|8FX����6��~����>�S��}L}�%��-l�җ䤄!!�0�Lן[>��1�٤���d^���t�`e�х�EE�"s��?�X3vءv�n'��>+F#�}�k�~���6��Ė��zm��u�/�	�%���]̞�@�z�r0�DtSL?���nǦ&H�s�K�Y�Ư�LFE��(s�6���(WlfM(��hO���?�3u�,#j*���������1VeJ�E�u� S2~C�������R����AX[Z�e�#�g��V�=${�3I���e"/DY�n$[�����(�ȘwZĬ��5A㮔�=���l�L=n�}���&��2��pL�tJ�d��%�e7k�j:��t�}�o#��4e��V�S,��)�ZQ@�Fp��KC��S�(��(A7eo��߹��$?���o�}d���L�偍�4�
��AÖ̃N�['�,0g~
�6M�^%P �=�\T��(8�߻�L��]d�|Z'��G�L�	��ێ}.<x(o.�#r�gG*��ڛ9
՚	�Ta�I��@�f��㌳9��I��7�1����s��J{]�t���;}�uA�&&�o���F����@3R�"�-!$q�.<���z3Ц8����(���/r34�Y֊KN�L�w`���FW�M���N��ׯ�wx��6<F m�pP�)vޱ<-8@&� ��� ^�e$�=�^p�X���nd�a�n,��YAT8!��@XF�E۱rc�}?�C(55Œ���3�tR��y�ٖ �)ɚkܾ����I�����W�]b�0L󓵿��b�4�p6��	����B�� �
)D���p�Rd^¼��u����^ߖD9�7��NU��������`�/)���~�[�u�S�:静&BՕV��#Ɂ��J��5��f����|;-ϲ�����W>ƀ������C��@�S���*�L�3����e.Mw�0l�{}lo��::[`g�쇘\}��{��5�#�3��:�1}o��Ɗ�~�$�&�.3.��ڭ>����K���3�G���E�ā�Vf_���@�\o�SN��5Qf����`n &g�\6?��h�~�`?�&Q!ѓV'�F��ԑ�Mg�h��8P��V,N�zۅ;�eW^�=x�m�1g��s�@�K�
�O9;G��4_�XN�[�0�g۩[l�>��N�CjEW�~h�����L��d�+Q�m%OWQ!����0)���F�5U��s��<:/!Q�L&_)�F�!�1�ϡ�	x���.Ö?|��ٝj�3�� �'�u� ���&v�Z���F�@u���6�Rx:	��k�jxS��������tjʌa�U���M~?�h(?��(|�]�����Y�ƅ�]1����~@g Ȳ�o���IȆ=�:O	�<���|��R^��zN|J� �NO�d�9�;�6"�*ͥeu�t�o��ZjG��u^Y��^���bt�&��Q%�a�k}�8Vc�@�U���~ߎ�	�q庵�y��U�I�`́��X���t�� �7/��.�����/l
�� ü�U�#����K,7r���#�@:��	AU���l.+s�H́�;��YL�IW�ґӚ��Rk~<%b���l�5�H@��g G�c\����P��+'�8���}�cK�����3����D��BWq��/���",)�E	3�F����-�?P%�L���J���	DL<>2?ڌc�
�1Ct��)!�?����4J���w�3U|���DG5�^!q\�]����Me�pW����T^U�D>R�CS��<��s��OB9��b�첧��m�LM��(��Ȅ���Ho��,�&	�P�)
k�������[�6�d������&�_��>B�1k�	�_�Ff1=��5�텖A���%��6�'D(}#a�@���&
hj�ǨayB�Lk�oA�Pt�5�1�<��."��k(�l�z-
k/�oM6���&݆sC��Hl7�z�.C��O[�S)=�ջ�K7�[��{@TFCT9���AS�;1[�)�X8�����wc(�{ lU�Z^�c��6�7?H�����Mքb�Q1
�R?��@SvUy�����d�J�K,��~�n��(i����U`[�<�	�f�.��g��d��1bUh;�2�����}8��Xj���Vy5঳�����`!r��@G��fl�-?�v�m���hU�n5��˦5k�7�8�cJj�����.Ȓsa7��� V�v� ?�E[6р���;heK}��R�9�B��C�h�sC�hڷ�@��H�M�O ���$�z��ۺ���h�G�/�RJ�OYKx-M�٧1�oq���zNO-%sh�F�Q�2!p}�o��~�U�Zy]�D����, ���Dm��Z;�
��SBޥ���c�Æo�y ��eGx}�7����w ��o��x�6E��A�0"B����RGm�a �b%D��-	��(�s��.UQ��{"���Mr�ФVױP ��g��n������oQdA�_8�f���'��6�LU;��EB��bbu��� 9M�]1���VEڍ�ٸ<ʄ)ʭ�n"������x��N�ul���������DV��(����d���Q{�Ѳ����OY�����wP%�գ��V����I�ab�j�^П�M�%�Qe�2�����|j�i�I�� l��.ڈI� Lў��&O�^�+ j�2k1���L�����f}֔/�ޔ�Q�e̳)"f���o�O5x�f��r��j^��VKϬg�!�3:���mE�*[h����`G"�ǲ�@��]���?n�m�7�Rv:>��8��r�W����/.��8��n7�] �1|����b��=�'ݓej8R'�xX�L�A�/�µ�Ɓe]�������o\v̤p��0`^�ܚ��E�X���@�1S��ͳ���Ȯ�2d`ƥtPˊ��-�;�faX������QV������!��:Wx
�-��8���-UK�aS�Dn�@���U�	�ٛ
P��B��W�	�Nl!��Yaa�c(���ާWw�gڂ���˪0�H��������33?kP��:\���KH���V�,��3�'c ��w�i��NM~�����������p{ڱ���D��fǌ���rvDA��ܯ��4�U���`��i<�m���s��@�W�1f�"��D�#��9�AY����"p��{Z9��CpI���p�]%{�v�a=~v�%3�+播�����Y�d��QD�k,��(��?C����&�	��Y�㳥w�"��%�g�~sv�S�����1f���X��H1�=mVҶ�b�L��v�0��H�Q�����$�xM�h>\�� &華�e�alK�㢟�n��ѽ֚���PH�����Z�$�s�@�����6we��J��kț<i�1����w��+]8�N2��J����@�%������Khd^�ZB�o���>9�GH��#���~�m1_͌##�K�Լ�{��1q���tg�&���/�h��*�J#a�PCaq�R
5��:�o\��cM��|�.��%��m�kTHA"�&G_���wB`�Ը��(2q݂��33���B��&i���mޏV1���
�NsH��*�b3�&�7�p�M��(�'P�J�yA��Z≾���� 3O��>�����J���ѱ�YO��M_0(!L��X����^dj\_PdY ��Ҷ���4�4-0g�t��:T#�I�����Ϙ2u��~�XH$�޶XI��?��"�ǉ�*/u��+���$��8 ��#�%����yUP�3�sB�K�(�Iu]j�p��.�m�+��6��x�)�'�;������`0�ҵU�`����<���#�E6\^"Kdg���e�Y8-�@H�e�~���2��g�~\"��S���N����I�ؼ����4��e�
,�)IEB2�^�P��!�ځ1�X�jA���anvy�γ�3%�U��&��x5v^�+�n�S5�r�*O���J2��B�'ԛ����dt�?�fW�<�άE;��>�osTFw��o�P2��E�`$t�{�f�m[�ZM*���0��_�P�Xx>�A"�hÖܭ�N�Q�rE,.k�8��wƓ2��W���y� �1�b��v�BL|�����H��:��D4x���e >L��-�ߥwM���a�OM+���K�yG���Y�8a���ǰ����`pI��f!%��
���C�
"
�Cz�X��ڐ#���}�XP��k����L�u���0]���73����\cG�s�m��3���p�fĚ�ٰ�O��GzS�M���uU!��3���T��E���k]�< Z.r@�h����0�s%���і�'v͐\�jc�(�)1o��l�-oX���4�dE���۞�ф8����_����@��%ɳ�3*x��/�8<���5{��b��T鉝Q�^��K^��Ƽ�*�s1d�8�������zy���,���~�o0�N儑�leۀ�^)v����1��j���UD�uŕ�U)�^��(��2߁}}�4J�7��L��bo��4q���k��}�����6�m��%������ �$Z�E�&F�쎎�αT{1Rram'�"$��	�#�aC�D�{�y��)�46,�f���n_�:s�����Z7��@�/���X�=�v�`0�+�>�=�MY��M=s���׶�A�F�t���EK�~��i�q\���c���hq�ethdf&�2�a�I�vuԼ&���F��k���\��b(����Z]<Pe�'��Ӕ5@�"
>:j1J@ׄ�S�̬�,��ݧ~b,�T!I�o;'��A���Bs=d;����Sl�'@$?�$Jl*���U�m_�����9��# ��h���X����ʹ�58�4AI���&d��4}���}��D ���d��׶A�,�K���S]��L���4������[!�~�_�����Q�-���u5��?��5_o֢�|��B��ŨN��$��q��sc�0�`����2�B8��-Z����Ǵ�|�䣟��Z0�T�y�8/0�'�(���Fz�D��O*�B�����l�#&lP�t���pZ�Ovcnt�x�d�8�	�"��`��#;d/4Ȋ���u!'w��{�ܽ:�6o�Ӽ��XYsn����R�+�E��	���#���w���F%c�`Ą/�A���P�a�HzN1L��E��IF����q�����*7�3خ�P���;����� ��0��0���U&�r+��o'H����-K �V�DƆ~�>�-�?l��,c�wΝ#�w�����X�CL���ռ�+ގ�<V�m(��|5�����m~4��vn|�*�x�:%1�{�RfVD���Y���58Ѻd���*�B5:>��ʙ���_�HI|�ә�`���0��[�==�I���֙&N�P&���?����<L�f���?���R�$;��s�ڈx�P���_��o��h�,S9�q���b�AJt����K ����T �*",��`k�}��Z鯵4� �fa�����������Xg]��B����;��iG�����@NNas�-��@L���''iv��)�3N>\zn�ЉL_�*�07�)�.~�]�����7E��r3�-->3Q��2E��p���="�]�^/i6� ��!���Nb��IY���$�X�0is��DD����"s���#����JZK���&�	}-���Ւ??���YLXL��Ex�/��!ԃ�s+Z`$m�%���Ek`�/�,W�����?��Pܐ����0��"#<2ZgRwvր���2S��I2{̘F���mF��F�CU]�)|:�"����1T���I#���i���ږ���I�D�С���7.��:.	[���Tz��߶�8���0�\2_�7 ~?N�=��f��Z���JFŇ�5��rcz�|R��U/���/�
l�y��L�r��!����8��\aJ���z�*�:[�vZ�W���6��[>W�uĚh���yQ�R�J8�A+���c7"��tWK�G����� f��'���jQ[�+5�;�C�%\��}B �`���-���-�5��L����x���1u0�Q�cj^��_`W?J1k��<-��-��I���99l�|�nZR��3����`_�ڜ�X���lt^ا�{lF���?�¬I�!���g� *�>�O8b�F��=��f<�_Kt�A�ǰ�c����f'���
I��D̀�d؊ze���ٿy��ҡ��z
KENAJ�^��3�:,��q�v\A̘:P�&&a�l@ym"�K�=��ג@�+_�<ȣe��,�O}��)F�j���2�@`���5��3�w�GuSP��R��'������Zj� �-��ݔ�[]# ��B��3�_��j��T¡�(������s��P�W=|��WW����s���wo��R��<(�Y������ ꐢ/�L	;`�t�_>9ҽ�9��N���׾�7��]�ۈ�J�!�����9H3����@��SM!1��gX�h���P���U21;�u��G�J�rz+te_����Hɚ=Q	>P�N��1��(�*>�Ȃ�<z�"B����۶xY�4\T!ơ���O��Ye��bN<'Iz��*[w�.�вL�ZW�H�ʎ���S0��z4f�S�TrfC�^<��sP44:]:�J/"(M���z�e�C��;�28��g������%�,��\�4[��c�W4��i2CU�Mp���>��ry�sA֛�@:�:q�l�k�H��-L���!�ސ���9xs���)��[PH��M��0�,w
�����Ҁ��T`�z�?��a6͂"D��`ƺr��)�l�-O*�E ��Q�|c�lhk��D��&�w�yu�(	G���,%��qR���u�^��Qk��an�@��{�\�=�o�l��̫E��/`j8�)dik�D��A�Q�����)�9#�h�D=�����r�V��5����o'"��	7��y�4@�ks�d*�5�WGN	�y�=���|DA��/�h��Yy�Ey�VPZK�2ћ�R���o��kBڂ�D�[ �΅�հ�u҆�'��yYƺ�X��uH,P}*#��
Ԃ�R�����Xi>�8�|���܉���TBvɈ��f����L��[�OՖ/9���棹l�HkH⑨�C�o(�r�%4r�	��q���Z#�[�J<\m��'�sO&������Ƭ>L�Z�����@w�y�l�'Z���f�p�.�>Nn&�]@g�q��f�O��$N�u�D�`��{x��N��}ѹ �K��厠�]��k
}���`�X؞y�y/:B�ɬ���@��G�2�7�G��F#�`�;S�u���h�����ė �z�;';�Ѷ]������\�X��Cj�>�59�z u�����Z>���Sd�t��7;*;
��0�q]4K�/��©J`��Q�h���̤�m��
�6. �yK�*�:��%��t���f��K���
/0 `b�\v�`-��� *�X�7R�� �o�-|R������mD���ە��<qzz��g�V��,��"�zwT5!�\����i՚�fa����ɱE�����H����$�G�?L��cуM���xM}pW���Ǌ����D������X�Δ=�qN�\��@A>�,䤴�>�Ex����F���-4ks��t�#D��=��rE��$fi��A&1j���,@IX�]}�SbR駘�,��	����^/�.�Po�����S�39F5�̡�N�:�D-%�
�H�Po�m�*�:����κ6|���!��D#M�4Q�Y� Dv ܪ�Wڠ��ϵ��E�߮�K�����g�U�ɉ�A��x����/��GR`�.D	� Jy%�Zd��YN�Os�S���@���x��|�����g��Ns����z�層pj@��Pj�Y�G0�^��s�� `?��F�����YH�W`8ѩ��R \ ����/8	b�x�����h8_����I��;Oӌ**t1��|�{���';ڱpD�}���M���;��)L��nJ� �x��k�P�cr�`0z�k��_�
S�����>�����ߕ�$��i@l%��杍sm��ˁX�@�֌�A(�w�uK= �ۍ;�XM�����P+c�����X4B�x?�xm��e҅�x�1����P���ڊ�k�j� ��)nj7/K�gH��U���J=������8�o�
��#��Q��ȋ��#٣L��.��p�C�g%:\�c����k-0�H �+��oH�N�4��٪FZ��f�<�DXή���Hz��Ņ�9e`���":Tk���'��QGS��(r)3��nX-�������u��[���n��mg� *�W��/������XN�����J�42P��ި{V�s/e#�f���xĺf3��ANw:d^Rn���bҰ��������9����c�M�@g�C�y��g�k��؎�\�d���%#q����qE�d��T6.��\�zF�*�j���v/.�l�v�`[���x1�Q��GXn�~���-V.�[\�@��H��i���g_Ǯ������:䉱iE�cf�N��Q8�*��	�-cc/�=rn��?�x�+L>fM�X��ד�Á+h�|H� �Lo�La?��S�a�/*[U4`��T�*���(tp,b��9��v�}�M&��a����	���'R�ٞH1�<9��Y�CCy�ǔ��;5l� �t(���so�̏r5����+l[�����n+֘��D������w.'3Zf}�13�v 9�z�%'�x��^�w������Uz)I���a�H��'��8<Z\�����>NSŬ��/ԡZS�ࢷ�!ro�,�X�<\�@#qJ"�~?�PG�9�D�Z��z]��t��X�R��.	�����>��U��C��|���i2�A��F�ʦ�~���J-��G=��r�P=�s�v�[���꽷}�A�*�aڥ}�?n9f$Ks��V��<�'��Pg��P���l�}u$Q�|"?���Ɏ��/#d��d{͟�up��Ua%�!���S�'X�-�
�Դ�Ѓ��Zםw��
�o���8��w�<�-U ���Iα�����#ɦPrE��i�����y�`����g쩮^ �N�>�D��#j�(]��U��b�&̃T�qw�C�r͑�	�_޴�'�+5���g�q���h�!k�b3W�����T�A)]�u��,h�A�aA%\�������ݿ}��Ũ�'N��/.PY`6j��R�<J�_���Ơ8��Bu���9د�S�LN蜴Л1�q �>Ԇ�:!cS��,%�حq�{z�4�a7{K?�"�y���4�-��O#�\�B���N�P7Ϧ\�3ok�X�Cn�`�69� �y#X|��O�|E�,������(������E;U���GU�~=��g3��b�N��}�{~���;��I�H��?����s�e��/�x�%rQ=����+�cs��z���K:��P:;����>��5b����آ�Y�oh��pa��}bg�^�4��H�t���v�ņ|S�P��K������IIuS&q���u����6�\��]�a�%��Ϥ��ա�ͧ@�M�l���r>� v@8  �Z�ؽ��ԗ����q��է��ÁV��?�d[����v1*b���ᗐ	�"�i?�?T%�(������We&?^��B�2�Xh�Lڞ}���^<Yz����~�3s�}g�#}����>?��O`>z���)�3&��[�:�@�!Sk^O�A��:�"!>����-����%#IӉ���]�A����Ɗ�d<2ý���'�'f[��lHKo7� �.����l�y�����t\|H��~swO�:5�>�-GUuf�n*��S���c��e� �v�A�6ױL��{��pjTf�e��E�4�B�ۂ�>
K�6��f��x7��]Q�4�n��i��=w�+��p�ށ}��
�@�Ăq�NƕͫMd�M4�P4M���q/L7���:\9�Կ��Eq�B�|~�,�ri������0��o��ID�A����@��|�H����M�0����|�sc�%6���ߎ-�G��I�+��[?�
��j���NC���ޑU�$�a��_�ٚ�wƛW�9�_�}��R�m_@c�Gh�?>�cV?Ď��"7���/K�(�{�&��]�~�s׭����1�12A�P�X�H��NS��h�'������f���
���V��
UK�>�7B�F���O�j�����6+�����W�j�geO�ʈ��.g����K�Hv�f��>
!
���l#��5pS�|z��߫�s�%~�/��#W�2�������>�`n��!��:� �ճ��]fB�T@�έ֖���)�98x��A7{^�^	�����i���rHRR�1^�����	9�V����8?�s���$�=�8A�������c6 	-H~}B�s ����龳��$:����]�qơ���j�����K��l�m����d��땵�X�cN��į���V���V����|��WA������BPg�D�����D ����e���V�݄�jPՖ[͛�X���U����5U	�����e�r�IqO}g��k{V���F@0�kk[�h�����7���em��y��a�I2�m��v�9�GK']��?�4iD�9�.ST��������Sx�L�$Um��8V��,d>5P����E�pD����UP���{g?7��y��o��^5��2����N�%VK�я�怌����Dk1�� �f$��׭R�k�IM{��~����������w>`	$u���.�m��H��
�0��!g ��>�8,��e�F2_2��H��K��Y� P�ҙ��t�L��\�r�?�$v�P;L3��.�:uScݵ_*�X�΢�㼕IuT"���FL�
�9��q�������<���u��5�X�Y�A�7t�Qk��9I��7�9���b��x�߈�E�����r�"��Kؘ$-z_�'����$����C��Y�BR���>�E.,��4�K��1&�#�eE�S��K��~���Gra�l��17�).d�ئ���3(=�/uI�r�����$��Ze�ffA�?���n2RP��hi}���mE*Y�\2�3��z�J�%_�����PD=RKn�uaI
 _����D��|n"$SrDcEo���Xd�	�?o��,q�<�vG�"#N��Q��]_������*H(�����N�2}��b !��)�/���HĤ��4�L^�k'�˦�>���5��O��ig/,.�MP��4m��nڴc�8��j�L�[��k����V��u!
��<;��s�)�4UV�L�%9W��EXE�}|����!I\�~Z���`_��}�sBu���_O&�-�B@������#ar��|=C�Ag��k5T���jĞ`�頊ȩN���5���"�A����Emʇ��=[���"�vN(6�����ZM�����>�_���9��Uo���5ċp��� x0lS1�	y���j�ʖa�t���6����˯��RI�6)w�_'E�1e��-�I����y���{H&	�k@&��x�ͽ^)5ߙ,ڔ\��g�i��t>��������܍������"� ̵��r�E����ɹ��.��0}+��8:�^�<�a�d��)�� ��Ȟ�F�i���{�vfh��K��%KgԬ��@u��f�M�o$��R��Fc���<��&��kq�7�K�2�~U�NH|b.��o��}Cx�`�T�O�	W��9�>?�"�k20��Iq�Km� ��gѱ�4�Z���Jua����{ �&&"�~T3�k�d��n�f�Zߺ�i~��Sw�[u��ə�%l4Џ']_{�Q����B'8ֺ0���^W�H�o��&��+_뜗��7���	0.�h�Bi8�k�S+~L�(J
��������L�+< �~|�!)t�McI����@��2�
�Vu�B-%�T@�&�o[+��B��N4�JVX%�W?A����a�L�d��c6�CZ��?o�+R
��U��1�!5I2��y��4�v%u���+Z"W�U��#�+�~���T����Hа ��hO?x�튿lc��k�=7欇/Od���"f���5n6��I�n�����S6�bh�]�̭dE'N���ȶɇeo�,����ԝ�j䞝��3�T���8J��|��b}�C.1�X6u��gYZ5΋eE�~���fn�H{�����o�%D���zZjK��o��OΠ8x��!���.7�b]�5�Ŀ�A�o�����Dv��������./#x�mPM�p⠶ж��O��"�/P��;��8�����PN��~!�W�WA�Q��V�4� |�w]��VGuq�i���-�)86�f�{�H�j�r4:�譜 	�Jǵ�(W(��~�nTNȬ7t3{���x��̢d�8�=�B7�Jz��ZyǠ�2g|��#L� b�J� r�z���N��n����;�U��2-Xkn�7�p՝y���p�VX��b�mJ:J�q�@jL��|ʳ�Z�{��M�v�����3���*'�#~����%��,A���Q��,sp�?�%@�ޅ��t�)���T491G"]U��u�	>�I����?�Y>ě^�ڬf]^��s�'O;�+?cQduC�� �N����B�_��^�:@k�(59���r{���Dt�:V�a�+d5|Ɯ�=� Α�JNu7)ON����7t���9"etc�n����]�"_lK��2�:�<&��I!x��K��t��q��,���t�u,���l�k����T�W1ɼ0$݀�UP8ua�s�F�x;�S���&F�o��N�Ji7w���}��*4`��0�����&^�M����+���½C+��{�D��S$i_�r�G	�I
�Gґ��e\ ��@tC�j��U?��3�n�'\��f�s	����=0��
�O΁��p�e��'8q�с�
�2�>Gp�l]�v%���`?�IZ��W6�<1���� ]B��5�H8��
�h���=<8����Wg��n�\L1�䠽&�+ؼ�q�	[�,���PJ�p��I~o��E�G:��Ů�c�|_���Q@_��FE�ꨞ�Y�=�9Q�Frp�1���;aپ�n�y��)(>ZW��drq�yve=x�3�/�w*���g[�U�6Gi�	��[�z����d��iĝ`:�\Mx��6��K�1P����ا��P^L	!�9]?z�9�=���c�|�L�3p_�nب�,�:�-2�&������
������~�8Fmӿ�5� �<*A��Jc;�ף�P��U5~��ɎЃt�KJ컡��<�a9�hdv��C�ɚ��a���R�����/�l7q��x�Pb �f��	�3`tmf��!���<��{��D:��E��]$��M&�9Ŷ�n���	q8gD�ܐu}�tNF�
p�I.}u��uRLpɪ�S�i3�V�>��	�&B���u���@��i��Vr�H1!k\$�[����4�6��
� ��ɺ��k&�_8Y��]�_b/R���P񰱈�)��*�p���~��c+pw[���`��{�7��0n�ۮcQx�O�m��9�ow<	�&�h�qV�i���8!>,�T��2��ȦQ��>R���0\�Pߤ��`�&|�w'�� �^�$֌3x����
`En�) ������	!�ÚnGIי��ƺ:��y��t`��k��N�~%G<|<�����ً��_֖��d��z=FT�r��,F��o/����]@0`�DS��l4�z��Q5�"�W�2p�p!O�N��ج�D��R�B`� l"�ܶ�G�~R�&|ы)���W#�}z���lN_/�(,s�#���j���[��0�PWe�dz�!��x�����:*
���e���3m�P��AX���wmr4�sE[�c���G�ySunD�3V�5��N\m.��R�r+���*G����{΢�Hh��-��R�X\�y�mX�͡�Oz����YI�;�b�զD�?v���5thiS��^(:���>l���H��	��=�����.���"��Iːv�:�����W��*h�
�f��x���_) v_՟�r�g��
ԥb��κq�������(z*�$��ݹW[�����U������]�H0{X-J��V�]�FT��q�@�E.Հ�,�j3��
�������A�Oh����Su�3~�D������wJ؁��3��j��#��c����K���e#K�N�����"��_n��
�d]�y�;C���oϞ6�32|z£E)����y�l+����ί���Y)��Yk/l����.^��� �1��}�Y$0 b�?�<���dU� �����Wϧ}�c"v���o[)VF��$�2M��zp�{zTlY|!�C�C��8��S���?ݵӫ���-�T-�8��G�%����E���0�Q7�Na�B"Q,nK���i�l;�zk�QGZ���G��,)�X@��pk�֝���:]�"�=:�R��ԋ�k	cXO�L?~���)�PI���)�b4�ww��[�ⱓm�����%,%c�InZ�76<M�f�80"�Xn����0��wIk8��b�`����0�.�u���c��X�޾��*���.t�l<}f@0�f�ټ��n��?�&!���\؀��	L��j�h��m�-�c�S�k�9�l��gS�C���MW��ul�#�2pT'��$A)Z�s�"^
��@2��Y��]\ �����5�6�S�&n^6�<	�lP�]��ᜬ�<Ͻ�a>�J}&��@>��Iw�E����㨍��<�@����F�3�_�l�
�|����Se+�M�ɔz�01Wl��nū�43늫ԃ��g��6�P�t0����
<���g��,�=�4�j�� &�t�J�J"�i�b{m��
Qǿ�E@y�g���T�0�1U�� �`��~���
�	c���pϮ�z�U��Y�.��p$kMy��yh��d�p��;�O�Ϋ���w״x�6kh�����n��K,���꘳+|�4B��S�i=8F1�fi�0��ׂB!	�g�5�&}��=5�՗5��m�?�����c���w&���B%��޷��5���y�OR��I��<�pJ���ni6���5�/H[eMb��WV��]�,5��J [�+A&�����8�.dx9âY���������K>�3��f�,�lq��{������s=����O��LQ��d�s����VO�]�7Зd��Aה�ǜ����B�w�
��$S�7'����R��CZ<����&e�?̄S�W;PC��r�H�ʃ�oZ�a�� .�"�@�*�%��
�#�bᲉX��yl/���!kC�`�+���	�>�r�MR�5�;��B��b@2pcxq$7�?�9�}��rjf����L0cČ�#�m�#�`�Q��~[V@����s$�!T�ز��Oʦ�84��aA=HQQ��h1e��5�^[�e����]Qv*,����'JG ���w-���f�zڷV(�F��L��w����R�M�S���4R�,;�}�?W��/}�2ԑ�6�I��P�w#��x)E9�7V64%M�N�c�^Ex���$�� ��X��o�J%/f`�{]~p�L��ș���%G�l���0�!j\b�w݋ی�CH!?B����`�	[��2
��K�L�|��Q�Sڛ-w��
��ϒh��>X����s��|�,� �8�*�ӈ4���-�x��� �7����"�m�iao��!PX����PJZmݰ��i��;Zrl�uǿ�b�Y:�.��w��CO=6��>�I���&;O�x�`�X�G���C��)Ҏ�ϩ�,�ԣ��-I��M�G�����`3�V�M6���yfv�1�q��9!]��V�]�+ւ����R���'DY�'�:�K����v°`ҙ<����+��gU���^�*�}BqLɊ��>�6�[���0e�D7)e��+����-V���m<=FM���ɀr=Xb�2�Q\&O�����������p��݃)@���(���b�	S2n[�{��4����7D���l庉6�FLޤOV����j�;�-�OV��M�]kN]Gy���I���v4	�?�ф7+C����ʩ��w��$W_�B��@�EZ�q���֌���hMu��l�@��:�ݺ�;��:����Q�餰�V�u�*_���ِX����T���i��&�e��1O¹xXǵ�����N��@)O?2���𰜻M�Dٲ�!IŮ���|����I�?�q9���P�|�/R���&,�oRQz��p*
/�u���T�TacGڥ/��7�h�}@�`�����9ĉ 5=J TbkH���"
ԅ�ʓb���@J�d_Yп����C�yeS�7����x\�P�&��$:B���-aM��k���`�1;�G��,ĺr����84�O֭���4kfrӲ�ғ��O�>/��K��P5�7��l�p���'и�߿�Q/u(^XL�����z�`�(���)4�~��*j�8��e	�Q��r�Mx^Ͷ����Rb�lL�Kٍh��/���;�)�\��=S�+p�'��tz���nC���g�&��6��_B����|M�Y#������c�Zy\a~^�&=�b.�XOkǶ��3^Y��aָ��<pZ�r��~�S3 0�����ytd��L���;]�!wa=a4�?j0�2n6_X���?	]z��MT�ǋB�l�l���#V���j7vc�h	s����(cGQcbf �4�d��a���Q:w�ۜ6i6����$^��$����F&X�3G�(�ӎ�⍤�S!����9��s�D���>0�볨4a��k���DxO߫�`p��s̬a�boV"�725~�J�g!H�O�����pT�/��<N�6���'������q��^i�YFn�F����W�&����X��yΗ4�Q��	^%�vc�c������ i��>���T�@� E�jCی/m���>%�G���Pqȸ�%��b���I~����ٯk{Ǻ9t�W�7]bb �A�����`w�@7�bY���"a!BU�����d}�*�Ȝ�\�~X�����>j<P|��,�'��F旂�&��Ә�_�Y�aP��wCܐ�G�.(��a��fd�]A��s&��%�Mh��GUE%UG~mp��E�!q#X����_�1���}�u�9�`��D���Λ��o����MN�z��	k�%~����e�6��Gh8C�hȎ�����q���?��`Y��y>��2snb�r�>�C�e�o���w�xBw��}$O}1��f7����y�,�z&;W���Q����n�*<�zV�����ߤP>�c�DC4w`���j-X�	(�1��cA����:�y���KM3�4"��t�����R&춯y�B��s��Oi�m�]��E^�+�̢Zš����S���A�˄�&|'Fk��K|��,Q�^žAE�4�X�ĉs9�v<&J�ymD��י^8"ސ��8Mz���m&��4��k|Y�c�;˅����@��(_�f=����Z!+D7KL=#~a>v�Q2�d���ǵ}�JR��,��>d�ÐF���wg]��[?�<��&8��9�s\�w�l�07l	(�[�����R<|��h��]�wF�����_�G�vm���w��*�,_�,��q!�h��w �m�H�-Tb�
��͛�p��)�lg,W��?��$�83�i��������$�fs��e�NӂW�.����$d�f�i$c��6L�2������/�F��c��/լ��#�����!\�ds��Q�RƓ�W�Ca(���ު�Y�=���=�G�����y�5�p����D�(V�@7^�6#$��Y"K���pc�-i���2hv���j ��yN�O�#�D:e����r7��߄�Nԇ31��|s��bh�|KUŎ���݀Ġ�=��R�V��1�N�М���i|���_����$W�������kd8(�����I��]��V�v�PR�XA�@�;r4��4�!�W?y�|���;.bG�nt}짧Y�b;O�5ΙbtOq�E�O�d
���2bT{E�8�B�ʘT�1+_�!v1h�M��%̝�j�w�g\�+���<Vr�ugOol]i=�7<��nb�R)�f�l��`����`�J�0'�1�D[���վ�Tf�a�{3���_Ɏ���]�m��!��Vm����`���[ᚈoU��M�֖��b���X>��5�"0nk�ms�HoM�T��E�I VE�s}v;���!1ʭ'���A�C�~�x��2�?2a�]��#`�sqtGJJ7#�����Y�������~�5g�m��'�7g獀g�2�F������N}�:�B8D �i ��LZ��d�n�RE9��!��$`�l.�t�a��9>�K����յ6����'�P�p<�_+�n������5�[n����(�~{�2����@e�����bU
h��)���˽3�S�Y>VjW���b�t��9^��ϧ��?Oj2���%���]���MQIv��?�DO;+O�Y�N������4J,9ɇ{�
OG�?�#z\e/jf�
L�KN+.t+c���W��'տ;�\�/�P�Ŧ6����Se_�Ⱦ^�f<���"|E�y*C�8��	I$�K�(�aO�C��E��J�@"�`�	�(��v6_:�1|��Ʌ��=��m���ܡ���[�[�O_K��-Fk�g�g'XM˼0�m+���
�y�3
@��#�BqN+�j�RU�2[�t�" �2;���!p����!pG�{���l��N9W7�\(� c�IґN;N� ���3�2>�����`�X�F�L��a��!a�<%�(j�%��ʭ�\���oW��������V{Ն�d��g�I�OH2?��Z��9ǣ"�"�8�a+
�Dt�Q!��������ݩ����=ux�#������[_<w/T�瞆&1��X_T��fϟ&A�j�&���V9gA��!L��!u��"��'��C}������PSi�G�0�
��q�?�4���ϫeE���c� =ɵH>�3� ?��P�HRq���;� (E,LX +Nne�u)�e�˙�ء�~�X@�|� p^�L�j;u���܅�ߐO�p�zŠWVI}�������|1�3�fm�hz��x˽D5���I�a��Y}8f��úEB�L�s�td���G ��u,~��x��!5 ��ѱ���s���� ���ݾ�����p����XKaф$�hb��hOb�ҧ�0z!"t�96:�!Sh���Hк*��L�=*)a�t]��q|���M�M����?B,����^��W*�4~�v�dC7,1{"�7^��� 3it4�x���~c�LI�ρ�<��bM`?܍���ֻEԄ���Y�Y|m�,����W�z�~���H�e�x�>���nל���h�~
�ǵiD9V�!/�sW���H�ً���8��g�MB|Q�X�F�.�G�-1ۚ���A_���>�c<誸u�@1O����q���V��Y4�ǎC�u�;,��-��=�c2)��Q�g_�{]�7)̎�%^���4�H��籦���ס��#M�>���&^b�oOKߨ���f%�b DҨ�N38򂩧LIZM���2�I��z�b;Z'�Hyb6�gDZ�Uq� �|4�y�#��O��x�����.��	i5���}m
�Q��~�o$�RF$`�[�#G�y(����tq�B"��V�;�.�/\�At��_�t�	eI��w*ݶ��;�~Qc��W� %H��ߩc�e^
�n��h�0� �ݪX��1�Vn���ax���	d����<�a�s�q�)F�u�"wk�@���Z���B���}��'�H�;���TB�q&�z��\%�D�Q4 պ
��ig�+o7��q^x�gCY��8�'�+�M}ף ����<U�hDwi�{t��>�D-�P�~��K=ЭfW8�4��z]���⦡i���Y�rv�gz6N���4@��.+�ч@mB!�:9/����*�ϥ� ����u0�������u��8-/���2$ǘ)[+�I��"�*���Id�oˆٮ�S��˨9rP�����x֘H!�����-�	q���
z����m��<IR���I�nO��<�����s[^�m+o¿SҎּI�w�KGuZ_�&��͇���&'S4~#니�#0w��g��W8�ɩ;�y'��z���m�����{U��3���P~�������9�,	l������87�bZ��%�����G X��'�:FI���i7'Y��];OEM+4VڎhK1��rF�Ț�%��h����=	'��Ua�6hآm:������`8)��\�������5�5HiI����z�,�s�/�}E�2���g3���˫�4�&l3Gɒ�^�3.,��ن}M���+�������tx-�JV�9
*r�aޫ�|yP�Zk�q�keu
Lظ�1��bw���&r���UDa[mfF,��M�^��S�m��s�7�ip�>���5��G3��Z#Z���Ƒ��E!�R�+�/���=6%���륽'S���ǵhv)\��X��O�FN�@�1[�#y�Dzb�:����+��g�-��,"Hb[�zͷ��S�g���jI�iJ*� rf��~1h��z��-��䏦�EL��mw��h:�E[�qة���n^�Z
��	��D})~����S�$�^nL*�B����o�J�@���A�&	:������lm��q&�>��/7i���t݋������a��lČ�JX��nB
0�!~k��$D���$��yX������Kr�s?g����,�RX-]�����cU�F�@����t�	,ՠ���RUD�����>�]���zo�b�N�^��<�V�~X� �@ʗ2�p��&:�����oWyM-[�DX�b'SI�+��ˈ�5V��r�`.9����A~���x���Yh!
���Bvҩ\U��#����h��n���N&�����Ea�_���� �_�a��Q󁕠�L��8"��^f/q���%�v�% �g��:��������HC�$<=Y���{��8����������	4$��,mۍ��274��N����a��}r�����R�2���Us	j+8���IZ��W&_kA^=_<>�U,�o{0�<��Z~a����ϛ��� "[d�lrX�f|Ag�6E�݌�X@ߘ,"%¦Z�?�5����hP��-f����xG�V(l�'N�"L>/����b.��f��p������]]�F8�Ө�*�R5b�P��I;�a�>�U��M�6����C�+F�ݴu�B���6������N��9��V1N�(aQWǴ;�;D#���Ɨ����%��b7X1g�QK�!���xR��8�����=�P�� �}5?����k���b���$�8}��Ee�L�.���yt`�D�N�68���V�d����{K̉���Cqڿك�M9Xy{Y�0�3���|C���C�s=X)���huS��$�(O�f8������t&�X�?��"dL���{�� �t���EeS4Sr�^И���$��t6rC-���A�ɋ1�Ŗ�4�����ښ����!���^�uV�1�e��ƛ�Wp�L��E�8�^���q�'y�}}�9������t=A=�v����lj�����to�^u֥�S�a�G����2 *v��]���l6�_	Hi'��>�e[D�j�����&�]�%�c��a���or� Q�����{-���Ms�X�X�=�=`�(�G6��M����32H=�v<Mʗ��j�1m�\� (�;��m��UL�_u@�?����,L�5��]yv�ԽV�V���m�����n���(�����b�ov���y��ʴA�؜|Y
�󉋍f����a����E.�O��_�Ϧ�n*L�kk��Yd
};;
�`�8�@�x�&.-����(�w�a;�o���#|�)�˜�����5���#W}��5��K_4��ͦd8�Ճ�,����,��d6�F��iV��wR��:�^*8DVX:��n��Gg�{o4>|�%`8�R:{:����U�Ā��S9�A����;��q)D!e|����U��y̣�|W�G��Bu4m�Y���<;��<d�a��P]�]���ɸ��[�^h꾆�k��(X�{����VY��|| �!�'#I��[8+T�=!)t�elK�Tj�����ŜצUo9�i-�7���<W�E��ŹC��^����wC��qe�\w�� �\*zsд�ϗ.^/���V�ip��*��I*qڒ	��tX*l1I�y8�j��>�;yr�F'��5@Y a��(Jԫ��D�#4s��<��8��h#=c���Z�L��)�6��m֙�����F�lӥ#=~o�ယ.��S�*�&/��o%ۦDN�G�$��8?�w[�[���V:=�2HG�����Hc��2M=�0��<�Ο:? �TfA:[1�ٳ����7����VI/�>R�?A����!3��a"�����������su�;~�@*�v�R���ho9M`�V���\�5T>P�9GF.!�����Qޘ��~1�,/�%�4����N�5ï:�ZD׫�@���>�w�X !Ĩ�=��P�z����N�u�^ ̧�dEC�8[�G�*~�_rG"k%��n������;�V���9oش��Z~kAD?�9���������z��x�ߘ���(�a��W �8�;�&�ì�9./����&�!�Rk"b�`!"d��!W�9�e(+*Y��>Z�X��N�w�@��)wͰ��JmV��
jz���������Q�Q@��]�黣#{g���*��Q�3_v�Q�l�t�f�X\Н��������mH��ʆ����G.(�LP�%�#5����*�Pq���D�����G�C���$����g�c!��}|�k?l\�h\ b�4Hh��ӡM��^?iuoO?����S��!���j���$6�B���ZU�ԆQ�m;��h��*�R����Y�e\_�CO�$*F���z�NT�!�T��$\����>�2��K*�k�LU���������{[(uϝ������t&<�RM̰���х.o�+C+d�u�kˌ8�R����H�g�s��:�؎�������9z��dF
��1�@#	"ț$F�UGP4G����/�z�$~=%q���oY���S*�oOc��v^7�iB�D�w�j�%&Q�ֳ�)�x,��G�1��<��A�C�l���6���i<-��de�36��Y*g#�q���mk��z��&z��ʺ��	F�@Ș��V����R�޷�F�-�#时m�5��q�jyX �-1�I����MI���n����;,K��s�QU�Łv��~T���4a;o2~�}����ZX�+����5�n9���-�����]����F&�
D��w�0r�q��w0U��VE�����l.��I�?�^ ��Zz�7�њE7k��Ss��_�D)�̎,1�$;幾�(�O�
KQ7Ul�Bea�o�ۭtg�5���^C�}�n�u5΢%l���p�z4�'��_e�i}�R��\�Q���S��	����3�9��*��w(��uNd��g�q������R35��s 5���M!,hXh+�<1�8��{�����d
�?�Yu�p� y�J��ʘ��|#�����k5�8=i�8�ޮ��Ñ�pg>k��N�:�s�Q�_��ݔ=�ߦo�!"`�Oy�zN�u�+�a��Y��>���`V�X�c/6�:@9���w������ ���^\2� �t�g��X���ct���kӛ�V���� uc fG����i�6��(�� EeHU�x����0z(�']!3)����5���`4�w����
*O��B��ř���FG�Q�i��qy�6�h&�ar]����q�W��s�
��;�p��~C��ab��AZH���\�vf�Q&�P�[m�Ć��C_��'o2���P��p�)f�>��~C��D�^�]�����\�-�+$p�w����!G�e�jy1Nd��P�KT`�����2Q����n-�p�ժli�60;o�p7.t^d��Z��jA!�_K2n���^h�+9�����1���?,��_)|z�f���ui���%i�@�2�"�Jŗ�|�g-v�yl(��S0��*޶F����rrX��yNvl#�Gb�Jk�����qq��2����I>oԖyn�*���2�yz¾�ߚX���}[PF�2��Ҧ�f@�@1�7?�Vi�����Joq&�^������{�z����#c�a�jKn�v�~�5\�9�!�����x���A�����[�����B��D�&g�j��lZ؈���m���HH�qV��2׳D~$J�3�XE]�oT/�:��U���՚�m��Y����֓�q��gP~�~>@k�Q�;.��x���3	O���a�9y*�|� ٽ��>dIfj�d=R�^j��
Q/�a���(�1�e>��Ӡ{~��I��:lR���}Ni]���v�Xɀ��|qEg+T�;�����l�Apz�.��_��~�C�Xag��!���by6�J�%��͕A2����.j���oZ{��Q�K�$ "?Ё��zY$	�1@��#FT��]�[UD��J������CZt����Z���"U��{l=s���K��`w�Y����Έ!
�4�����φ��54���Wun�bO�����K�28�!Ysa��Y���SE��c��F���]լ�����K���r�&~�j��6��g��T����"=	�����S���q�o�/U7����r�g��X-1�I�H���=_�Ө��ͱW ��&���Q���J8��$Đ��yh��o���^<gh��۰��M�������:{&O��H9Z)H,���Zpۂn�ڸ晇8�s�N�yz+"�	���/�F�dr�Z3���K��~�j�2�=�1�u6��޻tp�FiȂ��6�Y���0�R�-w�|_.����H��Pb���Òػ�����/�\��6�<J�q��-��k�3�|%��(Z�� �[f�����5-���^GD�hAg���^M���o�����C�v�{�qD�{	(!���6�|MN��U��׹d-�ʹ]�mf����^��A+�M���
r�3�YZ��s�)����?c3�Ǐ��u�F!!܃o&���'o(?�\k�O�|�-��lJt"[p���s�,܆ T����-	'�[��q�ؔo�?����V.ݭWd��Ӳ�����>����_��0��"��qxS�@Tp�D��{4Ty��B���s������,P3��]Đ�Y�n��~2S��?�)�i�@sQ���[��v*�z�!JY䶥ac�ۧsc��M!a]Ij)���#ݵ���Q���M|'�n�Q�[�`�Y��l]D��D�S�T�\�,_�L�T�Z=;ğl�~i5�#K��d,H�t
��H���v�N?����>�����tW�|����嚧Vrۃ����	9u�2&v\�F�+�d�ڊ.��Z]݂�HIL�&���j�1옉4�Kɰ�we��� �ěr���d��3"ζ|K�*)�I�b0�[�F>��b�	�ӿ\R֤�k��߾�tF[a�M�U�I�t�� ���}��:�RƐ&5r��Y���\S�NJ��;�
���^�<_I��)�6��A��@X��JMA�tG6�ē;(q
�OK����}rH]͂_��ä��O�s�dP0��Kˮ}ے�ʹ����^w���mR6�87í��	�N*EOm�IEt\|Vʼ~�X�/�� 8���̻��Y|O�N��g'u�c�X�C�����������H��b_�7��edI��Y���V��)
�lo���!�r��f���+�f�Tw��tkv���m��H�+�4��q�a�p��d��;{R�|���c�A&K  (��#!&FL�*�F6=Q�hYkCą1��'���u��}��^�SӐ���N>"N���ʕ������q=�揎`������9�Ld��/�?�'�x��i��-U\�swFEt��`�~Z���hw�R��� ��<u�^��K@0����E��?�Z�1��/���~�C���wڝoB﹉�4 3�]����N7"�fE�=��$u"��[gڍ*Z�� [�96>�d_C�~#��Ӵ�X��~ҁݻ��jQ�@�B�}E�M��'ی�������YD�����y�kϟ^�S.��U`��d�8LG%T���H:М#�l����k�Aƈ84�탌y��*
&f�yZ���e�Nג�,�uI0�͠���؉#��؄:�Jٱ9(I��IBb�Y�ls�+�9'���q�+�}�l���uT����/�	�e��|TİP@������񳏛h��E��"�e�]_�P'LV|q6��6�k��jg9>6��޳ٶaj��g�p��"`oY�԰C��p>2�9�.��2�es�H�g�l��E�4+�U҃`��GR.dN�����(����:wbQ �����<�/PZA��,W@�ͪ5|(�ep=�_�h�h+�g��cFDl���ۀ���Hs�J4E��� t�/.{���[�9Xfy�v�����?����M�Ct����y>����+��&h�I�Q�Չr�GF��U��*!��MQ���@�*8ov(��*@F%�?r�S�<dj���!�Bg�ӛ"z����� -�>&�^ ���u��Z�H�8���˨h�!�$z	�����b�R��M�:�����AH� ί�JC�ѽ��rn�]о�lE��*\���=
��E�¼��@D+z��҅-"��P�'��30��J��`����D��fvk�a�7������q�?X%�1�p0t%u,�2�i����X�������y�S ���|*;w�Wْ<}��)p2! �������G4C*�Mº�Sl5��S���i_�Q(pW�����9�����O/'��Hқɾ���Y7{���[�妍ߋ�O`����W�B�zH�gm��������������P�*�_RP��7E,�)���2�u7��p���9�ƴ�������rkb6�cpm���QMh�b1?�穠�J�� �"1��I�i�D��A=���ѐ�����v�Q�O>=K��R��8��:L����S��t����Ԏ4��Sb��,�> f���%��$�3�_�����	|i��`rhZ����1]��B��8�5Π~H��עI�:3d�/����}I۾�fG�	��#��s��ˍ�d���EZ-�#�Ԝ�S��p��=y���'�`��"��z�8,M�0>�`(`s"S��c���
�r�4Ei��O��cz򊂞�3��'���`�=��
ZM~���Jcs���0;^�D���*eb�^+iVˏRt%Ȁ��h��j�'����jL����J�4=8ܬA���ʝ�@��� �,�QtC�;&���*�X-�^����(E�C��f��I�=���&�N^(�2\͙��$���>#��C7T���-� ��6��dS�3�/�H��U��#hBkK���R�Yn�$�}��5�$́� �Y��M��o���일��������Ph�2%\;���
J�%�E�lw�t��q-��W�����;a��¾��S��oA.y F��Ҿ���C���)I˛���W��r��Q����qK4�Xv��.K�M��L������?�-婱Ke����)zt�9����OB�;
̴�����q�D�^sn#���]�$��yw�c�ZtT�Q) I8������z��NL.�u2�>lsE�Um�3�9��!��L�Th�MbJȲ�8
���TߌC���D0���^��)�$��R�z�LҖr��F�I f�~���{��"D�E[V�\Z˲@C~��=�#f<������x�(01�������ͦ���AGʇ�I �>=v��^�Űa��.��_~���~�n�8y�0^=j
��|�������-�(p飆v�g��u{)_�������Ex³�b'�0����P*9�xi��U��\���{���g�'��G�P�,]�q�\Q����:jW�au%�-h˴^9�֘0�)��g��8-���k���hx��ʾ~�Ǭ��H���n��d�4����$=�j}��V�%��$O��Or�m�f��p�	�w��ڈ�p�:�a���A�=�-C� �����&peU����":;E��RndF��F�%��YU��[j7.����QR(����
����GP����:5Ug����nN^5���Rb���V��h��������z-J3V3��:Jk�#�	V;���8!G��٢���.(f�d��f�&G��?M|Gz���":�)��}b��i�`���#��ß���z8�I�D�n��?ϬNC�&Ǡ�ZW)��?RM�S����vk)��ܺ�ר�kq�W�/��21���Sv�`��L WH�b�ou��|�5FȻ��l���8���Y��a��F�F�΢�	#Kit��
w��D��z!qd5Q&�� GЈ����'�`mT��W��˩��j�&5�\��k,ȱ���,P��L'Z,IV	1٬e.I8�(ߊ�LG�xI��@-�p��֬b��M�L�ZU����HV�^�~��PH`��+����v!�lS�J���JwI''�� T~B��t�->MU���>���F@>�!l���5�ȑ2(���GT�%MۯNUU��X�����>�W1�@���+gH9,Z�[��Ar�Jv���eE��~�W�m'���0�:����8Ba����s�=wxo�_�	���t��~C{�Ҋ�r��
�zҾ7�z�2'e1���s�ו���ߕإ�]:s!�������q�9t�N�����ѥ������� C_�@4�Te�g�������&�*�G|�8f(�Qa.FP!�����[�.��J�,5�'K��/���`��y��t;U�f9d����J3������]�#
xZ��w!��6��>4X��m��A%f�C+5��A�_�1�׶�b�����M8��v���I1L���LEW�A� GF��
��ba�����,u�El�]0@�y@�/d6� 0�*z��-�ݢ�����k�m�j�K�D7�6����IǠ�$�B�>��<~}n0�����共_��c�$��sY�Ùc�fn@u��|����$��ٍ�Y�޵�wm2eLx��@2���*	��u��ʅ̳���5����8�̇#�� ��T���8�!��������J�|���������
 �2\ۆ8�R�$X��u��3��%D��{D�D>P�b�l~op�{�.��P�	g)�-�(��TAu��Ҿ���sU�!���P��YE��+��59�mq���IZ^?��3Fc*da"}p���Q,
����U��]�p���[I4���\1�q�����ӽ���yH������Z�(�2��Db�ն�TI�io�od���G�9����Z�m����:>2	M7"�KlF���l�xQM��jTQ_{a�$IB#C���=q��e܆K(^`䔛sP�>��aKl�_���%�V��N�{��w2L5�������e:>/ѫ�Hk�6+��a����n�$��wԯ�fKrd�o,�r�O�r
`R���X��w��s����_���7��%^ �Vq�������
6��WDW���`�$�Z��!87�k|>���!W��r&=Y��S6Oc::�'ѧ���ݵ0(?3|X;���i�&E��:C��NC�8f���!�s���0�ܖ����:��0:�V\�� y�|����޽�G\�L�܆���Y^������,=r�7S7�+����"�m��M����w��i�������t�h#�m���*���/�n�����}�����a�3�o^�.��4�{��v��~�M��`C���1����wU�9�Yu)�'On�i��v����p���5tf*(NW:	<t!7~��-�T|D��]8���̋�O�o>_eDoC8�X+��<P�����m-y�:f�؄��};�����ʣqNb�dy�:�Ewݯ�cc�1�6=�ܬse�(s��y!���u�[����;s#��v�UQP	�5Zb^F��u�U�>,k틩���^�a�OE�H0I=�޹�ENѻ�S��[��5�H�֗h�I)�xJ��.�Ȅ��u��dl?���j|�\��@V��cɜ�ф�;o�]Ѿ��t�?�������%
��t������q��i9�y{zq^��WG�1ƜG[*C����p/u@�%(�;��������I��U	�V�}�]�c������h#��i\�wqγ�ތ ��BT����7���`�4<c~��E0�X��������g����~�9�����nO�r�*�2U�]MB"f�P�S ��Pq/�B��e��m2����'n�������mp	o��B���ZUD�(�[��_.�W�����&�8M���%�Ɍ{m
��(�Z7�)�v	���|1T����nJ���W��aķ�t1k�&�)8��38��������[�9�ѡ�dg»��G"6EC����?�ev(���A�'G����D�l-�^)5"��d	�����Q�����.&�=�{�Wt�<��tB8��CD���E[HX_jZ�Eli�xa_�����w~j+�C02����4�����<�`oV��*Q��7r�w1�A�[,I~B�����Qfn9�e{��#V]	O��;�2~�5��S��>��W����O�M���xa����\�!^� ѠY&b47��_����!),�;�B����H�����Ø�y\g]��$��#�I"s@ �s,�E3t����1�Dx#Hw�k���z����ч��f��h�$+�SSD_���.�w�!ĿI:�y�p�͛	�F]�f�].�~	*�>�,NJ>�'��v��;)mWo��H���G4�b����/Or�>�� �I�b�t8w ��a;U�HF	3��%}��@�������aj�̌Ռ7�<�d����9y�x��Y��2��^��9��y�4�.|6	�OX,(��6�`��X*+�PR��6�[���	��i��>��w���o���@ ��m����>F��Ħ;�g�,=��$k��QA%��JI^!��Pw�lv���h��ʯ��4M��1������������=���"��,?B��������Et^���:M���X���W����F�0�6��.�T]�^
�ޛE?�b�t�0˙��n��1���4��8Ϳ؆��q߁f��-i����$I����#w/م�I��f���V�I+��{`�|�z���kHDm�avZ�ȬaP��J
���� k��+�^��Wvi��Kr��꬘�O�lHr�ok@2���s�3�y�� �8ڍ��WG��o@�� �CpNC ���Y��Y�h��[\^`��s�����ğ�?��$�.�PmR�9F����~R"*AbU�����]I,zh!��*���w��`��2�T�d�𕈐V��#���)�L"Rs���7B ����~!���^�nx�(�Y�J�ֿ��Z=���n���~
l���5C��']z��u�ŝ}����i(W6x�\,��Ɏ�=~���&7O�c�FIX���"Ǔ��k�`bg�p����ݬ�75H�p���bs�b��;�[����;͙ڣ_;�L�Y.���� up@��_4�bY��lՁJ�u%�S;����"g�3�����y/�k���e�(�!Uc�9�I�PU2F$1"���,��n�[�WO~" �E�f����D�\Y�wypOR��{��kb `W�X&+��5������������2]-5��7� !��o�f��t!�	���P�|Z��Y���U��6V�R�����j2�ڑP���(c���>g#�>����q�3-Q+b�
S牘J��(���Vhӧ�3�����ye*���~m��=��܆�U`��/ؕ��`h~���q�%������?>�әb��4IF��F`������Y4cE�6�F�yL��̞Fo�����qN��#�O�6�l����;9�O��8Z�����8|�x_y�3}6����2&����:J0/�\��:i5��_3-�N��	���]�v'Y;�}1��c��{��t��C!@Sx��t�;L����_��$2�ɣ]-�x1F�3��Ȼ��K����Z���N;�Ka�Q�n�$3�ۙ�̗�۪�9�a�z��fM5��z����c�#lG�˪UX�Z;�he�J�o��v1�s��^Z��E>$����/F�*M� iR�?#�_��� (7�iD��U�@�Ͱh���m�6L<������HH���S�?�ϖe��� [�ǜ�^옣��mM}L��,�+� ��d���l�W��qor��B�V�_u'Q��&]���$��ǁ��h��녮��(d�oj;�2�^M� QE�9�@����Q!B��+�i	1��C�C;� �Z)��s2g�X��tMm��E��p���zV����/�jM?*Gr�Xx�"���b�Eǔ��e�w�2"�0ܬ�=��c��,�z��� ��$�z��B7:�v�A�$B('~O9��Y�*��G������A�!��߫��G���)��B�:
�!���;�޵ݫ�� �[**�o�����`If�'��7,]](|_���4nUa�-�0xVR3��葛Rw��"c��N@�oeM���<� �x��jH;ػ^����~�#��~���ٲ��d��5xm;Рg|���A&e���_g�2!�y�J#V��]�g��,����=ճ�����V(N ��֟�iԤ�6����(�(����Z48��]4�h�ǹ���Q1��cV��j�V�I��W:2�Wޕ>�X�����@��'Q�5(ܥ�4��P7�z�(k����6�K����N��Ex<��o�APmb�pϷ�	c�V��p�øO�5�\i����ps̭#�R�u[�r#��ͷv��m���0�&se����G+X�6��-%���h��{O6|��� v�C~�2�>ky�J�TS&D�N䜝���������0DN7����9���$i��!�奫�/>�R>�(U�򷳿��c�؛I����uT��?�%��Z�2���<�m����qv�����4� 6���;{H��*��'�Z��9��1��\]�2���mE�B���T����	�_į�L� V��B�纵�̲,���OШ�Zah���B��QR� ��Ʈil���O~;�"�3=+hꭲ�2I����OƸf������z��Rǚ٨���?p��n<��24u��W�JB��c�?��3�"mO���EO�{��|�J���K�9BUmT���f��s(������(+m��E��-)'���kj n�&98������+a@��):q@�eac����@>�����=�U���q���x��zA�=D*̘k���k*/�Iy6��h.�*H�BK-g�����޺fL�q�E��:�(�N`��τ�'h"�׳�D��4	�&
'�g}�H�#]�ʜ�/:~{��p�2�1jda�U����Ufz��K?�ҬN���X��Sk���m������5{<,X.�nE��;�Q���G��ĩO��w> m�_?�d�:��sH9y��e�D
�t̘�G9O�]Kqɓ�--�e�c0#��L���%��B�Nd�ΎP0�%�w��գ��g]6B�ǘO���Q�l'�����"�*zC��*'Er	�$������.���HKJ�,4�2�%:��p2�Z�;��d��`�)�����8Oj��hwnF�.�h(�ߌ�WԶ Z^v�>l��.�T�F��/��
*�i�t�!��A��ۦ*�3\"�XT�A_��9y�+���AJ��a.I�Y�C
�ĥDy�K@�%��
����0��ySy��_��*qg��'A�m����v��H��r�����)��U�|Xm�x� �\+�߷j��`s�3�➯nZ�t?�D�"�Y�Dg1<��&�{������s@��6�:!^�����!a���b����6K%�{'� }a�2�����l5����I*DBKMl����/���` �a��'$z�T0�S��yV�������Td��V�\򓛓'Npa�X�!+=4���5�C���~��b�I���c
�,J�H7s&E������<������3|�.���o���ƀb��]C�4C�{O�a�L�2����+jq�e��E����ѿ� ��ı�]���� ��h�&��'>���l�����?�֊�hʽ�X�YSKɦ����Q³���U���Sa�F���J�j7/�O�V��E��Xx ��wDOl(������Z�>%${-����h��%>�5)}�h�@�R�����d��l鉴�c���]��ƭ_Q�@�-B�^�ko8�h�Tِ������7A�*��IC̑
��˼ю���;)oY�r��}�O�\�5�m��:�Fr�k3������݊���\��OVΜL��E�}�J3���r_��A�a��q�X�y��������*]���S6&����q���ϑ���}��6pP�>R���S��:M!��=���r�ƏA�.b���J�vƀЁ��>E�Oܡ���:�eN�+���2����� r|b2�(�O�-�0\zv���������K�Y�KA_'{p����;������H?�.=ĸ_b8���g&�Jċ>���z��S���^#��/4�bu��� �]�S�:<���h�F�'�U��F�|��gc(��{궿9�����.���Vi�cZ�oK�R����㮎/"l��s��{z���9��XN<\)  !dq[~�s���_����i�W�e9tߋD�s�q,�K����	e����@G����6{�JX<���j��r�+M�x��xls����͢�����I�fV
��/eX�6BH.B�p��l��A�EA���+���t���uͰ�$Lr�Ön��Sm�J�ڻZ��/Ǿ��q�14���w�2�ԙ�m�:RdfP�ݑ�r��`ڡ�D%ZE:r� f���� fH� ʄ��#N9�d�Զջ��ؓ�Q6i����� p�� 4��+@Y\�ش)�J9�h��v7��
��y�(�� ֦�w�/v �p0/�T"��Z
]�n��rc�����]��gXp�\>��y�B�]ۋ��|h4�	/ԆGg��;��75�3��Af��
�:�e|�q��~jg��#�v/�acsS.o2K�j$�2�{�ˏP�op�l���h�*hW|t�L�X!�b�=))��I�m�+J�f95!�W�,���*땖�-)�V�����A��o+b�,M�M��I���\}����9j{��A��,bi_U�Mm��l����9���~�K3#Ce�T1�;c=P���3�']SK���x���hdW�\���څ�D�}T3���x�gX[��L�)��z�S�xHb�^Nm�����@\^^E-M�hD��k�N1���X1B,b-�
�;?I�!����×���gV�cr��8����D��U~�55����bj�h��={�l3R (d֪<�c�ܮh}�9��1���O�y��c��Hz�ԬQ^)H�mr�9(q�1�{ ݳ9�;z�V�i.[Y�T������l_i��� t�E"��<��pK��o����f��	n��:���f��'����"���	
WOw�2}��K����+���hZ�x� [؎�.l�Ŀ�ǡ(d��ލ8�� 2A�R�9�:��H��F�8:�a)E�Z��:�O��t�s*��Su��P3�Q2\�T���-2��8��FN�ı{�d}�F���*�����h2��T�E��vd�kN\l��
0@Z��7-�J,��8(�����+!MJ���AG��9�9���~��ޅ�Y1%�9fF4�iOD�Ya��ߘ��~�"R+t���E��Z*�!⓫td�>���d��|;�][����E���x>=^�[)�U���aU�7$��KJ���4�~�Tp���G�Wl�%R"T\O��dn�����i+�/y�<���S&� �a*ɜ�*x^��9���m9=8J��Y��}+��^�Wı�5K	�w@60��s�a�|Q���	�~$V��n%L��Gx���\�5o�	��{p�`���<�����g(�CX�d����*�_
�ϛ78u;��i8��L�Z����>\��2�~�h���Iw������D�<_�\�O�O��4R��̐��v�����v�<��v��Q^[���]6/)���c����8s�)bA�W��"p�$*	F	}��d	߂���鸁�$��'R@Ds�l��p<�i�֗�_�Q�t��/ $u0�X"�rnZ�O+�����:WI	��{sO(�|E���}2_î��\���<���]Y�W���&_\��o.�,�郟�a�A�B�<T7���eNF��3�7wK�J������|H����O�noɡ�a���-@ys��,�o�4�_����S�qc7�A�~>p�v���{���d�.�,�i4ir�Q��#*��'򥊟Gx*`�47�hR/��h�4�����k���v��z��f�H��O���]�2u��_����l����R��G�#��@b���P��΀��;�a#�]�3�����-ͭt�;)C⎡P6�9�"�c��e� �c*��JQ�XeGV0Sm,��ßE���	MW�%(�ܬx�[x�m��,eJ>��y~�+��Fg�G��ө���j��a�+T�16�K�7Pt��d	��E��3!U�!%�;��_;?`���F��N�f�����E�Y@~%��k��J"�ԑ�upG̀wum�Ǣ8Oy }�ل��^ViO:@e�P�֊/���q���$]VV�J!\�Q������2�{�@?��h�<W�\�͈8z_CAz�
|��.�����qE��EL���%K�:iR��м���رX½�h��1B��b:T��s�kH��/�������*Уu|��P�Y̩�����=:ݾf�b�.@q߿�p8G��#�K��xU��_A>$����c�M�rw�m�ƅ���[���(%X���h}̎�"��3;�a0�Ils�t��r��ZHCH$�Q0�%��5Z�$c��V�f�ͅ�j����"t`P�'���*{--�Vjh��w�H��
@U�RzVT%2�H��4J rp�P5� ��4�.���o���m���1]R������Ub�a��O��*�j7��2:,�kj��J�5��X)����XfJr��d-��?�����w��a��$�����[�b>��u�!�OND��J��%B���S�#�����J���a�"C��yq� ���f��puܵ.r�y�V�����%��`E�(YC�J�9l�1F`�W�ad�sU�U��ˑw79�5(�7��ID��*�������n!�q�� �><$Ĥޯ�i[�+����KU(v��$��RM�aj�~X��|��]ʹ�q@�0jLX ��~��kf 8]_��1m^�-��b�����j`�Is�7گ�bo#���)VM0�����J5vߧ�`!��7�����!�g���J�-#Ԑ�E�l����z<����\`�������b��*�A� ��F�/4�·�	��a�&�O��}���[尬�N(KW�AA���K�c:��7U���{*�E�ix|�|uv3�N�u(@���|{g�x��
0n�a�∞~8�c�W��:��de���${��+�}I��d�a��|�#����=DH��*ꎇzu	 ����b�Dm9y��y��G���P:QԖv�@���C�969:�2/�t9���ɭv�y��ܝ懖RR1���"��.� 0�cC��t��R�-��"G���+&�FAA���æ�uU�"�Z�yASP�qJ\�xuo��Ӏ
���C�h���IpD��@I��J 4�Bv����q?z��͘x��c�q�Z-(T�ق)�_�$��9�3�a̫�c�^'ŧ��q���ag���o.���Q?@�{��#8����xevTu�0v�#�oL�wը_f.�~,wf�W�̃J��wj����[�#,3���&�f44��|�}���W�d]�|�7�{�.RĢ�� [�����=Fz�s����G0�
�*�q�@=�)�{dWqm�&Y�h!���8ña��*��U����gv��nV�k���	�:<)׳�o/k�S�H�FtU�.D�)����ϩ.��9�F�7 劄kfŊ��MS2,]j��5�8`�v��l�H7�EBCySZ|��(�2[>�^��@�>{VQP��>tr�?�>x��N�>�=t�-l��a d�t�rs���0�/��j�ΈOʘ�Č��c�h�_�Q�^˒�
�	vn�mN�P�Le�a/ǆd��g�	�d;��(N��+=GN�z�g�8B����B٤�O9�I�?��I#څ�����{�H/�'+�8�5w�D���2�����ғ/�,H�wg�������a(nf��(ʸ�9�w��D�/��lz�"�z�	*�5�?@�K�Z�����Hf,ߖP���q:�����9dc'�˦����J��4����m�8�Te'<bߖ�0�?\�u�%E[�
� ڵ�z��+
�1&y;�.EM.2��g-���}��in�w�V|Ks�i�Y�
�f���h�c{�4�j����һM�x�f˯i��f�a��~�8+d�N�.�p+D��/�����C6O��O���es=��]�ξZ���w����	�����A�J�σb��w����>��v�b9�IkZ��l(|�R�{��9ͷh�2̊�b�5N���Q�o�x^�kL
�,�c�J����@�{K̹��u `�0���z�(�P�ؙ�xo���՘~:���h�uM~a	%>�rЁ�FO�m��4�J�*tbJ�]S��N�ݒ~O��ml���/����߷Ȋ^s�ShU�kͩ%��߾�t���9�D�Uޝ����a���m>t[����ᨷC�Ӵc#6��1������^��~���ف"���{��k�8Ue�z�V�G ;s�Z{�7'�p�����(L
g`��ٺ��j�ت0l� ��>1�6��-mdv���{�����Y7
 ��)��s3��V���j6�����䞈n�󓠩�f���?Ш�cX��)A���J�S9��(�m��v����C�1�N��۝�EGaK��	��W���䟩4Y*����ä�".P�$�RY�V:'�c��Y�1>Α_/�ˊu EK)��iC��w�fN���)=Z-���yԴ��f8՝R���&��}[2>j�d��2Eb��y�I��X?n��5�TM�̄sC��Íg�⯲=x(�a��f|��,���l��L��H'm�O�@Ty��Z��'�����%��ڕ,�h��.�Z�6�C¼�.�WZ::!����	%�wI⢿�_���%�h��� �u&:��ōT�չ/z�$����w�1��V$/:12��r�4wAX���o.F�T���@4t�wR��+�$�dB	%�mgӋ�3
˸�l�A+Pŵ�K���oK&<��n������sm��r�C��	��W�x��=�a�eU5���"kG���j>�;����U�2��uD$��;Y��;�ڼ�w�t�ƫ#g�0"��qn�����ױN!����w�?�ߪ�z��Gt=� j((?��y���g�V�ڬ
��[:��*�]oj�,�}�B�����\�"�`�j�H� ���lnݻ�v��M��e�.&@�!2���8]d(giqi����$ iJ�J����������qYJ3�o���BP:�7�������M'�Q� J�����¢-���Of�{�+'�����ZQ�27� �Ј����Qd��=�"����/ �Z�&����
�Ӷ��@��iY7�0�<8����?����UL�/Q4�/�	���爫oJ���< �>q��h��;E ���2�q,���� �:+X��i�СR���
�쵔م�PB��fs�+ z(S�_<i�q�J�D��yY	�4kN)�q�`�K��Ƃ���rHS��h���ݠ[B<A�%R�9Q�V�1/u�����I�]�Q��V�Dr�5���[M$B�A�b�#�x�V��� ���6H�4<��C䶘�ǜ���n�`��I���0q:�\?1�'�����%�e�v/=�&��)�*^�vB�.�ZYiq�IdD�>����Y&��A�3wq>g@���L���K��W;,�|� ��;�Qvb���N��tI>�	aທF�`��MziX%�Wԅ8N��])��kL1�֖�vzvL�Kgֈ�}~�����\�!��0�����a?M��FLV���ȭ��V��R�(�*�N��f|�.�`x��
���$f��5�Y��Y&h�9�N��5G�:d!D*M<(-�ى#E�s[���&G�:jFzs�&����nw���F�[w���8^��6���n�q��V�(0�4i����Q��E͐�A���ZRkLu%ߔ98�P����+�p�LhD��N=�2f� �)���(���I�(����A�	�AY_\����G��ᴰ�]�S����e6P���U�N�޻DF@WIt�x�!���5�F�������h0�JV�q�������^Ӣ�b��N�1�%S�B�J~L޼"���Q�b�?�l� ����!���cVd ��/PJ��A(�H�A�#�:�}6�W�=w���ב�Ok�d-����7]��Ұ~.�^�L�;�yځ�L�#ҏf��4�a��4�s�_^�z��e:�3����j\(_�J@��e�H��u�p��$A�`f��I���D�C/�e�G���n���������Mt']��A({2�c�Wu4�jE�w�x��)_km[��]�4�T�Ӭ7��H��lJ;i��m��Ѡ^���E�1Q�[��P��s�:���ޢ�k3��~�֔���%!D)`�\�;c��W��M=ۃߴV���p�ٿ$�	*�b������bi����!���6��X�ړ�ڪ͸@�ZgmakB�r�B*� #
y-F����8�L9|��c�4�I���c��K*1Yp�fՙ/�̞!DPoh.}~Bk�	�1	�� G��2��r���Τ�񚮥�ɯ\�{Q���I���"��f��ގ�@T��Qh�틤�|�P?7����Ox��%:���]�H�T�щ
����T��ʕ�/yky�ȳ��f�~H6����$�ϢlZ1�_ׄXEE��i�;5�]DT�vn���x ��<y�+O:���$�2+������Y�B"\^�S��}PD�1�w�Nfي�>�Vn;/IH��3$~�Lf�� �ʉ����"/Tl����C@��~6fPMU����A�]�dܩ)��I�5׃b_֮��ե�*��u�$���7��]�A�����/0�'Țأ�he<?��^�&<ux�އQ�d��n:���f�J�6Bj�����~_�I�w��#C{�X�]u�iHi� ȧ��#�Q�QoiL� �$�Y�F���\L<��1�e7O#��BNJk���yq8���n��ǿK(l^}�fRW�(�`�v��hQ\�4��Z���1�4e>=vdi	���ZU��Ĳ�>TO��Hu���V+'��W.�癄��٧C�7NK-�.�����k|��ٵ\v[$�{���J)���g��{#�<,�c{�z	T����o�b�������j�=ֶ����U;�V�nB@�٠��i�x8W��0=V�q8����?��\�M�ɢ�3��W� ,j�k(�����D��s�nU�C�ɟ�;���-)�U	U�t�����L���io�a#��剼���=��A;Z��o��.�:W���ﳴ!<&q�����`tp����Ŵ�9	=�Z���m���Q`ȆL"��Je���o�e gx�8>_�vZ��W������o1}4��Ή������#Ɨ����Ӡ��s!$���T�v�#9<:>~������������q�(x�I��)�p�P]0�$�1nv��F��B��9���8dR��E�:H����Q*e_T��b5�O$�-
�����*�:������%���f��[�!�oB�@k_�l�� +�T�N~/F⅐��2���,8w�[�����be��y�Tj�	�澥�������+�T�m���A�͟/'X�C�(�H	9"���y�8��bhn<�ݡ���s�����x�EW�G����)�	w�g��]) �)J9���\)�;WP-������xt�E�v[�c{�VxNW��_3Ӻ*93�>(I��
�2K?�
+�=`HrQ8��M3�[v>Y��؍\j8�Z��ۄ���J�����):�y�j$ޖ����zykx�)E咅Ӈ�	]i.�ЊIl�l�;M��5M�2��a����^�oE��t����1_������:f�A�'1�iZ�S
_Z�E���aP�u;�i�O� �}4ը�m�ML���D�wy�V���]2"7H��Y"!Ske9>�&��+p�y�BG\Ǭ�>��[��~��'P\N��l�?���B��V��, �m�v�9�MCO�U��nMB�#�h�?(�Ƀ�-֖�:Z��$��#� �kW����R�XN�a���bw��#x=T�c=�B�˞v��Ӧq�`ƴ���E��n���1S\];Q��Ly�����؛y���Ar �I��+��F���T�cЂ���ji�7d��֬��e|��۔d?�\9��q��ɡ� h%>O�����Z�T��w���O_)�g������ꉷ�'w����
���b��<:���[�(��m������i�������H�?����G�Ϲ6}�I�u��j��J��4`M ���t���~p`e��[�u�
q[���0��4�-e�J��\��P����yan�.g�K�ȋX��tԖ~B��gJ')�C�Q~{d% %SŽT�VD�e���B����4�^�b�7����)�Syu�r�2�?��
��D =�a �`8�1_��ա�7�o+&�`((G�e)�sV��u/��Z�K0��
}���m�j�R'`WUlx~G���G�p3p@�-?���7������x3���U�Qh�؞��Ǽ��Z n_@U@�QO(I���q.xS�*��
���7�q�.��4�`�Ǻ���	�#UU �鈝�����5b���@�'���-����E�H#��{"2���JI�ad�(Ne�����.���Z�a�����g���Z���m��P ��6G�2�u5�`�V)tM�+%I)�q	�	�nA�����#�C_��x�0���X��$Ӌp��ߗ?���xK3�R�h"#P��{�j���9Z�+*�(C���Ϣ̩_�Ȳ��ijI֍�`0g{� Xù�\s^��RXYVވ��H��~㥕W��u����>��U#�$Tid\�n+�:>��j�g�:b���f�5���?�n@��Z?�����Rx81.ԹGe�eّc���2�&�TiN$��>�ݏI�G���ΞAiCOe#,���PZh!��Ք~��.�5/ْ.��*Uh���cXcy̊a%�(ݷ�۬�W8��.-�� �%�U�W�
1C�j��I�a�z��3��~P�ܬ]�� ڳ`�_d�KVD�VP��rݘ� ���hr=Za%�zs�r{s5XQ-b=!:?>$s���������*�[����`Yt�}�3}��e�N�����Ƀ&pn���%����}e��|�V��T�����$MI�VF�oP�ҕ!��2:h�����R�('	Л��`32�aM@��Ǧ*���#�N�j��=�񘿐��Y'�ܓ��z���3�p�4�G���s�����uD�����w����AZd�ONoV��+%�B$����9g8����|�pJ�x�4]D9��6��կ_�$��} ���x�-	��δ����������~��ցmF&���A��.Yf>���/�sY��Ru�`u)^�aѷ��������g���؎�rkd�1�ۯ}\�~S	!o `�	NJ	�"'5׻3�9���� nȺ.d\\"2��Oc�p�+;�h�����>�=KH�$Kϓw0F}	r��������B#�*��;����_�|E:���zu%�l���T���:�Lܩvu�oZ#޽1��gl	Y\�Sp�ju�(����I��ʋ�~����5!�E�/ZrPY-�B�U{�+T��k�F�͂����L-{�Ch�+j5������=J&�5�=���g*��_�1N�ˇ� �1�2u��u��D8�{��AZ��OM�=*�z��O���ݤ�)3_�=(��Z� �#J8.w�4:����Ŷ�z�w�j#]Dxf��U��+�S������{M$�Y��`���zr�r9�6��q,�.�r_�%'"6=O�p��A<jۦ�$����
�.�D�J�D�i�P���>��8O8JF`�m�5���c(� R��! ���t��	���b��x��`�}����ׄ�ӗM܄~��,���f�L�!	�5��F_W�B��E�B#�곿����S�˃F�L qs��F�wGv5����:�R\�"��
�G*!D��n�3O�~���~�W�P�qc,]=~��z4�Z��X���{%1�Ё/���>���F���$�)C�[�fd�i]�<��T#p�'Iv�����3[��T��m͒���/E5��T�:�;o��(�����gF=�s�G)ɮq>�(�"���e����GTk$�1!<�ۨ�^MS蕱z�s�� xO��p�(�O�\���ț�_�{�Pa��,3P8������a2�{�ŤEx��R�;����{�W�ؔYN�V$l��N��X�2�$�����n�

S����jP�1�Zw��E�o�K�ՋPм"Up)�]6�ҙ"+7���G�%��ϰ}N����hl�~K��x]�V�9"�&pݨ��K9fd�� �L}'i����p0Xf��WYX-'�����i�Xْ���[�$���N{�ݟ�\)�veL4�v`(�!��ҵ��C�(r�ٜ\}�_қ�o�s a���7X^ܗ��@X�m�e�Ji\ӈ����^�2m=8�/$�dv�Fl�/)�ǯ�?ff3,�߇@�7"*�[���1P[�?�cR�>��V<j��]����T�ȴ�D]3#ۯ'/����A����.�v�/8�R�4��xh��U褔~��7����R��.�{�&�~S@w.S�L��`����,��=ɐ�ֿY�����Y
�@lI^M�<���e�[�o�5��B T��ɽ�~P�!2t�ye��:Tw��:�u��Cf:��f4���f�+{�ױ��؇�J{sߙ����V�^8�M<�8W�P1�7 �!ɯ��U˓��L�z�����S%��̕6�֧Lg�
��>G格QCc��$�5�����=:�i18ǶP����s�MӜ��\/$}'��ٳ���
ی�9�����)�����Z�ϴA�t:�Z��S�\C�?��Q��F�,�An
�r�ר������^qC!�-��Й�+��mO�:=��߯_	���`���#�w��!�<����9t�1�I�A$��h���$�wV��W\����c�)U(G��?��[���?c��W\[4KP�_�E��!��<Fj���D�7�w՛NO�|��
���hӫ��Ļ��"�a���ǂ��U
��:�֪��D��g��<rJI'u�`�6��@{�������\h�3��znQ�ΰ�sjp�O�׬�6����-�U!9Z;9YD.��{2�LͱQKH�X=װ)r�7>�&xi�tΦ+h��=oMz���F��ig;}��w�����P��L���C3ñE�7���B����0*Z&X�%��u39ЍհǱ�T;����/����q�v%w���_�
/�K2�M=�2`�6� -A[ȼ������x<��V��n����r+��Û�LĨ)G�B���Z1#����=�^��h�y�-�jv���%c)����f��IC	\��X���/�jd;��C�4Z�x�g?�U��^�ξ��d=ݦˮ�h�$<��` �]Y�H����ɂ7��&M�`�wbz�A�V�AY��?���Ad����B��
\X�)�a��Au��;	I�KT�����ܞ��9��#�^g/a�����*y�����&�)� N�h]&�>l�Ì.�N��"۞�%��s���S��T?����RRs��V� ��V�����8�k�N�ۥ�"����M�j��ED�~�
�޺l۾��=�ť��h98ڰ�4��"0q?�4[?���q��/m2�� ����� �\�53TJ�ש������;��G5ʓ�[��+!C���b����>J��ܮB%Og��z"�s"�}��$J�D�+o ��F��n>���iv�����&��ֻ{:��݊xޞW:������{�X,"��˨ @$����Xi�"V��k9T������3�(��U���"��d�Ǉ�`ɪm!�j5�"+�*�U�T��]� =Ob�������L�EO��_j��Qi�J<� <؁�j�<Rї�S�<��!�F�cN�3c�,�n�J�z3�W>���"���4�V��L�`�C$�0�ꛢPL����E�1��b�GMS82�����K�a����]%������ʘ[��ښ_:6H(�]a�Vh{�{�')�A
 `qt�l���S�0��W�p��|1�Hn��/qQ"��%��}լ@�ʡ�g̖ؗ���,�����Sk���C:�����Fd���Ӂ�0Q�r�����qB����@�Ҟ�F^�X�g.��f�7B`4~���Z"���j=��'�=OM�w(��`��^d�ǐ@F��Jsk6�r}E�6�|W����m(�^���v�|����a<��U�k�ʭ�t#ȷ�j���۽��w���H��hJ`�<�>b�	L�lG2�����.Л�&Q�G��o�;���V�%>�"	x,����K/�� ��_]���Gh`΄�^�����$;o휪8́��3��ԟ������Z�w!I�^�wV@��®G�OM���0�)%���6�X��NC
��哄R<i;D?9a-�����!�\��W��~,�����2���MBXT`5"������hz���v�dg���A`�xY�]ʌɗ��S��Q4J���8�JW��� �Ư���X��pg�E�/JETh��I��\2���+�t�c��I9SS�:�T^b��g�G�ۢ>�s扮G�=�Ͳ��"�$5m���W�|։gX���W
Vd�)>U�gM
T�%5��#�I�?��SQ��m@�&?C�7V��x��I�D�G��J?H`�Ρ�]��H���pwG�S��^��������!���[�����z���%����i���d���_b���F]��6j� *�����/j�R*t~�Wi�^Y�qw@�G۠��Ѯ�^�>~�����
��<�H�4�tA.�ԡ=42�����IlR��[[0����cl#!��|k濝����)�RhU��A8�Ϸ!n�,*AU�%Vl�`U-vc4��>��<��Y��'M(�ʐ�2����Qj�>fכ��:>�vّZ%�W��[t�O�Q� rN=F��R�<�K���>�;���Py��9#!.ś?u2,�q)��h�#E��{ '�̰v�̽7C�.n�EX�6LG�6p.R$�du�:�K���U�!%�&J����iuX��w��) �Iܫ+�[�$�U:��q�Bjh_R����8��95�
����؋	2����:8rw���8���~�X�kHB����O��(^�x�->|4.ڻ	����!?�k�c�[�
Q�w���s�O7�������$Tl��'Sʖ��X?�ڐ����0F�`3Sk�&FQ�>�|�~��4��j�&���!3��V���O����/}5c�����#��5_�HB!�A��wÔ�H�[��NKo�@c�H�����ZB�V{�8&ӛ*"�(�s��YKE���{+CA#�Ś8��]�b` �&��WQU�F��D����Y����?x��[{
�ƞ�;�f=:0�&CV���Sp�C��a�L�-��O�7cl�<�(4�Z	�*��PVLQ�����L��l4V��V��`�Bk���ڥK�����h�H�{e�OG�떴����uz!��ݕ��A��Il�^4��`R�V�EL��O��%s������;��g�w�v�mR��8:��yȔ1U��~�:^����l�+{���'+:V��;h�Yl�MP�=x1n���}���*�Ur�^�)th<�Bȸ��yi6�Y)V�Eq96�?6Z�� �x~����,�XK7X��9���anu�F#�sW��A˝cB�Ht�s��]���d�u����H�8��J���$`%�tl����(�a���>71��s�դ�+<K ��v�L ����
�60�#jm\A7jF+x����f��>Y�N�N¯:�PF��_���$�_(?�+��Uۑc�>g��_l���.��m
<�b�)_#ܐ]� (������`��ide��D�Œ�� ]0�����u��.��`$�o+=�D��A�f�Uz� ��nMU,H��Y>y��@v�X����-!Λ��֒2�%u'�-�t�mL���@�M���e��^�d�uA�J�@>{���0Y���Ε��f3Q�p]q*�g���<C�P_�X��Pv��	��y����F(J���wD�{��}%�v�u%��T��y��na�H���
�^L@�X�f����P�H6 �=�G���ɺL �>T}�l ���'}���;|��S�n��dl&"Y�9����X�|q��;2�W�z��ϼ��a,��`� C�7�9��x�Tc��%����o���s�D���+���\�r:��Ϙ�w֣��E	?z9��g���2+�������|���YtC�Ҫ>����^)�$�]�f�2Nb> ����oFY���L2W�Ү����f[r����MzW	v��{���rC����*���r�R곖����C8�:̀����-�OD+Ik2��s�hL�V�Ka��*O씐:b��;`��!��`��h��y銟ρ���KJ9�D�6�0 kM��WMji���z�t���_�o]6"�x]�_n���D�+AVf('H�kr�Fy���@�� �@�\E�͙GY��/�"�x�~��H�N�i����K�^E�}�*D�������"���j�����r�D|��&}<����[�˭�b^�,�$�b��<�n�B�	S3� ý�x�����Tz8�,@������Z��P�]�K�C'�^�6�"?�*��ݖ���$`�|9�sT��
���4C|J�T�KM��Q�i���z�Nw��&8�����Ry�	m�2�!$xQ��
��f���L��o��`�@h��~�B��C+��Ρ�����fs��\�C/͈ƀ��A4y�*��I�����%�j�N��G"h�:R�?��.�m��S�B�aO���Г�����vA| ���QM	{�5�r�~O�_u�������e]m'P��k����?ɲ�1?��چ��R��"�����2Eo���-�j>�N��"���8�r�?B�����7�B�B���ހi�R�bˊӍ9�䍩W�Vmh�G0�A��m8Xu�`=;Ok.���W�_�"K��$��`�F�&Ǹ+����ﻟ�Z�{�O4[�b�wg�a��͜�_�_ڨ�ٸ:2���Y�J��d"����3��.HsܩZ��Ev�B��=��_��k�,��(q:xT�����(�*≅s�<YO��k��,��f �`l�'�i����k�1�
~*�Z�ml[��z�iz��,�X����g�/5-i����
J�Я�3i��l���?u�� �H]��^8~[fL�P��xZ&�|x��X��π��k_�9>��<(/o�%r��^ �4�"�>�t�=gEz�_l���30]�ۗ|<�R�9gû8�!���	%��%�޻�G�g+�q;��/�sf�?���A�XN>M !<�G���g
��<����P�^������$t�3v�bK�Z��L΄� mـ^���M����CЪ}<A�x"���5<����
�����7mՙ�q̋t��z��bNJ��0%�����oD�=�'ц� P0������=�~� �t��D9�1S|�X��'#yp ?����o��˧>Yѵ����S�gQp�k�����f���y7-}��g�EX�=րBW9?�P~�c ��^Ɲ�<�
����L.wNV��0[����Ɯc�A�A,M'kqh�͍aJ@\����iQM?�U롧~N�FlZ���C�@��X�ԝ;��Ĳ��i���$ka�A���+j�H�j	\�y���m^EN-�A9����!a��K�G����E�����]#�c>�S�RS�0I��U�o,h{j�"��*���ŕ$<��j�'#�������s|x ����o:�]ꚉ/z��X�`)�q.�����N����Ao���3�^�<b�<<��c��ƤҖ3c�9X��ʄH0��)q�qH��n��6�7��v�F4����$��l:�#��
4�rѽ]����F�kô�iyY0�Ğj��#��*u��VC�����t7�s��?ΏL�B�Hg֊�C���g�AJ:{��~��4ό�Θß��m؋Y��ּ�n�P�!N�;?%�*���~�!P�IM�0S
��i�|��Zz���M��3�����n�Y��3Xc3 ���݌�R�p�N����^66�w����u*��4�X3&�������,to$��8=����C� /6�/�������s�����<x`Tޡ������gl ���)�o(Ш�܌	����ػr~��s-�ϊ��U����Ʃ$�7�����|N�L�q W�$]�U��7����i�%"O̖�VZ]���[|���"~�2��Q����DE�"�yS�ȗ(��p�R�������Jk���2�к�� �T9�9Z,���3x8�Vj�=5���nBa<	,!�A9+ S����3i���W]���}�(�5�8`�=��I{S�S���4�^�B �����`k�J@���V�%go�+z�ϼWE3 [�h4屆~���o����V.����;�2ʞ��0֗7
�vY"`��l����'a�r�t>kH�$W�4c~�k��Q���G�s�sv�S�� 4l5��ln��PY]�8~�U%����'8��A�ugM�L����(�	��JLxA��>�?��e&r5'�1Op�FST�s/��Ui�vU$��k@a�X��_e��3"���!iCW��5��e�����(K�]B,4��J����6O��}߉oTSq�,+Z�X��uw2n'��?�S.�Y�4�>�n{��9��,#p�_L���B�|�d�<A���]G�n�D*�%���˚�S� �0�u��j�����.�7D�����.h�7�r9C^�=�����5�̹�w��?/Ȏ�=�J?��:Xe�.���'�w��1��R��"�~&�z�\����H���W&��,���}����n����b��ʁ���n��ݢ:����L��G�`�BX��[�K�R��J8��4+=A �*�pJwqE�L�n��H������I.��6�U��F�z���a��`@�JP����8_!:��h<VkV{PN�ـ�}�e6�����h�i���]�j�5���ȰPܘ� ���ڳ�$���܇e(mt�fT/�T��Y����Ϧ���v]W��:��x��q�p��2��|�cGW����Q�l	(<�b��(�ϊ@z��|��{����̙reW��%C���O�L|;I_���{_�1������Cd��q+�%�9u�Q��,r%j�PC ��%D�9��Aԡ��GI2qR��C!`��=őB��� 6c�D��YLurD�7)S��x��J��"����8������j���f����y�}�\�\bf� J�0��w���BU�I7 �)<���)!�H�g�mX��)�D��\�A�j���,���5�J4�&A��rs���1>��W8�|�����03�h]��d=�
jڟ�7���6j6����2�3�E����S�}P�2`�Ov=�<�W6@pV�yL�`�z t;��ԫC;����A��c\����6��� ��q����c�Ӕ�K��2�������n���8h*�\]S��+	�"��p32�NiY��Ѩ���?0ʈܳ�)_�n87��A|"\��;b/2�
���./k�ҭ?�4c���9�yKhl-�Ӻ������"�D����:�ܯ��t�wT*U3M�)����G�S��ӊj�F�C[�q�-��~�\OA<��e��	���Nг{�!�f�*�T�U�"�x�;voM����qO�����R(�����|��NYz6���?=�G�:�'��h� u��p`}���*��%6߼�/��f� �H�BS<p����H������n3�n�c/]��&�3 ���X����^?�}��Vg>���E��wfЇ��_��D�H&\]���Tgq��ft�o ~w��8A�b�`l+��
C ��V�1󒨆U'���r���������[��,Y�iy���_�1�@�,)�Y*	t�u�� ��Ó������4�ƥ�9.�@���3Z0��B'\�N�'�d��-��؝R����DR�P�)�O2�MmU���1�0��'gQ��&��>�f�&�e��w��[���l�ƛ��U�}��	%���?p����g�}4 �� À����#mn�3B�Qk61!hx���!��d4��U�.�C␒"��8��X�U�t�I���֎�qt�@wX��s��c�D4$S� t#�5����ك���H��.ˍ�ؗ��t*�e7U�i�cmk.�oh\S�1�a2���*��w�t�!9�F+���~i�`j=�����~�^)G�� �k�/��RV!��F���(�]�yK��YT`5�?p���naK$�v{Fkٵ�l����"�em
	�M6?��B	N
�|H��4�*+���E�[��F�^|��c��e&���,��82_TR�~QyY�����~�^��� �:�;�ٝl]?ϸ�n�b�O$nawX&�������l��U<m(���;+f3�Oh�{�����xe���jy�װ��}w��_��X��Ƙv8id��"�����gV���L5)��<s���$S�/��=++$�y�ZB��:12)3"�US��^���߿Y	����X����7@L��̍'�q�r���g�?��2PMHD�F�S^ԅV B���ɮo�W��gm��pm�:jz����V�_B�L:��� B⩤���ް6r�W�#8��3��%p���"V'+L�)�]>���o��ޫ{��A�,�Ȁ"��}���,�uu?yk3%T&��A/}Nn$go�'9~?r}.���*�'�����>��B1�6.ce� �A|�S������)�b�&+�u�d�0ڐ�(���8����Ip��GQL���})�1��"��c�?�����=`D�E��a�a���d�;lp�������q�$Q�I�e�Hȑ:���Ud�_���"�
�\%=��ԆRh�tt� �p[H�ÛN�Hí�$U�WZ�$�Թdl��
�;���7oc9�ʳEy�30��Œ�r����!,O�ܡx���4cQ�9����uv~�b��}��ú����"�2��u �lGQhн�/6�=X�}���j0AZ���$��a��3Ȝݸ�胗�I�8q���?���˖ů���<�<V�U(�]�ۋ@��3��)����Cc���\�f���o�Zp��8r�,�A`HÈG(��>�-�!�Yd��<T�q��_�G�=�v7�D���M�e��رp�~;L�����T-0�fAtY�Ҧ����V�f��o�w<���}�M�r��?��	�1�,*���N�$|��P�?�xNW��0���1ݺ�?���6|�]&G���v>U?A����ct��_��r�_��Td�����5�b�6#�-+�ٔ����[&M���	e$�r��}�(ڸ�b&���m�(�|����g���McR�քp�p<]ϣRsf���y��Ei$<�N���n��\^�F"�I0���������*�
NO@	N�,�y��Jۭ(�q���9���:/����,(�K2[�͉E�6}m��K�r�tO	Z��kB�FY��r�/����Xc��KbL��5�)�,��>f��'g�wzVV�j<�Jp�G�P��ۡ��Jq2ڵ3�0D>�]�Wq�o����b!'�9�����ƃ��n�4&�� ���ڼ�֔��S�Fɢt��0h����KC�F��mы�G
��7?Y*��E�0�Ѫ���3��΀�?^�;>Ƚ*@��� W�'�)?��Ya�,�-������u��Q�F"3��e�1ޘr������6�o\9�JL8�*���=�]R�#�pή���,�?J����ށKz�+��h\+Wc�+�8~�j�Z�
oep�S�1�h&�B����*��λMve�n�8���}n2{@P�O3uk�g2���E��	L�{ڑ��{�a�����'�p�|K�G�C
_k���{�_��`��j�ob�ZzL�(M��y 5�=u��*�P���:�4���৵��'���e���N7|B�3���6E7y;1��.�7�v��7���r�C�L�,��I�R�\�<�_�)Gw�RȋA!���8j��g>9:�M$X!G�_`s��'Ҋw�K|�$�	4���n��+e���w$0�"6 K�`����3ԙY��Ro(�e�R���?�GEO���"Sr�݃Iˢj�"̐�s9��p���G)�0y�B6�[��V<6M�q4���s�s�{@9~@����D"%��n97��qg�0s _K%8��oG�
q��W���`,9q�y�ۢ�����e�n���_%"TH5�_������ɝm����>v�U�SnU|��p�&V�`4�'D��S�䩃��8�xZ��VY���?,�f���)���]O�
bK��S��[�|O������k�u��v,�!�.]�O��X����lN8��	�"��ї��w��M]v��.���,wwS��(�4���p�iN��ӹLjj�}�7�wiy\�{�:�Mb5 ��j����a��J���L|�n��~�ѣw���Z��*"��om������j4�PL��'�ۈbIa�l�9�[�c�v�ع?p��r���c$Ҭ( �n�)6�����`HIcSP����l�&�����4+s�4��ʳ���rh�a�#��Vqk��P-ʜa�_���g���z	�%Q�m�h��8��є|��t�Z5�X�9��w�?�PV:g�N��E�>?�K� �Fz��L��y�)��Q��c�*����j��K��u���A�9DW�5�l�?%b������i�},�i�D�X`�O�EB҄o�.$Nf����jlT6���o�K��O �˅��zŢH@�o����6��h��~HĽo�R��c'gnmK��eC��'�p�,�s��3Y����6�~� �ek� j
d]���dp
B
âv@S؁�v�">����u��{�z���&��y���+ͫVk����a��Vt����H�wZ�x�&����%Y��15��t�t��@$�{F�U�� ��nzW;����W���B���d@��q�\�j���������
Q3o��w΀�cJ�ȓ��Lt�ԕ���R��'=Ԛ_�d1�����@�g�i����a'H6ۭ����.3Иb�G�<��;��3#S�.y�Jꆎ�"Zo����H#> �l�(V�O��= c�"�?��o�y�\���bau]��}`,.�̻�F.N{�(@Z=�(p�h��!LӌL/gԦ��JӤ�v��T�H��=��Gb��}����.^�6T=p�ZL<�H ��^�!J���+���Rs;o�����;���ێ��5y�	�ow7xDe�������#_��?�v�������KϨN~���n��!�3��.��]��iRk�Nt.3��?1|f2��C��Ӓ~:~��/����rt��u[&a=�,��] |x/�.���ڻ�Ƹ��%G�H�����;Cx�"�r闘Q�w��X=U=�G�f�k,?�A���o'h��	i�Td��D�?ɯ�.-Z�$TmKz��U6ԅ���u��42��e�fY�% U�X/Ϊa��}~�/��#�Iz|_�Tl�OA�]��h�j��S8U*ύ��_<ݥ��6%���yߟꥄ�
s�Z�;j�c���U�Ad).��6da�������d���lUs�f���N�D�ٽ�l~�=��}t /�
��%Ύ��C�����ݤ�]�x�+h�)��WD��g��t�7�)g�q7���v_k�B��.�.� ��ѝh�ol�����v _ncY�pY.�h��i�ds�K�J������R��[��"๞ia�si�%��M�KD�����a�)� ��N�<� j�����u#������y|2����yC�p�rk1�s(��	R���u���B����Ͱ(_�Q�Q_�u���"�N�)�kWy��k���4C6Mq�(_�ߒ���A 6��{�nVA]��%v�����'u���X-(���O�q�u^@6XD����jNX������h?'0�|D=OD>��7kr9�򊪑ܴ����v��噍V� {xC�f�������-W ��")Z�F6 ��]��n��$D=!����"�������sqX�)���Ǣ���|+�#(9E��? Z���5��;������d�l�M�=��ۋ�����ix�8�Ǒ��?��9NT�f<-MU����S�@:���qQ�8��G��g$����K���.u�*�o����$��FKE�b�<ck�K}�!K������Ed3�h(�Z*7ұ�3��aZ��Y����:�3'%��=?s���v6ҿ�1�8���-?iͧK_���)m�pc6*��._a6r��[�ʖ���>:L	w��-d��ךI�JJ�u��ۖ���L�4�����<k�Q7vQ��cj]?+C����q���j���E���8f��AD9����u4� j@f�\R���G��.�p`S
;�(+e�gӋĈ܇�dui�L�md����4v!�z~�R�]�m��@L���6O(r��V=���(O�O��pt{�K�KP7F���K�����w�$�{����,ͼ�)��{p/ �c#�ʹO�&a����k���T Y�!M���bc8<�5p���Q�\�����^��,�ROV8�n�|��.#a������Zc��_쐀�@歀ʅ�Bs�W�e�$6miˉ	�iy�
��U�76}�~z׀���U��������O����M�dh=%ĥ��˝͝;�O��Z��dT�#�0�ߞ���*TDj�:Z��u�P����W?���Cf�BO��3��%v�u�Bןsi��А~��۪���[�{B�ޯ��s=F|����kuD��B�(?�H|�JLK��՞���l�|�U\n��_�l��t��Eă���M�Q��\|�i��c�I��ES��04��1�w������3�5��8Q�\AL'p���-��Hպ��&kI�h���:|�F:<�D��K�����*����D�����͜�+.�ϙ��$\�%�v������,/�Y��L����>��ӝ��y�[���OL���O���T��Ȧ"�i�r��3��Q%ǭ�:�Z#+Cr@yd<����>UC�G�����z�v7#��N�Sj"xŖ�J��w;�������:nw}��_���4��U���S�d>��I|�g��H�~��k֑�M�IU�/�cŗ�����
��(3�<��*��_|��L���7���j�y�X���k���%���f\��eW7(a��m�8`e�+�fL�2�J�I�bBD+����������1p~m�H)��������0���뵕�{5��
x��Z��	~�;,)nH�-d@u���c�Y��B*��5���vE?��:y�v�����[Ǒ�B2D+��#���#�G��H}vG�gZV!:>z�~>�]�e��vr�� ʞ�{k"�D��q{ �`���܂?��� �6j�����c�S��Y�x�؉�tm�blT;���N��ҥ[㙏rA�oU�_�{��G��>3�~���� ����ű�A�Z4R�q��잌n<�	���Cu�v5ya�;'1ஈ5��������Q���s r���B����j�2h3~Ox'd�.~�P���w��.�^�QF�g�P��X���B碡�_+��}Pn4���d+��½B����v�F2��j}���Z_�%�+�'}qr�P� 	�)��?B<	�������{��B;Ó�,���t{��MtR�q��h�F'c��ʶ:��z|��d{m+���7i-�����-*c9�����ި�E-*8pGh�/	_)
m4:j.����,9c ����
�g�3FoD2�S�L��e`0� ��.� d3�/CH���� ������m�W�EaM���?����ঋ6`����p�r�����������2!�@�|7�j���D�e���Fd��_�����@?�	����K�s�2ձ�	b`�gߝKr����L����6�9g�4��r�)���j�:%�8�B�r�!���[�����7����f6E�����a�eO4�1쫙H�N5��_� g�ȓf�NH&&��B�����0� V�ɒ��K���f_�	�l�T!Ԭ�C�=.F-���9n�A9�%�����c^H���v�T��Q�P&�ReZ$��]G�|lzs�0}&?(�רW�P��	V\�����%��s���yc.�;㧚���~�Z�%d���xp极b�B��#�Ջ$W�5J�� �9.�2���zq)UA(�mj�ҍ�,��|�QZ��O�X���91�Naa�
/,|�7�A�~�ˍ�<lᏰ'����?},�I�N"�c.J�ȼ�N�QK�"�5��� o��7*oal\c]~??��,��G@�Hf��~\��q�{��yx.ZFӄ����N�ٟ,��:��v�\G����j>M��}|M�~L��g5��+ya|�!��sA�;p!������A]�m; �.��̺�����o|\wL����}~%����&a<����}�Es���)!O�?fm�N�g���up�{;�8�|+� �̯m�	�fH�bA�4�8:�gn��'4�GR܅����z ^�b[�)1@go��
�W`�x�R�7�����6Q<�ۺ-(�n���I�B�,��p�����N5h��R}M]��c�$����D��li�����U$c�(�z"��G��rI�޺F��J�"�<�f�U��W����7`�΀�P� ��q%�{V���M��͹ɤy���s�^��2�����M�Z���(^#ed.b�?����Ӣ֒#�S&✤���V�Fr�U��e�a>���c���Tcl�U��l�Y�!�Im}�����ER�:�x��������Z���٬�`S���_�fq����J����	C�*�7��ި3�ͺϹ��z��Ҋ���yh��|�I��Jʺ5׀��h��}�/��Ϋ�o�a����X��Cg��CUP��8bSV9k�� �V)�Ij���'g�^���^Ni,m/�����I��˼KS$�5� �X[�Ff7��r�B}�Xu�)�`y�&���WfNa�{�2���m�T��-��K�!��v/�D�B�����&�Ne�����Ks�e4����hC�AkA�ᛙI����4�:���qn0cAS�J�F���^��Gj��z���H�w몞<�p�����>l}u^�g�e-]��R�U��ަlA��G�0����<c�k~�l!�W��H�u��B9�ͤӯx�,l�P���hN#�V�=Ӹ{�K�o�H-��)��W	پ�,iw�{pc��L�;���Z����?^��0Kq�#������;ޛ*پ|��c3&�S��O���K�
_�����UJ?�<FX�^��!1���e�h�:�}�rQ�>z�_x�ǭ�`܅"�����8iȍ�?�	��L�����=oS�r�"	���.A�P�����̓r-���xkP7�����#�/���3�3f��>/㗰x���!�*w>49�����)|�ʆ���b�EN��"Ϗ�%�h�'�#�/���x�Nn��I�c�T����z1��RH�$��鉗�Շt�Ǟ���E̓����
�)��@ia�Z���H�;	���"�&y���	�������ɰ�ִ^Ŕ
���&\�Hx���G@��-"�$�5=�p�� ��i�䁜�ZP�D�&D񸈣��zuO�@'%3��	��n�V��REL'�ĪA�s�������Ϭ<3Ċ�PP�ūT�Z�le�<*xp�7�����E��] �VAmu���ƍ���ﵤ"��%_��?6�U�3����I��[�
�j�li�R���aFo�*S�5�i����-KB��`�c�0�iw��]C����"���yuC�ج���RJ���[�����9��uj}B�:�ת��1�tty�y(��?����U�:Ǒ�sē�v�D.�/}�O|�;'	|���'�
�ѱ8`(Feh�ʦx26̽���U�Ш���Z�5Y�揁_�������E�:\��M�-)A�<�-o~���4�l�Sf\�aQ���+���F�a��݋� �h���C��&��_�X�\6�&$�f�۵X��1K�6+��Z�?Џ`-^�kC}��u3Ƣ��	�؂B�Y���P��������j+�1+Nn^�#���"U��y$&dА��+-�����wK�B%/K�&w������\�z2C9�c�^Yi$�X�eL�?뷭�ۉ����oj2�ʫ��u5��:÷���f�_����w9?4����~���� ���p3<퐙���h�c=B����1�wvW��mf��s���~rė�!Q&"-�O����{�=aI�fƴ ��l���Q��u��\�D
�P�!"�3;G���@Pê>mh���s�t�]�xb׳���>#Py�z�RjY�����d��5xc"��J�"���ǵ�#C�0��#�,T�h�)$��ljI��;h�^9��]γ�2C9X��N��� �\�{i�R|��\u�0l�B���U�
"���}�n������)BYA,h�-D���Z�������lfgI4u�C�@CJ�����U���%&�`�(�C\�Y<��h,�r���������������8�$M�b������I[i_��%F���u`��!5�D�"=[4��l�^L�/gT"y�� �T���u����'�����<�9�� �)��=$�Ak�������V�.J�AE<��f�A��P��/'�(��qٞg��Dy�Vў
��X~SLE|�V���L/�&Y��T��3���*׊���L'{�n87KdQ�9ل2�w��D��w�Y5��_T7>��,	��ْ̡B�ӹ������
�]8�>�1�(��%ī��j��O~�R��# 3;��$�=�1��s�u7��Xh̈�t&������Ҏ�����{�	u 1�@	�W���{WC-
�Q�0nf�t��-�\'�w0��Ĭ(rU�vgݾ�S����u����������]E����g��\��忾��7�3��ª8�ux.'�&z-���rT�z2�����l"�|�ȩc"�4Y�b{40�E�cHNx�mQ�LB�K�kS�������i\$���-C�x-�,tւ�.J�f�\��L8 �]�1�������J��m��Ԍ826��N����UǴ�~��z�
yz�R3��	�P}>����cP��.�=!�&Y�:[����Ty3��?��o���5�(8�^��8-߬�hd0e<#�QS�qO�q0o���ļ+K�J}�9�Y ��p.� �
����:��u�6�%M���Bg�$��ˁ�nw��U���/Q?���ral|2��=�Y�����Lש�K��+�QtEȲ��M�"5��c��0]9���Az��⇜蒵ōkaJ�tW�CZW���6���Q;Xpg����O�M��&0']
v�e����V���<ۃ��J�;��֬��u�|��jI����E��UP%����U�Ζ̴	���6�c��3F�~68��� �яu-�-̿)�)�Sz;��U;�l�_�Ah����*"��[��9^�������m�5��`M�P1��1N>M� >f�Dw7�乌M�F�'ה�v9=���"���Q�=�w1������`9~���QW�1~\�������#N ��/lב{o�g"���JU���M�B��v�9��3��k5"^P	�B���۱�&*˒��I����D� �8�6c��'Q�����A���X*,S��������]W�J�8�,���)P�{�Ϲ� �?~�fˉL� ��E���h��Z#QΓ���]�!�,jEm�[-����T�� ���8
'U��܉7����7��L�܁K�M�"�R�h����Z������IKe���$�X>�Cŉ�P�u�����|g%��������1!y�C��\�R�ePz�L{���_�#n'a���*YdV8��S+����v�6��	j�
sX�G tW�r_�;��M����氭	'���kP��[b�~��W"�lX�����Y�R�f�����sj�$z�_K�\ c����R����W�pPYH_�6� �����
���x��1T�E��b.������!��K9��I�D��.��|��7�1VB�I¨>9?c�˫�1)#�s|��⪥��C���iVl�nlr*���z
P����~v?�	�v�����w�x��5�D�D����w�~z�K�@ �W~=�\��Z�C�IU��Qi� �H�C���܀`�
��� S�6�����~������7���l�}�P<>O�I� �J;��"��V��,�A���W�G�"9P鬵�$�p� ߛ@���{8#�4�����a�ŷP?���0U�!뵯5���M3��������!���-TgT������S�0Ylk��'L1�����jaɅ�)_�M���j|PS�N%���ƃ6�E۪O��%�PL��yi\^	��^h���;BA��x��vi���(�HRj�ԤqE\'�/W�iA|�Z��o6(���:��ڝO�c/���N W�����Kjk�u���8#�L�!2�-��٘S�����W��;@��L�/?t���i��W��4c���QL�����p2�H 7�u�]�����}��|^�n.��e�:J�+k����_O�	
�ސ-��+w:٘�
�ȨϿ ࠭/�	��(�{���?��$6y�2��[�I�ԫ��O-���vs�P�h�o��Ơ���bX4�����(���C��$괽���'r�M�#��E��),�OA�a��g5�<S0ГG���e�y�%���(NG��T�h�"	���X���ֶx��5�U��(�s��I%7����\A�\�)��IIуf�sj�Cɶ�-LtҖ�
��1OW�+\��Rb�eӼ�y�HB�q��?Lr˜R�O���<�����������=��<+��u��&�,�kE(�uVW�;�J��<к@F�d�F��i�@|�}=(����z�hҠ7b�O %ޱ��yM���-�ז�a�?
L�Z�")��)�j�&SUu��Hκ2�+
s����2�8�M!�F���$����u���M#[]^/�� 6M�~��]<�	\2�]7�{�[}��!jI3�|�:8������hlk��Q���?~W�`�SC{��E0D���#y�à���ٺ�G�l�8�&�w����"b^�y=�z�@u8�g������\�����kKE�/zڂ���R�u�7"ֆ��/�N�]�gYn��b�U6�=��ˤJ�G� �М�t��4��PR��6�+��{,BԺ�J���qa���/���~���πn�v�?�l�BfrT>��T�>��kصw�E_sb]����H���2b21+�$�@�.��*)mA|�ƺ����@l�6e� E9��8�1"��u��Yw���#����6���ɐ�}��F��[��5�u�-�@աq33�j����J{�.�=�q!��b�= ��E��oF42��	�u����^�\�L*}X�Y�)Q�Z\�:m��D��#��cp����Qnme~
�1`���?b<��N�u붤�QkJ�7��.f���/���a��ٷ�,�I�`N�j�p���pt������N)��S��Y������t\��Ȱ6��4�����J�mN*�;^d��v�ʳP{Y8{�)�dX�ʞDe��x���WJ�w��p�O��-��%�|Qm�����@���>�N!�a���3��D;�DR�R���3ȯM78ݠ�V��`H2m����g��z!1�.*1ŀL������9�_.��+��vϪ���X�qtΘA4��ex
���y5zW�Bq��;QM��Mlq��)�t����?����j�*�9S�����g��sF��4�;I' "Ob��F�3�"or|�X ��$C�[Ir|*Q�g]{��+E�v-��"b??��6��Do�l��5�<��tn��2��ɲ���-�p�����W�u��@Y�{V���"�F��j�j�((���8!F-�9x���AG���e8� ��͘B�ܖDfR�[���(�Ŝ��z�����t�؊�]<P/iY`x�*�W�K�����z�����4��)ƭw�.8�z/	j*�L섗x����P48y*���JdJ���W�?����Y��5� �f�r��0���z�EO�Ɂ|�� �%���j-��� �*Qڹ��^o}�Ɉ�r��D��}�;\�B'�P�3�������lCrk������[Ϡ�'��z�X$�,L�/��C[�b�Axt��j����c�li(����H�!�koL
�/�*ɢz� ���Gt?��7�%��!c�ޡ{6I��#Ĭ�o}N��4��+��k���$x��Z�������Ae�S�VO`������-g�;G�3⣴��������8��Ҏ(1�@ܘѸȀ�����g���`���x���5*"�*v��yp�,��ryZ�A��O�� *-���тJ���;�K��Y�e�eAk.ؚ�67o���T2����ŲJS�9��I*c����M���ǖ�Q�H��Y$p��<]�M&�ʧJ�|��q���%�aӇ��0?�Z̈���!��$\���%x #�A3�@`9~��IR��X��4����O�51�\^&^�EA���nڵ�xc���x�,q3%&�82�"��t�~Q���P^2�_/66��b�}���%��1����T��Ðz�"_2�o��ƴ��k�����O`�i���C���{�DG�Ǯ�$\6�f�A�]U*[�-5Ǯn�<��<�N]u�=ی�)騺��@bȍ����E�cs��jo����t`�Wq@H�ݸ��Y������4:z���<7c����#�:u�2w �<���m�J@]/�/��mT򘤿0M�?�:&�0�]�L�R��vTF����iM7���G��n6���!�ꓔ��,X%�}��E$��>:�����}J:�<A��t�7��|��E�"1	cѷ��h�J��5"�I��P���@)-�g6�ɜknNl�*�G`�+%��p��HY;!wS�.��dNq�Ui�ڸ5���s�!�����*q0=�A��s���iLu�ߟE�Z��Jf��7����O�y���e [�"΂x/X���9~S�!k�{��jhi��U��M�+صWu%*�o�,�rd`MNZ{����E����颴�7D��$�֛�Hkm�y
q����T���ӯ�x�A(�i���A�	1�.D��{!D�
 q�g@�&0���~:�xm�[��j��HhQ(�85zӽk6@��:�A`�%liz�cA6�t$i�ɿ�t+�f�<@��������]��n��#���Ӱ��@�؈����R��������4�|,s�A�Se�U�W�iկ&��ƀ��������=��%���Q�rٶ %������OVZ�p�50��o�2#;��+�O�x�م�����[��R���s��H��ܖ��(� ܃�=�}��3'�׀��D�bZ\��n�#��΃ޡ[pV�	vMx��c��&s�*H:h���)�yf/|���dՈ��zK�^1�ʡ���tu���UCJh��j"��`�D�
A��H���W�\ђ�?d�+!�x1�!Sϖ����nRC�/B��wAǀ�څ᧧�E�	�Qg��|̭�蒖�L��h떱��"Vj��0*��j^�5b�KG�G�g)ʯ��� ��Ϝ��HU�h�7�ήE2�#��ш5-'�u]��Ln��j��Z܄E�
��|�һ���S�f�{	�X�y��t��CS(�-;c�.�*Oh��i/a����x�%�U0�y���X`����p�v<N�.��Z
�J�gW�C�1���~���Rc�LoV�%K��ƧB��~Ml6�92����k�iѠuw'K�s`�^�ʮ2q`�ǒV U�D��^�fN#�Y����ߏ���rni���^�>L���=���8gC$�Rt,�C������1��T��E��y�m�r�"�K��t�N!OK�?�)�Y`��,�W���cg���8�ΐ#�&i�o������]�a��r�Q����+2�A���%t<���&H�dG
���	r�0�_�ȑ�^'����xЛ��I��m$�/�e<�� �]�|�ѓ�3%1��`��M��\CY��D%�"Z(I"q=���j%��)���'�'?��4'�����_ۡ՞���8�\��m�Ԅ۬>���d��Und��ju
6�gz0Sϖ��?�V�`�Ȼ���gv�=� ��^%i �})�` >Oj	�p��)�p���N@�
993F����\|?g��g�jmp�t�#k �s^�,P`� ��k#D����]y� ���Q%�T���ćT�������C��^4��낮�`�'�#�;��<�4�~z�2���%�
;\� 䇸��?�"M������լ�!�~+(�)^U���gd'�'�<�6��(ʒ�Asl1C���7i���`{�������i��EQ�uu)�#7v���v�d��/�<���&mz�-G��@u��N�3�����p�5�����/X�D��Jk	�G���c�N�]�J��O>�-۳����l��U�hj���։YmX�5*9�SQZ�ܪރ�Ⱦ=�4^R�᎓i���-�V�	'3�B�b��t7"8�p�&����sD�s��v��@�L��CrHQ!m�#���w;Ej�g���w6����e������B�{��Js��W�W���DLۑ\T5��q�:��~]
vBw��=gm5^��SO�a�ݞ��fU���D�Td�g�pa�Y��s!U�5�T���\�?�q��:�����Yd�-�a�U&��ՠҠZRhmJ�jy|�ḗ�+�@�[b�ۧ��7���B&(�yqD��G(��Q��LەPS�Yq��/�xp䜒�Q|�D׸v�$v���dU�'
$�#�w��+O��K���J:|�R�<,�x����"�}�qA|��;M�@���!?;��rpWϼƹ�tsR���Bkc'A�^�Fۭ���$W_�)(}5��<�	dP����[.v�-:oFI�{����ip�L���5$���#�ʃ�l�iNc�>8BZ�@��ũ�H n٥��(��z�Jw)����E=�Vy�.����@�I-,���'��H�� D�r~�&l(t�Z;��Q��B�L�Z�ò��u%��޼I��so��E/n*�h�%-�����,ѻm���~�6���������iȯ6�JNٲ��L1xVc�{�Yq�>��f��d����h�Y�ҊO䥹h����"�� ��\iT�.�6.ٜMhɇo���<㏩�D����F<K*P�.��6d�6�n�f���dgN/>�u�(�0��$\P[����£�>#�K�uF7�^�-t��k��9�$��,2w9�,}J����tVߎt�$]���[5b������Ԋ�_�������T���� ��yp'|wzH���)^�h�wd����c=FO��q��}oM4-eW�,����h�����
��\Xu,�m��{�V��� 9C�|/>^�EI��i|4���`�GУA,�ד>�o�����=a�S�tj
�=�`�Xݕ�K`�]�ϔ_��t�~n��T���L��Čۮ�G�k����^�b����׌�-ڇǆJJ���K�_�F-!U��$�g�VA5���8V��ّ&��8�{�:˴�X�z�<�-�0�E��0sۘ�:r4�O�h7AO����eojD�W�؋�B�٤R�t���V� ɾ|�]�wj��r9�@�h,6�F�1Ez`]x�%{�l��>��� �V�&N.l�S�*��󛅽�a�Q�~�ĩB�ڙ��cu�fP����m>F�_AĀ)���6��6��E�V:|�l�wJ�b�xb/Y�?�7����m;B�f
d˵�dY��_���'�z�Dr|4>"��*��Be���\N�'���P}���fn��]�������P��j�O1P���L�k[�r=~�,�/ch��]ڙ��TѬ��06]<`ݺJUR�vN`C0�#��r�M]�e�z�\�51~�wC.U~��#C[�z�0�ض&&�lE�[#>D�������E�Z��N>�������3�*hUè!���ԣ"H`�߽@��7f["�֣��z;n6��n|�&m����}p]�-��ޛIb���bd�����~���� ��u����!60��>��	��]��w�������yF?"1�e�r��Z)��$Z&?�X�!�<]��b�&Ly(����Y��&�.���Ϛ�!�臤ׂnd�T�Sv��W!��*H8�M;�Q�p?�Cｨ;M@`ư�6���������
�w)���$Nk��%�?8_��;���7������!��O�����n,��f�_[�����s��tU`o`|�wc
��:�%���� �.G�QaJ. 8r>h���9_�Ut�JEd���q��� Yx �6���t%�Ax�ٺGF=B ȟK��6 ��Jr�C�p�۱eS]��n��ܝ�Ĩz=��#Y}�o�NB)�g��묭
�س���o}ES�1 &Hw+��z:p���Hӈ�լ�����ok+�=��r�BW{`��<��Pތ	P�W��5�	v�c�N���r����-Q$��|[w�h�R=�f*��P-Qb\�݆��K/�v�e��tLi�Zt��n��8�_M�x���D2��=J�>[]z�:��Pq�N��^'_������vP���Xj5Q7ƴ�h	�9�ܫ��z�6E���N������$^�������%+]زbV'Ff����y�&w0[���4<��LM���H�D��';]l�e(�*�h��F6�*v���Y\����^q.�Z$~��a�}�#������l�~s5d�61ui钒�K�ͬ���&�:7�mg�]=��9r�(���^���J��*@>],��)5먣�U�SK9�J�'�J,����4eTJ��DebK�&/�MM8��5�����n�&򅑦5x$t�>��� �����]��CB��\��<<�H����ߧ�t���4-aK#�{C<�A�vj����U�.�r���z�.R	ޥa='譾���E<�k&��nϖ���]g?Ш�1��s�K"������M�g�/�� ���xF�K���	2��� �����Ķ��tT)�1_$��O!`���K��1�n}qȉ�྆t�G�c�pG!�\�ǹ���I�ApD���'�N�y{n�_�R�K��5���8�ב��������>���7W�[�E3�H�5�p�8��p֩��8+��!l*����Z:PͰ7�{�N*G"�P<٥������aअ�D369�8\{7XE�Nz�S�M��O�.��H���[�6
��j�嶙�}{�����W~�v!��dHo:���������u��=X��haT�2%��o�"=�}�� ɽHO�_��Q�� �������[�e�G\�~ώ2[BAD�Ͼ�!r��kR�t�2_9��|����g}ۻ� �|�M����teވ�G��)��!��u�M�5>�����0�6މ����V���K\�$>Tl�f���,�̩�\�:X����*��;��*Gj
�1���@Q�`��3��2�*lK��2pXX3�T�siF�(������u�g�0E;1�q�}v�+I���)��JS>�׆��3{��<I�
�FU�D�x���oR��eQ]Ji*B��ls'~��m$��i����a�V[Q���b>�<'s7|�p�<Vr�bd��C�ƪl哅"�{�~��o^��4��dyE
�-2)��ZD�WT���W��J�AM܆��?���C��rt4ݿ?�R#�dX�%Z���Ъ�*voH�G�ʧ���P�i]�V��d���9�;���Sr\"��T)婄�Ү��x�k�;�͏�*v�o*�����T��i/�5��}���5
�ek��F?�E.mr�J�����<�cQ"N��(�ܕ֜�{D/ ԆHiͥz�F4�N� �B.�n6s��z��[��G���$F.dTbՈP��77wfJݓ](啾��]����7;Y�@��b�)H��`T���{��iĺ�A��(?6�d�T9X����^B�f`v��0Z,9���Z�[wE�[�uam��voם5峋�
�.��S�i�*|v�q:0	�Ӯ�~"��k��+�N�RI��@yL���/� Ō��i�Ӣ�&_R��]՗W�x]Z0��W~�2�:����+v·�	�zV�(�	��{�_��;8��n�!	w����E>���,�t��O�F�|зƲJD`14=42�l�+��n��R����:~��Ӄ�aK��t/�J�qPBS�ˎA���<�p��!�͸�uݘ������r���l:6�t��T�$���=?����R��Gi��u>!4��P7��Pm�Go�l�IXLqB�N'���$�ٰ�����o�A�-��*�f�)�尘H�w��F�BX��>�;�.�$U�c�d�x 5�ӮlO(�����?U�h��u��%���V���7y�'!��<\z�\�a�����!�8�����$d� Aņ�l/�8D����[/����}����5!�T�n?4������j6:TTp�Tf��Хq�b�&����f��i�z&d�!��\?����M��OX��	'eX��p�{�B3k���Eq�zE�~�����Vص$�B��Q��-�1fPJasv��7��b&<an�Y3� 
)/4O�f�"��O ��-A!j�n=ސ���@��v�� 0/]gķ^+��tfK�KL�n~�	IA���EFW�vb| �x�Z(( sn�	͵Bs����H	�=�}[�Y�A�$~@ߨ2ڢ�uH���r^��X�ׄ���I�DY�^��Sz�8/��r��F���΍���Qs٤�+�fM���8��bw6������W���D �F�9����C�F�j'0�<�d��`�u_j�v����ׄl�6����[�%.M��Y��z�K���%P��� ���4u�k���5�a�K|�-
$k*�ͻ4u9�����!��g�p߶����<��TK����C��YaO1�mկ������T�=����\Mz�@�	Łppe��%To��׮p�}�uf:([g��z=!b���~��.
ъ/"�tVP��m���^�hh��_��y-�V7DS/����qW�ڒ4*<���
�KAyu{7]f[���ɠ�TԺ���z��km[����5O���'GJ��F8���=iU�;��`-��⒚���((ܡ�%G{��j�e�^OBB���wPt��l���c@%���:�N�֚��cy�~�_{=����w� �A�ӧR;��O���7	��[�է*t	EBdǿ"�����`.�>�e��G��{Nĺx��y#G�^�Mr5D���q�w-d�T��V��/���ͤ�Ģb�=���|�`���5�o#�G9��N���t{Y� �;�g�����6����a�w�C��[� m!��oZ�+f��M�,���#�3�d�8A]>�����Ң"d�;~IAwXo��̭>��� ���J������b�v���(�o4��c(������*�:	qC�V�loi�������	��f��TvL0Zb�E<����})f8C��H�<T��rQw��Y쁸�mfU6������l�T8z^�(�����������\�2� �|��9�! !�삺R��n�jy�ܡ�3F��W��VX����R&���~[����/a�����ff�Y���g�P�,��]���j�}�r����gY�:��c�[��p<~���۽m)����p�vϭɒ��Z��M.<���������rJ�w����d��tH�r�i�H�q*7/���8W2���?G��g��G�����G��\S ��V���9$�t�t��>3h8�/7�+>���,J8�-�j�s�8�Z5�W���C�,�o&�0�%_L�vO��~��w��X�?����v�bX����
�X��e\%�lq�}���i�ݘoϾ�3t ���V����xa��NR�7@�8���P�\|l�W�f�T	�g ���0օ��K�� Z�H����A�H �K��u�ϲ��M�GB�<1��� t��,�ll_��Q-oT�5�IW�>��)ISr�Mq�AGB���7�r�>������,��I!O�����UC���h�h��W^��.�@�Y�d9���˷8'����]+ض:��%���u+Aʠ~���'J�rA�����(�D̾����c)���������X�ɾ������&^	�V?��^#�?�J�A��N;0�钦w�ܚ���K��C�%��\(��	�,�Sօ���'�D�8�)�;���=<��SG���u�&gV�qy��G�˯?��{�x���:�C�C����V�W(8qO��mQl�O�Ik�۞N�m��t\��*�m'���ԓ�>��_�B¨�=F>"���O2��5�;xIB�����w��l�J�v~W�n�)�9C������#���놀���'��3.x|i�����\jDwm�^�g�˗M�����_T\P�| ���L}-Rn��V�n�m�Qyvp�$'���&�H����m^����f�(/j�S\���E�l��~�ߎ����ta�E�ψ�h�����$��a��+�_X�1���4FH�,��|�*��]�E������sUB�:�[<�f�����BE;�߼�ɍ�R$����
A��1��`�=g�/ZI,%5�jX�ziDL+�曡6+U1�R3t���z ��z?�5+y�%1����y� �>ko���I�^��F��/�w�-%"���t�u[�Q֢d����:�_�8�}��2��8E��:>C��<1���:�*�@c�'�[wX�'No�~q�	X; C���Zf�i�'��Ȏ�-_���z����L67�����q�*�!S��FHz��Ǟ�����n�z��j��bU�5�Y�.h�gi �_ܢ�E.��i��A����|Ęr}�=W���0�FU";\H���?`�֛9�v9���J���0YD��7����W*`2��ZK��g����*��i�l�*��z������1���6���'f�B	���
� z�Y��v�R����Y'����-i���F���Z�t.UD�[%~��"���.%~���]v�c����mץ�=)٨�c}u�a�6�4c���2�=��ؑ�Ђ�*\��d}%O!��\���/�ؐ!��.b /�����҂��)IU-�����73��	0;����`���cU3䙬B��.��� �u5h���Q��䮯h�x��w>y�.U���˿K�j"F��h��}�D�o�]����hE!�|�ǸY��Rt��p߁%Q p?2��&��e��7"VU�_�^�,����p��A����Ɣ�p+vdS��[�ra�Ũ�I͈��anÃ��Z��F�\8x�8�\��-�>�u����5aGڈ�X��_	)W�cH嵔kw&r���*�-��Pw�w	�e[n�f��a�k���A���;J��p@4M��̏��u=u�t{G'��eo��Ru8qG������\��EF���<��ڔl	�e���y���SS�먿D(lc0s'Mo�7�]�����p���*I����B���{Y&��P�NAr�m�1PV3�8I�E��P7�v33}x��ܙ�w�"���%}�#�e������%�4k��
����%�,�7�}ftM���	u �xJ@Ĝn���Qx���^(�O�jJ1���@��{���U9�δ/4�Jv�uc)��Y ���lV�>��@�������Xg��)��<p	9+:�f��b%P���BB��x��ޫ �Ke�~�& '9�&��C_�ON�S�P�-V�%���Qc�S�%|���I;��Ї1�4�xa|���lk2�ËL�f��.�	m�Q��d q����<�S[,�(��3��#%?r6��[��IN��r��Q��W6/�b3BF�������)��L�3n[���͸Ym�&^��a���J��kZm��V�&���nc!�u|��Y���� �����5]hSm������2F7S��F�C�j%�:�	��N����a�����
X���mDs�r��Ww��X�i��E�ժe�h�:�J��E�i����\PZ����Ϙ" hR]��i��3#2i dE��4u�`R8����:,��j,�?���"0S���1ӣ������җW��I���bkz��#��
�"EQHȑ�#�F�}�&��~97ET�[�>c�g*�o��A��I!�	��r���^���:d �'=�O�iݘ/j^Љ�D���JT6em<Ļr��ԳZB�T]y�a�5�}��є��B�,�~�M�k�ē|�ĕ�Nݼ̫qh��4�!�s$PnH5<E�p��aዝt�ʃ_�ǭ������������!�r��=�Z�aN���<A��@ ��:Ә@}M�ֹ�JE%\s�O�'�(��Q���	+����I�OI�<���f��J�`?,<g����D��T<�5��Fq�N��61b���ͤ?k������4*�M�p	c��Y��F]. <d)x�Y�	&��T���2��ӓ+g��#�,Z!C_`M�R5�5��!f�j�?�co4T�E�[d�44��DxO���Ι��24�;p�g�7w�g/�%PRY4��Z8m�3c�4}�¾�ԉ��U�-����iD.(�&��=9�l�]�RG�������,�H�1�GS��2���������'*0��#|��p�e�H�����НT���+�%U�a��&7���tZ5�$�J����[C���d倎Β@��\�F���jƮ甮��8��@��H)�-Ux�|����"y��S!��O=y2��|V@���.fӚ�废�2f��1�e��9�|z>`t�<�6��}��]f��	.�f,RVl��
��f&�Q&��:�f n�9vC��>��i�1nK����n�⛿}_D��[�a��_��׋Y{�����Q�Dd��F�*�H��)�pחt{�P��U�4B@v|��W�&%Gk$�ƂY`2��q����O���Xt��3�M�/��^���7=ܨ#T�=ɶԵ�KL�*X�
�d�_(�C\��r�u;�s�t�a�=��B��D:ۖP+{�Z�eJ@�����c\��E���)ڼ��bf=���N�	b��S�Ȅ.�Iq�����
&��rM�H�ȔY�^����尊n�TRv)�$V�!�;�����v̼��4MB��FG	@A$K��~<V���8Wt�é+��j�.�%C�Xͧ��ۊj_*�}oH%<dK3���աp�E��N��Z��R�J�����R���6�v���6��&�-��}o�0�P� L*�R��t![��70ѭC�VjE��y��1ke��Ł�LA����&rR��7�B�P��{�x52�B�>]��T�]/)'��Hg�ʶ t��Zx�b@k��b� Đ�l��y�/�N�ꋰ���:T�� ����(?���0%��՞t��X��&C�9;1g�T\x�}��7^�w����?dBz�ȴ�L�z��fopEl�L<��%;�c��`r�b����I���p(������I[A�m=@*��v�/��XF)�������;$cu�UJ�Q<�_� �}r�1�[UǳFo2�y�0f	��H%+�;�8�*:4��4�����ȳ�$q�lu��UT�ey~ܪ �+7����H���mq3+�;���С��it�½&5 �>ۨ�an������㐘���l^�W"~F�}�(N����ʁ��qM�ئ�2�N�aH�U�uV�.�ѕ� ��� F��I�n����Y��u��	3@!U*�2}w�0��IFQ]�;��X�jӫ'0�aw2.$ǭ�����GH�h�����(��}^����hdAh@>�_�y����?	�kA�Z�U��Rs����n�e�yê�	
?�R>�������3gi��������shzĻaB7֪q�pzԇ��z&ɿ��ZD�W��f���9��w�JX/`�rA��@�dFd�bi�
�pօ�˜x���i�fτ	�p�P
���h^a�H*��p�{L��c�����yT+I*�8����t����f$��,�6Y��>W�7��V��|��'c�^O`}B��Ԍ���)�0� ��iA����a����-���L$�j�g�mE�T(�B,���
��d��Lv�=Ŏ�.Z4ހPt��LBx�Gx��e�jD��*��J&\2��-)���bmyS�.OA^6�	����k#��cT�(
�����»�"�ȏ6����= q%g����Y���f�x.F�£		��i^�l>���n~�{a��e[�R��g��>��	��u*���6 e.
�F�xCN,�zWG�4���($��o�T�ނ��u
�F�9��q��R�D���Be/��l�j*b�iPM�m&��P�Ӥ+��rxdL�y���Y��V�J�(+s�Lh�&jV�������1|�������m��o�6b"�tuK.v�EF$�wX��>��I�VEW�C�΅8ҺoP6�ЀB_S����i����(i����Ts�4����$}��Ӛ����(6�$���!�[�'d#�nՌ`�+g�5!�چ?0����om�k��Nc��Pm��Ny�4l�U�d��H�)�j`��WӢ �-���"KЈ(����_�l�r��k
�i���?��_�<I�L��Ѿx0����D���U#'���6q\|�]�3n�H'@��d܆_�%Γ�_3�����m12Ee�]�E���Җ��lO�E�̑~�����E|�a��B)�o����˘$~uJ�4�T��I�n���gx��_�jR䇱�k�e�7&z-�1B@�3q���*�| '��i�`A<��^~���� ��V	�8ر�Ҽ�l��>5��� ��rS�=M.[x��%�æq"���8ߓ��,e �L+�a���_W��SȲ0��F�����l`V�Y/;��t�M�؜#����v��/C��Ϡ���0����h���CV�z+Cޞ���>e�f�8��t\�^\���a�;��U��Y�nF�]�ȑ���q��n�6b����e1-X Zβ A�{�?q�9���?"���wF�6=�^@����G�r,�ƒ�x[�S�t�����ô�RL�hun����$;�R��H�� �QDo���M�_ ѱ�zu�׏@��z|# 7|��vr)���|��Gp�/~� ׹�B����H�.͠��RM����=n���3����\�E��A5|�U?Wz�$��~p��nR�\e_�JF�{j+�i_��Nį?˺nlD�<|��T�J�NeD�û+�.�mlǷ��)a���Я_�X^,w-)M�ɬ�YL�p��xg.�Hl���N�q���4��x��E���Rj��tY��U(���,�۶8��Ɔ���>�,�%�^~��|!�����8�PhՇӸ�Ė+�Q�C��EG���2W7'DY���q��A��"E�3 ����?9vb;�I��Aˠ�pr>��y)��D�<.2q���&;ݖ�1G1f�9
?�ɗ��� ,��^*'Ռ��3m*� @=ɏ�ŧ���$0S���R�~�\�)�q��pM<VlZk(J����P���8��-H�3��Lz%P���� F�r������h[q��P�ҏ➽y�#:1��������N��X����A�ŗ	L�b�Yu	�P�Ed�M@(�����?�ܳ�}�t}v�+U< �IOG�����F��#>%b�h��rMڈTٮ7Ո���/.4��wT�n��QV�fm5v`�13Yb[��M9g~����̋ q����ն<�n�c�T���(9�]�P�I$��RۦW�\���xݾ����m��g�¥ۂ�۱��H�����ox�i����ZC7v3�I��Şm�u]��� g?����QІ�K5p,l�>Olܧ���ɐ��M�n	=A�	���{ql����"P�3����G����i&N�!���Y\#�G^'^�ʾ��©����j;M�!_��'�����S��,���,q�4i�P��_o��(�cx^"�7��
W�Ϋ�CT���`r��G������,�:c�S�a��茇K	,���Q�ٙ��S��ͦ�W��%f�A��׷Y�q��
 b�6ګ���i4��h��9���-H_���3��b��
�l�+`2�=�-1Ⱦ_��:��b�n�����V;8��I�Y�Q\���M�h�2�5�(�5��gG������ �1*PQ$DJ�rW�I�*z,.�/S	L��q<ѯ�iӌ�Cm_��p�N*m�|�eH	�]%g���@Ӄ�_���j?�J�v)ÇST��2�.d�Y�@���V>�z�pr�SF���ʨ#O(�p��QG�j��-F^armW��]"3�6��AAU3<�+z&������o�dB��l����3�t�v�r�W���o�!���{C�k�x�Ǒ25t�����WƐ��N-��Ѭ�!Nz�5�ޘ�D�yI]ubQq�O_�~Q<oMf��BMG�ab�L�9�R[X���u�����ZS6%j�+�[�e���a�BO���x���i�ȡ��B?�C)m7�Y���M3�a]��D�.��K�����\i�K��NrWf�����0� O���}���[�>�Y��Z�}ޔ���Cj�N0��g	F�U����ہ�6���S��6��P@�Y��8�. ��+�N�Ș�q�����S��b"�lxQg{!�=+W����iH���֘��)y�}��?�8a^�JDo����*#�5ylc��,�-�(癦1P����	$p˿c�g{>d�-k��E��m�Nu��嶔�:iÿE�VC�LA��Ռ7mK�Sd:��0���h��'�Vű�ѣ^&neB��f����o��g��!���"��?Yx}M�h)f����k�vI�R�M3pm�C���GUž��$4)��D'	�ӕNT&��0bP�6+Z7_5b}��ks�a��b	}7]X9�<��!��k�)����36�!�����f0�x�b��IG�9���B���zs��C�yXi�0E2;.�_�G�B����cǯ|OGN���lo1�p���es8��y�j���BVm��CN�
�g���3�Km�(A$�`5�G�eT��2�=M�k���b�)_!6�����M����.��`oR�i�����Ņr���k���Ss<��/Gg�
�{I��z$B|�-�c!<pɁ�0e���]�.�s��
�:���]�:q�Tk���zմيؖY��v��T�i�7r����aL{�~��m	���V���K� ��}��� F�A�U1w�%"U��)��ac̹#'�����'?�">����L�y�Y�p����ƃ��zҌO��\���X�+*.Pr4j*��!�..1 ��{M�eA�TԾ@W�
5JJth:Bs��Ԗ0(��*�`��̷9�D���G�uA���8�D�È�m��.�/��^Y�8�F�E7`��X�8ݼ����I�R<1�Z�dP��sZt9�F�`�9���sA�F.Fd*_���ȡ���(�⺇���@u�؍6K�,�ِ��6P�����bft眑.-nfD\�l���I&�mO�,�Χ�T�[	�_ؤzz�F��}5����J�Մ+��V 1"`�ْ�]�"�����[���I_��t	�.�ȕ�ay��ʭ����!��_�� ��[��t��`_�w��bL�[�|i�P����,�B�g*���﹀	 ���`*��Kϱ
�Wi�\�A��V��-��˥�Oj9�Hh�&����*&�e(���Y��ӈC�X^�;�[&&�v�E֎e~�.�;��4����8>�Ұ�ZON�^��·(�j���o��^_�4�d��N;@��%��k;
âYr{��-~"Ж
�(덋�|�̦�K�{Y��[�#f���s��3�_T���9��C.��V�`��/�FZqB�Q�7{���mA����m�1dx�ϩ�y-g��?��a82����5.$�1����Ġ1=־у��1$��Sɾ;'���$��Vߑ�����D�*��ENH������i��c7�#��<s��=D��ugoU�����frB�s�r:��-)���_TFr��2q�k�Q�%�v�������Q2�Nk��3�R��&��"ov��P�� tc��yv�$&O�%r�T� �:��ۯk�d3@3k�P�np����[��F��jj
�eV+����]����~B�s�4�\I�Y{������_;��SsU�Qx�W��)�����U����e�Ǻ�b��N�cc�RY6����W��x�r��=QX�}7����������@��\'*r���"�V+�|s�;:�8d-�a��n�e`Iyٷ*O��Z�$+��%4��K����h�5MnH�uΩ�l`��G�U��S>�9��AN�|I�.F7?�ܺ���E�4pw�rōXI�BG���)�dHZ�-��3Q��c�3��}U\G��:���侃#����;�O�"�^��#L"�G��x'��h�q{v�.=���Т����x�B	���Q���ޱKI"��-��6��XZTu�7�:��&I��n�FD<�93�0���o{���PA��5��b��[��,���ba��$�7���:��x�I�e�����v�����6�� 0��~;L��7?+��J�p<���PO�ܥ�����I9�c��k:ý��8���3?�g���hl#�t��r�g m�;%�FYV��'��gr;�1�ez�s�/�IO��Nw�	3�,uLv"�Lu>�	 Ÿ��$lOqE�z���h��i���KʮUQJF!�d�b�n��:FJ�����x��v�uZ�0Fh�K=��=�g��P���L1`�{�WH�h2��]�Xӟ�O_8��VB�!|�&r�WMM��P�{{w��F%;0���/&���9U��e�e=���#���N[@�=\�O=<������&��`ӻ<!��v����0��m$6�1��."�ޒ_���4��f����6�4�2��D���_�3j�:F���$+���H��"����i�E66���DJf(��2���7r�Z�r`?2r�z�&`�/�g�Sv�@	�c�M����6���2J�OC�w�w�Q�e� �U��n��>�^K�d书�Gl��n�31��Ro����<'ո�%�mRo�}�bL}WHm4��E�m�ni�M��椭n��K���8	�XP�E.Ӧ�Z�Cr(��ꂞ�ؗ��1T%7D�m��@k�{&C��c�։U���M#�����\@��P;a���`*r��V��umw�!�ll`Dݛ���iAh��ԩ\��6�8Z�������Īsq�c_��BT���I ;A������	:/
�mz_��t��\�eF�y`ȝ�Lˢ��݀�^�5��
���ð��g�q�� �b?�m���:U_�k���dz;yM}l�8E��#�x���3�A������X���1���}�(!p<����-����:�G��9D�
$����P�DvN���䚨���O��<�c��W/K������p��+���>���K0������`p+\��_-,{#�D~��䭙�h���̣hy|����ك�f�P��\��NO�gj^X�u^
x¸m�$�{���{j
�ri������ ����=��9*�+��;)�&Ϝ�3�0AA棿')#�fԤj8�����l��I鵑��M�������SIJ�a��<�p�8㈼d8^/�1� \>�V�iy�OK|���f2��F���FqBC&Ǚ�
�zQ!��3%R^u�VLcd��a�h���/��[�d�t��<�O���Xv�Lz���K��G
�E�֑�/�𯪂�B�t�ϕǣB��}TR�,,b�K����Z&0a�)%�RD�b��F�ƛ��� �?$�og<J��kھ;�g Y�[��t��h=��Ð�;�Ǎ-���^}T�O��@��'��q�v�Y�'�`%�(U�hk��7�;��aЇXogy�(!�'z�m�ʠ#ɨ!A�E��w���Vd��՝o��1��Z���'X'	H
c��3���S�J�l�&�p�0O"��4қ$��m�)���2��Q>7b�ߥх�D����H� ��q�3l��S�Uп|��5�rP����MI�6s|���.�*6��]�?���IԿW{O���n%�CZLO��B[ I��ՑR?uS���U���26W7����hXF�IXRr�\C���:+e�B�@[j0��0�j��Y�9�j�͡x���?I_���4��֜��#�!D�-4�C�ZZ�ӡ���B�2�֡��*���|�NJЇٌ@$z��g��;-�:�`���{ε����?�ˏK�<4|�����e�)��;|��[�c@�9D-�"�M��z�<ew�L+��mydz�ut_S\HO�c�Y�'��La��Uċ(%��!#Q?h�x&�T>����U<r��U����]��K Ǵn�Jt��S��b��:��� ����SD��#;��`�ͪ�7^ͣ�W�>(]Eq:�L�����%vy~���Fl,K��W���$Kڸtҿ�
Gic{�rX����Z g�Қ���C��e������^WT��U��V�Ւk��Fx �Co^J#Y�� ��#��[H�zO@K�$�cK�*Ž5`P�j�̬K8�>h/�Zu;��EES��s��qן��%���i�IB�v#J��u�ΰʼ;�9�%��i,�E���5}W�4M�v�p^`>p(^��v��uK�k�����cuc��ň�f;�����i��s�����S�M=5d��P[U��K�`3��ߝ�%���}=�s�̮����G�/����_<Wn�!��G"3zpb(�L�w�)�VMS�����K7!�,�%6v�.�Am��@�MB��otq���~�뜶�f&#)�:B�莠���O�X.�Yhp�����;�=��#����#u��!z�Y��D��f��\�`�<I�U��s���tgv���D� �t%�t��-?UT��"B�R��)���������$$\���h��Rht�=WX������P�L�K��tu���P�{I݄ZzPz[E��w�酣�,�Ś�C�D��t�Z�1^�wA�Hs�e��A��
��]q��y�f�`�Z�>�޽-���,��a��7:*�#)P�,�<R���Q����q"�ai�r]A!#������V�NVkZi�1I)�|[ʝ�F�&�h��9����g̪�#b��O����t�,�����A�����
�������S���V �$��!l��տ��3(�!�4�.B�ޔ�(�l2�F�-sH�]��~��~�M�i6�]9Sx����������kF���'فI�Iĳ��[~@��Ah�@�pIpѹA�nt��^q�"�P"*��%M\:c���Sh,2##�4�o��-8�G����q��w��d�{NTv������祐�������@2����Q�������C(���!f���.��	:�4]����+tM�J��R����)D�d� �M�EY���eih���s%�J�sؒ���O!�(}�R;���F�ܲKi��e` �@ I���E;�N"h�Hµ��b�i+F�3+�0/9ZÁ/���Al���qO���sĥJ�ȟ�8"Z;�.dXPn��ie�s��w�g�JpȄ��ꝧ�߼�/c��g�E6��fr��Ғ��]��*�J
^�˚�%"[; 3�"�,C�~��zb�G��&�L��B���7Q���6�l|�<րk���Ѱ��M2\:��؂�E�6�����x�s�o�jq���U�޷m��^�:GئA�ׂ�n�#�z(�HRΤ���(e6 �(���8���p^��U�
"�n(Y��9#�0���s�l=~dc��g�95�jO����E'*��q�C�(z��\���b�%괙2ųげ�g���jrP|o�c��j��Z	��#Z����5w�gh��+zE� ���^�x���N>��s��^.�\�]�Q��=9�Џ�Z�3&�ւUc5G�h�Xz��qfܜ��ЂY�jSd{���QR��1 ���-"姓tA�r�cz�_0�P�pj]!aK��_!������r&)���/�1p����'рN��)�,Ϣ�X���}��s��B�b#����]���G�E#�2�P붎�-���.oK�"	l���s��Z�r��JP���|���e�k��%��ٯ�@�.�������pH���%�U�b��M����a����$A����⿽�WS��B�mA|"��%�����{�3%�ګܬ�J8���iO�2�f�n��� +XS-n�&�Д}�_�
%M=����ϵ
&Q���B��P�(�kC�8)q;��V������qv��+_��_�|bM 9��i��GN����Ix��n'��q0�z�|�ܱ�:�Icc���e�8����f���6���6���k�z/���@�$<A�K�J"H���Te	��)֣���;�j�ow���%4C������;�|P��2���)�׽���qη{ߨ� N�,��q橀*��m����m�b"�ko<l��J?��p	�̚��^X�e&S�4�]�:��7��	H���/e#�9I���;6P�r����_0cw��trS�n�ti ���1�̯�6��2-�����Ր�s0aF�^�R���~s��_��ʻ�U�s���(s�\qp�]�������-��/�,j�%@�[��9����d�W����a(�#R�s�<-ӛ)�'�I�E�R##6:�����Q���
�����ִ�w��fٸ�c��R�'u��׎:����KY���N��)r�:Pҟ�o��/ *��?Q^&��5UD'�~�zm�0fz� �8�x/�]:������|�(7;vT�]|�:���/�u���$�tX{c\Z����kM��c0D��]�C��T��p1�V�~⡦]ޗd�� �(;(Za�7\hM� �A�
�h�wV�b��(����:�����?��dE�X�,9 ��5�ᬙ2�G��Y�P�-A|��Cȇ&��Ī�a�U��gn��wv]5])��46>�UN%�|$���Hu�~��G\�)g(�U�����x��N	�2��R�h��BG�hD��a��JZg%�PEGĄm��%�W��n����0�6r�����ףT�b,�rd�\�t���W��I��*E�5��ch�e8��X�R�m:MX�C��-�Ŏ�~K��,�L�C҂t�yϤv��jsz��J{�\QUI�pة3H�B�a�.�3Y��x�vp���	�Zo�,�{�����o���&�I�0'�M%�@��ވ�I�N�uű��G�� i�y� X��`:���6�������Ë�@$� E�W$<��k�1y4[���Fm+�P�'i��1�3��Ëϸ���v��W�+����2�BH��	Y煰w2�XNP�p�.��׀H�1��n���#��F����G3���j�!݅�L�8�;�ٸAW[�H��'�x��oU5X�'􊐻\� ���;��W&{���x�(������R4
���N=N�jB8T�Z]5���0����_=��G�ţ��a5d���qf��_]�2��e<]��;���؞��l �}���W�G.�nz�r,��p���.��k![������ɅB��rД�f�7~ ܻ2�&���8f���d1M@4��ʃ�|a��9 ���;ٲy� ��/�#,�c��=UofK"�@慱ߙ$��z��=�ڐ����YD��/�0`-��2;/Rkyii;u�*�q��"����?��+�zo���r|�h�b~v������Y(���C-�\&*��#�I�{�Ϙ������<�Dz�O����sF��`
�o�H�KʩE��4ވk��܂bT'G_�&�(*�Y��R�E�	N�z�BO�I��k��L�d���h'N6�J��O���e&�)l|��l B�ZSR\���(-��%(Jw���;�;K�}��lԿ)=x5t8�}	]�������I��Y�+ⴐ|���Ŕ��G��o>��Y��X�����A�u�֓�0e�3@yl��}�B�ȠtN�+c�ڠJuP��j�i=W�Jy쾍�|�'���bC֗�iKap��,�m�`d(-9���?���#/�1�@���D�>e�ڌ�%����_L���}n_�:�S(E��� V1X�_�'i�җ9���L(�~-��v��+		rh�ֻɶ�C����N��\������ �w�a���AE �kYy��� h��pC'�k�iK�Y]�\�o�&��Op�&�S�/��{�~̽�g��wUJR]V������;�)��UN�MyND�tMm8�(Ƚ�ǱN���E�τq��D��3������xV,�Z�\[�'���G>��<��.ϱ��C�$�J6�-���?jU��q�YX_�M��xU��yT��0�s~�߸�:���Ř���|��h�dÝ��w���Zն��qd�����t�m~��g��>�Ĥ�t�� ��6���5�g�j$��|Q�Z��L���c[{w�kf�\�C��K=!�@�[����.�R�Û9Fw��5}*r��E⓫���>��:4+B���^(��-C�l��X�k�X!����"&C�tbd?gL"�?���.BM+;5Es*�J�hV�R�WSdk�7lې%��'�M�;,N1l0�V#�r��sϝ�m��Z������F�뉹��R9)���ɺ�I��eE�H�e��<&����5��*d���6�1zRyk�ӿ���u��U|s{th�7�e���E��{�����t4\O�`Âc���8��5�t�g_�t2$v���9�=��!�p�q�C��F�`�S���ζ�O��{��*'SA�t�dq��t��o��
u�F�gO��$O�DWjj���Z� �۾3	��[LaY��4�I��� �%���%U��<�`߆�\a�������W�N��^��Q-q�����ƫ�����_v��#�^���Z>��[t�
B�V���������SXg$�CDԱ�t
� tH,E��=���j���6��R�!�n�l�;�慕�*���v� 8zy�R���J�|�Fv�-F��*!�.p�=K�UTz�';�F����|XAn�=�rhl�E �Z>z��$t�da��_߼�ƍ�mϣ���ӿ���e>)߼k���"\ð�Ӌ�<h��lu�&��y���=��f�6�dS�a�Ǒ�3�cK^�"� %�#�׾��)%���Ah_�|ZŁ��=ztxnJa:�r���j#ԋ���8��j��eR��/�Ŧ�*�E�Y�����{�s�I�7T�◷��(�����5p�\96v&�}����`8�%�+��G+�"�P��{|ѵ�r����q�L��
6),�6�i�#'�3Q��Z�o�,���R�yk��zx�{�O ����=���]؇�y��}��65�p���]+��ղ�����Ƴ�������2�0�>�aX�[ٟ��	(퓍��-Z�0S ��#]�k3E�]�[ʹ_�5��텴/�d��X��Fr3�ֵ��ļ^�"�����r(,�9��O���r�4���Y���S Cw-s0�w_%`=Oi�)/�i� G��n�k�:�G޷���1-�Cve��p5��A�����-N���K�z�(�[���yF�Dt�譯;��ܔڑ���F��Ғ"�eFJp	#��P"u����É���  ��V�5���� �@\��zމ�a�-���Q8�����S�b�2*�ڒ
`i�dIxb)i' �B���25�L�f�����I��$"�f=�����]߲7����bÈ"9Ͽ��j�dK�T��
뎪0��A��<��oVQ����J|Ì&�d& 9�F
M�U r8P"�xB)���ˤ߮�3 V�nd}a�}��IM9�\v��6���l8:=�X\R���j�٤�#H�;�?$�L ��	���-p��Ĭ���ivKt�Տ���w
�傾MAn��xI�F�IszS����xw��2��u�g��3���d�c&63u��]�0��H����am����b�]�A��I
r�^��(\<᝭���#�v��<b�"B~����a����(9�5jm3�NJpq	�6G����03���H��,��^\�h��!�����,�GQ��s���wK�!�5=���������&.��ZQk�F>�֪�<1�]3�;Ǆ���5�$��$M������;2�����]oͽEB��VI�	�KՕ�~��v��{/�0P���9)�(���ud���e���6(�N�.�����H��=�� '6�|l�?��08,�~K(�}���{3�S�(QѮ�r�aQ�t��M�fϣ���i&��Ǜy7��i�j8B�4HŽs�~���}O}�,����f��.U�\y�7#/�c.�[�>���?����v�k_&�}!���H04�����t�	z�c��Y7�_<��n^j�4iK�(��_t�("û�
��h2�=Mu7��hB��������W�8�a�n㌱k�;a���}�(\N� �υ9����Q}����x�%�����*o�VP�
D��a�tr�:F��@�F[�NǱW�Z�^�9���~9��e-���֨�䍼��j$�c�l>�����+�ÝSW���{x��&����֊:�|�5~�+2�U�k���{�-���򳶽���"}��=8s��u�[���A~;���41X� ��6�<�o �3���n�0ϻ�ĝ�"����.ِ`e9������ w�F��m��	��k�]Du����Q�n_(�,�I{�HG���]��OM�����Z�MP��q��=)����RF����'[y��ƺe����B
��x/{X����ן7�tn����$�@��O�(���ǘe3n�!��-��Ռ�e�Ѩ3ϴ������5���M]��E�'�>\�>����{��)ҹY�P�$9}�����9��ǜ�g�V{Q(iM�Q�>��}��qgޔ9�/�Oh��Եv��,�Ƥz ���&�e��N��c�|����n�WS7y&Q�|�,�sZi	��nrK�ނ"�ϻ��Q���؈���E�ep$��b��ge���J�qf:�-A}R�ܤ��Z�^���4�~�;@5Nm���	8C�pT�=R�v1�k�m�&9�HT��cNTɣHjʝ'�3l��ɆD�N�c��޴K�]��{�iO��j,0���)���<r� {�j_bk �����ֹ��ܞVÚG�C��o4����>(�OT{q�2�'�Dk�ΊEڴ��QcD*��t�	t���j���,X�r9���z��yH�	�DAN3���H�D9j3p�@�UFB�ٙ�c�}5~$���ܶ�o`v�
x��sߣ0(x��Ȥ3����A�(����c%��Ci�W�Bd�*�,����H�V�������}��
�������Fb��+�WE�`��`n�~�ъC㗕)"�_�Rh�qBpO���j=-���'o��� ��eM����&>��3�[<�
\�� �D��ےw/'P�l}�N=�����|kظ�ϸ;y2�t7�{���N��$�� ��$b��*��É"�����r�"�B�[�KjzF* f��:Ɵ�T�*�f�1`��{�u��c5ڢ��k;ϡ�t^��I����۬��j0T���N9Kl�[?��)��ǥ��kq5�GF����!����O''�V$��T���%9�l�1����?��4П2��C�s��)��1{��a��K������#D���MSf�]���I����~��FF�˝��>�>R����O�Y�H�j{��7B,��;���mi�PV���7V�� 6K���3ʲ6�;ĝ5�7�u��Εx��'ݪ�硴'8���SIY���،�*�s��)��A�����p�U��V����EdJ�dw��s��L�p��X�_=m��3�����Oe�#��\�>����?�u��;���ݷ�D��}�m:9�c��� �����O��^�.�J�������z�!(�����/����I09�4�ٓK5�P��:��7]�.�4��%U����'�x7[-�5���y�� L-<s�s��t8�So�4�!uq���Ɵ��i�]�W��TľX �f5����T'�ZX�N`����Q�I�L�󄬡�I���ž�	�"�'bq�L�ïe�V�&���Ji��%Z���ǂ��ڰ?4�:������v/������߽�29dWvК�X'�Z9�#w�C�����f��8��kGؿ#��?)Jﮝ܄��}[��x�&�=�Y�@s��6vEm7*��F���$L�Ms��Xe,�fu��XJ�Z*���*?����8��-"UTIɲǲ��rwl�X�����ˑ����F�lx��2b�v�NH�� G�i��b䙤c�
���y]#���[|�J�
�8�J��zB��n3�����B:��r�u&�C���MO2j�EXwiGN�ܹ�?4hb�԰�B':8���_B����= �=����q#@*�	�������^g�?AJ�ifo��b�E�A��]'���ˉ�a��Q�b�D\�I�Z�Lu�+Y��*(��A��jp�h	�S�3N����m%�<� ���ɦ9�}r�p�R��O*B�PH���l�����H�~$mЖ#ȯϏZ���Ki����<�����[ J�M�t�����̳!{/�jZ�HJ�$ޕ+�`����r���>I/5�&蟏l�<�Ҭ���F:�	R�S��Eu(�xo�քdL������J|3�^%����C����u_G@�����0c����?D���Ԣ��-�X��=�dn�/Sx��Ã?���K�| �xt&�To�N�:N�؀���W�,��# ���=���T�;6�a��T�L�(���$��g9c��4	D�y���܆P����3��G���(���s��K�OT�X�k'��6)�r��͍@��
��ǭl90��:V>�R��"�q��U�:��U������;+���V�6b�z�	�7�o$n���֞vrb�z������aY� 0�%�������� ���5ܒ}���t�3��C�7���F��T]�!��ń�[����t�Uy��\�\�|Ԍq����$������N�������S^����({�v��]���	�ŧ5n2[]]3��^	W�}��&�8��ؑ���@B�\�l��-���^�j��0@����/��;j��eH�� � �d<2�>o��4bA��B�PQ�0x�~�:�J��Z�1!T�a���lG�Q��9�_�}�Y�M�"�@Q]P[p�N_qLa�60S�;T;�c�#᯹��0�`^���t_�)n2Ӳ�N��y�Nq9�0�����l<7΂�����;-+~�
���t	�g�̊�O��C�غ��b(sa�5�D�'<������0,��H�](�>��M�j�N��5c���C$Lַt3�]�r_�+���=���1Y�h� �|���!�E̟T]*�l����b��[��ڸ�x!)C��/L�6�憙��T��2��T��O
&N|���p�?¸���Π�Ӱ4�����~�Ogk#n�Sv���N�=Qx��T�<� *��%�\�[�^�»�2�Ս�빢�MI���2�z������nt�zl5;�0Tΰ����d��Y"�ѧ&�+��q�Zc�KZ�n_�g]Y2,B�@�G, >��C�&�T���|�j[ �|fb-�!<��q�w��a4���c��\��0����̚��?}l)B�1o࠼̙8u��Z��G'`��5�fa҆��R<�u����So�@��xL6�{���)�j��	����2z����@�C��Ᏸ%`��Qi�p�i�l�e��l8u�064�1\�hNV7>V�{�ִeY�6���C���T�D�lurp@��c��9�v?R�|��
i�Z�ܫ� �a���7�aI��G��(m�z'���]��[!��*��FE_$�^�z�����?����t��ok�_��AH(�9�=��+�U�%�9�Qp��:�;['J��^6J�4N�<]Ld�R�X-�Ea+�m��]�p�ăD�!��/�E<k2�4r��v�b)#�QD�O��xnX��I���h��֐�
�"��ud%Q��E��K,uu��o��^���JP�N)J]wȖ�H����	ӂ�xa�쇞�ܽ��u�׭9�����0�S3�]�t�W�xY���y{���3}ֹyz<�Nӗ���9嵁 ��Mhv��V���? &<^r�	�O[�OǇ���F35M>)a�9)���6���O���Q�k~?n�j�1����o�Mv�I���Nt�%T�7�Jϔ��r*�Qz8����q]��V�%JN`��v ]a�D��٢�!��ز�B���0��.%d���7wv??�p�?�.ޟ�gP�<^hW��ڰn\ަ��@%8�R�����ӫ0��|_Wߩ��Wt~DB��'|�G����|�Y�s2	8��d��a��,@�ϳҝ�6ƚe�S�5�o]������u6�����p*!�x��;����J�j��~N�6��Y��
��=B�WN`�P4���Ğ��]�r^��Դ��G1�{[�p{AAp�J�WY�O�.҆��L+ ��+��w�$��q���NF:=�=���TZti�cu^餆v)� d�)|5�{/��W��q�[p�΅���&C�'�p�+��1�V��B^���C����7��6� ����\b��J�Ѫ&?xع:�417��aJ�G��A���� �#S�?_
gJ}X)�H�����IG�!��,od�(���!j\ԯ��?A���K��s�x���\-��C�F[�c��| {�#����v�����VƸM4�W��|/%-f���
�$F�gj:;�������s�0��S��Ą#e%ْ�B�-�$����e4�nn%�b��h����m"�أz#���aL��zx_��Nx��J���'����h��߳��(Idv�Hǣw:����j�i>bՃ�{!�(� ����OUo
�Rd9��)hO�P�{�ʋd`g.eu�s+U����]��2��t�i�ol�����8z��6�]�3�
��$��}��w64S�/�[��N�ռ;��dM��yP������Rzٟ��¯ouuM������n��YHs�L��J����pY�����z�e�h���O�=	\�8����6�꺳����@�g~d��|1(Je��mQ�@�\���Ƀ���񠟖�ƭ�׼�x#B �%�6�V�,Ą����K���!���Z�
D��V�p�-�IZ�?b@�Y���;+�>��ĕ�U�-���yM�%���L&�#����	�������O�C���G�eNl
�X�-����5����Ȟ�DZ�0`qF����4�GP�
�؇�凮��i�{f!^���yx<�Ig�n?��ӭ�S�M���]���pvh�HhӨ�ʨj� ck�Ɏ/���'|A�ZG�um�f�)S�_z�O����6��j9�{�u�P���>��e˕/�)F��	 %��.!�Ȅ6�)�n:<�{�+��M�� =�o��`=�%������x��xX]�?߄ Y�Ce-��gnsb^��j�RT�=Y	����	����|X,ҡ�h�J��czFS��Gr�PM�Sf=��_%�CITU����e��c��eC>_��﷞�������h1�zfMN0��J�%��ދO����.���~��Ե��2{�L�j�;_����C�|���o�VM���W�]��k��^et�BO�H��V"�!�-�(#�U�08|A�p}
&�֛�H�)����̺b�����n+�:�T���ڒ��%Nf?�Nn�`*������)�)�)�/>`M�Q<��h��%R�:�JR�$����ǊaY���"�	��SCAX���֎��1�d�>��8�?�k'� �D���"~�k�U�d����z���&�H�QPQ��
��et���<��lb�33߄xvR�{�O�É#�����A��e�ۅ j�����=���dԅ��Yʐjt-4�"n����Jo�$P���l�:��-���:
T�T�+:[�(ɧ�&�fF�J����
�\�Z�X{K�-u����1�I��ŌN���v���ʆXɸ����J����0P�ǒ��g�����V�o�޼9����U���0$�ّ9�)�i�+��E�]Q���(j��g�(/_���2z�i��Cԟ�3܉��^|y��;�m2O�V��4\�R|�}B�$;��ཝ�b�N~;Q�=G� ��WK�1}K7�Z1U~�dه�u�hA�ۘ��ӫ\>iؚqy����1z<�����}�W
�ʣ��><k-�����0�nVY�%�`?�E�'}�9��|t�5�s��1^v�g�_<��uT���"D0�́�:�t���@�~�;`$�k�-Cݒ�����ƿBq(XX�s�g�B���.i��_�����ǃR�P'c*������ֹ<����h�S���R�BW�=50E��d������fB�i��"�|�, �&EO�����[�~̐�����
�X*����!�F3��X�%�[�OM���><^�+�:��� �H�6�IW�!��3�$�G})C��oD�D���_�{|T������lw��� �?]m�}�<g/����p\��SRPf������#E�@.�Q�Ѱ�`�W^�W�| ������Y��V=�KN �@G����eG�x�|�FT��8e�P-�)�r¶
{;JJ%^�7"����u�==/��t��&�.p�8�fK6R���DX����l�?_���B?��E(������Gy)ؐ}��p�d���`u�yuFZ0�֠�O�|W\��lY�X5(���-�S��0y���7�tm��yȥKۮ)y��O�#��<��Hn��h��1�W��dk��-�~�l,]P`�,��]*@.ԇ^\�u�'L�l1dy �q�_���8;�l_)[��|k�4/͝��L����*XG��I� ���F'���:��f];����+0J%��{������'D�d��w��f�� �N�� mѐI�K3��Q�V�����/�_"���:�dV��p��<���i;�>(�X��)�(�6�ԣ�5��f�C�(����/���#�,�TMϫ��<��'�X2h�%(~%�>s*ب)�J�l�6c��V"�&f&�!޷��5�e)�,{����De~J�L�R���ΰw�rm�b��t�p�t{��EO-8�$��Yj�D�����z�ƫ��[��[���;^��.$�~��2M�
o��e!/�CH�->qp�Ɠo߄��ŉ5,�Qy9y��؏KV[_�����,>��m?s�h:7yN�_��o<�E�rҗ�Oc���ľ�����B"U@�Y,� �^�*ݼ�l��M��p�:�B�5�)��4��w�M@����	V���u0S�N����B����X,8d���&#b/���j"����2��1�|^[P.�"^��b�	h�1e��*�"i4�V��*BY�����,�y�)�;7J>ۗ�� ���6�� N�*��G?{�N �6�Eq/��Y|˔z�9��o�E��ڼ��d0����>���%]�}�V�"ߺ����R�FV��pj��m��`P!�*��G�B��g�6O��E�T	�=]���tH.e IHM�J���8��'d!��M�n�x&7ӣ:��b3�����Ӥ�;����7�䯫A�A���X���\�ޭ��9��m�L�=��%%�H�Ƙ鿵�� �D�Y����o����~ɟ�p"���a6� G��b��7`Y^��&�v(�0c1eX��0(�9F&�C5��/�[c���{�(%��l%��8��ɷQ'EJ�f��L&v$�QQ��T�w��F���=tO�F+5!Ob��LJZ����:��'"y�V#">�,��H�����_'�B64����,�,��̝�e11�@G�J�d	u#�i�l~*��\�a��C���y�%I��ce����r?����"��_���rCD��&�  K��^\U\S�-�%�֧��$mF�0��b���m�*l�K�����`>�У� �b�\@3����l�R�IVg�~I�:��$�ugd�r�o
�B�T��G��U�@�N�/P��^�i�+m�k����ٝ<�B�L��n+�I��+�W����}�j:W#�r��-� d�zQ|q,v��nE��nф�
�q߻[D�v�GZ�:,��k�߳)lY�.+9��I�]�r���@V��\�
x����']�;����B��|�װ�fm�hϷT�G�)�Y9*�Ha�ȑ��3��qD�x�G�5�����y.�cK�.���u� ���B�3�����o��5rc��Y���H��G�86���\�����u�&up��Â�����{���y���w�G�{��ܝݟ=R�Z�X�Ԣw6���=�v��f����٠�!K��ĭ�ِ�'M�3N��&�\*�u���N��dF7�=�Q�i2ؙj:p_��Ȅ�����3_Z"5is�5jݍu�w�(��7�.+�^A"��㼌����R-�&��7���F�9�0s{q!�,��ž��ORT��T�*d�lo�7*����x���8�@�;����9	�����:@i�B�E��Wh�ۄ<j`Kq�T�Ӈ
#?d�(�Ѐ:I����WXu8��5]�<��{�K�,��oM6��S	�C�����^=��o��� ��qF80���ft./���JI���ɳ��5�g5�qF����ߨ˻G�-�������cx� ��u�Q�@wZ��d�uJ���S~Yw[BS�mP2��I��O�Z+J�gM[�!��C�/�Q�U���rž�~�}6<�ho1�����O�����Y�<ŤC|l��sx�m�������0(�YY"V��K����� gW2�ӛE�p��dSAҝf|	}�M�7�"*������Cn>�X�9��'�8��U{�U��tN��6�[/�&-�v�E���hj��z0���9{�T��|
c�\�~�	;	����U�;}��_�`gΘ3�p���y0��>+fQi�����}�#�� �ێk|���<6O��i15>j*]w�s����>�׊�˳��K���vz9s��*� �N*N
�	��:E�����>��f떓F��r8َ���Cr��<��+cE��w�j�����/c9\�}���֟�N*>���[�Y�0���H�T��II�rW���)����e�@�4�T��X8BE_���5��R�*�,' ���NZ��P6���V)ՌUHӉD��"�(5�~\�?)�_����u�66[����(_� �K�=�.f�jZ�2KVY�Bg��@���Z-6��da���f���g�WM��W���6����
W#���w�$[��)��}߬�B�Tg��*�9Cg�4�L��*�J�;Ȃj��4D:�p� �A���E�}�<�������p�bGj��H����	�%�y8|��i8`D�)+TWꎃqф�d��,�7����*9�|�M"�=3������3,���2X��_Q
�7]���C�#q��=1Ǒ���=1��F� ^�eR_y�:�CA�)�b\g�m�����-���� '�E_S�N����;��q3o����}�}݁P���&$���D�989�J	�^W���n��������ኾ���īZ{�3�\@X���?\IԱQG��R��^w����'�1�Z�4a7�u�S�B���?��|Z��K`1��8e�>���9���93�����zt��p,��U��-u��ϻ��~ʉ�r�����裸���G�V��z+b~������3
#|�4O���q���{�kM���r���{��R.��
����\�Hi����,��=��wY
p�LR�C�X�Г=#��Z~��������E�*�
gv�=�aJ�k̖�O"n�&9?��7,MEwD19n�>�������A��o)8��eCt���lBO�X��������,Г���*��D+�&N�4�.�(7C��؞�]���\��xYq�:#�r��As愅�R3���mQO¬ޜ�=3y�������+}�­��d'U�Bo�d�mD6l�	�fN��d|kOר�G?�l������5�#c
�;@8vG�^6�V!�ZV��%�F�F��U�Sڼ��jSS�|��=ƫA:�-ͻJ ��c�Y��ye�N���:�`:"O>��5EA�)Q��*m�rKUwd�LOR#���0�x��?�G'#�\z9U����	U��*K|�S�^�*4̨���?���H�x�q�5 �E�T�/o�B����"�����A���kgh?�ju�*������i
9#+�OF�(��2e^���ZV6/�V���bA��Hq.��R�_a,:7���� �3R���s�
�禎���IFeh[er����J��5i��h<��M����"iSs+؈κR�ct�=P����u��esJ�#�C/������K1���W�B� �3bqf|?^��(D=��*_���I�.����� ���T�oĺ
�h�oW}≭�	��8sQ�ʥib@+����a�^��ițIF&6O�sc����
w��h�F.��N��sj��)�J���qF�%� *��:um�33"b��_�v~!��A�^�K�f�o�;_�$:cG*u��t�����K6LP������RZ�R
־����?��.q�/����O���H��qT:���7�zmj�4SU�[�&��-N�}�-Vgǐ�ZR�|0�Zo7���yũ,�*%#�@A~�1��Z�о�e�Yjb���]u��&�$$z�l�<y�<�����
V��o���-_���$�ϟ:46^f�	H�x��G`��U������p����ޫ��W� n]7b�.�"<K�m���S8F���2�ƙu�ݺ���%DE���DO�����{����WVyĊ�� �g�G�t��3Z�L��XnR�ܴ�j�9��O�'�L\W
u�a�M�M�d��4s�
�Hgr�~�Ӌ�]QQ���&�p�!�fh4gK ���2��ݹ����tJ*� �娌��R�^SK�|�/����+��A��oQ��<�=����70&!(��t|=|����F��@%P�5z�Xnۥ�{_iŬ�4�{-�ō;TI�'���j@�&&zb�Taڝ�9{hƉ	b�P=="�_$��H6��{���fQ@R_ڴ�P!L�Q�g�K���$�3&qe��ׂ[��b����H��������MB��8BtBd@�z�b��Ƕ�!t��F}?t0.�d]��_�a����|�}�.���g�Q+@�"L�f�-�g{"1]cw�no��H,.���_4��j(�����oL����	2���:��1��65���N~$�|�vH7�mb�^(�RA����3E���'ev9�s����I���.B��2������1&_3��Y��jZ����6�&�tL�~d���:�ilL�z����4f�����4���3��I��� s0��{��f�N�5��b�m�w|�j�hr4׈��m���I���Y��A�Y�,�|^I�95�-�߀E�Z�w�*�yŮ=�6U�����4ϝo����s�<�Y�- �-��7G�B�ː;��}Ȗ!�fe���u�9r�=]Wl���q����XB���_<X��e�0r������(����k�ZK����V��fV*D����i�Q:_�$�a�s���~���d.S�jM~�
�Ul�Ɨ�ף��2'�M͎�6&T&�(�(io������j2^���7k�N�7��BX��a'9���@��e�$J.��wmF�'���^(ȅ�]�o��"�f�M�����[
_+ d-�!	\��n�]W��;���@��'�oY�Fz�9 �^�\g�ǰ��R��[̈��RIW��	"#�Gք��؎9�2�}�p�W#��!l��f�0T�x�Y��Z=J+W�n�*{HRҬ���]^�UI+��_r+�����vȀ�e�y��>@��L��G�'A�!|��i�FTf�S)��=ܥtO�9o1)�&<a���ԽrX��.!jYy�gu�q�Q�{�m�|���{	�Lv�_�k���G�Z�����(*�6�����_����zX�H���<�� ܔx;�]� ݌OQdt�ҏ]��ř�)��	[~�����b^Ｐ{3-+ϒ	̞�x��v@�Ίa��������x���dU_���Ȱ����fF���,>�:'��#���6X�d���Ll�
w�Q����~ ��R0���"&УU�n_�YO�����L�9�ZM\�p��&���@��?�B��3��Q�L�kFkK�("m&��|�l0���x�Ʒ�TU�"
ڂ�e2�W;��IHN�h#��1�;�� �	ĞzB��l�/5�ӷ�֮Q�7����v����h���4�pP!oO��I��dA�1�2$�B=H��!���ì�)��fcP� R����v4�泱��pO�6.ہ��?������X�c1���S␖C~��q^�3�f��9Y�WɈEM�i�t�����l��]g �.Oz�>�-Cs���g�xYW��R�ԑ�����P\���	�N�<3g)��vg���E_p�>V5��	vU��c�	�YͭiE��$-0���K�xP�O����j�@$�8n�!;��F�ڭ�h����'Nw�:;��\l(��V��ӛ|���q�4��4���5�}��G�`"�:��&��:�t�Iy�Wc�:�XB���s٩\pM���jh��i���%�+ٗ��"G ���:7�