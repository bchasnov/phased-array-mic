��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\����q�?��e�I8�b�Ǽ$��"����ׯ1�V0���C��J�"7���_��p[�� �*�G�j��Ñ�#��}�S}��B����q�g��F�?�̡��^�.�W\�P������w��jφ� A.˞�AH5��n��MV�����W�#�l�owܛK�J��@2�
�?M�3H��
��y���8��2�����0�1p7�w~9����M;����jI)�O�^��~F�_�����W�]u��0�kc~�hr;�LW.E�Jj轧s�&�.`��iRp�.�:�cI�#��f\���]{���:'GhYwE��I��1��W����K���0����m�k����4R�ʻv/D�`�!��Dׁ��� !�'ҩ�!���^Z'����ɶ:W���<<%�{�M���*�q�L�L�6SQ�_WU������2<���g=��g���Dc��A ����-aW�~�f�U����17dX��Ϥ�'d�� Z_]pډ~�$x��ʖY�ʟ��_�����ˢ)H��W�ul�����ܗ���U����v�:<�5<q7;��q+򜑌�&�;(�M\�=�~��i���S�?Cz*�m�p!x������U��Y�p}A������v�CG�u��j�#B^Ԡ4�zR�Y���2�E�0��7�i�E�BJ�t��#JY�R�6�/)0�G
�_
�lN�8�z���ѝ�8��V�y�]���<��@���?����ń��{�����ۅ:���)x$u5N�=��c�8~���D��c��n��'&Yk�C+y��׮a7�Lj=�EC�@�=��c�%��,osHu6�jУ�H���f�~�[�D��_�P�
s~���I��:@��n�Y�5g�����Z�Ԏ|dޕvq�J�K�׃#�3�+B�" �:�\?��.G��B���r�����pY�3���.��:˼z�v[c��e2ƛ��d�Y�b��� �;eo`y��73l���������,�'��4O9�v���1s��yѼ��.K�sj|G�un�@O�O07;��[F�>8����;"��q-�A���R8/���ȇ� Y��u�O�0�z�P����wk��[���9��SYr*o�2����U�R ���`Z=�Q��s�&c�C�1�F���������%�������)凨^?ިgm�BQ6r4�t��@�q9t��(��]>�}a�<��}�g�!/s_x��R�*":��e�ڔ�=���	�T�EO�{YTl0٨r�y;߂=����Mdx��]��>�%A�PWu���������]ߑ��D�I4@K]��Pp.���W`�>��o��7P��B���te[y[�T����0Y�F��l0���3���N!��kj��?Dެ����7��/�6�#�y���;\�ju�smg����uE�X�vA�)��͚q���ǣ9���5��Zu�!gM�T٩J�.�ʃ��i@��h{��OH��&�h�η)ݳ�}�R��
Y�l�n�d����y>��^�g��ab.)�̸�'�&���z��#ؼ���Kw#�$�������������8�t�V�&�o�"h�A�24P΄��\�����񙪷�q�'[�\��<����s.GG�E瘐�V���u(j"���9�	=��s&�'x���Գ�O?�`��H�ӻ ��'�DZ2�r��m�h�� ^��7z��SXC�F��/�}f:Y-�l�=���qUu�X��mH�Lb���V��]�w ���f���U�4'g� ����Ӏ�a�=X �	=�hv�#�̊!���K� ��,��>��y/�p��͟�x^�m[�R��R��1�DtП���M16�䡒����b�#����0�ڸ{z��<���p6E9�qN#X-4;Q&�?adSN�%��XHv�jDZh�����`�pğ���@�c:��1"�Av��1ޜ��?$�U��O!���L���囲w�(���i���=M�i�K|�n�@��o�Nn�4ws8�eN�F�+���;�o֒=�V\]�O/��>��z�n��}3�0�ނN�Y�Zz�|2������O�힃�I�c�:%�J�`�[�Qȍ$]��Y��k��W��}�6��uh�m��W�s��Nin,��s��O��_�Y<+�FL0�����So��`�h���pVb�6�U��u�4�@|Aߥ��ecq�� it�9��#�,�fE�]Y��H�o�HYm���E����i�fu+|ߦ�;�4��q���n�Уܚ������'�W{���Ny��.a�Y}��_�`�Rt��MY�K�kEN}���S���U}	_���K�k Xۻ\X�g�$�}bՓ� H_/T�aF�]����mw�df��j��� ���x���ٺ�N�BW���L�4ڙr��oH�2"�.���K#�:sV|Q�<^M`$���~�������#�LT.:FXK2)1> T��~rI���
�x�����n�b�A�+0��ަ^���a1U�������㻫Z,9YdF{���14=�ʫ+�xÍ�LU>Hq���O7�ڤ���]w����%�6��y�������-�q�$�'*�(?�O���'�r ��*[�`��-��>�q	D)�Q5#��
vk���uGKI��7�;�wU��Z���7Q���O�������f*�Y�[�F�O�,�6i�D�BH^T�G�y��مq���
�\J���0ā���em]z��G�.{p�|>�k�yr@% �W�H���)6�!<H�R�ٶea_�AՖ#!Lʔ��n
���ή헼��d,mt;�:�C��dX2r�6��q��X%�j��n)Y�������r9� h����}-C�x?>�l�`o���)�n��Α��YݲI��p���>���9!r�N�-��u��$�o�����ul;��3��P1:�Z2�KOW�%ۢ�ꬣ�?u]
��}kF��Q�w�"��\XP\��� �ɉ^�L�����R�T;5Ј_8�:������ �~AU1�*�"��.����稿�wO�dQ���@]l"�Pcc��f��$��R:}f���6מ�c�Kr&�d2ˇ+�y���:/�f�"�omJj������mAۣ��~#�Q�J���NM���f`4GA�$_�]��R��y�#v�+�:���H�@�%g$/5�_�)[̀�+kβҽ�Ͳ�UP����»�#�w�f3^u�3�@�9�X���弑�rNvjZ�J\��U|B�-�����S� �ˡQ�f��{��M��$O�}\��=^������Ӄ��jD�e���W(���"�d6�'R�m��k����.C�3���p@T����;�V��`JU�XZ2�!+����Ԧ����>���G�����yh�(0���SE�m��(��{�?����]0���Jڳ|�a�Ǒ�9F�ݷ~Q���y-�齷h�X������.��l!s��r ���UZ�N�$�B��݀��[Ԡ�����]�R/����g!cX�W�
p����?Z�f��O��2f��P�ܝ�F��9
9�Q��]b�/8�O��*%�R�4�] �/N?��פ�GT���n9�J�%<1"�dw�4S�+��[�����5���a���d?���RJ���.ž8A|^�T��㴟�1�k��7W�69ܴ ^�w1N�%W�.5��P�w𝖓���i��q����d���>��O�
��2.�hL4ue�[���!p�ȶ�x-@t
�@s]̼��Ƥ*&�\�3V�6ҏ��ڧ*��2�U��~���0�b����]��F4��M��������y tz/�'7�E��^az��D�h0�ϫ���(K{����G���2�e����[05X&��B��)c���@뙜��/k����4e��	4������h�<�� ׿z�0��&P/�i�s��͐EI����,��Tĉ_Ñ�Ar��k����N�M��!^e��;��ş�����$5�T9�F�ȟ:��.y��V��JB�<'s\�:�2h�,:O]��m�+b1'��y�S#�������Z�������`i�y�я�%k��~߯K��DA&�I�#e��Q�Z�~bNl���z����Q���]�(Õŋ���pa�
�>B�+�t����LR�����߄a�doiF����<\n�w��g�*YA�W��7�s@,���T�b!*�d�/���?����/+_ي�_J�eѮ(��z�Z+���2��wy��,��[2�%����?U����_�rS�m�*xK�\�v��d�����L����Ò�&�P��N�m>.���"j�rre������b����O�ap�
�Z2���լ��`*z����'��{ۢ�(��.]��eH��=h��-���x�w2_D�>CD1:h��,"ө͛��|�ގic�B��ܛ���YЭ��\��<�`t�cf��Cn}��A���Нi
����a����4類u� ��x�$i����ƿ�S�S��Oj�[�OJ 3j��:}�Pc��p��F5�@�q���l��*����.7��P�5Ψ�␴fbK��0p_��UHqժ�W7�S��
��<��~�y�Gh����D;��fn=��J�x�'1�@��:��U@$�MVp��Tƈ����<%�5��.��
��v�-���Nm�(�(r���1�%�e��+J\s��6z4J���Z���䣠�A2��eZjeY�[=$K�|�\i<&V{�h$�nMj��L�:�uLbS��g,��܅N�v�7n�ԓu��8���	���ok��ԗ>��D�vi{\�j��2K�+��Ӊ��q1��h�Z�L��!�ؓ�:�.sRg�S8�	�s�:���8��7T��]d�W���Q�Z�S"�S���Qv&z V�)�9�a7�Fԑ��F�Ou�������/� �o���k�w|��6�t��8�.j�?+�<�0� ��g�ϟ����^rYG�g4�&�����Ĕ(\fϽ9J�ұ����C��W)��/Fc��G����8��h��HD�)��|a���k()�߰�<���2��~�z$��"b$�V@�2i�?��_-p3��0��Nf,Z�I5�Μ".��Ї�x!���hs�gA:�%j�6 ����T���a��[
�$��!lu*�-��Z��z�
5�5�"�M8��t�x�X�$+�Snc�C����`\�J��iNx�Tu���+�:�҂㖽"�������n�^Ra�-�]���ϱ{6�Jz�A��(�5�?=���St�S�����JR��`�<��Uŧ���k?�j̩f��:����M17��,��$#��y��ִm. I��Y��}@�4C���L�X�Zið�	A�#lǕI
r't���I7������`��W��,$hl����j�f��n)�\ƍ/@P��u-w�ӽѮ�N#"U�,䨯_��g�+Ą�԰�m��7f�lYk_i\5O�:0]3��W�N�R��zJ���A���,�"��S��6̑M��emL��-�/v�8�7}����f1��6D���9�}��V����ˮU ��T]���l �N��܎}\Z�*�U]d��[B�+K@��y����2Q*�v�:r��
@	g���Җ~C�.�-��Lx/ӑx����*5E���}
q�Ɉ#���w+Xܦ���6�$`�|g�C��}��Z�ʱN��pT��F��L�� �Oh�!��G�)���?�W�@A���}@\�w��	��>KH�:�X�ڟ�W���8��Ƙ�N(��ޥ)�m�y�Gj%J~����/�TH�qnT�m�5�a��*��m�J	D'2��\9�wS,��5�� @n&�N�"�F\�U#��JF�s���i{������`���~����'��1(�\��V֒a �=aO5���e ��a���ɚ�g��a3�(x��6�LG^v�	s�s8e�,*0
�KD��DK��d����W��Z��/?�cyV���YNܖ�]�3��v=N3Y-z&Ux��,��� �u7(a�q�!��������Y��lW�����	�c�(,����]��̥
Ҍ��E����z������J�w�-���b��&"�Xm���4��U�..��uֹ-�M���F}d2��n�i�ɏ��2�*���N�s�G=X���.$�b;�w�
vi��IT
����eW��B�k�4)�ے^^����=6x�O��Ӗ&�ӗ��/�a�Jk�4
�z�`vj����T��j|C"���^�O�=⚆.3%#C�Dµ�Y�Ԟ5�ϡ���$ŧ7�cj�{_'�[򏶹<�o��1wd�yP1�{ߧY����@�(�?�\�����_�\��)����9 ��:%R�7Gw	�8�xU��cذ�ӆ�><E�=Ţv�%�{�C�l�o�
Jj�����0��-viE��x�����g�����{Yi ���Tu39��@�-�63�r�pB�h�p=	0�����B�ɸ��}�2�?�Gs
O7��W��a�°)O7|-=ڜ�G�#�S��8ߢ�o-�#B��:
���H#t�C(�5��ӹ�i�@{�������Wb�M�/#l6�٫LJ'���$x�h��״,����
���c.	hۈ�W����KMt�i@�.;+DI8�%���Y��@�eP��s��?�\��T��K.	!Ē��O�= /�^������2�E�UE�p���W�7e�9�o�ԁZcLGY���"?�D�C��̕!��A��9^\5�Lo��g$���Z��B-/���4�g�xlrR�o�E�;�?F�0e��z���Bt�m5vu���JQ�En-�/�19�SLX�K�3I�����q��3RٖxӪ������trFG�7�O���F����U�����H)��G�1T�g���Q���cX��0`Ӫ���+|�< �a�c�q��ȯ���s`%������,#5'��zJ(l�i�6�˘,\��	������9'͋�����&AF���l!�[����p�f�;�y�����Ɔ�s��yQ�rq�N+��Lr�_�A�r�%N땸�ō��X��-�,k �������߲ꦷ��e2D�C���t���pw� ���(Z�&B��<��F�p?��Ӷ��'zD����/"X�"��o����ƻ�߂�C�6�yV���OI��nDWLW� �Z7�E��}��k�Bs�����x�Z�v1y=�<�{24�pzy�S��K��屬��ܻ���/p�˅��0�̜�D����v�i�1ʇB���Ho3�Kʾ��#��EBT:oε2�sL�4\�+B�>Ēi#���� �VZ?�H%"�贶|+�ã��w�ӱ��;�!�&�cJ��B���d���\jqD~q��p��� �z�d�a�1��c�G�I~FFn�X;�WA��%�c���u%��0��L$tl�b6r�8�eMv�7YtG�����==��R�}έD��@�FCg��>^$���~ZN'tk�/����qYw���%���T -b�xuo����f*d��&۳�M���D)~�(䋦n{~S��u��nLLHR-	L}��:��^"��a�.��.\�5���J�
���c�WG���x�-D����-9%���7��`�Z��1��ʄ������`̑�tkH|��1�v�g�Z�|�����7�;���x�VV��!��ԻlK+̿/PR�q��Ś����b����#<�p�s�NA���\3*t�:.ȟj
�\|ja|*R�v4R=z.���V h�	+�K�Г�Ie�{�S (�IK��dNOM�\���-]d
ë�_�z�l?�%
  ~��(�Fw4�y�)46&C��N@P�A���V�1 ���C7��lo��3J2��Hg�1����9�� "V�Q?��m�+"�
�٘'�����i��$�f�#d�'*�d�!;X�8��L=}�9q�U����K�@%�������W|>�� �K#����!"B� �\m�jH��w.˘gf��.p홗�3k�6������*��~�N���1�Dfwf=�F���|�Ps�e�=5p�uH��>��������4/��a���^��.�*��I�RO�p�{@9u=��Om)v= {7�ҭ�O�_�\y/0 �1��[�
2NS�x=	�x򦐡���xa���S���#ۘ��m��ԑ�둼�aE�#|�S�/���\=�dd�[g�k(��~ˑ���L��D��Ajk����"�6T܄���j� ��z��j�:�漍�d�'� �Y�ScR�C�o��"�+��Xx��u D]��O�\�!٦-���\�[7nQcn��*�,����q�m��(�5i���7=��Tz�Y�4-���M���O��ߺ��(����<�T������o8L
g�L[�-����E�}���i�zxk*�Py��-���Zi�f5`	$�򕌼6�'ز�v�;Ma��o�6ބ܂��:Kw/y]�N��_.L�����z�{�o�}Ǆ'����3`���e�VG��Jh��!�I��A!�Feôk��~h�_�Ώ�ܐ���}Cu����W�{fpQ�C��B�m��d����3千�@���H����'0jjß����F=�f�ؚ�mo: �b<۷mye�I�B/'%���Xc��5� `y�oeș4����m̱r����2�S�B4��w�m���}7	�����w�$�)_�;P��qzmK��b>�1�xm�8�b�Rܖ�˩�D\���=%(��q=.�_m��K\@�b�z@y"}��n�5y�f�^[�;�+��Q�{P��h���ꉧ0k�}�H�ы��`��.��O�#)��g����q�^�(�?OLF$�uL�e�W�w��\&�2z�'i����>��|R���4y	$ׂ������K�tZ��`Nƕc4���I�WY��/�!�Y�cmE����,�3ķ���@��ߎ8�X\��=\�F�sE�U��z�1���y�'f���W�%6F7bv�M�A��k*�R��U�٨���v-iQJ�"�rT4��wnM_~5�1b���tZBKu4���sI_����!��xX㕋�#�Pߴ^�M����ͅ�N�����.��>�n�0�e��΍����Ae��7�]8�����
a��@����ojC�j�8��0�Gҹ�RҿS�d�7r\���;#��z/���X�d��v�������J��؀ML#{~���K\�:i�o�@3n�m'�ݤ�YI�NQa�L���1gPh�y�[��CI�$糺�K)=gWY	�FoH2�hg)J$x�wr��P��P�4�:~0�R �ȵX�_��k�b=ws��[H����𿸳E��6�	)��o±·��-��]�<�Aù��:��lm�\�K������C����A��˞�^'�C&I��c҃�E�e�v#i�-enO�\��"��H����$(�r��8�� ��&7�)j#k<��U��� �6~�!k��nc���eg���b����~g̸͆���x��#�^Ѳv���Iq]����D)Ў$�V{��6��y��<@��<e��Z�pH���B���(*!�))�_�)�X���7f���F�`�4��jn�/���\)i��&�6��48����MP�I�b7����i��T�9���=�_�&['�+V6N퍭j������"O����
�;��Z�.л�0��ޓ�O�d��_'���Üܫ�T��.y~��kvܟZ��pN��z�6�5o�{�MY��=����'TL�xu��Q�8<�L�V���j���PګΚ|��IU�w��t[���J�E����7S<��GHEe�<��9�R}�����#/V���vB&�& �ēS����m�:E��ϐ5.�W��M��)C�	u� x�h��s̓nrԔ'�T�"*���Җz :�n��b�iL�^���W�����U�"\'��O�,
0?x2��yNN�C��!b�����������cDޠ�WXH��i��\�A߸\�{{mq��Ft���>����J('��8�V#�P���۰�a���${M����i����߅�Lq���m��xj�)2̥�u���}I�Mv��-)�j���={̭��%��!C�O'���š��AT��>~� ЮN���	t�A)��VX���9v��8\=�űq����a������)��o����X����ط:���ڣ�3��o�ó�\`�uRz�	@z�^X��V���[�Z�t�����eL$��������do�U
�)�x�|K
^_h��ŗ���t���!�/>#��c�R �9B=���W��=��pf�:O=�R����Ȗ���S����n�V�þ�d���1������� z���]N"?��`�3��i�f{9P@����kJb�����g�<�L�\y A;G��D���:2��B�TC����x��G�i�*�H'����W�O��錒�mꐄ�h� q��X�hҌ�v��@n�k����9�����ϴ~�\�CJ�,���ܞ�}�v˽�1 C�;��k#5�Y�U']���	��!J�C���l�Df[K(ۿ���QC�� ��4.����A��%I��z�lᇔ�@t���!�NBe�`YZX���iF�4�j�cǃ��` G��'1��^U���l��oQ�:ԣ,`�^]�=�)k���j��O�/4�`�
1�G��f%���{�qcJ9�AS���
�뇠$1�su�eI7r��f�䜗�� �l��Z��b��>T߻.�3���=I����ݹ$I��u�fQz7�LZ��ʗ�$���J��xr��'�3�~Ka �E����y�q�WG�G���E�eA���h�+�sceA�^9T�ۮ�b�_��̍�_����i��wI�l���~�������/??�{
`�
z#|�~w�uzǸ)�F�h*pQ�$~�?W��M��FN�Ȣ'���hc�Ѕ�uc~!߰��=ǦM3*�vB,衭�A֎�� ��
i����u��1�h��v#ƾ4o�pJ�8!̄X�lѸ��,Պ1� ���Z�3~Ekǹ���1��n��@��P��LP�b	'�@�b3�9AO𴣅@��׏M���+�z�.s��Z+g�o�'��y��c�[�N�y5F���8wx}�N��C��Qg��� g`��ҕ���(���՗����ڸ'��$���5ؐ)?���pK7=S|+�f
:�N�'��Xz7N��o&=Sy���e~D:�A-%�2e�9�j�3��>x���a>����~����\�uR~�b��A���V��NSЮ�W5�LL8���/1�J�&\�!�R��eBSȕ��Y��7pb���[��q����']t�y�����T��L��)>�kǏ�5?��ӣS�Q�<��e�h�T_C�q��Ԯ�K#�Ȣ!�+ʥ��CZ�����g�@i+�5R����%2�"fl�؏d�	�������d�c5��.cW�V�%|߉�ڮLO�d `?�ű�c����l���	 �D ���#G�@A�A0�Q�S��J����Ծ�I�����r�_͍y�d֍ì��,� �V�8�K����1-^�-J��q���Jix9��&�,|�[Ҧ�<��	�kϷ�Ѝ���8`<FtKnρ8xSs}��X?�es�Q�鞘�&Q�� �?���B������4��Dt��U�n�Y�-�r ��ȿ����ڡ���|234Q�s֔�n�5�W+��`=K*�~���
m\����F���O�"�Ȋd��u�P�Ş�S�������T��c�N�Kov�a�`s'-79����'��<�U���6"9�������N�5���&%x��+
�+ՄWu���!��A$��y�g; 5u��r��0�?��� 'q�4s���R���Sc�DYy��&�H�g���n����Mt,&�����{P)��������쵖D�g�E���D,�~w�A"t�����G�����?��q.|���*�e��P"\���F6����^�K@{(8��C�'>2���skic����7���w��[��a;Y��J�=�l�n�hGipo�B�0�\�h��!��HoI�Y'�BNZ�#�<˟d�+�[���1%�BN4��9UR��]��F�[Ggm��yD0���n ��]��|2�utYٴ&3��z|�s��P � YVBh� �m5<jWm��mYx��^=�h#�9�!
��<��[Q���f�sS-�O���Wx~�2`���ŕ����Fޱ��9s~�!AU|spM�K�߯��jy�����ӣ�[��MWaE���t��
^Ca��qD���KnnBu<x�}.�j�&=��I�i�����?(��e"���yT��D�1W�b���v^��?F��� ��K°H1����͢��$�K�h���x�n��P�����`���<�a_�c���׹d,9�}�{~_��F$r�D+w�QfW`�����o|u�ϙ�\?���%����Ն�7d�_o#�%��~�KL���D<d��(�Q	�3q�ma�K��E�m�90]�Ѩ����Ьw�Z�:�d�4���2��$bAr�H>��Π�� ��>W[	�y���W�8��\�%���+۷��+���-8�L����2��p���-=Y��Q�?ی�R���DEɾZ]�L3��VIJ�V�<�HyV�uH�,bgSJ-��� �D���o��K�kj9&�!�y���V��ϭ)�3���={��7�+b�� ��'�H��)�Ad�G�#��.���'����2��BIo�$�����D�淠jG���3�����W�t>	�4�l�S�} cT��:h� �]�_E�iU��v�j�d�+��ɿ%�卓�C�B �0��9��PHj�9։����M��Ϸ=�]��tɪ���U�f��R���vĎ��lF6z��)��$#H�w1a!ٌ%zh!Y8�ydrn�cm��Z��ɛoI��ʣ�<8$��p:-.E��{Gg`�i����ˣ%��v���5/Sz\��:)1xoo�����1��,�"��Ң�c� m��dMh"�͘V�f9�m�jI�Mim!�B�_�!�z
Li�ژ�I�[��ǋo�hd�?r��J�XbjԚ[8��O�̘-6tyw�C[�#>�	��-4t���@��D
��9��+�f��R�NI����u�;�)0<�2��j�Ξ�-Ў8^X<�!���"-W!�L�|Z��_o��7W�T<(�5̵���k��d,e/L`��=�^� ���tJ{[�"�f���D$�8��Z��m �v'�F��$5�fͮ)��(upAc� �)g� �jN�����t����4���� h6����DN�ө������h�~c����U��d��g-q����<%`9�X�%.08]�Iѱ��/䤁[P?�ͳ�J�QU0�ΊF��� ����*[�<�{13�>}%�[��GP���)`n����Q�Z�y����G�m� 8p,zDA�UWn���?�I������q ���Ĳ`�Y�����h�؃w:������A�a�GL+A����7��z�,�/)��ƒ%�H�F�31�OB���� �������Dk(�BĨuF)�H�W�p������Ѹ��)R�-E�����PNY�Ӎ>x!����#�G��5�گ��73v2+ax��PCV�7HG�x;��k*�]��f��b�
r�	<�ؤR��p�j��8\�Q����/��X1	w�YC ��nۀ�H>D��F�uB>�]����n��7����}�5��i��k[�:�����W�0�@I�����v5�y֭1�`]�Y�(r��a2?�~�X� ˊ,����F��/�aς�6O�I?/��1`(�g,�iE�̥�l���4�� G%�%<x�!�\�ui�YBdu�%u���/<�O�F���*�5Mm��0^Q��k�6��]ø��Ĺ|C$Bw� �=aIq5�9*���ӣ�(NuA'I�!<�r���(:��*��	3�&�`����:u���A��z"�D$������.1�`7��C^����OI	�]&QX������8�Z�8� K�-��~�6��_dl 8��=�l�\_�;[��s�@���t&�O�{�`�B�~<�}ՎE���|:�`Ωö?�v�H_�ws��ݹ��\#n���l'������!8������|�&�)�U��yrϢT]13������L^<u�*}&`����_�S�'��T��P^�kҠ=Z���ՑaS�Ac�\�A�اE��jF�`�H�z���f��^G1I�L`D�d�����ۃRCsm���*o��.b��P�@v_bu�IǑ�I{��v����j���FH��K:R�M�d�\E�%�~�w����P�	,����r�� ~��l'�f2B&������!�C���MM]�l2�}���X��i��W0�s����@���3F�u,S�M�	^nu�tz�^�8��MR��j��QRh�4��0����G #gSb��u��D�U��ǉ�N�z��������k�`1K�������5M>5i!��y��`U�@�Ї�3�)h�*�h��.����7y��*����"�@��ordg�w �g��Pqz��7�&��H��;���غ\"��#4��8-Z��9��*k<�9c�-cZ�4ztߝJ8�3i���>���{�fvN��F\�E����a�P�VM��h���'l��R���0N��R�]9����E)��[u J����g��4b;,[W	�
�h�T�һV���N@���s&����8ƪ)-��.#�D�T����.�U����;D4AT���}�~���#�ti�.��%�?'K�ĢE�OU��Z2����p���t;r��۵ν�8;F�Q��6��V�j�`����F8�e9Ny��HZ�״�{f�2-aC�$������x6��g,����LEO,X?�Y���'O�"{�hh�%�ECVM� zRu���5�[(�y�!a"O�~Ur��Wm��T�F20�P����/,�X@`e�B��������fp�TW"� ��̉o��	�/�@��2�#��"�s�'�g�)�\z?����w�n4Q5lW���$�)�,p��V����#�7�֭?ln��I1�R?p��*\��׎Y���!r�C���8m�T�z�X��ƹ}���/Qc���H����� ��P��Ɲ�Oj7�����#�A�-8JrG�f��yѼ˲��aWHE1H�o���*L(�n��N�Y�uΚ��[o�u�����څHZ�J+�m~b�&nzֽ�z���wPۢ�� �>���R�Е�剶��[�H��]z���/9!�Q�|�%=��`�F�D֗`�HZ�6ߴY�fJ-\e1X����X�IMT�U�0�0|�r���	+��^����MUŏʪ�;�@����c.LM��R��md����q%V�0ԡ�`8E��;�e�
L˪~��M�ࣣl� fD�v��o@6Ѝ����_	�81� �ݲb�9�Ӕ	oI�WxA0����6G��9�x{�Y��d�H��t�0�؂���A6>�^��4o%�Y�U���z4��M��<��'jV��+��T�K9H��E�L2];�"H��q眪�YK�Q�=��֝i4�H���հSF�׿*�`i?K ��%@N��˥W�khr
�{�E���YӺ\֌�>�S�;�x���m ��f�R;H{�[fC#E��}\3!wshE�����r�->
���q�~E�:��!)(#�y�l�y� _�Ϭ�kӰ�NT�ш%.�o���&���@��9�yg�`���	uVpy��ǩ��~�nEkC(5)�+�ҁ��Jn�Y���Fp�=�����"8��Eƀ$L<�j�=ʲ��E���d�#������G�?���0գx�=���Jc�A�0�߅Z�J���;z���ovd���h��t5�f��&g�p�*'��'���\�o�/�v�^Qj,o����C�zg� +B���r���ذ������؇+)*v��[�,=[s�S)��A�~�'�W'��X�/����Y�����<�6��]"YELH��txWC��5�����G��y?f#��_s��;�n�d<"�� �O0��X���9��d9Q�Z�V���L/��������F06�]g�<Σ�˽�ג ��Z0����o}��,fm������E���ۢkr3B0�j�V�:��n���/���R�ch�
��ڿ���P����֏��g/�
GR��5}��%%U�b�yq/����Y��J+2�_C����>� e?T�؁	E����w�!6,J�ЌE)�S��4���/7��_ȋ3*�l��'��	d噟"
#����&�&�W���>��ì�JN�B���KIVW���$n�tN򯒁Z(S�v�D[��xށ�)�6��,��%a�oq:|����'ɽg��� ������.�X����)§�����O�Pz\���C�v1q9x؎��Uɖ����k5�%yuk
��U�]���|V�����1�Wġ����8j8�Z������=�>Ѫ���/��R:10X�O��$��aW{ğH�s>���pW-�)��h���I�c���4Hq�Uu5�VwXv_�J��h�o������J�!3��	�r��gҟ�m�_\��|��s�=�%�@�CL8ш��Y������Y���־`);�[v^B��������8`ѿ����� +�~U��@��Б�K�����֖o��L�l]���[G�b~�.�u���r�z5�VR�^ϕP�q�u� �?ֵ�@�i2X��Rb=��;�(h�<���A����_�|Ŝ�-���B�j)!I�2f޾�nQ��YְK`�'�����+�ܛ�Alwt��+����9/e��2�����e�~!�1yl�+��7�lCY����|n���?�qR���g��J��u�K���>#��"Y��;F0�Q`ƕ�ꪄ�%�É؊��
;ާ!�F�'0��R���Z�nQ����ڑ�뷺Pn���.I���~�z<@*�Ϧ�z�ӓ�=B���g�WQFQl'��3j�'����A���oq�N

�M��L���	���`�s��xӈ��#C���ɐ޺�ٖ�>��̽� |�S�%⨤�冝�MN��3x��Lf��$���ij��k�G�闪x��:�>�h�Y-�oz����j�ST2�|�^>KZ�#��p��Riɶ��ͻj�T��2��}{�g��&q�wK�x{7�������ZT&j��0H����1�x�_�{ݢ(�2$_y+n����-�&~���))��Cy�����-C�Gv��Л3ߚ�lO�"E���L�����ĩ�0�/���O����DZ�Ju4���U "�^���Ik��Bcc�E���d�yQ;��YgT���9LM��U7zZ"�s��⋭����X�=s��n`�X����w�Uvc��cŞ�ա�r���)�k�6jd{�A��\�e/�D�Qv%�t��_kbxj���^ޜ��W2F8S0�N��u����C^k������K��4�wj�N&	�V����bɕ0����������Zs6@w�L���"~KTĝ3�!�<ҁD���nq����'�r��N8X�bv)� �����Z��B�ib�?��8qY!t�4�H�ZT����|��j�4B��ޙ���|�Eab�J�ڧ#�)�h��fW�����j. A��Zlĳ�|C2�(��c�S��_���ҡ�<�2ү.���]�r֮Q��&����qǡ�spoq��r؏���s�N�O6�;���ARN+o�H���Zme�����-���4�i�G��ys�����$P!2mR����}<H�ik�Y��#<��Vk��w��t�zK��<'D�|�v!��⸭�_����/�,��Ѳv��a�d�= ��Ϭ��g�RGv]_o��rHe�l����Y�倇"�`Q�U/n�;�<P���@����:?��(�C���,����+�����'��{Hdw޲snQoE/y���А���$sV�i�[��*�B,�3����$E�c�z�(�&��X<�lX����E�3<�v�Hx�5 �y�tl�̫E&@A���p��P�V1��6����~eh�)ʯ��2��IA��mN�!I�����z���Rh+�ȣ��J<&�yx�om㆞�J�{��(;A�� o����� �мz�kC��Fnp-5"w*��\X��n��(�����
(�Ežt��K��g2��ImH�>�33���C�֑ -��6	4E��z%4�GA�lq-4�H-����Y8�mA�!�Q�� ��t�RRZ+�y�WR�߯2��0�W4��B
�^��� ��`ƫ�EN�|[�M�t��y­�8���Yc���<���S��H�f�M4cK=ls��Ps0��C�8ןZe��UH#.'��#�&��IO�<Q���OF#�cJ�91@ѕ��ۢ���n��M�F3`��}��i�ڈ�}����f�.�F@�&���o�g�6v�^�$lʑ��=�\2�?.�O{����Ѽ��W���JqeC��<f��J`��k@+tQ(�PB�u�ȽXV-%�[���n��;���=���&@>��/ie�J�7�\��&�W*\�F�`�)�\��T\�U�Pc��U�M6�5��R)''H��Y��`�UğI}���ri�a����:"W��m��� ���S�s��y��-hoݖ�k�
݌g��-��0��	���3�si�����X+��?��彋~��⻉�L�<FCѴ�[�H���<�y�f�?�yh���h���
�8-�Rn?o��0rc�T��e�
t����DoC�B�֒N:M*�]�#S#��U�A0H�
�!L~&Ͼ�����FkȤ�Q�:����pHU*�9
܎��N��˚�=.f���p����wꩱ�e5�ES�ĿwGX@ͭV\l�(��������&�k �[U�i��Q��a^��^6�E64�n�fd!:*�Ί�\�9^�Q��"Ҵ����5	�V���R�(au�^�>P�$�Y
:/���+^����0��Z�]���5���;.�	���Ż1�����h�~�����0������X^�	�Dɹq�knt�j��)��:x��K��k�QG*�}E���!��>��&��Q�6%a���+ɶR����B�FM�����F&{C��K�j/o"�[�$�J>�#I?>&��\�\i�Bm�k\E����{�X|��3:M>1��3�A�m1�6����n�fP�Ő�1	���s7:�!\��B)&aH��o�q�|g����i���_��i���f95�3e#J�\���S�\� �̽Ѡ8yD�m�d�?��@1�9�\��N�AH����B!)��8�=_��x��7"sƊ���^�L�A�Alx��[^s�,�pm֑XgI Fm�'�&����#QM�ٺ��v��	��������\Y<G������V�OA�E�g:!u������.�6\���'Wb��E�����E�4���#ĥ���r�G�X��hVV�e���`'q4Y��P��Px8g՚�K|�]���
>c~~ +I�uq��$���~���a��H���F5r!�i�?�h���E�T2�|�m9U�EO����.�L�[�?��P0�����0ɮ�2�С�#��)�i'�u���VI5}�$���u)�_x�×s�`��n<�[
t���Dw���3����IMAe���]��U����O9��2����hO���d���,Ue�EpLf�_P��t�L�-�C�?��t����&��f����~㙽�ױ2�?�g����;n�F����:d*2�2���t�,�{֨Z5��'SR^���p�u��I�K�~������<�����袕��$���h�tC���Gh�x�#? @���8�mZ�?��i�DA�t����##ˉ��Ɋ�Qp�o.���{�-W����������x�"��Zd�'������]�$qyh��7��^�?[]ň^�ל!�����;2j�İ�۔J��L����$��T����h�G
D�s����4�ڮ�_&�<�x$�2>(�Q���\�FdY�"���۴����t��8�ňms��
?��1��M:�a��A�]f�ȵ��*n�>�Gt 	�gΩI����򠟃3����v\�I	�.�nc͸Lϓ��~?��5�`��u��ƌ�x����I�Tr���N9����䶎p�����&IE�����U� yZ4��mw��r=:x0�xc>s�e*w�5�)�W=+�0���̊�_�U~�]�$}N���ODAߨ�ME��������M��1��ÿ��**M`)f/����������g��� X�[|�s��Wڐ�Qg��82p/vm�a��R\��t�/��=~�"� Zb�y=x3+ �ο$�`ZYY�@�C�+?h���o�`H�A�
h��'��,�SkP��Į7��r�uČ�h�������oNk�G��;��3@�7��ՀdrD88=������4�j�j��͹�l�2���ۻFF!mLd���?�̤{t4
t�FI2�|t�u*�\�_K�T�� �R��:�D�ר����@4(��ۭ�'u;v�n
��v՛�E�$zŭ�@�`�3�	�jf����G�������K���p�V��.������<	��@��h��H�yV��n�E+�P�GS�)��=X����㹯c��yG>�g/·"�����E8@'B�`�Vs�e�K��##��S{!��a7�v�'G�-߭<�D"�2J��R��"�O�^!��U��
q�P�⯜/���do�y��R&��PW�l��Re�c�$YJn�a�F�K��>/�'vWf�E�)�.�
*�Dc�TZ ��d�a���O����6�iX�>3L��wȤս�e,.%����{�3l�q�7| -���3�KJ�]�\-Ң�܈X���̙+��{F]�ߙ�g��TR���1��XPW+�G�B\��t���P	���=J�|7эK���~)��� I��z�bT�f�> �`�A��,�3�:|��ɖoa��k�dK������sF_�+/��At���,�]{�h~�B��y]yl�		���WO��j�3/xz�����[Y�x�K�ۮ�e�!�.p����H����V�j�����/Ȣ��I��p��;[���+�f���<3b�7���^\�k45! ������4��JbEȇ_��@�E�%]����뵿�9�ڭ���.�?��Ќ��.͞�;�$�Pl	��,��"k'%�]�a8*B�R/��J��K�y���䰿ՐP����k����=��r�IN��8&�5v��G��3�i�7j�ZbId��q��c��EB��e��ǃcg�Ke������nq�;E�s�,F7R#Px͆���6�%ς	�TU��i���D y�o��f2�-�Z������"H)��w������R��:�1�T$���r��J	Vd��z�:�==DrП����+����A�
:/�h��= �wu��3uݓ��7s�12r:]b�yh��14��-���]>����3D�SS6�ۂ�p`����^�d1�xć���	�ZI[da�4{l�"N&:e/��m���}����+P��b��,c��-Q���p����B�UE�6�=����b�� =p�>�'gxƊ��XS���ȥ�7
��3���&���k4��b!�?ߢ���I$ɞm5V��䧘lS���B}n���3�l�"��x���ņ婢�� r�-
�H'����Z^�f�=��[�����U~S{���R��1�����)O<�a��s��m���Y�H�<�&�l�	�πuz	��22̿��D�u]������j��@�.V7$L��`���Hʿ�<���F����R�ԭ{�X��L!���CAR�{+��U%d�%��p��0��j2��m��?<[]Ql�{�yK� 66��+��OXd;,3@s��OP�O���\͠�b��tNsM{k���г^�, 4�y�*��u�Kja}'��ΙH�,�|�z�ʵX��y�b�c它�q�c�`Ҭ��jq��_���Ûtn�����H���G��M��걼Q)i�9_gTCߗ�=�X��-&�#
�S Ʌ�^ORK�����י�!���D�ǜ��9��@VK�:iF>�!��b�o	o��%�]����x5I��e]��d8�lw���~b�X�����7�ܕ����N����YT�)�J�Z�j����
6ّ�u|�<�T�xn�H|=�|�]�����d���#���v�����c��������2�������)�+	o�P�m�����V�[����#m�=2�)1�K̹�C?.��k��d�Fa6� �/r�3��cE\/�cs����*��D��K�oxY�`�"���x~@� ѹ
���>S2�@���P�ƦG����>�yjy��(��$=�G�=����L�k^�/�����x"�[�X^��px�JeW�����A��S�������%U����a�6�D��S�t�bs��'CH��e	_�������g�	d�]؃�Yҡ+Űe@�Y��Iz�P��kũ�y��[��U�)�����Z���? J;�x��Q/p��Ip��()@
�����|�iO�*�I�S����ŪMۤO�8���AjЙl�<x̣'Y�"���3�-�8��-��]�Wv�7V��N��)��C�j(DT�k���&x�%a�
C$ǡr��m�����ժ�?������h��ܷ}>�q<�Sh�^9޲=>��j���2Wp�\�c�w�A����縣�C��$g���5�)�G1Ȕ(fC_��Vs�joX�`�����Ƨ_�"�BM��EII^h`f��K��h�"��������]��>؈�<���9��F�2!�N�;F�UJ[�I`FDe�G�?@e�I�unz�N�'G/Q 9�
����S|����4���[�'�5/^�7�����d��2=��T�����؃���a�/v������%
5>�7^���df�趥!,v�ՠ��!P�_b�;�B,���nJ�,���ik\>�!�XG�+sU�E �?���#h����B��햴����툘�AǭN"s�ЬO-����������-�%w�TU#$�<iV�H��h��r�\�����0tÄ�r�U�(ܚN�&5 ���J�����	y� �.q#�~��5v��_���̫y��a���Sr�pY��V�x�F�"�Ǔ���d�!�
���ѓj�c��UK"�fn�J~�m��֔���g����(r�O`��\$U�vOwa���ϧ�)a�ߧ�T�3�'���������?N���ű�A^;�R_�\p}Mg��n���L�3�6я����n�S���9fm���J�b	Q
��TG։_��вB#��k���7�a���	��a��eޯ���`�^r~� 7DL�[�Q�S�7�#߯!ӄƂ��х�o���Y�>d��ta��* !�z��ڊ�[���"׆�����H�,A�H�f�N�="�'!.:� �R;ݳ>_�6S[�V��Z���x�3�dwz�g�������f�U���t�Nّ�]���N����#{��Z��~O�Y��%i�؋��a����!]��
��N�[à>m��PYePoCG�kE���,(�`���pK�^��y��u���7?���ވ��)I\H��'��QJ1���Z��4|��f7%�)������[X�A��f���b��3���I[6�";�b@X4
��`�c�}�o�.�Ts:�d_Z���!�Ք���4��{8�}E�*��j��+�B�M��� �%�L!��v}Ī�g ��N_�'f(��P��KJ`"������:��`7z5�u��vڏJя�j(�̩	)�/��� 5G�06�v��q�;��B��:P}���͏��'��b��y�w�����l�����O�!�+��*x_w��=0PPu��4�6q�������m7�XN8a���|��!h���2�KC܊x"�T½miP�1J&�W�I�Ĥ��O�}9}�L��+a��it��|FT	���(m�1�G!������T��~��$�׏:�$oQ�ލ+�Z6�K�z3ƅ�6N*r82BKP��jaN��C��_ R��ϼ�!���"���Z��������|�w���Ŀ-֨	5��#�&} ���^+�r��x���9��3D �>��f�~zسZ����|������R `��D�� �uݴ@v�5x��\z0u�����şUx=�EJ����XXm(�u�U�-
Aoس_���j�օD���z?�:9ߑ�;���8N٥��"��*;�k�iM������"��s#�=���C�6�A�3��E�����Ƿa�J6�Z�v���k<p�>a��!qqN X�Wd� �i}�Rbk��{�eF�Y�)��W-޴����^� ��'ߝ��XB�z�ב�t��!T����۝��4v5[qw'ʖ��8�I���>�q}f��R��I�w�f"�O��j ���$���Z(ox��)�	��ݕ�Z@<��=s6���[�u��:�k�o�i0IN�ۥ�zzح�̎�F�L��Ԣ�9m=NBR�(4��:Eh���f�8���̹�d��;\\��snMo+2	o�1�3�U��&Νu��%j>���HLfŲĒe�>���_i؉,\��Ή��(_Λ)$����IKyō0��y��f#"F;��ܫgDȭ1��M�)�lAD�.e����ҽta�w����n�w���S^,E�Y;}��H/!hf
t]�F�rV�*^�}���q�,T�.��4����Qj�)���m�7]�vD��̳t,bEd���`�~�W�p��+M�G3�?Ѩ:�0��X�~l�V$ܕڢ+�������$=\���CLU�#k�yqG����l�+ �y
�M�	/�'��~8�w"��!��'�� ���%!�ZkJ"�ٮ��K���EYFB�v�0 �.�3��mw�rr�PL�_n���/T���E����_��Tٹ^�$��3��
 <��޽�t\��TX�]��㷖��36�L��O-<BF�U���!�L��]]Q�4�+蠃�mw�:��߲�e��I��i�q5�F���rj�ofd)�s�?$��|w�A��r#�
?�m�'T���7P�܎+��E"F�"�)�Ч�j�y�	,���M� ��f�>�>����zU0�4s�0���՗�L���(���9'�5�������x�/��&׾Tg!F����N�T'P:E��\=[즬�4�б��Œ<��$�"]d�&6Yo��PR;f�F��~Aõ����bbd��=�������f� �)l��{D������^m���J3��Md�ͷ���{�/`�G�-a��jcZgAA��~.HFP���z)��3�&'����u,��sk�*J��Ȱ��.�N#Ǟ����FTZ!���l1�ՕB��헙��k�O\(��&|�^���:׹�H��1J�w��ҷ�-&jQ�u�ݟ
bq6dP��:�[G�C��z��ho�#!�gH�vq��M.���)s�o���i�51@��EVL�#����v4]�"��ue�d�L��d��S]��v��>��;'27���"��X���Is�g�/�B�.:�p�~�>G�AJb�
�pU�9]�R�����T�a�[� H\C&R@�����^�kJ � (󣙠�T~FJ��r�9���Mq��g�W'"�ol%$�:���׷ ��Bʋ��uO���R)k��KȘ�G���v�o�#-u�F��4�[�t�r�M��O�0q�H�`T'��ҦҶ�B���}Ыx�$[g�[�C��o�8'}�ؗCN�$}����V�}��Tٵ~�����Z9,Mv)�<t���RgJ(�\৛����j=�7Y8�{d�;+e#t_�3$��r2��&�h"� ���آ�Wi��ߣȱ�/f���|�VE�u�`��?��U)���i��/�M�B��'��'޸E�(���f��:up
d�9�?N��ѧ�������*���m�*Z~�t�<��Q�bJ�3�R��rb6�4X�m�y�x`��&�'��ebS�d��.ic����`��r8��� ��%	�I�,EV���A7?�M(;1��`e�#dRY�$�]�ܽ���AX:�C/;;�G#)P#9����O%���6*]?{9�H�>����Q5֞.ᘸ���a/7�KgP9b�46���w]={���^�M�nN�?o�cѧ�ʮq�Q��J��'��pj� ����¯��4*�.Y,M;���>zt��zzt%vd�a|x��F�4
Ʉ����'��+Ğ��AjYpdRf�L��+����j��	�j��a��3^7y�Im�����F����}�WCK���<��`�g51<��@ӫ��Ά8G����;!�鍉�������Z�+W`8fE�a�@S���ˁg�xJ|��3������JK:�][e9��˅����E�k�~��t3i�:=B�8�5�X���NW� ���<��&JxD;��-o�ҥ~8�a�Lt0�����p����P����s\����>��t�ѓgC��i@R�*�Ǖ'U�SeJۭ�t���Z1��ik7�u���q�xK�k�
�2?D��/w��o:����(JQ[�NC�������px�צ��M�ӱق,�d!��UEh�Ȓ�U���	Ѭ�,gT��i:�C9x����L�u`�/��|G�_�k���ۚ���KG�,�>�_*|��G(�{�p?�Cs;U'M�WM��p)f5�$��P���#EʼKj��A���~�~qg�ih�:38j}ֆ�ynp��%�o����\T����������h��V3�3tV}��S3�5�<b �!�JP<��2՟��,����~�=z�kv���'��fB�g��ݬc���
�Z�(��xC=����{��  s�3t=uʎ$p���������Q�ᬊ�r'��M�*�J�1���p��-������ �2�J�&g,�Hݹt�iG��K���"w�I��_���&����׏�4�LI�Z6<q2^�2)��l,��y'E:yk��7vR�� �� C�F1ɧ����;t���LE�Z�j&��T��ۯ;�Lҙ�iG6]�Kc�刉H�″D,P�~��$;W���<��~m!��Xe�{G9�m�E��+ͦU�qy�v8[uߕc�V��Kw��p#6�g?�KP�*em�ӪG�$NW� ��$~>(邍W*v��%�6�ƅ��+���{M�w��~���Z���חٔ��涫Z0p��+{��������h�FMo[Bվ
�p�<5����R��y�{m	�Z���/��C>� *T�W� �u�����5��W���	K���o�Λ�YL��P{֬eC�تJe*Sy��]��\�u�JS#J�I��������<dҳ|��u�yU�w��e��:�"�ĸ� �-b�۝�jњ�|�M)�hװ�P �CA��cw,n���@UĭS~���Y����hG�RD4y�mu� b�Tob|f8�/��_��Ѯ0�		3<�kgɲ�c��=�X��Y���+�A ����������fi���U�gY�
4��5~����bڰ��HTw�#����	�	�A�&��VE{�Yͬ�iž�?��N����l��Xg�b��E_����&Jh�"6c]4X_�]6�����YG��B��_!�.0܌�*K�ᣣ��j@~�-�~z������sޅ����C��ԟ35����;]�nn�Nb;�-Φ�7���|G�ϟ��3y�9&6�����WX�Fk�M1h��AT��['|���[]6��b��(c��	������f��#դ6&�v@R��[�㐜ݧ��|�-�Bɳ*��I8�}@P9.W"��~�����^ϱ��C*Y����,�B��J�(�=H aIR?Ǎ�ET`��ÙY��!+��]�5��lu�]*��t��R�v�FT$r�`!�e�z��|&�Ӵ�Ķ"'�ӆ_A"tg�D��X�|΂����/�!?]�-8z�����
@�ech���(!c- Κȱ��} ��v���U��h-�����f������ybRZ%���硟g� �;��Z�H�*c��ʪq!/�gW���/��f��(G/��c�1�]����g��8��=��H�lE��`uX�I7��
�T��<���*A�[{;Y�z��E�5�:��@�&f�]����[-����0?���z�5L&i��J���ɩ��s���n:��a�ň\���*2�j��!ފ;5k;B!�Kr\�����|���6{�\��X&��w����fI*����}��g9����6�����{�����H<�O�յ�2��}��h���^��Ɖ?9���R�w����o�?J��[��F�'^�����[>Q�Tω�U�M=ă�3:�qa�����oK�z"A>��Z�t�1���4��#ܐ�-��(����������ɋnZv��[ځ��S�-�B��I:f�#�P��'������r|�M�� �K�^�� ��� Y;�SAN�^����)kg���Smp�6�˵X/݀��(����ሀ�I�-ї��lP���!���RX����/�Ё��c5f�	�=̍�9�e��X�r9����+��7��9���a)%?�	�b�Q[��؃��5Y-���*U�������~;D4�	��GȈ�?2%䚴��16�\�oe�j�@��i��tbLD~��lO7�~�Ԉ-HZqY��wO4��l�j'���FǮƔ���ȡ���1J5bg�!>�[@�w���1��\�ɶ��z�PWڼ[�C�|��������!&<�nh?��#ߞ���q���W�`+���p���ES�zM\�W�4���)�������_�DMG��x���t�d
EЌA��H�^+��i��vqtҤ,�\Z���˯%���-,r�!*�'NI��/m���<<��r��<���էNƤ�� )���a*�(��S��y�Hʦ�Ӄ�Վ��"%,|]�'0"��-�Y?!�#`�E�F�V���
*��q�:bWۂ�}Z�^hBA��h鄙�E;?;���1`�p���י[^p��)l��,^�b�0��|�����Z%T�����u֐�l)2�����k�~y�EG�<�%g�֟x�sTg�cx��D�t�<U�[��_?=�V�V��w���?��2VY�z��]W��1d���f�������$��n��^�T�! ��q⫩�36����b6����Y�Li[L �?�1DP�$�e"Ϳ�@rQd�T��(Swqc0>QV.�
��|ʞo���_'�(K�n��}�#�O�8�o�p��r�����y��^�Н6['�֑u���[&Nk�6X�!5=q �?�� tJ��7m�O�vj�ӊN��F{�^�y�@F(����Kt�D�/��4r\r�x���ƽ'�@)��=�I� � �r��(v���5���3o�Q�I�Z�0rT��<��]�f�^��_�Ĩ�������Y5�s�S
{�������������䄻�/>
�k�^$�B����;	�=���9qu��P�������y}_����I^>N�=�g�O�ӨQ��0�=:rw�*���DA/�'���C���&y���6·i���kS�8T;n7>ٚ붆�f8j�oYE�ݝQ�%Ӯ���'3�ʁ����܈�z���.9}��dC�:y���<7��#y�rl��ZI(3�G�8�c4���cA���i��;�u"�)a8s��9EJ7=j����� >^fj�˱��@�E�Ics4��T�U�-%��PN��δc(��ڤ	�7��2����Z����5�_��]L� ��T8����@D;��[l�mS����**/{i.��b��m͎���J�b��cJ;�^3��%�(ү�>[�NE��}�{>�����ЃG��jV8�נ���8����,B����GݶHFl���
���n����q��/�<h�qfז�u��'���[r]5r`1�z"��4�F�|��͑Q�1.���q�jUcA	L�KR�mQ�N���x�a��y�q�����KS3��S��%r9+��4U=Ѹ��Y�\{�G�u)V_c��p�ʣȶ�f��]�9B읮F�U��b��ND�݌!��f��4�1�1I4Hr�Tw����vB�0f� �&*��FE�%�̓Ҥ�8��Ks4�b֊`�\0sr�p�_�;�\�i*�� �y}�z/��'���l��9�	��EWL�U����z���]�X��n,���qyt���3��ں�}*+���ړg����c�@�V�QS%:,�0�̄�1!H{?Gw��dR�^��+(8	��e \�����K��s7	(��(�-�ŷP�;�Fz���.������K�r�åT����H�IZԻ>�hb�޲zH6U�p:@�����u�r�y�P���}����	c 5���b��&���{I�<���͸f����:���Ctڝ��h#���is��!���;z5O+�;��r;e���d�ڽ!i�F����3d4�Ȣ�ԅ5��?T�ņ�ɭ@>�XRo�ҚN��ƪ�z�ew�`�5��W�3<�U�t�q��w�gb�G�Iό���чs3j�QH�\��~u�O �����]C�/��3R�j:l��'����q�p��i޼.�J|ܥ��c�v��(��(<c�s����W���p{��-h����:B@Jt%`�/�c��C�yR1�fJ�k&N��C�x?^E$n��I)�w|"�*�r~N�&��?D�K������ӣͬ������8�w)���,���غU�h����M3��WR����V�(<f��N�ǒÔ������x����Z��ᔫ�U"���zS C�9�wG0C�>�xD�iY�t5��#���׃8���Tܷ�2�g�\�tx8K�!Ă��'���M�j����:j�sU~�=������s�E-�m��>�[����I`z�CC/I�T)���*0yT���u����6t����0������)�1� ~n�1�W)溭�A��5�+[,[y�1�b�MS���c��	i�Р�����J���"��D�c��@2������N4�cM�Ҳ�m���1O��į���P���Ni����Փ�N�Z}n]8ED}�b4��Y�5hF������s�5N�0�|Yo}d�t�;����X!jC��a�3��z�<U?������5!i]��#���Τ�iBs�{@T�Qy�v�l�x��[�ENg&~�������o��+���gNwp./��Q���4�C��_��\���J�ƱU-H���ể���]�֕�`��[�&֙��c��q?��H�~lB� ���,J=�r�qI��]��E+���i%}$N(Ê��FZl2K�=Ѯڙ9jo�&r�du���������@�1��Л#� Hgl�X�����P>K��훳;P~Ƃ�Hs3幁8��5����u{�	B�f�ׁ� |�*�j�'�Q`����T�j�cY֨�S+2������V��}d�gČL8� �`�����9�O�$�M1Jך����[o�r��q�q�P���K�p������3ܗ���U��>3P��� ˟RH��|'@��r9�Z���kNZؘ�&?�m#�H(/��V[Td��TE��u�κb�syv{6���B��@�?a=k��?ee^w϶dF؃d?���Wo��:���Ϝ�e��k�>W�x*��7���}�Y3"���� �۷z K:�Pjb�����/þ�����������ɟG�ź��U:����MP�0`;S)�G�D;%]X�q�����ނ9]��a�d�V�1Y�_��`�rR��b �o���v���^��tg]6�"�o�H.�H络toҦ�D?�b�wI�.�']�;�{� �gX��ͧoDL���|��{*	������A�}[Z6o�jĖ�k/(껵~m�)�q���u3��T"���X�����!� �"�G*���He���5\���w���:KU��7�e��2m��!��Bc�����(�o��RJ?b�"�^���
���˂�XU���8Î��j�	�0$�I�(.n��|�e�T}d��߾�"�EU� A�`�+�+�������r7k�	绯�N7SO�~��m�Q��'�냹�&M�ɭƗ�t�枏�_l׌�ߑFL�+B�Jam�,���@���ɹK6��22����@�|��WU[j��P}s@'@�"\����?�/����I$��ad�S����ҍ���q����%�|��M��R�	?*i� 6����9�`2�zy;�]�$2��������XI���*����C��G�����6{�l	�X<�$��X+�՘4�u�pۚ��
��Wt�c�w�w�W�݆g�H\r��J��=��&����u���T_�;�0��3G���[����5z���i�����d|���f�-N��/9�G6f�W���J�t}��"^��v�������+�*�.}.�\'��m��n�ۓ��Ἂ��Wlt��o�1$0H�f��W������1���؄F�kDfl�T���34K�Tm�;ܗ����˖΂��Ծ���$��4[�	����}j"�J��Ue���������_���o�F�@�t�5�����=s~pw�=�mƩE0��T|q�iW��hNďJMU"�Z<|d�9����e��n�%��.�b��D�O���z��]��)�{Г���O��m��#�x�ضX�S]�ֺ9�D3���'c�@���������uLņ(��+x��5W�U8�%H�L�JU1�?��P�y��1u��3�s�r������<��R�|[6u}��ϦͮQ��v2��(V��c����4�M�O��|�T���j��¿XO[�k�����A�{�g�Ƨz,K��2t�A*��L����"����8I����c��L	�]a�[���v�����Y��D�� 2�v��x�b��q'����ø|�%��䞑.~�/� �����F��0�P�Ĕc�1���K�M�IH����MA��W�Gy��v��J�Dy$m�z�`h�Z��-�gg*t�I�A�v~K;9z`�-�-�O��6�O~@a3	���z�D:M���R�3�[���;]��}������sf�ԯME*���0�Nxr�<h>7cֻ�lL�M7��WYw��"�>���MY�̞��x�0�i���p-�u�(�}�J�6����_/ե��̎�l Ҁ@*�'ݱ��%�Zdf�.��g��Z�����k�Ƶ��ߕ�9�����7.6�8���!5��O`_��~�I�K�0�'1�劸��N�K��L������	wp��+�e8�Q��"Ey�t�A2�pq����������Iy���W��1[=�4p��Q�=X�z�l���B6�̈́�a�
V}m= �d�o��V����z���_�u�g���Y�%�3�e,��8o�����g.���z�L�	$,��ϓ>�;����ڽ<�K?/�[���Z��?��5��!m�`�4�B�b	ֵĦP�On�s4Y�9��Z�Qe�ef�����O_�mQ5?S��=�̛�@���C��rLY���"i@E�^��#�<�)��	���O�>+�ʹE��G;��'��;���Ùr�&G���E�-c\�(��~�8^U�;	�Əݤ�A8�+�q�71�Lx�
 Y]40��M/dɂ�6]FY�>�`��im��d5k���
�D�N�#~�nM�mހ	n<��÷�����c����
\��Z��/����U6�u��^�̰�\K�0.5��Q�!v|����aW�����<>�����ߝU���qh�����F�tc�;��d��{����8����h�FYָ��c����Y��1m�#i@_CH�g��j��ς�9|M�'`Ȋ=�
�����U����^�mk�U�a6T
67aa�8�3�nD-���W0�����K����8^��	D�Ԓ���e�)z�G�jH&��[��K'̷��z�c*n�|�1�ed��Ź���*��$�v�]�r�=��&��X����p��|@'�pc;i���g>�[OT��o˦�G��C�fS_^Re�� �]Z��D�tbYy-���nE��J�q;P���S�8K�L���̊۰7��f��?��@/�	w��GI�����7�G�������£�.P�m�>�ဆ+.��_͘P�U��1�2��X��D �l$�m\<�Ӣ}�
�?�᳈���4����9� ����d2Ƿ��$O�拓����ێy��2�b37�N���yI�BW]�LqH��0cؗ�>WD�]t_���9�mA�ϫ9֧K����ƛ.�$Frs��C-f�c�V�o	��Vs[0L+�0�1E�lkz�W>�!p��5a�~L���J�[��2�,T��q��FAjhI���ج�`��u��Q �N�wz&·�[$����M�L�VDH��ſ��>U��G;u��4Ϡ�3Ă?�#�_9��>�  Fg/�7lS�%d� N��(�V�d|���*�(�%G^��ྶ�K���M{�8��g�izB���_ā��qs��9�ÅJ�Y]�"�eT!v��Ċ��fHy��c�3��.K�����p��x� >-^�2���7�o�']��t|��GyD�6��0�=����z������D4��e����x���i�� wI٩;�}C����q����Sr�,.�=�	��e��0$-n��<pr��s w؇#����A���Q�c�T����5х��Rj I�q�ڡJ<g��;�@^:��� -g/�h��4w2�f$駓����ݗ��֔`__�	�H1ͼ1ҝ���$�
j��@e;�cސz�l�}1(�0�{S��o5�����g����d��[X�M�
SN[&��Ȟ�Y��<hw�B��aoХ�lv���;���X�����A(�u+f���U�t�d�q9=k�=L��7��J2 Ӝ4a�|h������b���-j���r�� D����y��KnƋ)0��е�����Vr��g�J�;���_�$ﱐ,AмQ�)�z��K9�ߐ>�+���Q?�JdJiU!���̗o+.X�?O޾1UE\����8�6�����KL�VE�q���mB���0kZ2���vr,n�����X�^�.���LN��rV6��uW�ߝg�t��hF[� *�n� �پ�w�=]X8T��KR�lׅ��H���z��Qv����lX��r��_����� l�&�K#)��-�i�2W<9�kJQNN+�]�9��-k%Ҟb��v֞)����x�G�U���(d�n����	�0�j��	S�>BjyU �}�i]3y}}�\9��\(`}9��b�4��d��۳`�L�:��j��}?�3���^�#kxk1EG	�	����Bͱ��,Q��mU4]��G�}wD0��H�s���ƨ����Q�n,�/+6�B��{��2H����E�yoh�?�4= ���EZw��M���AX։>�ę��.�Qd�qӬ۷3�!#�ģB���Gi��b)8\�e���|;u�� �!�f����L��
V;�A���ߤ��m�Wҳ�>�5CwBq$}�*L�
-���q-����0pd]9�G�!S�$�v� `��ە��J#!��W�T��
� ��d-_�T��|�C�T��y�Ȫ��#�I�i���� ��d("��]��s4�*�9��l�!O�4a��ˇa��;`�s2�Y�d[�r��������5��k+���,�..�Wrﭺ�KY��|�0�ZT(�@v_k)��n=^YX<���s3#��Y�;��E�uԥ�D?;��5�=/>�'��4Y�o@�!}Bs��Ao4�TOmU%��Vdyc@�ϨO^(UH���	�˥pjJ�� M��o���xq㡉��v��u_"u�G
{�	���VQr���S(ڭʱo�@}[�Hw!��~�X!�wpo�X�҇@������=X?n3���ϕ\�h�Ogq��-}���#c�-��m�ÚL�@��98=o�Yk�'S�h>�4��,�;.t�rQ�I��w=G��IPD�<r�G�b{fe�G�+rW/������X:�A��M�aM"ܒ�_�~--�Y,�rr��}�I���`�ޮx������^;�Y�u|����+��*ruh3����Ǫ��3�$����EM��R����#5�BJ�fdzL&_�	D*��xׂ��1��.2ɲ:��Y�J�Z�7����W.B�y�&�?��*�R�E$�9���KwnS���5x�Gچ8V�pG�$�������5�=���[F��/�X4R�]t�6�L�{2�$���eLA�EK��ۍI뿎Hi_oB����u.$�<U�tv#��%%���`�fvP��K>�?��
���֤�_���z-5��c1��5�Jk1��\Z�������닓=..���8�Ʌ���g��d@G���U�N�r�y'<���|�d�[�5�c�À�mBe��!�d�J���:Y���@��'1%�u��Lnm+���	~ѱ]͑��`+�Y�K�'`�������/E����H�Y�VqX�҉rq�'l��H*���]E(+.cq�+�^)W,ͨ��ft��
Z����U*��>�S���V���	�����lxP������%��EC�B�pj����xlw�c�O*�Z�iwųm���^�i�q��Dsgր��������-����zˡԚ�0����#��;D-��DP���u��O�HvJ�p��/A-��=K�$���)~�G�+�sn���5�p��><�y�Z~o�ްu����d��9�ɱ0���綴M��F��^,P������ez	9���z/��~m	�Ż:�	*�\��2���G��+��3�ȏ��b�O�OXJj���y�'x�!���5�֑��*��r�T _��x�m�BԮ+�-�`�O㢠�l�0�z��#�4�N�n))Lnx��z4�,���>��'<sJ�闡D�^���7����selZ��<<�#pat z#�����n���
I�_���5����^T������y���E&��������f�諒�5a�'Iߒ��<��"r�JU�^WNxB3}��ߖ_˦�dx���^A����d	?������n`�J����1��!p�:��=	퓩P�:���Nx]8�$��ܻ���*Ye;y�p��-5�f&=7c��Z^�b?ۄ�Ѫ[S���&�b�`��-���!L0]���� ����v��nf�q��Yj�h���r.x j��J+n
oj4G�����l-*�>��YG��Ϝ���[��3p*1Bi$v��M�Tt��z��3p��V��ߥE4�Ԣ_$q�)!4��5�c�IQ�����q1YS���4R��#�
n�ЋM�>xb��q���\�U�*�Q'�A����p>�P��o�����H4c�)�?��]������Y�ϭ��C��:��V;Qk��?-3�&q���VO���pT w7?�f� �6ً�}"���@�M�?V��f=J�8�̫���7|��`G��9�,d)
H��gقI�V{�@�Y���c�^�WG�َ��qXWl�C�/I�}In+N�ϴn��7�e�Z���Nf��(��8�x�*��0�]0��'(�3H�f����0��X�p�y���!k�@�u�xQ��n�%F���j��G�yFy��+$>�����%����Ybq�t��O�f܍��I�B�p��2�wLi��ѓn,�� ��㰨��ρa��ǔ:
�0i�D�/�q�0�!�F���ܡ��~:���-�c�ӟ�ق͘BJ47��v��� ����H��MQ�^B��7o�-Н*6i6�z�jjȖ�Xu�/���	B9^fx[�xzX��.�ժm�rV��}�X�p��=`������݅a��q��$E�$�5��{WlO��2�k�����!)7�O=��%�K�o@��\�j�o�����M�Ҏ�sm��ຝ�K8�˻�e�ϏO���ŕ�|@7�4��� �*N�t�Txo�*K�@�hiN���/ݕ'/o���FɄH��I� ]3L�{��-#�%��
dNYDIGq��-� �/�:l�(##����޵p��(����u��1��@����Xl���];R^��#觲��w��m��[���;��]Wx�M��}(�)����i}�2y*�����f$M3=(g�̑���'č���OZ��
3+U�?�xp�
󩿺z:O��6WS�:tL����D��eR�$Pnٺ�6�����G���>"�� �=�X���޹�?ϛ)�?^�b�j�.
.jx��H��H�t�(r3�a�*&K]EO��)5@Cg�h�6?a�y�0�E%�oK`��A�p�I�����?������0H�����a�G'[)�(�ga��i�[��0Er�K���ն�-ɖ��1$����������c���8�Y��>�\��y'��.�����ncJ�=_2�޿��
�h�y��L�uv��}`�Z�V!SЍ-�H:�X��d�>�����06����[c�5��䵬�\Cܦ�G�f N��'���&L�Qep�o!�G}�(-.�	#�T��zE�[�8��� h��	�hK��t̑h�@�4��9Ѵ���
����ѭ���!W�۟�85`c�P਑��LG�L[|SƲ�2T��� G ���u�Gxs�2?VňT=G�UH[�5�ii��JfN=ڮR-�/���5k&�?Q':���d��l���g��\r{sz Tr7�L,�ں(�P�4wb�},�Z����fQv���J۞�K�Q�_i����7�(��㫬��]��t���[#$A�����hv$A��1�f�a��(��<�$z*���ܷe��l�����&K�S̻�[ߓ_��(���3O~��\z�A�^��R��F�Ut��̘T��"pVA^=��vo�;�\kvrJ �lE͋� n�����&���3u?T���͠��L��4M�? S���w�yz�a;'�v�K�� c�|�J��`���� ��󠖣�V"�<��d�>߱	�`ц�jr�#���焋��@N�')��>A���@4q������F%��1ꫣN]�-.��-��#��p<"1��N��A@�w�}M#�b��<�y
�@0x���S�Gd��4�(���1Ȥ�G��[5Fq��>{��JX?�ˋC��6�bE�:e���"�7���7���VY��4�a�����ɤTk�EW�N���&���?�(H�8����$�N���3W��cР�5��m�s��������������M�!!����Зe�s�o��`���ZꜢ?@���״:`2g�Tc����Ƭ�TM��<Ў��Y�q/��4�`�]u��^"�^�c�o;Xk���@��:,x]�{}�a	�4�;��W`G� A%���"�"��H��������)b~U�lH]�R���c�z�@�T�̌űM��䫫�q�O.��6l��~ف��=�>u��5;�9��pqHd��x}E-�����ֱ�nX�,�9�y"��������}��{V'�.����4Q�����c��;�����\��M�є״�h+e.�{�n�>��E�D���LՓ��8�q�{�+�8bQ�Tf�9��ȕt�ieƩW�(������sy���]���#IQv�[�^S����������jQ�l�*e���[psFTF���O�vH�஫�'�1���al"�n��C�:�\y ��!��C�.�Ӵ��蘙�.w�iv��dQk��n�ˀ.��GP����ʓ�N1)����!���ע6���L�W�I�ugtB�9.����:�[d.�Z%$��8�,��꾛9��ԅ{1���X��!�w(��Щ�KءG��&�sUIEp�;�mM�����]��U���2���Y�\��Ӛu;�fs:��i��D�����<�'��˿��~�eҶ�<8V9�4��.t��>�
�9�ՄXi%2���f���'�{4�C� �^z��0)����h��m�߃l�{�$拻#�����B5����;0
�ߐɾ�4l%�u-�@��6��^����9V����Y�+��)*7܏<�a��.im�c��/i�a	$7V����u(Q�I�['`�7B�`}
M�>=�ƛ6���w		�W)~�0h�H�_��Z�I:��܇dΰ.T;C9��
�1*�"MUz��T^�Dӻ�YS���Ւlˠ�Zޠ%g?n��B�~_�OJZ�f�W�w�Gmx7SbL榮�Ѥ|J�I@P6:�i��&��Zy��ǃH�]�hE�]�r��̐��M�RP-;O �;>S�73D�75�(��'�ϓA�C�R��G`z�d�7���Ͳ�(�}�C@�t W�c�$x�xOF�?(଄=��<!��Hę�g��?�}f2;4^*r8���&Z\�7L,����
x�ݾ����/�$�,��S.����e�u3�;��CAw�a���N����l�^@R�#�7{2ƒ�"�d���юS�y�[l����/x�1�X�Gt�i/�$پl7�{}��Rtcj����.�h7�w�J��=���?���U�����q0��a�7��[f��a��C�������ZS,��չ� iIll�f���k��N�:�n���)'i���4�`��#�1���� �����Y��X���� >��~��}����jFT�$���g� ��:<#��䌮���t]l
,��Md�������ﱥV�vv�^��m��Y���f!�._��8˩ړ���}KS(a�y���̪�0<��so@u��)Q�����d�=��Pg�]���c]uE+䌨BoNU�q���Ѐ����o�E.�ג�eG��Ȓ0Mw9p�h��C�v��;�p��X��F��9���C��y�`H�~ީB����j�h'ڧ�y�3�fXO�ъ� +u���c�z9EO��:R���m�p��,v��R��08ߪ^�k�7{�����?d3qq�xk*SO����t�D�_���ܠw9��S?n�ә�sO5|���/�������pQ��[�TZ%XW�,k�����*C��U������J�i�")�A*����ظ�MŖd`���m�Qk���Ut3��Cr�I:�M�u?������W\��9Gn�0q7�,nz�UԤ8���������K���\"�8=
 ����]�N?�[Pͮ��N
����-��ݾ6���^�5�l'%O��� ����H|ƕ&�X�Q��P�f�8��;\~R�ؗ!ˤ	"�PU4�������O�l�{<�Su�����5���ta�	d�^��O��+*o@�Ùd��������k�}ı�T���[�^[�}X��X �B�:́�*�mL�4���!�S~����(��O�qW�n�d�b��	�8=�*�%x%�
�����V��*٩ �z^~�[{�;�	�`�ޅ�I?�Ø�D�)|���z����ŀ�>q
�$��֡-Ʀ?�N�CY�"ݚ��g�-�r'S��^��7��ʕ�i�ϱf<�2I�rm�����N����w�p���@��+�:���jюPѴ���]�#p�?s&}���*�UW�;�6�:5�N!J0�DN�I�����H�.tp�Z=��	g��9"	��9��챑� �T�%D!yc���x~���V��f�4��* g�Ԗ�>��%���l�=t���È%��N����¿K�"]���T��6���h�{\�A��%�F# �|��ec�o�QǨK�C��~�����;��=���13���~�F�"��T�݂:"��}X�TXA�ȓ%o���qτD�ceWh�$p�nya�%�
80`"FJTO_���8J�9X�W��ȅ�'���m�&�Eb���j��B/%�m�}��,ђ����k��F*4��o����'��71��&�?�ׯ�2o�F�[8��JEk��r���ͭT�[���k/�4��J2���kNjq�G#%{=I�|���<idF�t��>S,(�Ǌ���
>.߻jGAy���~���1���M��R[=[ݩ9V�|��A<��9�'��R���%㷮Ю#^X��m�" �)0�ɰ���m��-~��[��P��WB����w$f6��b53����9����GT��pC���hw�(%�����������KvƠ\�=�96LCܹ	��]M(�{R
�vO��[o�G/��ۼ� E�E�<1Uy.0��ո{X5(z��)�)�Z��-�LC��g�񗖉��J���/h|��m��L�1j�X�*C�Q�����S�� Ƿ��p j(kG�;}�>�gD"�ݩ�C?Vs&����8R\�����^�ߐқ�n���'լ�[�\'��Q��3�ѱ�Q��i���p��W=Es�8���i�~��X�AU�s�A���K�ѻ���g��&)A�?�܉���uX��Hͱ�`ӑv���NO��f�囔ъ}�S�{���j�[oz�o�m<��f��?�iO>L�H�?��[1�/g��9L~72�\o����υ{�������J��`�x��U�M���,�/_*��緇?��t����ʳ�2J�]�jp&�9YRPT�;q!�T�)��lQ%���N,��b}6����{[���Mam#���N����5��\�6�{��w�e�W�(ܕ�y7Y�zoٮ�O���Z�?��Y�%��C@�/*���oQ����ʷ{TɆ���-x�Ƃ"st��>YQu����X�1Ynm7��):��Pi�Yv^X��	��#~W�U�Vz����d1�k�|V�щ�����5�&�eI-��p���.��ɽ���`�\�������o��K|�IhUdox�1{!L���
2`��|��B\��E���hsXw�<o�?��i*3q�2$��C�0ir��$�M���A�����(���g[�͖�<=��o	#C��>�Fi��|�L��q�u���]���8h�A������Ij�%
}��-tK= �@U�ɋ3����K�-��Zq��z,���d��.`O���K޲'p���`C�l���v�c�Q�+P7X��E$|"gm��( ��������k;�&:9Պ��|���;h-B��۴����[4�(��,˚�t8�1R�%���hC�"-��4/��=}���9\�QI�ڠ	>2T�"���q���O�о�M�o�UOۄ�*N<+Y�K�y�d���>!ƻ�ɍ���J8)�H�Q����Y�}˕��2�i�D��ל3pP���L�a��_��vwI��X�.a��s�ot�o	@���n\�z�Qf����v����Ӑs���N�~�n|U&���Z�u=�xu�1�[��po4w����P��	c��1���W������4�#�M�ew�)dk5�aS�<>30鹶���J;���ͻ��)�bz/g��3�3������*7�(���uJ��{�A<�s���a��,:Co�8��NiӞժ���x�g���� ��7R7�EO7��a���|�n�o���Be��*�Lot �� +��g�W��>��Q���:����Dؠ�^�o�E�;A�;H���&���81��Ѷ��Z�Vu7��˳4�Kw�h�Z��l�c�CկF���_y��1��C���$��38���k@w��(��xP�mݔ盈{�[��\ �!֋-w���T��:�(hȥ��گ�{��қǭ,����d��	�Q��L���lV����Y��3g�W����9�H�9�$��:��N�bϚת�}�a!�峏6�Ĭ���s��~i��Pܕ�J��&�k�w�	��H�w��h�/�h�n�'���:�C����;+���ڔĆ�+T����QRS���lG.]�����Vl�i+'&��d�[���k��aX�R��j�E��6H_c�Bw��D�^▬��R���Ncz��2ѡ[bm���9���bϪ������a�uJ��uG@�|8�ӻ#E�����7�
�
mPxe�mPcE�R��ض<�tbe�>�S�"�}�x����	B(� (-�f a�i^�W�X�G&�R�b�~+�+���'f�f9>��SOJ���n��y�nQ�5H���ø'��vh�w:�9#'���c!��U�q��3(u�"�+q��s��P���|��5�e$n^C%��o���Z��n�'E����mJ��1c[���Yc��M�^�m{����O~%�(��Pi$����VYm^;�U�0�+�<�����#N�C��0�4P�,H��ֶ<D���v�K����8TJ��y^,�ӱ�S���C��h�`�6�_�þ��2�mg��o��%\�bck}�钽%"�@���'���o���w��ߕ� �S2��Ǔ�� �J�I��uR;�Ym�IQ�_��=��T���̸��%Z2�|��\�X�JL�ۤRe$0�_�������Z��U�>Ɵȇ�L��91פ~�.֋��`� Ѩ"b�o_�HǙ��
���.��DVb��H�p��%��B+��q
��O��0&�HMdR���×�IB\b����lcퟏ�Vϛ�����h�_Su���/E�*�MH2�;�o�H4�%m�SƲT�yo�oSW-x#V�؍Z�M�W��"�Ux��r�T~�RS��-'+�����ر��#�^<TR��4٢��dD�>��3;����]�g�5��$y5��'FMbK\B0b|�p�c�p8A��r��٘�ip�8�>����5=F߸9�}\���ĭ����JZx&���E�"fa���"p���#x��?CM�M����Y`��y�Y.���Tv�s�N�WWKD?6�3�m[Y��n%1Gi�o��R����X���G8q1:`W��b.�x�⏇o���>�; �ⷙH��a�*o2%<�h�z&֭�`���O�h�Θ�;���m8�P��6D�r.nl-�ʠ��>����jb�d��t�Ie��g�y�_V���v]�q[���uV�W����rb=��ݎf,��8���l�?�o�yʔ)�s�'���洉�p��^o����8��˄��פ�:n8s5�X����1��}~�O�6G��Q#hJNy�!M�f�nQ[F��Rtn���4�h��uC��q��`��}���;���2�3-���]��/,9xު+ҡ���A
�8e��Sb����G�a�?Pѓ�KQaFx	�+p���ؐ�;(Y��������u��頋a�
ry���)vh�x!'s3)�h���J׺�lS��)"]�����t5��^Y���8x���#:��\���5��~��W��cn�e�����P�h�����m�d^���=.[�0�m5�B��|�4�ߋ�N�Y8C��;w�upR�4J�cU5��b~��3ȼ��{'��l����u�y\D.J�|f�p��*�����N��Մ|�{���?֚�2ŀ��z%����+滏�/v},��q�P\D�t�ʏF��zZc�%�A��9{�=iy������gm �U�v#s�jQ ~zȆޝM1�Dv,�y�t9�q��h���ֽ�K2�0���K�=��9H���Ր�/��:��@���o���k9p%���9� �B[�h"r`�T�F�J�+��+"�q3d�l�g�pʽJ���?²�+>��Ø�'����,� ���?aUo�r��6Dv��틚���d����s��\n���WD߀jbK�<HU;E����I@���7T��fb�ӓ��c�zAcgbC2�<�I
�y����.i����x���㿪�)��Qtz�p �@���\Q�8��5��(k�{֕�i����p�!� wZ�������V`l�����Ϸ������o)�VYk&(�~ZJ�B�*�RF؆��Tbf���v����ԩ������r=�hQ�����u���]�a׭��C�/=�F��y-_їi_��E!�c�i7c��&�c1f���?��y@�C��+r�����=�B(�D�3�d�7p��gm��,9�[��z�x�tV��'�J5��O�H���'#����o�lG���r�d�]{��̉�����֦K��1-����H}�9�Z?�#l^JDB��Î֩m��&��a%�m$s��l���M ��R�۠�ke�E:��@�)E��ޢ�(=��;[H�Μ��ꖭ��v�c�r���G��G��cڬ,�S&�X�k�TaRj���n���� ��N.��_��N��<�"�W���DΤٻ�G���^ϖ�W奔α��K+�ZF#�a���"+�H )�_���A`!��`�dQ+䏅F%��#�F��`�u�"N��^�2A�^�������
��6��
�Si��#�˳~.���h�����P�!���.���n/��v�릉BYղw����B+��!*F�Z|��L�����W�ܻ\��}-x�5?�bT��*Pʅ��+iR�:7bm�f�����3�"�;2���_߃XI�����(���6���;Tɐ"�H�v�S���}��٪Y�}u(�n��|��g���
�C��6�`o�X(�Vn�]���q��6�
�`z�@�����re�Ŝ5vV���K/�Y$�:��S��8:�����q{q�����1ʪ�>��^0�8xQv�|�VG|OLaf�+v�Q�o{� �k�3#��V�p�s&%Q��X��o-��H4.ʷ�b了wa7@u����]	��W=�\T���z�Dk�|�����#�x�@�h�ͅ5e�����_��(���F�E��K�g5�)���Y&�ʸ
l���d���W�;��L3����*���'ä1QCk�}�d����3L2���ڄ��N1�c��oq��*��S��>2w�,_����~���k�����9ʽѾ�+D7��n�'�>�8�-S��
�9�u����.A�Y�-C7�E���͓������<?��ԩ��ެ=����Q��6�X7�+S�FVz/K��bD��g��|��ΎZ_��
i����]�^zh}��>:�u~Z?y8�K���D)��k&8��.�*��_�	�:��JѦ7�~���I�!�i_&��3큂�
�;g䌈#7sB�w�mN��t�P��O�/�O��Z�N旮+
x����r�lX�����`�+�9٘=��+o�$x�J�v�F�Ш��K�%�Z�y:�.fD�t��Rm�c�Nj%���;��=�dJ��/"���+����2��Or�`�f)y2K;8
`�|)����f;�M�׭LX�oEpK)bJ��Ǥ�-U P��E�RhXY+_bD�O,�����v�jʲ�b�f�Ao�"q�>+n9�7M$�yUkX3m ���!I��\>�o$Lo.Y�^��c�������f��
LDgpHJDU�?�m�]&���|��0������q��5�m�a#q�6��K�l���T��A�׏�}TE"�����O�
8eJ?��^�d��%e��iC�����N�]��;7r0�ƕW8m��|e�tM�]Da�M�4q���SOR��;7�!BTEX�ۋEvl+�\ol8�RS�M�G�D
��9��	��?��"��!����OF��p��� �j� I��("�6���n!`��ŏ��2?/}��O�5R�W�F�l�<�|�K��P���5�'�6��W�(��� ���T�enEE����"�������un�\S�� a����S�s����iW��^�{+;��8�e�ޝ����袠<rJ�Z�=�B�J���	2�д�4T��T���i��p�F�Ui�0��lU�����m�)��� Mq���S<�v�h�w�s�43!x7-���+56�W�$̨�N%������Uf����!��>��q�y�b�ya?�@���)��F�Be	�܉b����XL�\,�b;g|G����ݧ�Y��M��_{�Z�8�#5e�<��Ó��G����<�^Z��K�8�f-&O��5�D�'��兀b�%a�
�x�V�\YFM=�2^��o�c�u��¬��P��U�$a<YѬY9�E࠼��X�i��b��g� ��~$Vm�;Y P~N�q@���Bd���C�����̏�hѩ�k �.���)D_�J�{��T��a�������Q�ts����_�J��<�Yx2�3!p��;�3��I�B�N���ޔ&XԵ�� �u��[�,"��x�!
��4{o �3y�k��벆����k7��vkU%�.��o�a6'�
�Ksוֹ�����X2��9��l����ϻ8��>
�Wį�28�"�Ы^�!�A��NK�~���pb!r^8���DQS��D��m���(|(�
�\L5�Ŧ6>A^2���-2�����A+�6l��\y
����P�p�涕5�5֘���HT�{�*�o�L�mL}G`�>6J����U���_Pw�(L�ܱ��-��O�U/��:\�z!���P���
�I�X=;��A,��M��D�@���ve\��!"Y2�;�΢Dȹ����փ���k-xRP��7�������O�-WJ�<-/��TE~w��L���Υε`x0F6�}m~v�c��`�VJK�_��^��(f;��N�� ��S3��S��'�\B�ê޶���
;��Wʍ�H��I��N��$����,ݏ��e��w.���d_nfRx�l_Q�J��㳦n���MPIֵ��P���;�&�Q6!�Q����6=�<�#NO�e��F���Y7����s�[_X�&)Q�͢�K��O���+[�6�<s:��0�� �7=`�������~�.٘Mu�D��ԑn�qX��Ҿ���Ĕ,�z0�1�w�v7!Y2g��PB2B��c�zq�8Rp���!�:o���:�xuF�\n���b����V��7�V�H�*Dl �O���!�ë�wVAt`:��yO�&�|NϫH�j-�N�j�Q��\��]�H�a����C���K?5Ţaj��,Jb��@}*!��O��ؙTϥ��hp���<H�K����愐��s��"6cOK,��d��?��-)_��y4�9��N�]y��l����x����GwĘ���Іf��0S*PYd��d�-��pLu�G�Ä�"sk�$q��Ҡ"$��3]`�d���$#�,�y�?�jw*t�d ��BG����S"o�N�b����P�u�V9u��E$4#��(�v�T��tL(q0����Sp�0�Q@��꽟�^�����5Pw(9�j'aY>�P�E��6ͥ�Q�������+P	bia�h���I#�Rsyp����R-v 
�C���[@���i����L��T�=��|$�A�俘��i�~-cJ��6W9{@L*ѵeCj9�G�5����~n}["�{����Ҭjv�®>���g��GzVڑ��#��o�8⧼ ���G��}�%
��$�3�����eg������͏�uA���aN�Sc�����Vs�Y��w���&����L��H)Qo&T>~_���I�MJ����2U���tͱ:u#�?�G���572���8��(ٯ�s��	 e�x)=��B\�m���EKj���C��!����ˣ1�;�'{��ߣb��z]e}e�բև��yד}[���fmkU|�0����eDK�H����X�3Ⱥ�Q��#����:�Z�xU�>�
���5.O�u[wx��T�+mSJ�� ���>����!1h9�O�]|�������=���y��h�~��D�	\ܱڄy�Ɲ�]r��K|���_c�N�3�:%�����H�� _fv;R�p�8}2�ٞ�r��5��X8��)�\%Xm��SZ���s_��|��A/� ��� lmU�4�@p����!��v�i�>����%��9}F����K�2�:s�)*�<��D�E��.׈��W�|�1�5���%�?��v��N:������P����f�uwe��9�\B�	��U9B=�U��@,8xv�{�
2j�e$+L�tS�I6��I�����TKȮ��7+7�}�(.n�ňw�N��3�5�0��,��Ir��&�tc�
����))E
�MTD/2�Cc摶���k�T)�AB�����_E��,�W�?���}�	� v>�FϺt�V!ڂ�d�R�O,��|5��K�ٻLq6�W����k#�3(}�&�c��.e�
�l��>��D���s��*Xr����6�Ĝ���J8���1<0���M������G��@ωީ�̀`���T�ș-l�&��\}���*_RZ�<��/�T���Au~���2�^��;����N���͚M�~�$�d'���gM�'-Ǚ�Dxb[�s�$�s���Ĕ&�2B�Z#}vwyq�"�J`�)�ah���M��-y^'����2\��΂_~ހ���H��Y�j�w][ý&(���u|�G�r��4�y��epf�L��!�����:)�(��G6a&i*n9�uw��q���S'���ˢF��э����bR;-�^�L A2}b��19Ԥd1�dU�Պ�@ptJ*n����,�+�0�*�t����;�.���h��T@g�' �)'`�U�K�?������V�%��vym1��[O��x�'��o�+��1� -��bU��kr���l0���Y<��S\@�eq�I�tB��f�R?N� �Ĳ��VS�qۚ�p�c��aL����D�����#!��&J�c�C�D�`�+~�Z�&c�(������6u�QQ�p"P?67�/H\�Z���[����$ռ�	��+mW�����[������E���-M���z�K�/|�����*�����^�I���9�V5/�(TG�lË�;�k@O�]p2sT�#��I���L���R�\i�J�o��]���@���FZ��%b������LCc��1
��7��y::��w7Mw�Fw�����̎�ޕC�bh�0�"� A�$���E����()�x�ԯ�߃{�C'�7�����Q7���eA�Ը0�Gs�-s:"WZk|yscm�֮J�n407�`)��A���S{Ԅ�5��.�"�
[��{�o6�ٴŻԡ��+��%��l?#�(�x�����{h�j�������N��~�̫>(c�P�z����:�bV���y-d �1sys��sj�b-�G�`��<��]�w�2�� ��g1`����>T*}�����������,�it���(?a�m��b1�ސG����a����XU=�!C�΃�>��^Xվ��<����{�l:je�C�����6)y
�f����t5�/��g{�NF��W7����������pci�Qxɢ��y�q�J7���!1K��eJ�<��E�<~^m鷫�ϣ[�kЪ�605��{�M����Gv��DU�UNQK#C������ߺ}�V;!#���J�]%�K�yr��-sg}T"���j8�e�W]�8+u�jܫ~\�MpGk�Cw�S>����)q\�|&�<
�}$�]���g��nt��#s��%t�Q�ϲ�2��%u$�AA䴊:�o���U̚2�����ޫd�q-29LfH�`w{��ަt'���֜��Լ|>����<U���3��(�3q;�{��=R����l��vp��s�X��qr���T�I @Y�o������?�E�7Ctt��tXѪ�Pa�v,��	����!���$�:���X:��F���$n/�V���d����HmoU^�7z� ��܈�	�|\_z�
:���*�H��Y`F��˛3G��}��S,6s�x��x3E�`�IA֞{5��Ff�~���x�옛�`�40�����"�\�!/�9��wT����k�L�θQ�H)�r�n���P�s
JT�� u����ԐB�օ�N��L�X�e�$	��5���0����}@up���&RR6�-�\�@�2k��P(&����ɸN�Yy��R������&)p4K��1h�����g��]��|�T��Yw�\{�}_�0}K7"��P~dz���ٰl���sB��vPmzn|��	.��kQФ1|��{Ғ�ܴ��7���6ZsX��ĩ�;����!In����W���1B���X�����V��8�r��ΎW.��|/<���v���������h2Gx�f�y>�v�^�)���u��Ci���$̦=�v"�����c�T�Y�$2�P_m2�>B��q���z��Ō���X!&햢��
o,I���6��?�V�9X���/ʷ�~�U�0ηu��;4��\�.���{(C;:�&���⿩�B9O��-11}��>���1q�^c?\.�u�� �l�(����!�\.#�t<���>,�����[y������D�OQ�_R>���Do��d9��"�E��Ys-
�yFvu����!�����fп��dE�^��<tF��{���{!l	�I�7��?�;��G��@w�� �4�O�gʂ�����i�6�Jm��Yh7������͵����v���nf�Wz�FJ����Lgnc$i"l`'�D�b����l��2fl��@�ZkV��\�֗�l*`�;.���,7��}��Y5�՗����1诉������)ox�ǆ��%���,
H����E��@�f����Q��$I�\ b�m�$He�؊4J�f9i�R���Y �d��Gլ�(��]m�8���v뿄������=K=�E�����m;��ѯ�p�X��A��Z�/<��<H�X�V튎�"��m�A��q�4���ҠO"׬D�g[���h�D�BW��9ʪ�q���.I��D�P5��m��W�����bJ0-����\+�rؓY�>�h�����%ͳ*
���u
AP*8�������C}���듶���y����k��p��x�� 1JP
~�C�w�d~����pJ�zƾ�)� ��u����t�q�sIm��a��r�o[��		�Ic�ai��ؗi�1�܋�ߞ�S�i}�ZՑP��A��(a�{G���s�E��ú<g��i'��/�eB�
-�<�-��p8���Q���.�B��uЧ̸�U�B�Jw1�	�?�5Ioot	<���_���g�
r�d"���e�^l��I������F,h��g��5��]fB�Vn>�x���B��1h�l��q�xC�Sk�za�<���^�Z����q\}��;t�ՙ�r�ѕez�z�Yx�J޲!Ci�D�@�NqEyW�X�X[lY0��}�L%{���d*{6�cO[��9�(.!�ނ���}{ezesV4Em��O�'��B�%]��\�E�Γ-<���T� �$z����Mx�X�2c�mN&M�K�,��Dh AKG���+�����`jؤ�I/���{M��v�Bf�����fN���������y�'�1��0����E�X��E�k	�`�%�GM� ~XV���1�U�h7�T�G@�A�0��m�Kn�oA�&��`���+��N|�eÚGQ����Q0�	��U3.�ڄTWJd���t�^`��3��t���L�A�i��֖L��zP,$�}��ZPy[?#���xO9�׸H��h:;Rl�
��g78�%*�a9���H*�qC9:2La�=ÎL��x|0��Y��ܔ�U������~7�C��On*�]͛N�Q ��3.�ڗ��wG�����dm2}'ޖ���b�F���s�f&?�!�mp��n��f��Y�8ĳ��M�|ʮ�.K@Gf�l��8N"VMpKx��O��+��C�1	�42Y���q�&�Ԅr��4�b��N'�mI������@�K�QR��/5���=�|�+�K�nxqpq����ٍ??�DU#��C��0V×oY���4#����tǔ��yzd�rr�:6��a�zŴ6/���0Ň�=%��d��RT0�L���.$�ɺ� W۠��kTih&����lǐA�Y��䄕|��_�Q�[iX��uf��Ύz�t����Db�\be����TO�ϱ����x��A�ztzIc�@ ���@�}��:�b��=\Px�Z�{�+��cyQ�'��?�c��B��
�*�I�Ť�f�q��D���־��K#��2c(pTג�}�8��=��<�y� ����)�mj�"�Xi;ɬZ�Rә�ޛަ�M�k�4�)GO?��9�/_X�'�D�0_�>1׼�lEp��8歭������C扺Kt~ �& <̪�g7�R�F�ʚ�b�B�xJ��Ьe����`���5���B#c�L�]�ڲF5��A��b�^D���ς	�<�ӄ�7��hM��}�1�.�wD ����/�K��U�c�Fn�����^��)�j`	�[�(GtA;�ܡ-��i�H1�w��MU�{3��$Ԭze�R*�Ff}I���z����3��a�������4��E({����v�zL��=�N���#v����]��ӁY@AFG3S�
\��wc�Evm�dT�g	���=J\��&7,}[�s�b�����b��墷u��i���ī8͛�:�1[��ԛ¢T�<Dj��F�j�㙰�&OLLmpdp��W�j���'���+���	v4����s�P�~��>�3NFBF5��n��s��}K�<���P���*KY1\j�D_��pfW.�)Z��E^
�'�ߡ�n[�cCQ��>�;=X%���h}>�T�E�f�x���S��i��JϫXR�����d=)I׀ؤ�;�0��̍��b�uSu��	���R��c*;��b���϶*
�
�dv�UP*QXh��*��Ҷgf������:���bUFy&<Er���M>���6?p�$�q�o�(��7��� �ØW�{�r-�!S�'�dw�3��tm
_�0���7)iC	ZP�W��D������e�a ��ص�N����kJd�O�r�_X�~���l� 5��x��D��C�U���_h�?=�W�y��@�ޜ���e�ǀ�&!��"�N�N��}EU��*R6~�W��q���]��FDU�{�Z3ި�_��Ш��N�*Y\�ـ��wd����R�Ӏ���T2#�Q�
�����ʛ9L]�e�6��i��|�q�ƴ�!�VhfV���w�Gt��Sv\Rl�;kN�(b�6N �����5�C#7�{fG��ӂ��P�-�E���f�Ѱ"or"���ElIg�}�涔��ċ��K�Z;ɉ(���C�'�����Xj��m�N��9�� N�)��lh���&@EH��K$?㩣B�S�|��X`�Mu���v�XljH��A`C��qAH^e�n��y��=��D�6E_�1@޼�t#�� 3��l#!�Z�d�j��~�����r�IWpz��+�F��S0j0���
����1=6EV�W��A�،��>�iy�'W7�yq���A�A�%|7Cv�1?X�۟�p�6�p���ĵ�m� 8Ьm�����g+�Cx�L,���~%[|{Ĝ��h��o:?x1�"��5!`���L4:�M��zZp+��D/~���/�dUx��Jrۣ�MpOz�'g��s��K�/�
w�'f=�pL���4f��19vG_�c���Ě�ݙ��bȲ����\�(Ӄ��6���9-��A�����Վb�.ޣ֩5�<�@ ���G�\
���36]�ߖ%9�����%St���|J9��GKA׾?�;��2��r�~�6�7���P��5 u�f��0N�^�M9D�P3ؽ#9Q%O���v�
����E�ǖ\��)�C�9�����]��T$#m,�T�'$а��I���u��6�#"ͧ�E.:��Mو$"��_ө����`(Z�����ұW��0��]���T�� �����(&t�hk���P���5���O�޲
^诩u� ������	h3��a'D;a�����2�I@��7މ����U�j�$#���y���_l�#z���+�kA�o��Hچ}�n&����M��b6����
T>"Ip�D ���[Ї���,�D��GŐh�Z/���
�C���[s�%;��L�1V���X\�؅�
<p��6�2�<Dm$î��!R�x���SUo�ɚ������BI>��<�Ѕ� 7WùS�A�<0]4����fV��o������o(� ����X��u�;�C)ڐ��b�ŻYGX]]3�*Wy�V�"x�^GұX�l"i�����ל�{O���A��Ep%J�(���@q:8Q*�� ��v�����H�2g��+�C���c�����ȴpN�~$9u?�[�̓�l&��%�g�������>�}�H�������@Ra!j!I�
���=�Ҳ`4(K�V0�(�������zO���E2�����_e˕>w�}��j�Y"�sD$kZ�4��]����][���M�Q%ʔ�o'd�T�L�RO��h��?�%x/��4���X�3X4��:���:
��P��wZG�T���=kˮ0�MT�gʈ�	�Z�ܢ�O�����T�/��b�S�ws)QBF;�4���|��B�"����P�r.�2��/���jE�k��+
Ĉ��NH CV&	��_��ݴ��]
[i�%1����v��Y2S\��T<����bG�̫!��k�/G�ʒާ�⍂W}�86?����x� ��1mD�#:��7!���@�
�}��͒��t��Կ�d@�t�ۀ�)�U*�����5�:�Z=k>0 ��#�7�'��?�.|/u�T}�:@���Z�-�^��$s�ϡ]�ǮD��`x�6���6�;�ճ�>���:�Zd��%���n�U�EJ���[�]��ѣhĆd${^�^L�+���x
M.�p ^�E�	k�SZ���. ��G^)����z"e�襊��R�bjzd�����=�~�SLC���i;�I��3��k�e;w��]g-x����� ���iR&�T����=�f�_���C��*Z��!+I˗6� ��ב��=0D��i��Z�q�̄�	 �	`��#�.���<�?�Y�~E��n�b�$頳@f��R�|d�f�p��SN�AjZˣp=¬��2�o�^Ù��i� {P�Աn�;0{�����~�#� 7.c��w�	���y���d(YW�E'݌�u:�fw�VT�X�GE��PY���Q>o�J"�}�}�o�A�IR߰���x�����^�`�G��^rȃE�m>�g6����X;��:�p�� :2;�y7�&�u��D?$͝6�;�\Ɖ	�K]N�=ufc�Ř��c��ԴĸG�I�<��D�_J�ʻ+��D�
ڲ7�WL�>(���Y曑�9�5���0܋����'A^���\�8la:&8*h��U6��?�r�Ѣ]��Dr�n��t�X`����y?�جru]�īp<�W���`p��-F.�W=[�MyiG>J��D5�Ƕ��.�/�)��)W$NY�F�{Z�ND��ܛ@[.�
���؍��]z�̊]�Q����iYϼ����D��1
8�|_�~�A�o6��o���4�j)��<��?(��bh�Y�W����.`�9�b��t��KS�L�n�	���l���#
�.m:E�f��|���7wPj�WŽ��{�~���m>��Q��]ݔ�.�$�h���H<�=�����:�ʗ"�oO�n�G��x0pԻ̈́W��^��o����^��h7�M���H �Q���%���i90"e��FՉ�#��PoN͑�w�����Cl;*:�d7�~�n-q(/�3�	>��^�y��A<,8�'2('YzE:�3!�]Ǻ�W�:
�T���~����ܳ�C|#� Ĵ�S�:i���?���OFN��jI+�#�N��Vȴ���b� 5��W��g���w���c��D�4�"6���=j���,�\5� �z�h�1r��F�:Ŗ��Ϙl���h�\Fdyf�d
���}~���9�v)���������~�|��9�@Q�� �A���)�� ����8��ؔ͢�b��|Bȇe�����^I�s_�@�����.��~�g#��qt�4g�E�ZA�D��nJ��ڦ�a�|�K�/�`Z���n��1%.�f��W�i�_�>-b���Ɣb��B�!�y�l��x,��S�&w�7�d��	g�C��e���\a%'�y�t�Q�ؽ7�4��`34^���}��>�X󧝮��:Zʕ�Ƌ���&�z��C�g���>*�������f;׶T�*]#絩��bpbB����^�K.Ӫٔ��i"��0Kn�O�qݓ2\n����nRU�ұq�x��n� ���x6���
Q}5v���k�R���q��9^��Q�7|-�"鮖�\������0����a�fT�E�ZFN��.�*���x������`���wU��ei=�a��"�HT�oAj���4"��m<4^7O!=��"��$Ƌ&#��Ǣ�9 �E�n�)�zS����:�<v��u���4�X��=�{�k'���SyR��O���+i�[+�Xg�e3?�#x� 
���ts��)�3񟹤܍�Z�NT�w?v��V�?�*+�tbȳ��fM��<������N��@��Wy��F'��W���|k\5��:��������Ⱥ"j��V�Hn����#9X6�t�S��ۚÄ����Hxu�P�����v���J�R!�eK�3�EK_����|�	�֝����C����T�Mh=�݈��8z��"���i!�5E+g�[���~_����1c�9�����j�y�5�:R��hM�䕅��&Wѫ!LO�j�|eqF=h����ni۰�!���y��,V����f��ڠA="�?����|�"���}��w���_L��R����JR�oJ�H�7���꣉�=*W���+�]�>]Ώ:�H�!���jbl�ju����U�[ypAn4�GS�yU�5�4t����G��pgE9p��T#�gW3������8�%��O�l�~��q�����1�?���S�5%N���F��Sp"�C.�{�����1v��"����|D��������9|��)G��1A���?�.r�G?8�g:$��b�F��F��P�=A�F�������#H�@<ls��{(놠+ �EwXB`&=��l5@+��C9pm��W|� ��d���,0M�zj����y}��g��L�v�cN^jG��p��1�Sc=��>�nw�-aW!8#����]���tw����yy��2~���I���K ��#"����>��D_�|.p/o,��U�/g݌S��*�ޞT����[g�x�㾆{&��ΕHAADw�=��4J.jm�8.�����܄��/c�-t�lx�7��t���P�l���h�c�Y�#c�`#�J��K�ci��H�)�v�^�ǡ�'۞�8t�$�Di|�*yڝ�\f'I�0�UU��OC��hS�P]��^;P���Up�l��r�d/G��g�,�n-���GY�D$��y�W���_���~�?lT�����%�4Q�a����WO�56(��� w�2̧�H�<K��J�њ�̯����WW���"ق�b�/-W�X|�龿D͝ȫ���^�}آ��Rj��u.���N���V	�וo$��A��O��D�.T�[���+.�Ed[`��{q@��D�8k,q\l2+d퍺��3�� D����4�>�,-XwYg�~�r˜0�y���� ߋB����@E�4�[��|�oB���1���Bçx�+��D�s-qL�a���C��s���\־l�#���p�Z�vFOܡ�Y*P�:��xєg�n����m�A��c�{;ʜ$���G�Ƽ љ�$?�ŎE�0�s�hv��>�t#�@f�I^�Ȭ�@t�����A'�u�����'>�$Y=Z�
n2�<�^��<�)?��>�T�E{F��e(�_��I��KrW[�%V�)�u*�������K=ɝ(�����be���H��5B���w1 Щʉd,b�Fj�f�8���V��Y�u�iZے�{Ou�M��<D� ڵ3lK�DDD�k����Z��p��g3s
?X���h�Nq����Q���NW��Yz�F�>w5���Ar�.�4�L3��ʧ�_�{+E��#��^�*�9��bÅew�x͠�A+&������OYy�\`}~=���d��_a.�����E9%'C̄����qd���勅������i�K5^=cް[�#"6� �w��f�2��V�����/��S=~(V�V5�:A���v0LK���a#L b�&Q�K-!o�����Z5B�H��o)�֘x�t��7��m���ɯ-���LRZ.���X'8����_bp��S�'��9'� �k
�F���I�#���V�ډp92�G�D	Nʔ����>�/�!�Y+�E9��,���\��F=6=�4�]�4�g��V��1n��Ӽ�Y��'�{R�nI����Cn���E�oz�;��� �NV�(���V�H ��zf�/�5}��U�?yh)� �����i���8�p�����n��)'Q�WK{�w�y��u��Ą��N`���V���\���v�x$k�sB.�fio����\���g�S��˔+��x�9k-]kځ_r��Yi�rF��.�;g�k�!�q�f��M��V\^�����
Ԣ�MG�pfvl�{�p����%�H`�h��3�w�}�N�R݈��o/>���j*�c�$֮���(M�铿j����y1���k0��,|�1*>1(��g�+a���� /v9���K?~�(��
ՠ��d���X/���Y�����ٓ$�KJ��Z��������\�6�x�'&���E8��hKr�����=^N@�L��AD���В�;�?C��O��Iϒ̹S�7ڷv�׷3긭���W{)B�!:�Y'��� F�O�({Y,j�_��.�hϟ�����v`�aI\S�+/���3y�p�ӤS#�6�-x� ��Mx�CM>��X��2�Xt<�F����Ż|��}��k�9�I�B��#�4���j꿊�� ��F�i=�Ecuw+@oD�r���LJ���x�-}��g�@ �r?�|�<���*!zlzY`2E�h$�>�N�,o���Л;u��V�5��\�ߠ���&`�>�CB[�����Ћ��m��w�ITF#Sȶ#��d���΂	�YnﱉcT|�Ѭ�fE�K��"�J�\��v��V����S�U��\J�ִ��/<�A�&uIR�1�9;�] �g7��%���������5��KEں�I���b섧V;��Fv�tcR��<�#����I�Ճ/Z8�wC�(��1�E0�e�ū��q�GmoN�7
e\#3��(�ѷ; ����oC�p:�W
�^0s^.źnR<��U�̯2*痢ɿ4�B>T0��Iz�\`1�5�z�Bϒœ�Ɣ�+���/��M]w��T�V�����o#�'���W�A������������EO�A�6��%98�[{�\z���%�� �\V`x&v�|�z�gn���b��>�����{SjE�gx�b�	�8�U/F\� ��_�
�a�����[N`���f�J�M�Xx`B��P�Bx| 7�' u	D��轣�|��(���<(NM�?#���nT�Cn�]� �џ�m8�v1Y �n��1���t���Ϥl>����� �U���)sATnShl:�Jt��k�������w�xB��P��V�p1{z!">3��gں��EXa
�f�q�YN؝C�/*�f}�zem!���t���X%IAf�nR/�W����͒l��&�3�����4#��
�2�UL5�!-��~dr��!@�N U>��c$���ʼh�x�VF�h��kV�p�uTm�����̩�%�Q+jH�f��tL�M�_I��ъ�SP��=��/
�7�3�B�:K�����o�������1
�T&�ݑD���q0��H2	Y�O�<{�1�R��-��� ��F���;d7�
������u��, srT�&�5���"�y���P��y�/IT�Z�����<������8���vr�'H�W�au�Ga�tgM�fV��^A���̾I��X�L�.Ձ!h*>��
���=��k�D�5��ڋ���6?�(>�?��iǙ�£@������K��K���]�=�|fac��a��B\�sΖ
�΍����ߞ��@h�?,�,���u�1���f���	�Uj_>�q#���x-�=<K#�4�`�J-#����	ƶ�`�fp6��'��Q6���W�l��$�|@X>��a�k���!.�6O�o='Q$C�n�iK�����p��}w<�b(Q����,�C��O�.\`�n�Qq�z�݉�m�CwwuR��!��Z��X�*�D��C��Iű�զ�Er����gT�co$fI`sw�l�!��Tor4{-{��f�&O�| ��פ����<��+�^Y�8�6�2K,��Z�A�|���%L��S�33/�X�p�X������)��/��p���U��>�;�I�4V����f^�>����W�����K8�-���y�̚Kˁ|�uU�i�Q�V�n��ʪ�ӡ�!G`�Ljl 7A�CT����e�'�8�y9<�@�r` n���|���65�;2��,�~��5��rQ��g�%sg��E�P׸��Ts���#F�S9$��C�ʲ+*$p4�΋��oƦ.�P"�(���N/��-ivNX��7:��U��>��N���!�=���-R�dh�}�1is��"�$��rr����k����u�-o���i�R{v9�w%C���N
\wt��B��	�??e�O����̗MB�Y�bý�h�TJ��Yi���!�p~�C����ZF��
��Y�M��Ag���9������n�/a�j8�G)�Ѡ;�i��a!�/�t�F�1U����Ь��6
�}�����ڵqnձ���^�hfZ��㤥���[C�zKը�H���	���ha!U��dx�6�����m�VIs�x��X�8jQV�,;��l_�DWlD_1B�k��Q�γ���+�����\�~���`�����Q2۱ֻ�r�!'�'��FŻ:Y�<����{��Y��Hڿ��;,���d6={�� �����\�,p��@ћg��`�g�>�/Xv��۟Y��
Bn�8���y����a����n8O���6�����s��b�A��P�r�Ǝ܇�X�"/�3�*1M��;s�&���'���Z����Bٞ��v�Bӊ�V���C9�J�!�T�a����-�΅E]���g��[���n�R=1�"���TG�>�-G�e��PW)
���ǈ#�nv����t1p���$��fCVJ�$5^	ޛ���k�ʅ�;���1�����U�<�]=������~vE���� iԁ�޾�%g��;}z���;�pg���hT+��R�e�&f��A���?h���JD?��=Ѓ�"�0��5p@�thHWaJ���ѐ���ܝ�9cBZC������bG/TcWΣo�@��ض�A���c�?���*�M޼��"�$5�]��o��*��$Gz��Mdl�`�)Y�E`᮫���$B)�� @�i�_%�ꔀA�|<�~�w!dĊ)�M��Ձ:-�ZL��(3|��"�ܾϲ��]3i`-���!�;�;��ܾ��I��dti�5�|o4ݻ[-�ު�����r2�O��Λ�f���&���|;؅P>��9B��4���nz�)@��u :��4O�����ػ�G�<�?9�_�"�� ,a�A���J^����U#F�cj��
إ�<�_ 1uzZ��|8���i@�3A�@��\N'���)BVl��,�)�>��Qj�^P�/����2l����m=L��n��y���Z�&���Éq��#�7hD�hsf�04R�x���O��c100 �(�F�������v?c�]���:�g�u��j3���$ǵע��K$-ea��Y��
H[]C-����X�I�4#G�P-��"�\��#��UXG��ɼ^q��GC�Ϡ��/s�gy�1�B�硠���=�j��*��Y��������}D?��<���U�}�rP��'��G���'v6z�X?�r�=�����|3چ�{1"�&v�CR��A������K�V����8¯ج���w`���}�,��8�il�5��N���U��z!r� �刱xu��l����7P%{���sm3e�G��<"�k���Z�A�����N���h��#�Y�.U�麦��J*ſ�Q�^+�h}��8�h��Rr��p<��6���ya�a���O�3-����Σ��lN�t��vT����p�ҙ��O��s� ��o��?�>��#-Ǐ06�|�st����ͥ1|�~����?�w&��teU_:IN�b�}���{U g�Y�zI�?�jd�������ٲ��+Y����H��9�Q�B�4"�A!H&�#��O6��T;�n"�e-x�|���Ơ�D����A;��~���-��E`eoF�q��J��f�6�d�5D�Qw�9��T��y�௫��^�0^�>j�PRL4}d��7��NR--�!e ������P�?�3O���-��<y�&hg�/Z��[��xM��~6=ӏ�_,��֤3*�~s�\�����|᳅E���T$��|�6+�������2���+���_�tO�X"CD�S��2B�Sd�UF����3J�ݫ���l���x�������������b���G���̌���{��`pD��q1��==u)�O�R�줈�dP���rlñ��4%!�V��՗�+>��p�͇6s�N%?��!�K�����AY�/ɟr���T�����/? 7�w����8Ȩ"K�RJ����W2��q0B�H�3&�י��b�$��K��b0C�隘����5a�T� ����>�I�Mci��D�]"������c�l�/�n�м�y���XF��C"Ey%͎��4l��5��"�fG���"U�"+W�6v=?̝P)Z�, O6�F����o�=�_JP�ڸf��e��<{^���@
�P�B�fX���fjį� >���x1�,%��9�~]I�y\XqV2�&{�L�"lWW��2o�|��(U�9���
�U靉M-{fJLJ�,6��6F)��I���g�+$�N<\�?>UW,�
Rףu�[�9֣"ISO��-�ٓ]{|��&�)dF�������,�1�.pg�}�~�G����V-�V�� ��Wg1�5�
����N���K���^{�Tiζ�4':�dK�E&����Z����XӄRm��UtO���`��2��߰V�?�����]f�ܿ#Ldw)J��'3A���%�|��Y�S�Q�{���8�%Hֽn#�9ni,1�j���x��Y��ԭ�**�@�?bgP_���ҙ��)_�C��9�8KRv���S��m��:�d
��~W�Uh� "v�$���ź�6[k��u�l��>��M�~�Δ�����M�va���߂C���	���_[�@���aΊG#�@�<Ȯ�����c�t̀r��i�C�˥��R%0�q��^��� @��w>8�� �Z��[9�t*����zM8oT[Mi���v�~8�:hi�w�LT�Rcuk�'O/ 6�vѡD�)���}~|x�1���]>S>��� ��j���-������M� *<�|`�Pĵ3Aa����u_�� ��ҫ�>�rU�~��'9�J�W�}m?+�%KO��7�<�M`uAߪ� �"&߼������I�
�8AKt�$WF�A?ve[4��
ɺ�hu˹27њM���4�["���Q��Lá*��X����;Fў��6s���"	���nc���o->�t%"�.+�\ �|=����d�$;�t� �)XMa�gD�G�
�K�����[$���oC,g�ŧ��J&!p�Ve�t�,��0>b	�Ϗ}[�h/&&�っ^�yֱop*�ӵ�i;dy�,�#�ñ?RK�,��}u^�)Q9#�^:��D�ͪI2{�S),�D�YK�"��iL$����?T�LEP?�]V��I����.�!lFE&<�D��YO������ƞY�,,��Ug[y�p��ash���-�_S��ąMC�ɶV���Sn��������e}ok� �z%e%��6&x1D�蹮d���Q}����>���Գ����Ť�ޘ���x%���R,�1����Eۗ���2��M$e�C!5#�iQu�����(�i� ��(�m�0�f:^�(`�����OJ�+����DwJb���i�����*mO%QD���^3��1|1�ˠ��*`��'
d��!��61���]-�Y���;?ts�]�d�Ga�db2SM��B�K͛��K����; ���]�h�?�_\4VFk�2B�gK�w26nA�䉅�H�FC�O�8B�85��65�]ԝ�.��&�=nxb������>	��bw�dF�$he��cy�Ķ-������}�cz���5{"��|N��3��kb��3v���&m�c3W^�� �s+���`{cs|�s�eSʖ�#�A-�a�J�?�Zg?���oԢ�2wPd�h�H��l�mP'o�Jd�Y��v�9ϠG�;a�/�� u �%/��~}�@s�
�ݾ�&�#߄aΜ��l;�@��v�6�2̱�P"��E�������[H�i��31��(�q_�(k� R|�i��\�����W�h�P�]��ZV�q=ݧ�$\��WO,J��!�I�ȃ��m~��9��K�/O�MnI�Y�~*3���V?���$�,�z億�A�]X.�i
���^?+Ǹׂ}ϠH�DgY
K}�L�`9��06��Њ�3�@5�֤|��/Im�mU��vҟ8{v2�:��"eUQ�f;�ZQ�7o<Cpڌ���
�'�y��k@��-�M��R�9v��4�N�ap��~���g���G�V��7}�/1IR%�`9 pQ��$��y�� ��f1~S����LtW�m��\���­�j]�Á0Z��Pubʲ����b�����u��k���
o�j�:��cS'��X=��4#�� x��2XCσps�kTB�����Y��قP���i�x.�u�|K�_t���3x��O����x��+P���3�K @�ϮKXZKQ�Q�dj
����r�3a���EŨ���38:���i�*�7¨Sϡ�[�%ٿ�����iHܾ�"Nc�k��ߘ�'�o�8������$E�:�z������z��x�6���^ڇ�r�"8���c�e���uTD�B=>ԁq-LsthF�^:�y�
������']�io��N����PvF>���s�1���7�\=��)d��}�u�>�,��X��-2�	j6�<��?Ϯ��o��q�-���'g��$��NC�� �{|M����)���d�7��[�a�X�!~BC0/$��wH]B@tB0T�hEL� 2���R��ET�M;b��5�iAhϊ�����3�B�ʔ�
<�i�h�~�Y��n�. (¢Un���_F��*���C{>6�l9�jU��%3������*���3������d��^1U�֊��Τ5�a�a�����K��F�@����٘�	�U�߻.���l4;����U$R�d�N�l�,r���ڗ����H`�Ke��ˈ��S��U�_�=���!YfL���]/�ڣ!��ݸ��M�����v0��G�6w�JV�rhڐ^�e�K�&Zh�>�:�r�E�ک�T"�gT0+�s��H�Lts��Cp��_�![H���ϰB�k�D��%'��R2.M CM*K�Vo�*�-ty`T_��}�L3��fC�_�"N"���α�P��;Cy2�a�s��'n~�����r��3�,FQ�s�̔�Y��	����>>PD�Y>-rt*���[��F�R��a�"׫W�j+t�zs9 �+@I�� ٵ��!����n*�l�7sW���Z��L7M:DxBd��G%yd���0�yL�0����Y9��}���|�s%@]adE���1o�bx�t������ ���(A�y�V�F�rͳ߲�O�4Z(Be�v6�ρ�Q�w;�Lj��Or��=��9��Q'�ĩ�
����XM�;���?lIcjH�|�dbN/��3n�ZD7-0؀��7�f����|i����-d9�sL���9���5�SR��#Z�\�bt�9CP��g�UĞ�|oĮ��O䵾�P�[w�t�T��-<��D=��"���g�/Z]����df��Թh��|���� ׈�6�q8�~�D��#]l[�g�8�|H�!��
$H���l����e�yVc*Y&"�_����y�o��mB0�}� <}�6hI�U�!�-�8�9V�?.�p�u��p����a<�m�P�J����[w�"Deo�C�3��撕���7���3�8�I�o�%y�3�\����iطu�5Ɯ��3�V"��m@bl��d"R��4��ާ�
#�={+k��=�8uCl�S"�36�>�Я����nuI������G��B�J�����kg(q��68���b����̶���hr:l�$�DM���Ѐ�14�S�����h,)�yu�ovg7-W��B�A�5k�n;I�+�V������x�<?	�m�Ƞd��;�?yw��76�1�]�r�2E½MCO���)�B�k��L�?�&Њ��f���(x��{K}�T��DEq�K�e}�f��)��̓���Ԡ3Cf,G]�(2�����E�K�����(l�
�?0,+K4�99Rk�1���^c��j-�N����V�v�� �4I��?�b�}���:,%���]-n0�ZW�M��]i�v4���ù��Z��_y��k��B�=�D\A�}�� ����V�f�����$���5�P���C&��̻]��A���"ypt��KS\��D�U�w:��1NY��&��v����Yn�(��h�8��I��V�}Q$x&�җn�
Wb�F�RE�[~A
r�M�yK���!M�3�o�md�4]�B��C�TZo�cP&���~͹yV�B���=r��Ri���WI�k��n�� f�g��F�l�$u��yTJ�SC��9?ޱ��@��xO�D�N|�q}���_("؄T�1�mQ�j�O�P��B�~�A���/-��B����K�]���
i|���.$�~(�p��çE�.e���k�
5���k�,���Aa*�ۜ����]y1&N����f�u���'�����v7}zP��
S$���e	P�Y*w��Ѐb�׻H�{�1~�z�L�J�g�~�2��D؍#��U�ɲ��-x�p%�j����1G$ ���Sq���PC}H�p8�RLϮ�����n���3|c0��!yF�;V��{����d�:��d�oH+����c�
s��d�Y`����|��1�z9kip�����`��ԥ�NM�'���ZA�u3��e�tcPqt�[eس]�	�ݕܾ=�=u�߈�Mf`Og_���q�W��/\& ����0Nu+v.��t&W�{��t�Z�jC]�N��q�Ы_J(����w嶷���G�߃	��+���~�7�=h�B-�E�
�s�U3�ܭ���ܰ�_2����2�sv���Z��j�91@�@�F��of�&��nN�ůo�������/A�R�/@a�2� �y��t{�r_^�#�`?'7|Ҷ�9s��ܮ�����B����<�����"�	Q�L��4���O�r�G�������$#�z��E*�5��]?��Bgw��]���JZ ������������\� 6b�ez�m�T#�|.Z0�@R~<\��6��X~:8:5�C�:�Ap��xk6���+�T`�W'T�P�,��BJ=�c���ݓ!!P�Mmi���:������]n�������;�V���I���]�lV4��PKj����`�J������⬭+d�������bi�R���=�8�n*�c�M{u'M��*<'�kT�ApB�LvC>���l;���`WZ�U��6�4�����Q��X�X���b%�Ju`�w� ��dt��d��P�Q�-�-$.�S����9����.���2���b��g�.��:�������U�[������zatY�xw��<O��C*=��Sm�I�!����>&B'�!�gt�EC�����=�6L"���1mQMˑnְ�J�[z^�@Vs
:�<��B�j�Q����)t9�����v�ܕG�2��!ɃT�؎-o �dX�`���;�TLjPD�ũeQ.�2��ګ#N{Ͼ�T�bD�)��}�g@?��ſ� ag[�h?���yb�7']�Q�u���@�$��7�|�E�N�t`�)T[��V%��ybt��(+(�����8�nġ1no��\�0~� ��(�e爂��h ��� ��;B�Y��@M�H;U��]G���4&k���Y.܈���,! G�����iSa�W`@J�Y���B?B��@�ݩS��R�E�Ï�xzJj���=]�'̑ �2��]YQ`౞U��~���>���8d�X��e��+���,�8��]�d�8� [*@��l���PfrN�e�����b�]0�adc�9�+c����t�Xm��5"��b?�p�t����Dx��m�S���H@U����I�ؗLG��(�s�N�O���\�Hk��q;'�4�Xc�*N���^�J�/�#Z�Z�_0�	Zi���X��u�-���!zd���v�߮�f9�6'��WP�H� }��䪇2ݏa/�~�8J*�SB�S)��sv��8�\�{g3#�<�CLi��`���[/�����Ŵ1%x���Β�IKo21����)�w�h��}� ��=�ŰK�=������OQ�D��WQ0�xve��f,�:�3poX�$��m?M�b@N��[4a� �ʖ���5��"�����ȕ�C�;gҘ�2*0E��<�j|��r�$\)Y4k�I�D<Knn=�@����6�]Y��t��#�X�s�濷Q�մ�cG���Ic�\�4��$摦t2t/5�`�d_H���Z-�*Q���B@=|3�<׭f�ӆdk�~�ۙ���N��N�Y�ŴR]pe�����sߝ1OI`�)2-U����D�F���eH��c�����f�h�B}���|W�tO󹄂��h��U�e�f�?ϋ~G`#�R�My�/P<h{��U9��&vk��1�R��<�����O��*�̽����@ʥ�.7�d*��.�t��F&�N��~f��J�N���T����U���ܽy�8��W���d*���|=�V��@k���|��h���R2�?tv)F�b@V���\ ��ё3�� ,w��6�=�r�*����'��K�վ�����d�'�w(W��wj��gϲ�Dm��]��x�]��;��&O���X�R �1�2%�MVX|ٞ��~��EVWL�Z��]��+�}�\M��Q���\��53,~u`=W}���?�E�T�(�7H!j����d�R�(�f�j�ѵN��/�%�+����Pq��"����ͽ"��C�(z����4Bo�8�;�1a�<&�ԗ�5���|�3	m����VäShz��?�� h�lW]/��`֍B� �YfO�m��� �/dh���''i+<4bt�DR/½;>��(6Ӽq�C4���p�C��/Q�@k�%�P��Uf�����{CCzGe��6����:��JW��uÏ9��+�tM8"���}"��v�Ic�CgU��	��T���}� ��c�����M~���O��wrs��k���L��� (뇟o��D-��Cä��{T�$��[�-u�xw�J6��CnO�~�.�a�'gN��˻K�ϔ���{ �b�K�+��ͳւ����P�UoΡI��/|��*'�MS���5/F�e5��1��m��3��4�n�^�����?�\�B��x/Ii�������J��&�A�������b��_
�I3,*Q&9.�g~�TY�:a'�>&$������h�|ϱ�Aj%B������H��^<�H�~:�|:�|�U����>y�Q���
��s]c�rb[�nȃs<�BԴ�O���f�쟑frlǉ�Z���c�(侢Crvn��_�{5q�G�K;�?��>yz��5��UVk��S�YN���X�[W��-G.�Ⱦ�����hrS�l�U�>!S�_ԉ�D���1{��čL�%�_��<̮�ڗ�I¨�2y�_�$
e�ӹ�7����5�؟�0Z�2�Qn�ΔYS{���ψP�	��w�@2i�ɧ�d�X)��v�U�����S����)�?,�� |���KH�����֓l�4���*�|�M�D�C�J�)m���Yr�x�}gZ����Ց�}4��>��J����2l=8M��z;���C+�D�b��El}� t~�ŹR_���|���A�� Ú��j��c����#���2xC�jLE��$	"M��!��Y1�47�5�k����ݞ�b��P���� �㷰�l�?YT�HgDӆ���m�}2�_۽';���&K����? 8d^&A�[�`���?��[�@�$��F5=�������+F[':c^����JϘ$ >Ĺkrvv����wSUᶒ�J�
�ұ9�q>o�O�nG���s�O5牟������E��h[�C���v[��5�����;��;h
��SyVMٟ$��'K�&��R�e����򕨧�8t��L���A���@�����Y��>�0�t&����Ċ��e���X�l�e2�-e��;Wik��!�����x�]w2�|ւ
hФ�Uy��	��o�2,aL��Sn*,���Abq�#����6|�Y��4�}w�Ş|�e��P�.��6�"
�I9�-WH�Z ,����k$8���lZ[=S�����L?�~{��g7�����|p��������h���FdP	��X�'�0hՉ�5��z�/دYFm�)��HP�=�Ň	�3���ޚ�g�.:-���
w-�H��'mG]�m��3�:M�w���ڶ�x��C���Ɗx�]gU��/@]}z2���9>�.�qtP8�@����y���N{�\̿�_��%�0�$]Փ_�[��h��3�Jf�ZDQ�S���?�����^��a�n~ �"#�=���C4��f.j�87���Ə�}JӾ�knAM�������?�J�<���d��p��T\J��e|QD�7'l���}>W rj� �L�!|YEy�d�%h�sJ�j�f(�7��~rr�*ޢ����]w�}�.�+��g�H��e�U��Ji.�v�>��x���;�<�n�~��w��t�#h���,-�s7�m��ߍ�S(e�ب��L�Y�Pݲ{�֢�X��M��Qw�C�4`�;&9��n��w#���[�=��+=XOr+�H�`����YEgp�}2����s�\�0"t��U���H��!�� �}��Aħvb�_{������\�������>}�"��9, Z��|��/U�$�w�'�fz��1we�ps��.��0;Et^�L��چ����2�5&}�E��	�#�@��_PV����>4��iy�ay�k-Vf��{���EhjoOAPn��vk 㫟iӴa��Q�`�/\���!N�%8e��?~���.}a_��
~s��~~=�*6ʮ�)����~AųW#˚.OǞ~�e̋+S��t�`ƃ�|'$
��L�y��V��/���C�x�)���!M	��-�A��V��*�7qu���`ߤ�;2��S,@��_���`<i���z'N�x�_�j��\��t����CJ��PƵ!t�.X7���j!���"L��~G�|J��k���
��tk��&��6�*=���I>1���t���k߆p$��xWa���p��T�������l������0�rޫ�U'���JUp�~|	T@1�y��+��*�>ץ� ��ߡ���1�	��^n"�6H<	g���/~�{��4\�˿�� 
p'�5$2��躕�-Cmp[B#BT��Z<�����jC�1Kc�i,}�XLm2��:Q$t����s%iW�A�}�С4�s	�0���9�T��w��7���i��J�Ah��C6ޗ2�u�v5�O��@ݢUA�S m.8%{c�C���86���UZ��t�!S8q�X):
'��/�����X�p-Y/�F>�>`��S }�V���E��}(����m�X���Զ��mݬB��� ��O�j����
�=�H�b�C��ؿ~YVL���$�:�Q� ʗ��k��3Br� b��w7���{^b��p� �U�&��̜����+�a�\�{��K�����xGq�c@��	/0�e�U NMD7���c7�)5\~\+���Hj���ø0�@@3���kc�ڬk*	S������pW*6s;NA]�n��cy]~[}̓׸��UL��E�D�����D��L����WZ��������0O��lc��	Lx��I�ӡw�VD4*����h��^���tS�E!�����7qf]�_�%U�S��h"_��9�ʥ�R�r�5�ިai�̧�.�"@��{|�w}Z��]��Ÿ��G��k���D,�N�w�?���s��o�sV�i7�/�3V�P�6����L~� ?�^J�\�s�l���n�?C"��i!�}�Q��ĩ��������ov+�6b�'5nd�a*�+�X�UU��3��5�1��Q[ ������7��5�v�l�3�}���|��Z��$�l��ץ�i{�m�i�Ҥ��1>`dM�����~� �L��d���6I��Y5����Ŏ�d������I'"�+(��h!����T��} �6��L�V�dy~]~�*R�L=�4�ДY�ꈆ��Tt#�{�'K���*��"X��=�dˆ�y���ʇ�Rk�Y\@�� �+���X�{�u�v��P塶'$ϫ�a�y���������`��RU �q�J���~��������*���;���D�芦�9>�
+�ST|҇������/������)hXr�����-�fF�1t |o��J|������zɰ��#�<��=��ju�I��o*y$�U4T�R��mb�y�en��������w����zbmL�<1
��f�i��Bt1�M�C�j���և�E��!w�ʳ�Pf4e��J��b����&�a�=�g� �X�i��L���Ǘ{��jv�f-��n�Z�Z��n�����Cc�`=<����7�o-��!)�H�m��;�.JNS��M�PC�����$�LN�3r�p[;h�o�$I!-����@�s���J�}D�C�x���?i�h��l��j����o��G{D���P�����R��G:������1|O�!���  ��9F.$5p��zT$�I'���w�6�����e������E�EU K�A�{.y��#[���h����-ۼ�R� %���[*���ӆ|�VW=;T\����`!W�a����pƴ��I`�eC�Km>XE#��	l��� �ە�@��/�f�G�׳��C����V�'�S�U��q�N_J��17�Áiv���gF�wJ��P��l���\�!l,�(��]��z��Y��S��k��%�m`�P�2 D�Y��Bj��N9�����j��=�=�26*�Wh��e^��~Qi�_���H��1���ƚ����<1����s�ڣS�S^�^��u�x�]�4�������fɕ��?'�Z�'yQ{,[����Y	 hPıv��ꟹ���³��'4�=�)EOɎ�夏n8��t_nS�,(~�A� @�ߥ��&��x|��8�E3���[�J7J����Ai:��.��yL3�9^T�\Z]�ч���!�E���wTJ��;�K�Z�-�7���A�wl���E���/�K;M���X���=[v�����X'k�����+�FՑ��L���@����f�`�`Z_��_��.�)A#ij�����)ݘ(��!�_�|�"qJ��%�fz���;�F.��d�����h�:N6����!^^�<�A��K}���N���N�����Ҧa��� �Zrz�&�@(�Y�'L��өȋ�H��<5t���������Z&U�rR���P7��dp?=��f(����0�%����@"&æ0|4)k��i�Z�����p7F��"yGV�(Z�ȉ�Br�J������vWU�#�͈�l(���2��~+����*�E��Y�������¼0ׂx���R��t�J��u*���x���7��XoY&fR'������O��q��"x+M����thdH#*]Υ"rKfƌ��Z�hgqW���RNΔ{-��5m�EL���s���?�H�'vqE���6��X�ixB)���۞�H�0����N���*��f_��m~jD��?�í	�)7��ν�����Y[`@ O��.����DQA���J.~63k^���E��~ݥ�o��a6Væ.��#�"<�Q�e�Xp\/="]�'�`�]�j�3s��cvU7Bx����pK3p)�=�{�N�΄�2�vᾂ/����ӯy�I�^'#�ݴ�#U���G���֢��'�?�r�����V7�]DڼF�����I�~�D��E��qJ���XI<b�D�Z��#�Sǋr��Qf $�]
-��o%�-a���_Ϳ� �|̶�MTZ%���{oI���=cqv-c"Oݲ�\�<p��ݡ�k�$I,"II�:{�*<��~S)�r50�U�1��Ų�]x^(#�T��o���P?�G�~O�[�"{{�\�uL.֛��8b\��)kڡN
��kՐ�b:2�;��K��{$�pqL�bca�ћ�A	��h���}�X�Ws럙��w5�9g믧(sCLc;12NVAB��jӺq�>4�pӀ9��,�Z�t��+����DJ�Xa2$�yX"�c{�,zC��������*�t�ƪ���{g�)f���@ꊢ#�v�/�QRi+��$,e�Q�W�ƯZ���!�)Ӌ�A_�LWmw=���[�*c��K��|�胕-P�G��G��~�wA����w�׍A�CM��{�pV
��f�<{�3���B=G�5��j��j�/`uE����[{��?e��xQ�VF����kص����@U�h��>���0�ëk`\x=��7f�z1��x��qve��
�>&��9����i�kl?�>�r�yԞ���vC*�탌���-�\��(/���r���=�%���)����b�4����Y��\��SX��a�w����~˥��\�b�������+��<�P���5�o{��,(�`r",܁�Q�zΑ����V�C��P�'�aeKz�|����E��<�Nх�L[��K��s�
��HϨ���5<� �`��榝�C-Ul�-:��\��h�	/v��*��3@������]�����׸�t�K 6o��<��V��
�ST-D^�pޔ,�:�g�]�W��:� t������s/�6��*D��^��n��x������a2�tnL��Z�닜7`�1D�c#f��J����%S��q[�75���qN�#|��~�>��|rI�OΓSܡמ��H�e����KJGǴ��P�;�DD�/
gӥΓ����I�s�ڵI�=���C��:JvG���f6�������X�Xp�4Q��}��J��5M��Z|������!�$�t� y�^B����X=�u�g�U�A7���JF��$h��O�O��z��G7f�N"�a�����2��K5v,��zHH�	z�3�.Jt]��
Q���F�\�p�^�G�y�g�کn�@0�i�b��VBr�$��z��(�4��^:#��k�,�~0=�����h��u$o2�L}�",�5�����lFX�& ��@�ז��_������a�=kUQ� �<ِr��w���p�k��#焽Y�����-���!�y�,��v|F��a���� w��\(((�P���;vN�%]���R�*�ɂr�	n��������RC�D������Y���%�*l�&�t�����? ���-�����J�a�9�@�y�缋�ϋ�Yn���^Oa�m�\Q��Q1������|�i����$��ݨ�u�Tdik��|������=^�,�~��%���G��W5D8���Ug�����ص�(�U���� �x4�
�m�|.>�|`%����֝�,�G��A��Y�H���{�O�Bo��.����Lܶ�Mۀ{�mA���%���'?G|ဪ�#XG�����I�,���o�&L����B��7-
��>�vT�_��u;��t_v�_��(�9�nh���= 9@�t�K�I��
1S��;�+.{##
�C۱��ŷU�4L˒xc���58� y;�a$����ģ�F�x���J���_�ޕl�3���ӃtY��#-��� Ѥe�-����ww��S�'�r}�u���Ǿ�R/��
����-e��۴���Guɛ�������x��o�S"�7��)�U{�B�D�w��7a�&�o��X��<������vVGj��ݝ�Td�)���#,e���VE�Fت�('�_Lk����7\�n:��1	Ƙ�����$�:��0�y�����qЛ��Re��=�:����_���G�$ϣ�:��"W�Qk=�#�	��`��|�Yӫ��NQ&�\M��HT?:��qQɊ��u�%�r$j쵪�,�=��fŖ�����:�3jU܁�W}Ҹ(����:��O]~Ԯ�=����8�,��u"{�A᳏�e7S�)kg�f�[��Y΁I ������"/N�B����`�ȇ9������0`y�R+��(��ō��[~��a͏�=Sp�LX���Ư���G�� ��$����e�Ж���.�LA���w���Cc�a�s��C��)́Z�OY��U�t�(	o�x��k�e�X2��4�l=���7v�����	E��s>5�(U��P5ĸ��Z7�H�B6���Ϧ���1&[�j[B/!�gR�2?p�em!��o6��T.�I���n�`3����ѡɾ���#����$��
�ͥS��V�Q��;�����b��f�#��Ҕ��Ux���F��h�Cήc5�S;p��F�F���w��'��0)s
�pla�D��]�Cl�LX��fn^�'$s��*�t�b�[2�e
=�*�8_�%���]%�H��է ���A����]��A�ڌ��5�T"�0nַ.�`�3���=��}j1���.̅S
�.�"Q���Ӱ�gz�� �@�2�jԪs>�퉻9tU�%@��a���?BWa����!r:�r��]mߣ?�F8���F�^]��0h��p!4vWݤ�"����=ct����0�fA�!'E������f����,ݳw%$f��6s��%�����5�9��}�ܠ~�8Ȁ���uk�X��0/
�h���io=aco����� �a��	O/_!�[�⶜�+�+�`b�P@�3Nɛ}8����T�0��l��fY�2�k_�6K��'�Yi8����cY:����6��&�f���yn'��2�UMW���նg<h#����`��>�����X��Lq'��Y*��D�3X�	6N�Ew}����O�#�Ԥ�.DU �,%��c����r#���c߿hq�:����U�����
���c�;�E�Z�0j����P��a��(<�t�Ul�b9�{y(.��i����h���4�'�]xĠ�)��iP��3�3򃾛n�͵u�t[��rö.�T�]�tx��&:)E���v�cS��`�/�߲ا��_�]��-�E�d]�v�hV)�봼�(ay��y)Yv�����HFd����S� ����%tmn�@��ƣ� �G-Ҵ�muAk�P�;����o��/E��-�#��M?�|�}:�ڼD��+(�@e>P� q���!?��-;�>A o�*j���j�q�'��Z�+��[�S%X��Cd��?�Qu�~�|*��ӿ;;R��U,�`��/4�G2VU_:^�{��ar��i[L���o�E�W��f]'`y�v=�_ ��q��yq��֕17d�sM�\�7���Wh����(��yHN����J�|��ݗ��p���Rǘ�`匄#�k{(
��5�u������g�/C��)`���#��aEZ��X�?�߃ ���}7pĲXXx�	�D�#<�-`D�{l l{~�~3lE�b��M��U�k&�x;�7��ꐂ�g��3��=��*"X{m� �7�gt�.�W�[QG��f�у�m�^�뷍W�(]"7 ����y����MD��퉩���v�瘜c��2$�Թ�$�/s%8S��MW�7b?By��i_�y�gc߱
V����\װ��
�ϏA�E�p֐o1~��qw?B�L���l��J��!{����w���Kҿ�}�����^�!��4�NnP�5*�%���|,���-CQ�H_��tWM^�#ַ��Bw*^�9��7ި�0;)n�4���ܤ��°{EK�E����QI8"�ܤx�]ހ"��y�{��Q��y�V;�@l$���=�z�ц�X>�<96�	#O?U�����r��V�=B���|��D	ەޟZ@�A�_B�l:�?7�^58����M2B�r�j�������ME�����~W�\mP�"'�Lly
�p�6/ȴ�g�g�&�PM�a��i���_�|�l���D�Ιf(�_��VL��ʅ;������D(a���@m�m�\ah�ws"���gЅ�]��}Ĉ���^-T!b�H�{�Y]w��;�NP�嚳\��?�5�Gvx2�ѕ(?�Z9��e�*�K:8Ͼ�,��ժ��:ᎊ��?�OD��j_o{�^r��3�l��R�	cG,�5�_m��J�Dz����zpP�@=�!z������`!v�݆�Ċ�l׭w#����5aØ�W�L	���j����7�	,J�R=���8�$�l�����g3l^_Hf(e,8���'�a:����4�Î��b)	��xp��z�q.;����Ӥ@�γpƆ��='��~��$Js6�!�\{6�0[�W�`��G�lw��I��B�=���ƈn/�����L^���v��ղN�u���c�Q��`@m�N�B��KQl���B����h��c&e^�!9��{�H��

B*�lWH.��u]�-��c���{��1jْz�h�=����5�Xg�J�P_��f���_acR�4�E��>N�/����u�f0� Lu�<T�;���	��qߍʀť0��Ǥ�qhFJ��53nO�voި@Ma�� b�ZnUo�����.�ZV�K�#��!-�씬��m��"��F9;�PM����8\�$�1s��m��	a싖�9$0����	x��S�I�Gq@
i��
7�7ĚqqMs�>[���#k���Dzo86�ސfOG	Oٗ��J�M�\ܧh*d�V�R��=�x��^�bT���' �tK�l�g��i�p���f�i�-��	ѝ�p>�eBlh'�j1�rIAxt|�+�8�|��.ϕ����愫��1��Vc�dK�c��{�If�>���k�#/��mw�B,\/4G�r�@�qi��d�5����IXL�G�ٍ0�@��j��X&��9��yxl=J��"������ux}�=C��� ?�1-�!J���7�7�����I>�=<'�j�]�ܖ���ݛ"N�;c ��2�K��<!�^�Su��៚t�M=���v�A�@�k����gy��>���֛�>���!AӬ7��S�6 �{��C���jsPp쨷`ϯT�\�%�RYsWe�ڵr�/V`��W�`��b�.O��A�z&��S���^��3���ܐ�o�[;ݒ�RA]��(ȫ��h2�X�Q�����&���f�BJ�1��@T5��u�BgΛ�U����`�2&`�,|�Rb;#f���C?�Ϫm�i�|��P&�vG��?ݑ}��`����_hɸ2�T�y�
R� ��I��3Z;��BUb޳[0DͿܒ~�.e���$�{������+&KI�KV�w�?3�b�cru�q�P����b�*Lj��}��z�\]�,O��ewx�j����Md��Lt$�\�߮�Z����L�r=�|V��
�\U��D��r��p6��vlW�:7R�̘hi�����>ɲ,I���I%����e~E+�=��e�Uh�6��"�	����\ǻ"�b?^�L�2��t�=�*s�`2�kNy9K�j���l\��]2��BN{��K���9T#�|+�?M�o=K�5;VZC`�����Jo=�M���p��f�� g��8F�\�T$�4��e�Q����9vA@,`YjR�e�ơ��� <_������whk�`�Xb�ʺ)����l]
�JQ�i����cH�~,zs[.����J#7k��:k���	CZ�WZ��������1��Hپ��2V�GS����;��r���}k,=n|�_=j�?���oJbnb����3�F6�����z[x�1/]��f����F���L����RT�$���`� ���Z�R�l4R����}�T3'J�N��y�Y`���G��}�7�|��l�����'����"j�X�Dsiqi �'��*���M��� ����_���/5�+�/��UYY*-�j�f����ʈ~l.5����v���:{����I���q	��e��<�q���tz2h
���3��^������f�R4����o�O���3�
K����f����fF�{�,r�>�ԟ����nO�B�1 >V��=�
8i�[�x�_�T��f4���k�|�zlCj�"V��/�������K�<_x��v�(G�*�]�	^�f��0�U�҄����'�)�Sxa��z��Y���A*�<{4S�s-Id�=E��j99@DN�y9���E�b�[g�� Ό�bo�%�xN^ŭT5�$�p���z�<�)�d����l�p@Kc�da�<j����Na? ���KI>A~�A�?���đVZ5 ��:B�*��̩�Ga�n���������������GX�
�p��� ����a,J���'�
� �TӐ��9��C�U6�T.
�D�� N������sHw��6��$����������u��!��:���/����3�B��.�.�U��Z�f:g�r#R���׀W�k�P��7|�<��Iapz��P��.��n�b��Wj��t����8k&�4A�?N�n�&�V�3�
���rw#ŝo���?"*<e#�vf'����m����za��=�vM����A�s�$�JY�Iy�u�ʹ&
0z`s]���V�s��A¥>��M�j�O�W����x�3�s���@vA��~�Zʣ���I/��f�3i�lvq�A�I��H���P�N�d�ݷL�}:����/�%�m��.t����.˨�����	��+�jn�_�Y�_��� �7��Ủ�j�Wu��)�5��B�ſ7��n�.�aD ��h�s��T����rD`�}ѹ��K���'9��OB����W�&��+VD|�}��a�r2� ��4��2�����{���[����H���ߘ�c�Т�H�����@���'�Fn��H2Ɲ���询���'Bd�yp�f�$<�6��,���~ѝ�����8޺�?�OM�>��Ί��,Ⱦ�07�8���o�� ,.���;�}�3[LFu�Q_)L� �T�F�d��B��ŧY`��Ͱ-`�ƾ�@UR�/�W,`�Ƭ>�p	7ҽ;���zQ�k`�=�7�˝[��\(�ϓ���ܛ���c�*�h(�^���xF�g�J:�T�t;�ʓ�+yo��g���}K��j��?"a�l��;8q�I�rth�{Me1i���R��϶n�W�q:O����k�  EU[s��J����<u<����B����ngS�	@��i����� ���TwP�����~`�.����V;��W�0�Q��0
E�Ǫ%�g<t���=��b�Z�M}L_�g��Xi��XV������~���#%e���u#-�%��&���&�I����,�w�p��-)�j�����?���)g@�!^K���8T88D\Y�̱�����θsE��xd����X���6���K)�����g_��ә��/=��A�ן�ᡉ �{X��\��X։�:�s����{���Ip���:T�迓�t��i���V�܃�\�t��zR7�~Hu8��D( \|+���V@p��1���%���w��kR]r�ь�4����mk	rhC��r#�ơ��B�N�9<[s�`�ʵ��sD��c��O^��u�gekiT�LJC�,'W~��eI����t����TP��.R�#������$_`ˁ�8 �G�&��;���Y��KD|�E��U�f�dT��xՆ�r�tXBu�#��<��o�y�)ԟ��"!���Q�� �>JO�;"\���Z�u Ր���F��`Y�f�>-����&����V�u�8�[��Ry&.!!�h�SВ�C��,�����L<��f�
��%Ɏٓ��0TJB����EX����!���Z�@���unEi�h�J ��ni�X�z:��"֎ʘ�����K��=���&��$9y�U��~�Go(�J�V�9̴	��6���Ofst�M��"����e���O�`�^'d��k���*',��G�d�c&�&M����i�3��K�e�?�-�����8ܒ������=���ۛ5�Xt��� s������WBgg����ݸ%[�k�cڊhֶDQ�>�-
���n.Z�h����K����!hgQ"ۤ���6��fا�>O_���l��D���/�J{�����	�a��BB(sO,BH[R��'�^ù�)��%&��a:E�g�\�$�q�\���QAzv;�3�w����iN~�M��R��#��^�Ex�h���`Y�B/��G����dhU@�\EP˃^��M���y/�}D��}�+�f��!��*�RPL(͂$�5���Fl���Q���B<-���D�D��%�h��`*T<�X�f�~xq�'��!�t�	�A_�ڄ�=���|��c��A�/)���\��\-e@<�|s��O��oT牨=��]���n�H�T�'\�U1Vd�tb(���:u�4e�qO){�l@_�wTg��(��x�����X�M������B�#����$��<�_F�Eݾ���f�w��MåZ��4>ҵ�Bd�0r�W��Z�fin'��dԜ�a������{�𺠉C����n'�M	+���%'�'a���\6��&6�	�hː�n3vZ����Sx���@��!�9��e��W��P�%�Z.T�"�Gqӑ
m���Ĝ(ɮR*S��Pw�<.E��j�:1�9a b��>����Û�T�OV��XP����^��������8��w}伡�e�ǭ�!!��v���ɵA�־Q�,4şzݐoհ0����p�%���ړߘ��Kсi���JD�
Cp��]/$�U>Q�S�	�7\�hɆ��[U-`(-1�r
^o�	& |[����le�����퀐�Վ��n��*_���	
 ܕr��d,Φ�SG��zx͂���%�G�Pa���	c)�{	0=?X�=RF��k⮗k��E��d�@'�Ȧ���j�9JO+�'�qme;��8���*bY�"����a�
�MA@�{�rT���?�o��Zp���Ojϓ;D���Z]B�1��;8U
�UxK�I�}'��Oj8Q2��e�~	��x�7XWu�ߖ��q��V I=|>��Ճ$�=�g�X��m��u��N�9|�A�"ASu��kWu�ߗ��y%���C��|�f��&�F/~�0��P�ޤ�Z�63Ӆ.��� ]u'WG�)�9�G�HT8�4���$7��r��u�]�X�Wy����ŷ=P)�2���4;h��UP�G�[؀U���P�y����$�C6&rIW�"�3P6m�ѠB�	E�����H{�4��ESΘLu"�����
6X8xȗ?���@k �����%k����ު��;���1�L>X�؍�����8���mH�;�Ӓڈa!aS��-X=�A��J��"�~q�~�a�Rc�2����`�<;�N��1�I�t����㵯������Ӗ��gX�)��3?��BKz�h@��]�	-AX&^!�C!�9��2{�z��V��R<�z
�q3�4z#?�ԋY����$N�����r*	�@��jA��`t5�vɁ��,�>�Įl�(o�N0��K�x�(��ٸD?Wth�^@�3	E^�����
H���;F�xB����Sr͕0A��2����`݁�ARQ��)Х?��T��y����ʠ<���&z��t'������yR$G��d�݅�hm��	`�&���t�|�Q^�1��5c��D�m��x&�)�.f=�+���Dݷ��nl(� ��/1�˔F�;Ίkq����#ޙ�PeɈ��Rֈ�Azv���/g�/O��c�]�W�5��[���%��KxEa�c���d0�\Ba"�ѿ��ĩ��3��b�<ٟ�YP[�L��hp::l�c`�D2�TR��VU���B���=?�� ���y��Q�8��-a�fP�
v0}!�(�Zp��:ձ�6k�S��㡔B ��b�Js��L~�˓�Z���E����R\����Y�:%���ڟB9���0�q~�2�hw����Q�^���:a�b�"J��G�i�8x2qź��ER��ԥ�W��ff�gt=/���.���C��6s���;\�t�Tt�	��K���TC�&IW("�Ui�p�ݷ� @1���4
9^;���bB���f�z��U��n-vI�B׆�9[OD1	ï4wwZB������zy6/������Y!j�"qDͅW<t�߾���
Р�N��6+bcChrq�u�?m�1K��ŭ�7�s����pojyI}5'"��Cl���y+��gm�|�j0M�b���׉���%�P]$�~?V/���$�a��sܧ�D�Q_�rB-�3/����'��e�0�J6A*��v�y��5`#�j�AI��z�7�;��k��i2�`� ��r��`��
B�B"���&
��9�S�m�۔`��Xn4�iwj�u�Qe\:l��W!.D�k��*y�3"*g�Uw�\��i
$;l�J��)��Z��������@癗�5� Rʔr8�����7�����MG���Dg�X�j��K�2V��[���R��O�P�y��1er1I s���,�l8�Ti;��q|E&E��*w*<��(�i�P7�����ďǽm�R��:�1KǾ@�!��s�|K퓑�@��,0���t ��ORE�A-��e�Y��&�����<�Ή����S��!Wqz�B�������+�k8Dk#O�N��@�O�#��J��J�b���:i�j�TEh6�\����mǲ�Si�q�!�y�9ڣ\u���a�]bGV!H��{kf��$Y_,t���@�g��b��H���{e�uyхz�ҏ�G�\>�yX�#��*/{d�r�Y�b��n���tT�b�}4���T���� A�T'��Y!z� ь[����j=6��z�C
��U"u=+��R�����dqF�
`g ��^�Z�j,[���-,z�Zfqztw�an�Y�
�ÑK��uꀾ|h	h�e���g�)��N<drBx.�]�	#;�	o�5Ɣ2��}_�-+8����Y�P^�YP��R{�New���J���Z�'$8�M��"�^�p�m��3JgY��yB�?�����6�|[�a��_�j�ml�U�����N���T�o�"��\�uݙ�}��L�����;/8#$�d�H��1��`q��N����V`�^z����
.�5�����z&y$�{<�&es��BIK0����DIۂ2X1�t���2��vS��ړ<N���M5�&l�(�N�^��a5A���wU�b��e,j�]�zH3�QmlTGnΆ\����,�Ƿ?zOr��8+O�I����*�YL��w-8*���Q�M�:ys��84�M7?���^�4�s� <k��ރ&4	H��Ӭ�[���n�bɔ /� ��B\<�2���N��Ř��A8s?����-:'pf��q��o��
5��q�H��>̣�u!�0����I����6��\�Ʊ���|�^2D&w��7/?�/?����D#��� �dU}�Ǡ6l#�3�ݖ؟���M�+�Z+�h��б�~����&�����6�!��K%Hd"e�ql���c ]�V�qd�F�s�����;7#�Q�J�Z�
��+d��s�qP�'\	^n�B`>y8dX1�&�O*'��I<9�q���*z�НKy�sO�w>_���v��v$J{_`�<�S;�/�ݐEe֡<HF3���3/%�n
C	�R�vT2�>�����Z+��`%��z��]� �.VسZ��Ej|p�x)l��<�1U���.����|��j�{�����yt�	��:�(���j�8IC��TE��r5�g�m~��vɆ���]*)�%��`�X]θ���m����M�{౅��JؕllK�wb�Hc;
�À��+�zqp��m_6�<.H�{pCcl��g������6�<U?���a��Y�cq�i�gep*B��V����l�݋'P�(�{�l/p8�;	���*2G@�{ڞ��圛;=@
4�ʃ^v��{�A���ϚĐp���kGS����6����82�ǀ����í7f��y��ix�}�7�*(��{���nhfv��*Ge�hhUMj;���oAc8񮀞�w�"�#?�2��P��0MԖ*��ֱ6R�߰R����)��j�o ��Zg��)e[��%�Q��m�'T����)Bw��w=��c@sDz`|8��q���9LV����s�۰�*z���X����͗(��@�r��u��6�}B��b 7�X����x���*.һ���L �X����5A̲q�C��M0*�G��l�X��D�ψ�4���/zA@'�~�= 7Z�c#Q��%%��z��^�\Ə�⵰�Q�d��\�Ҡ�߮?�|��ʠk�������^�3�30g�āC��<���8�9�|>G:��g��{�V�Kͣf@ț���R$@`�.����S5����w�\��Hؑu��:{	z����f5S�l�%��re�?�Qy�xd���6)k�Ǘ_G��? "ڬ���v|*���N��8�Ag�l�[�y��o��9ݨ�p�m�
0݋&����Bj_�C�����X�?�%���;xc���O�~�(�[�I�Wu�zf�!��S?��p+�#��+Q'��B�7����˽��	��{��]����ߣ
���T�q�J�*�;a�L�	%��KTE�; �@�}�0=X-dJ��A/pΕՔ�#j�z�"ĉvx<����B�d8쭁�ԝM2��e���\��$Tbv~���R��	N��p��߻�Ľz}>bV��:��H�	�R�T�6�8V�t�L�v��8�sa�������<t��J�OI{p&��@�#��a�Ct$>�rd�;X�E����y޶�KnQ�V�<��gI�̀{Qw����ɸ$���c�Gֶ1[���adx���q�H���I��Y�Y��u�Iߺ+ps�O  �.�����GAn�BΞa'}�q�s}1$�1�|��튛���e�p:����? ҃w/��3�I�F}��i�nP� ��lA����0�j`Rl�����#X2
��N�������'	���FW�RJ/W*r1�q�5�[�b��p�D��O�B��k������:p�bv!kXM�G�����/�8����ޯ�I�	��m��t���
�4w���FF5@4ᗅ���&�A}�m���'M���<����ض���P��P`j���3{��g�T��x�UF��G�;)
�Go�Eř�l�s�ߝ���u�c���DH]"��Ò5J�D��T����@��/f"qUk�s~�etEiJo���5�q�$�5ޓ��5��l��/�)�n3B��T�b�Z.�ݗ-&��F:�G�]�Q$#�<�"�\�R�O�㬏lPR������6$�}�QZ�̉<.Vς&u��Q����p����B�-��:��a&��dL�鼊�o'�b5��/!kv�) 6���E�╕�q���[��b�y.�: WOB)��T���TSFK�$�)7�h�Ǒ�%�>�[#�s���n��T%MJW�%%d7���&@":�g���B����x�j窇�R�~@_Oߖ|�
�ָJ9*\���k���K����@��! �1ֲs-b�F�����^���ͷ/�Z�^����1i�M�W6�n7��]�j�9j���4Rį�)���:B���Uu���<e'��[O���,����Aէ0��9?S)#��`J���co��;�l�5�2#��01~/��H
R��ۚk�
Zd
�SI�Q`fp���Q!���W��)\!'�w1k�̈�~p�k��V\l��pX˪��dC�x+4U�������c=�}�O���B�?�
�Yc�UŜY	HFa��ٗ����x�N��| �����r�����G��vz|tӔi�^Q�����	����/��V��0�4
	��H��'L��ϓGhh�����"S�S�d��5��i����b���\��D�>�S�� �D��9���vN�����s�H�K��h;Ap[��1��� !W9~���>�F�?X� �rj��(�;%[�h�bD83��$Ќ���}[���6�%���ގ�{���U籅و�ܞ���.~����[+��T����J�q.~��Z^���$p�b����J�r��壣�V�M,0�z��h��
��{���󠑯��[#}�-�W+"d2��I��
S\��q�D��Y~F�4 � �r�d���CM�v�=f9��N]�qmo8y��ǂ]ChHr�B�g�q	V,Q_Tq#W��(T��K���[E������L���o�����W`w%�ޗ�#�����Q,<A�0��8XC*��Z�h3��� s�\M=��C��ut����y�;�BS��Vpe��w�W�ӗ��
�Fc�m�#�����������)�,�ǷixH�|�r�����Ҳ�2�W���j�d)�@��j�.ިgY^~2P�&�]X-q��Gp�l�t$�"��@���!DF�Z�T�z6\G��e喩���dI _��EM�;Xt���u%4PXu<���fϒIp��f>�9<����z\��"Ǯ&��M��A��Ղ��*�T~r���A_|�U��m!0��<L��9�WڅӠ����(Ƀ��Ji�U;wnPD�~����G����r���~�?��G��YԜ@{�6�4bO������EK�lC��ຕ+^���h�d��?�X.B�c�o�_H�x��Zf��*�g
���.��=�ѧ⥴�Ԟ`�?7$B��Q�p�2�M�{�r�V�'�5�v�V"B�K���/���6�f�K� �_Nȱ=]�����7�޷��F�jYR�>7-��1���}oU�����D��A�>#yI����E>�
C��T����N�g��Z�;���Cz:T)-�+0�D>3ך�54��pO�e���W���H��uZ�S�VL]���$AI�Hءv s6ז�
��h��՟JA��{�罃��������7RUS�:|�n���HH��`Cs�@�]ޯ�eD�V�T͚���H˛5b��:Ueȍ�7d��׵�f�����Y���R�7Kap?b�Q�8��Ž�"n ��Y�[T�UBY$���X �ϯ�hS\L&؊cC�o\4x$(m�}#�k�4��E�9D����y=j�=�4_*圴&�O��U���σ���Oz�,�DʗR�6������[�::�!�'t4���W\$�6q������;\�������{�Iw��T�nPz��$�z�[�'a�%M�R"�8߾����� � �fу{O��9��X�ҥ�pB��,��łR	�̞ě,a�,[�n�1lt����ck0��m{���S*�%�7η{�V���Sx�q�7���kE+@����xܔ�3�o�)V�I�L�����Ey��EMn��]n�!7��(}��t�[�)�&,^f�oG�EK"��{L�Vg��U"t�L%X�h-&^��\;0+燏ԣAlh�CK�W��>�����u��B���6��1��K�J{��s|�����W�=�KC�-K�`��m����8e
9�6���F���e4��L��8{7�C9�wR�Ӿ:�w��m\]��gv7�X�"�����Ժ΢�	���D�ϖe|m�F�v� ɔ�����Pc�U2De��3�u�\�@�m��X����o�O����k��'�`�)bIܥ����o��ce�p^��=��� ��39�VJ˻�ǨX#[�>��{k~X�輛�A�v���4�0����9�K��nZ�(���p![���E�?�����2t`":�5����o��`�v� U�և�	��E���\��� �T�%4:u.zL�d[~g��S�U�q)�%��������e��T�נe|Z��}���/h�ڏܱ;�I����C1{�@�v�p}�b�O�mya�C�L��>�u���{|��6�"�'�@��Ȇ�z��=��* ���ƯQ|�n%���*�b���8��p�>|�ڭw!�F�:����P��Wޑ�<H����☝��?s�,6�9x5�o�����_�����s�R��i�Y ����딁�	÷��Z�;��fAD�d���Yq>�bD�Cȯ�#|-A@Q�х���,`m���V�*^�(���Yӥ��� xB|I,�;a\,p䰻^�l	�_'�^��k���g������:(�Cn�-1@�h@��	P�h��+�$5���y��~���'�"�tz���ęIQ�c@$��nW�?/4eI�P `�����͢t�+VW���|+��ʢ�,�9^�˺��u����iīY�t:�/a`_u::]z7A	�,�0����:��AK��>�
�!�D+M�:Q�=[�jx�ᨽ�ԇ �2u^G��������zőP�4qZQ>���u�Z�ID(�Qu�����xL��m��id� !)��D&�r�dw��l���z��Gb�����P	��a��}䖤�G%�I��JXW�$qB �,�pG�E��o�H�P�#J�#X8N���
�2��D��Z�#k,��J���_��C�'��iMߗ��8�Se���`�Бd�vo��)9�<}�Cu���W�Q�%�_�Y���-{\.�o��$O�?>]	�K�],O�":z�tK+������iWJ��p�y���ʟa���?��r��-E���K�X~2}]��2)z�*�®��"F}Sɱ/��g����/�x� fcػ8�OeC�}�j��G�=�"�0=|�Pbӡ^��]�qP����׍cL�7���>j{�p|cŋ���А�(3�� �m:���'��ѯ�$Ta��W�$
�
���MR�*�&]��9
��w~��H��5�w�3=5���2H\�$'E����<�{��
�WI�{���h��H\)��[��
L��H�������%V���ՙi�Eo�B����������4B��)�x*b��>҆��_�� ?իKB��췭d`�>�*;h��۴��G1�A �T��C�y���*���@� ��{>!E�����"�ॊfV�	�\\�ɚ*�z�� t�"8J�T�����4����빥�fC%�-6�֔,�����*#OS0c�sx�޲wĞb�f��W�5}�%��rt���	7q�C������l��om��gFǬ�C�%�Z�@N�Z�)~�q��/�R�f��{0�ԞP���B������R��@'{*�U��W=��}<Ѝ���k�vw-�����ϙ�Y�=*�z��'SEw�~�t���@�9�X�44l.��V��R�6O���w�
�~ X�j �ި��g@e
n}m���t��8��2��L�tSҊ�bs�R�X��|���
2CRl��{��?��$�0�@�ք�k��S�@���6Cwq����N�V�F�>��O1}���[�.�d ��~Q ��4b���}�O��G�TJ>��B��|ʢ��M�w�9�pXO���~ڬMa�`�薔���QkI����
Y_�D�BItF��$Io�1Y1��ZK-Γ����=���C�z���Vb�]�hT
�y��2�v�R9�"���;0(�T$ws�U*�
n4�R��J�=+��Λ������٭N��]BC���^��R��p�?��G��u��	�5�\�u��1:X����}�s���e:��K�A�������3�>���� q-{�D?{���t���A׊��~J]uHˍ����VMO$3rxX烈�w����Or(��sm;��������=�ϫ*�Zcf ��c�t�r�ը85�l6���b>z=��mp�����3�����w�K��@˽Ac���<�qx�CP����\�Њ�x���?�`�m�	f�$y���}�%ԗ����Ore�Փ&,���!��H�dMn6�F��P������J� �[3ТS�e����%%���}�� =|o��z7���;�������ؼ�Ǻd�Fwp�k�����U��o��f�����[z�YJA�D����S��:���T�L���o��\����%�1?BU �̮��Yd�r�������+���i�cp�9[e7��˷���'c���U��	M
�?�Se|B2L�7�e#xv$D�� Nkhx����M&��=�9ey$�V��OFV�!�Wb��M��Ɨ�P�Ԕ0,+�ʟ4:�u��		j]��c�x������6���2CP�ͣV�)�LK�n.'����`!��eM4���<J:6���H[.ri�zQ+�[�$�+����')Ec�}I��3���h����7��њ��B�e䪦e��HK����v��u��}� ���V��'Z���������F���0!2�ل������>u����Y!�y+��QV��r��}!]��kp�	^?ȗL?c���uc.�OݪlR9�ŏcL2�络+��n�Fb,O�w8L�]��؆c�E���?����2/�"�L���d�?�{������`G�,��>E�
��!���&z�_e`$M����T�a�sāb��Hsw����Y9�4�+���x�E	��*�n2U+#�W=Q�/Vb�$����ږnB��64�t=_�p�R.��*�[mE��>O�+���D��k$�f �_�!�ϙ����7�Ú�ȇ��+ʀ�%m����]0���d2����{�Lx%�9�礙xk�
�a��i8ۡ�$m��˨�O(�e5�+u�]��},�a^�ò�(Mcm5��"x�'���;�U� _������Ʊ,��&��%W�	1�9�������`HV�L���7��=^0R/��ͣm��U�-�i�`�]Q��8.s����D\��r�e���r��bw	̍�Է����z8��s�Aj�
���d��r��v���=M���<!hL�r+y���?���{΋��Xʚ֞��F�NJX��B��;�#<t��B6_pzY!�yM��
2��W��hs�J�2��Ed�>�a:�@G
�q�ɀ}��>&�wD��=��#���fe��pS*���7?���	$��
j8!�a��KuG�z�5W!'��G�� 6�^��J�a:u�P���T#6Y���vtŕެm�1p`�'d7Z5��h�5������͚�$ʳ����s��pv���%�"�K����e��_��t�і:�q����H�qWb�h6�ezE�8òY�sɬEġ�l[0˿N��#03=���� ��`k���.b��%L���)��&�e:�D�	M��HmAEj�7HΎ:��,�N�q]��e,�rA�H&	wh�ɵ��?�3��6�MOalF��4U��>
��s���� �.��~�T�у�?�ጰ��w%�����S�IZ 4��XV8or�p�$���Z�)&�210�rK��jd� �%���$���'��/8g���(K���`k3{�P�n ��T���tRp�D����T6��6�0�1 a���[,A���m�N��Y�.�̈́J�P$��&ʧ5���.zs�յ�>�"�Ӂ����y�P맫!�'�~�A�΃���؜��%_

f�z���uM�2iqP�p�e��l�Uf~E��{@6�S��]����@�M�ph6���zq2\w�t�9!X
��ȩ���|����Wl�5�z�n4�%��`J�S[��
�g�<���=�Y�}��]*�[~Iy�uL�ZC�n��_���DuJQL���
��Կ1-#�n	шx��l
C�B	
l������$�r4��@���:||Uk���������YZ1{���O���m���N>�jw�F�A�XV�B��1{"��ϋ{J'f'��]\qt��羊���g!2]�AN���緻���f%nM�Mg�Y�fS�ʖ�㰳-P~��fڜ����<��F?�L������N�tᏓ��6��3��Hˤ��6�2��^��Y�۾Bɤ�q� �Ӳ�� y�NǦ2����X��{�h�����i���$_�6OIR�l�Q��@8�f^xGw	��wc��Y�y�K����\��~F�7��o�؜㬥Z|��L�@�8yI>�c�O�hD�f��b4�#M��Ʈ�T}
�Č�b��*FF�wEYm��z8w�{FF���ē�fs��p����.������(g8~V�2p�1s��Ch�;-����8�c��SI:q�]��A�����X=IT����-��Q	0m���N���(�"~���m�a����Z�e�9X�УI�@�B��2#�y$�r��LK� Zi%�oO'��Q0���E���5��~��-Sߊ�b����U<[�[[�r��Zg���1V���u�yÓZq:X+��3%��OC�ӥ��?�h�����a�~}�X`�❥�5�{��ZW�JG�A�����B��l�����ݘ�g&�m>�.�.��I�9��ᘏ'��f�Q`^�r�^w�����$�ܢ:���7����I-�f�Ȋ�ŏ����yfΩjܝ�j^�eh�x�!U�W��u��/p���6�.st�)����^y�lH$A/�:u��4�h�Djhp_�Z��?d]��$�@nO])�4�DI���.�����a��A�갧�2�lw��0ְA��9cͼ3	�f��ٴ���{7`E��"�\�Tm(��p���bn�^No���f�i_1�R�H+�/-x�$uH�l:5��խ�i]���?�2���Q1HbȬ����&����0��+�������.�3H�����H;�S�{�z��	��B�%4H�#}q��_��k�z�ln]��Q��Â_�YrĩP��d�G���n��l���!��`4=�?�q^U��y�݄�k-P���`� ��֞�J�~!a�$-�"^{�[��:��Y��V��B�(��셙�k�����3�ÁX��N����2�s�*Қȫj���!�i�38z'�k�P�πc]��-m0[������f���<�S�t���P�e w��W�������!wD8��\�@&&x]�D��^x%��.<s�|ˤ����=,�D�8�K�F�_k?�}t�m�0'�~*=u�>�4��t�;�ai�7n�4�(�b�=���v�
�^�M�\1}�����Ւc�������x����c+�:�{�����}y`�+��n?�~\ǜ�1�����WSL�_��[ЄG�A~�?l\p%EʹU�Z�[j[6$�՝��m`a!�f����D�-*^�B6I�P�{d���>�_� �h?&!�����Z���'��k� .�t�,�Ow}Mo��j���I���O	_� T`T� ����`@�D��iR����A��3�[�wَ�p��~ѡhH�g=��%D�S��mk���ܝ�W�eei%U�65�l%&��5�܀?5[�8/j�[(];p:�(��;q!h������}������G�dAC}zT�'oF�t?T�����Q�-�zH׵����'a��tq0��?q�w>;���J��K4�����s>	%�ѱ��U���`X�Zn�\���8"�1�`?��I����������r�Bvb���z�8��[�io��W��,m(G��m�*m掱����߶C��=��n�i�ӮE���̧���V�AJC򀸮�|��U������������C�4pބ����|O�%����Q/#�V�5\>F���Ψ(j���,F�<z���: ߼� w��
� ��rA]Ǹ~5n��^,_��n# 
�?8Y4@�qi�|��a�.�[w$�>���&�.O��n̺Q����z���NL%��c#(*@�B#�~sigb��MH*"Ĭ~�{�_kguY�b��]%]<^usUO�8Q}�]�g���Ѯ�1���3�n���K ��D�|�k|�|k� �)h��,w��?�������|`l��N�C�����f�D<�KQ�D���Dvt4k��#i[���š=Xi�йL��GS 9�WL��I�ˮ���
Np��*��
i�E�/4Z��S�l�fN|����J��H������N���i�Q_���hO}n�*�ف~���^���qǷ��
x����9�y�)+$�7��"d1:6XC�S���K�	���D����S�4L�]ź�qy������h��)���lJ�mi�k��������R	B����K�ɼ+���~�WN*�/*ׇ�ts4��h�)��h�sU�:���W��;�;Q=Mv��ǆ��=��]�pm��x���	��J�8O�D�h濤�[��!�Ǉǳ����*�������̗>��1 xL�<$�X����g�N�`���bg�ZvM�[��ۮꘐ�dz�;����q�ݎ�̰C٫�}�ֱ��KZڞ�}�a�������L��E��d����� I�c|�$�q�"�
y*��A]-����%%����\I����~�pQU�Q}�3q{�"9��	�� ��H.RO���\,G^B��t,#)q��Њ� &�Y�.�"�Eăz�Ih!?jEa�[�(eͼ�C���Iǫ����Li�d����
_��M��'�� �͈�u���$X�_�#[�u�&���5*�R`��ʰ,������w�ߪe�ݶ���9����{����n�����lN��<30Ҹ�C96�m�$≭\o��A*T&�k FXC;#F�������si0#��1 (����o�|�#�x?��-�M����eMU��q2BL.�#+� �?4�'!��\���g��8�Y�Dt�*X�r����;i&�-�#pa�F�2�.���H}��d,Bi�����Dz�ί��L^G��MrY�1B��e1�^��� �(d��Q�`�V.�&
ǶN@�ͳJ��J��'CTI
1�'�XH�����4�{��[9��m���K}�Y��u��[��Eh5��B/ڷ�3��ά�5�q���O$�*�3x; !y��dH{h��<JG7ܱ'1O�9��\�����hT4�C|L%j'v�����/���'�A�2a�YjOՎԐ����Ź��d{���Ŝ��B'ՙ�������ͺW���kp�Q��GÂT`��7��~�܎/���}�v��}K[5�9�$�A��۶{�.P̣ON�G��9U������w��	��9'5w�r�4y�s�e�d^�'qr���bk$�]�4B5�E{��5�����S�h㷧U�I7�������&<焂�1��4���������,1�WjY�N������ܺ>�]�5
o�i�UV�GΕ�+�w��qY�&C�&�/wt���ۅ��_68�D�ڸ�y]t8�%_6A�����ͅ�ú��^g.ѢO��40�K�h�T$���k����Kr�qfh�]��<�z�Q�
���Nֹ#3���{b΃��00W�t��st����;	�#\B�X��)-�5��_]��wj��D�!�����J#EMM4�H}k҈�~"��G��+�`�K*	L����(*%�\5��3�=�L#a��*�C�p�.}�{'�;$� dx�#��Ȓ�Х��{9�j�(��������.\�8��.���D�x�P0#�6��<��3�u�Q�͈&��6��>��`׈�
���^��曎�u�+��??�eȆG��[E� %b58�۲����t�~�.;����l�W�I����*C���r�~)�,{k�b��2��	���;-��Љ�����M��9��/�8��(3_&\
���4�p�FeNfu0p��MC���a��	�;�|'3�h�V��w�Ө.m���gc��/p�3���e󾑠�s��?�M/�=�I�g <(g�� ���k��`Uu�!1��O��,�mD�Z�+f����KV[�}�8yK���a���o�t�0����J�'+ʂ�%��T��C^m�������<`Q��e�pY�e_A��	��c���[�
��h��U��S�c�3���3�EyS��|�����c�"~x̝��~��q,es<����ȇ[�K@L�Z�@Ek��^�TTzhGځ������*���
1[/�:�e�^0��ݑ�/�����V�`[�3������ܣ9E�����aZ]c�b���`ۏ:I ��/���'�u��}��b��J���@�O��؋�eD��5�V�ٰ'��CÛMG���/�a*�+���U�	8F?���\,����x�A��!�H�&����M�A��?� `(�J�L��ǜ���\tv()�um<Uy� 7��>��jz=2�pR�ܐ?����ඃ��j]<Ag�6�J���_?�%I�@��z0����k�8i��(���I�-��D�R�H23g2q��@�J����$�£�+]�g�LݼB׵͡3)�eOm�r��`��xm�:�#(���|�~�}�R�̊�u�%��]9b��d���x�{�$��zqi��0�z~� V�#�B�BeJ��Ѩ1(e���y�9����/&g�J���2w�>Y�n-`�\�ev?EwH��1zL�s��5Eʜ�@_�E��ic4�ٚ�s������%0D��@��4�'
�s��T�C���c�ޑ�P�מ�&�����R���t��Ox#��D�zk0�kL� ���ч�>r����C3�t�Ix>�hN�<WKu�۶��+�j?��@�t��"غ5̸�Y��Mq�L�4p��T�fb�k�V�){m���6�߃�~F�樀z�u�gx K�)"�H4�
M�.�f�ʆ�/�1P{�:�� ���{@tK��Cv����f�b��K�tn���C.}�S79��E�w;��^��T���U�<��WP��Yx8v�ا{j!�"7a�m9P�x�u0r��m�R�ض�ӏ('U
�uN����.ф�^0�Li\��a��l9�@���ЎфA?�URw@�-�0����C�H�>S&��g|�9��`�=�sJx!����c��*� 4p�5��g�x'��׻������M2Fd�y�&W�$�2NAmm̛6�ƫ+ @��H0���M��*a�zL��'��U�U�i�mCĚ?��,��bM&����#,6@�R�񀰥�n��ńc���h��N^��``��3�n}b�U�35��D�o�J����K�F8���x=Hda�/w��e���ǰ|Lol�9�@�^��h�G�=y0�-��ui�&l�࣎�
��@S��� J�x{ gY���m7�t>�~ȹ�9��j��+vEξ�5�
��!�|cps~��ӓ�鏵a��@�u�p����8�ﴬ��t�ӯ���t�Z�%���=�{=��`�����uE-�
���S��MU��d[~3l7Z3�6����%�#�����f?����$T��3���YxI���۶yki�#'L����EK������o�P1���w9�l<O�q����K��;s@266� AB�{;JN�q_|��c��J�ʠ��*yX5Z��^�ʄ��83N�v8�ÛK=�N~�L�v"L��j1W��F�{�W��Jy�m)��.e�L�[e�1� �!�߻��F�yYHf�_*��0�c��+tivy�ۿG爆MOa	�cl��� ���y���v����(S)��11�O��	��d�(�@7"\	�W���
���#��A���������.�S�fέQ���b�v�8��v�'�E����`��ׇ*Pxϣ�@���"P��;_�+VZivZQ�r�C�#Ux��M��#���+�\���c]��?���f\uϙ�-��*�,!PJ��U�wQ ϓ���ؘy��E�'^�\� ����-n��/k�c�n'f���~D)�d�+*�R�w�D�r@(��*�Z��ؑl�ԗc>���EQe��7�}f�i�+��fJ�[ G�W�Ɍ{.W��Y���1�(���$IbK�7��D]F4�m=���_��A� ���^�T`Xy궐y��;�v�#V��'�h�±��ދq����_>�q%bnRa�:�a0J	��_e{��.ۡע|vH&�I��. yy:�����&iWID�א|�S��]��p���p����)�I`�'�� u�J;�W̹Vg]x�CT?�\77}#|A"�֛CObf�[�]������=F˱�-�i��g:x�����Zxڅ��xt|���~q�
�!��94���+��-�B�b�i�;A�I]���+��Z�v��f;����Y��1�x�&�Y��a&wU���Nt��\�z@-��q���0�Bp���]��u��Bm(�������E8DɂF^�U�ӓ���?�J�T���I��l��~����RR����C_%ד�2�32�c(����#L��y���?��^��L'RRU���$4R"��#���&���g���r����U��M�N��'k�y�1eb�-3�*EMs�~�hP��J瘕����0�BI"�D
����o=4Jc2]!2��aʟ��v�ɐ����遤6������YU\gz�����~���Z7���+�Ɉ/&�.\�J��-�3���o#t�@t��Z�-��D(�1kbA�!�BqNGơ���X<��=�}�x��h��δ����	-���"�DՎ�h=�;�iBI�{H��`^�/�,��]�
��_��!ą�F�c���u����0�bx'�^�o���h��0��G[�_��O��О:��X��"
���U^�㓕���"Ttl�K.��m�dgQAM�1���.� 	����Č��N��r���7���K`�a��O�R���*��O/�Ü�2�z��-��MХ����(���4ff�Z1�1p3\��j���;F��B�]kc��li��Ale�������ө�Y�{vU�=7�����>�6赇�vZ���w�vh��
�4��ͨ���x�́�l��ڴ���=�)��>�y�͗����O��V���g�ǽ�����>/̽6Ф�|����U)[�*p4=���A�mU�<ј'���ώkT�L����Pm��:+�&��n�:�W�l�ew���U�e��>���0�����7�d���5��|v0�:�����FW�>P���w�H�A��WW4�`1��q��4�ݼ�y1����%�10%��w��w:,�ʂ捑��C�s��ȩ!�i��Ҽ{C�����a5⎰�0������r9��#b^B��O��@��l��;��E}~�ob�=���U�Y͏�C�Ƅ�-�f9^�3��,D8\�-MM��~ŧ�w��ήx��#�[�޼sA��CEn��T,�Q�{a��
�a�> /Oأ�
��=�Du:��p� x��S1>��F�	�/=*�����ǝ�2�ȕ��{��"���}�$� qs�܊�^�2�yU0B���!��o:��v��E��<O��:#����N^�4�������"�gǨ�2Xo���EY2��o�s�rP�u�آD���^񛆞RߍRF�}Є���ȏ�W	� ����A_:dE���9�]/��@��i�!,m�+9b0���g��=d���8Ӽ-	�>���M!���|��I\�t�\Ij'%��OH|�1q��qj�n�V�-P#���u�댌rW��A���T���K.hnH��P~��3��B�!�t�4j޵*������0+�J�0w��t��f z�o�&ǆ5<��*��maJY7��e��wj�:�����g(<@��u�X��d<=�hu4����&��-�,B�ʻG�!���o�~��4y�dAڑs�Gfm3��/�������?0ւq��fpR��6 ����>a!^G�Etol�R�����e�03��Rkk���*��z�.k0koޱ��L0-T�՚���>�1M�Q�n��6�d<���/����<[A��������M���DOA8���4�NpA/սJ�tH#�}on.��;g4ܯ�.f�W��.�d p��5�b�~ G~"ة�]+�� 0$l8���
JI2�=9E�U3��s���κ׫�h�X�t!����Օ�j�`L_a�{�C�<W���M��e�+Ρ�j�w��?u�ѹfnʍ<��N����k���Et����?R(j[�7kL����)L:)Om�^��ej�{0�D�����;{�=uH6��/A -�X,�l�4�N�O��/rL|-w����r��\�W�e
Fue
��$b�A�4t�ug�q���u��  o;n�ovSFm`���3]HC0���#_�"�r���)��T��UwN�I�R8Z`���0�s�y��&l�Y�6��0(��p��vcV�K��w��:�E���2�ܵ�lh�]����9i�K��F!�Nz�O���.He��X��B�S��5�"�_�<�e�^0�R1��E-���b�Iv��N�``o�G���8��������:�m�26�c��9��Ċ x�U��D����m� �$��(��l
��AqQZ���B:�=���u|X!�R�+O\c��݂����ʥ[�8�S�et
����V�+���e>�aǸ^��߾h�3�3�=���i4��ny���Ò[龢�=�Mgw���y��?-Ye����)T ���M�<e࿙�I��B0Tigt��E�@,pIsb����N
Hf�L���Fjْ�9��xT�H��o��<���gP��$µ�����$:Ռi8_�:鐽,;�'�ߚ�D�
2�PId�	��H�	�ݑM؇M��������cp_tȬ��@�8��nE��l�������p�|��][>j�4͝�BY��(G-<�RB�eK�	u�6���y��*�ǹH��L���V��r2�&,]�pVz���T�QڢZJ 83q�녵c�g�[��'�(�'��6�z��D�O�mPô�t:k�|位�Ó�>�	�� (І�`�M#M��zc��}���7��9:.����zc����!�}���'�,�~�&ז�Y�^��pz�����~]���`	��?xI���d�a�1�jE ��X"iR8^Y"���/;�"pU����KK�l($��?���&�>�\��x7[�_t��v���|�����*���G/C_�<x�!7��Y^TN�0��?��҈\r��&��n>����)�����k赆Ӕ{j��L���Q��o(�0��ZByۦ��W
�dt�
�G�Z�(�u"/�xG��y�9�)c�
d7De<��*e�7M
�"L�����A� �?S���s�"�n���u�ȑ`{,Θ	�q��[���(�O�\8�G��)����E�5���7�+q��Ϩ����7m��X7<E�:�^��&�O?�c�Y��?��Y4,���kȷZ}�� �����@�y�#o���r�&í�hē��^�s�y�qD�@�W�Q����g:���W�RW'1��L-%�>���t=i� �y��_���ʌ|��qɋYsX��IFCTʜ�%�Z0:��Rg���r2N!�bf��z��C7�$�}Ew/����(�g�?�8~a9�tgy�Ԏ��|6���w��ަtゕuG��M��4	L�F��o�$��aZ]\�����P�j�u��ћo�,��E���[�n0�$�'1��bw�:�d������ 8x�#Aѯ��� �{S����v��b��#��Ir;�D�o!�%4G"=>�'Ǩ��z��j7G��"��u��e�L+������M��B�Y�"t>�'�k�@�Jo�ad�Q�����A�ԭI��]��M��J��?��O��Ƹ�ȳ)����܂5�5��ދ��U�ػ���)���J@�%��-������~��̿�9�47��>��Ir9��U��;vҥ?�= 2�>ƿ��72>��V�`mՀ�Fl1�A�V��P��cQ��S� &c�m��4��#�L�U��M���͛�����7J���c(� И���֋<F�M��ڕx
���S��./��vE}:�S¾]B���n��kU����`�0�G���F��s���`�#�2�9m�f����UY!0:`�oy$ȩm��Xd�"#�Y����3��n����-kn	{3��M����O�4�v�xN��ֹ�8.��WK�3@?
�����2�V>�3�	�ب|��4rx���ƔTE}�ky��}'ƈ������9q�'�1�S�֮ƫ�ZQ7=����+⼼�!`t��(&���j��$X��O�2��@w5X0�(m��ם�,�fC��J��DΉ'\r���!�uc���6�<Z`x���݃H휦+�D�V�2'��]5�����:�[��1�@/j{�7�/봼92���������ܚR�d8�&����g$�ֳ-o��p|:��P�  �Ց�Φ�k�g�7z�RK���yj���� �ƿ���?���6OB|@a(���~f*y��yЫ�'�������@�ڈ���Tj����:م;��j%g��m��g��>�7j7@|s�0�0O��zlH��F�tX�<tn>c&�*��J�Aͷʪ�c1���m�x�*5��&�j������qH�M�a	�I��� s�ٛ[�.
��ﾭ��ߴ�΋c��QU)^���"#h�C��[ߧThd�f,t �f�jS]CR"�$J Ю�Ff�`��s�S�"A\\V�H���|ʑh�2�B�am'=��,��F��l�.��R���r�bd�tp�%�1q!�0����B�L'Z���~���ٍ�^��*�R��(6���c�%ϟ�hޒM����h�4�iB�?��Q�Z����GB/\��}G"� "�䬝;�m&�5�{T�C+��<�#R1b�>�3��[�ȫlq�#= �-�szu�������������,�v��K�	��)y�[YL'i�6��4�!CQ��~�q!��M̙e�-)ِ�Iul�q�mݚF=2��5�!�ٞ��g$����ٽ�Y=0j|y�s�,�)r�=�U��To(���x}�۩HWJ��/O@*��Y������u�yj�(3j�C��u���p�ϻ[s,�|���=(M/[Z���*�*�T��Γk�j�2����!?+��9>tw�¡P�i�XV�ˬy��qO[֬t�E�!�`B=I/��@�w#�昳xQ���-�$����7������]\Ա�\t��FitU��M$7��6�d@��:���P�������@��7Z�J*�T�Ý��Y�Dj�UR��zL(�=Ȫ0zvl!z^����Nr9J�&�+��-�m�l5��m
`�[��i L|���d��7#��Vc�V��:�ilF� �ŏfX�E틶$~l2�Չ���o[�l27�|J�fme�9�"x������燧�ˌ6�%q��#��+[�nl���`����җM�98Y��]m"29G3���
f+�®������ �V���S�ޞ����d����{HD��1c6[�w��K��~�W�2쿋&d���M6{����*(7c֋RӃi�#�����6�B"��))�G�`)</'�>��L��a�Y%w���m�f�H�G�l�����$^S$�LO�4g^�bx2c>c���Di��/$�5����s5i8@5$�_	�|%�sg0��{0�9��UP�L���ay� -����P@���ۮ�������p�ο�ӝ${zv/�}��0�����"�;B|�{���Z����"z�ԠR���f�E��8!2f��js����������bF�p��G��sZS�p'�e �\�Mc���7� u=Ga�:*�Y�%��}i@5C�n�F��6�O�2C�%�ﯦ���u�M΍���!ϧp��)	4��}���:���:$�9�Ũ�ճf=5O�ڲ�=1�t͝�ڒ�q�~�j�A
�SB!�%���)�5N6?�����+J��Mܞ���X6I����&��d��K#skN0�p����;�q��<��ϐ�י��B�\x#��^RBǪ��ؑ1��?D��A���k����|g���(Q�j���� �\��f��59��☷jH��@�h�E0Lg嵣.��)#�c�wd8򤾙��w@S�}�|���W��`bw� G�L��Q-8��2��(�6z�G$E�%I]�ֺ{7�f��p�GG'��m#1��C����Bg��ʉ^ɤ��{BV��!�brj��ڣ+0pF)��L�O�5܏�`t��v2>���� Xy�����f��cDvV�!�V�Owf��Ej����~�q�G$�Z�FxW�-�_��~�DL/Fdt����a�ͮ"\V�w���� ���v�o۴�(�PX��h�x� z�K�<G�Ɩ��v�j�勳w
�Z`�d�]c�^놅2-�1H,��.����l��)8{Jr��S�"�"��B�,ᎩfW�*#2U����}���h�'���iF~_��Z��Em�������'a���;�z�J�59�	��`���L�P$��VTW�`�dןz�+��Ca����g���av<�qw�+r��%�֚����#�1��@d9��hd�U[��*�Pɑ���-q�6%�C*o=?ۄL��p��B�`�OUk��	:'C�v�i,��A����k`Έ5Op6-eD��a��b��de	���ǋ��Md<㷫����n>�S�~"�v�j��3�cS��K	�eg���{ɐsВ8KX[�@��ݒ�2�tʲP�^v�v�b�v���Ŗ�0}IsA��_���]<A���HA�R��P�'6)���(�y�M-�9��'�]���U�Q&3�	)��jy�_|���z�?�=��ß�K��<��^Q�پo*�$h��P�[vs�~/������4�]O��պ����eK�����a�u�b�L�&����~�F�Q��<��8@�a�<��ϕ2RCU�r?��0�-��D�c9��-�{x	&��GJ�>���<)j&:]�s ��9��3��»�x����*�}���~6�Gi.����5;m�V�逫 ڜh�+4������j��\RZHi�^����Ҭ�Jm���yFp��)�\�8%E��(0�y��v�~.��m��/��)2�68�A��F� 3����	�:�CS �wNҾ�D��̿��Yكa
�D��`\S����6&�5�'iBE!;	���"m\���f���Q�[����5��F? q��������3?���O�\%�$����ߩ"˒��o����zDx�
����Z:�(��V8X�P�r8e�,���0�q(����I�~���n�n��LO`aK�M���<qڙ`*��<I|ڑ�Ǫ�Uf��=֏z�ݾ5�O��JkY!*L,ڑ�i�V�����@��׈����?�88sƀ�|~���%����]r�H3�pm�w�SZ�̈́@S?��^�P�s�X)z7�
b���is�q��8�����\�xi��^�7g�(���*��:7�2 ��g�`�55�^�s:*`c+���Ik��Wa*d0�1�8���>R�R�����đwW}��ZHO�[7��Y�v:�������Z���Ny\�-���v�6��A-���ˮ��w�	���J�Y�R���/k�""8$��(�:@
0#_�[7Y��(�D� �Kx1M�&�Y&����n�)��;G�|}b�{q(|����@���<�_�C@�R�6���B���8�,I���C>�^�I]3R(K8+�U��렊��αb��H������>���M|�X�Y�WF��O�F�wS���v �в�p2TF���e�vV�et���yd����f�MW�3ߘ�|m�u��� � ���D})1D�����W�n]j�G�J�Ѽ�&���t� �./S��P�ٞ�59� z��rό.� ����j@�#��Ǣ�a�����9�H�NA��$�6g�A�c������ĝ��Twǟ��쉣��%{P�]͛�ǢH�q5[<0��$�&1���Ti(t^#IY�G���<7�RR���G)M]��t�w�'R���úN���"����gA�Ɨ�H�)��v�e=�Uتz �+#��W��}3�no;:�,��I��&�Y1�w�/�>:9���v��{vZM�;���XPGR=�&Ϛ����B�߿�{�zw<�X���b~�X����$>���[t�z%�6BźW�����C���)��<�v�i�s\4M�([�g���󅜞JJ~A��B��ћ͎���a1o��`�
]lg�ҙswT9��fa��(\l��=�-�pJ%��_��G������s�{���DEg�sCm�������^���gz�I�!Wii����ۉ�;�v�+/;�⁊��A��ɽC�}���$�UdS���\g���Q��>��mM�tbgj1�_���ԜvÍ?$�B�4����M !�Z��ߘ����Ф?�aU���w^���zHA������������qA��\�!��$lƚ����	䤒�HFpQliq�?B�sg�ieӥ�et�C����dH��M�b|Z�\�\V�_-˨�Xy�.���k&`�w�+��8�OC<@��L�T��BM禗�39�=�7�0��)::��b02���5��;�|�	�;���nf�"��R;�CI�!G��m��կ��H�r%y��J'�J<AO����;=��r���Σ���.�m#����r���+o�r��#v�{��9$Ɂ�ݡ�#��Y�oz���ٮF�˥U�G/xT��=�տ��������I����@�k�� ��l0r��&8�[qE#���~8�D�N��6���.t6�gzݔ@h� ]��Q*�TB���k)����4����m(qG���XkŲ� �v��nDj6�4H ������a���8�N*�����x�Z�������(���ؤ*���]��'��d�w���BqB�Ȣ}�-��OKPCįB��_� �Bw��'&�c!O[Vl ̚��ׂ�ߗ�a�kb��^�`d��Fy�5�?�RJ���Dxh@�J̆����X ގz����Xl94��_G,t�i��h�O�[Ԁ�ƞ}��ZY�0(��j�p �/����D�H���[��g#�{�8g����NҠ���
�U���+-�1>��<�Wj!��:���'YT��h=$��l3P�n��s���g�]�#���M���":t�������f�!�b!be>�|T�s�v���r��\Z:�ᴅ�WD6;{֤ �������
R�*s*��?i4����h����T,��W<�#��N_`�Ta�c�p,��i��$]3�����x��x��2"�P�:`�Y�pk�H x��%�U
6~~�3�Rϭ�d�0�S~�W"��gu�����<�[��/.~ZȨj�����XL'�e]@0�^XeO��|��ZEH�~ �_vA�����c��^ �{��RXf"�������W�S��A��|� ���l�5Q �a`뙏w���o��P�,:�E��:���͖gy�w�ީ�(�H�˧��:�o�N��t�O���@oN(m����5ڮ}�ﯳ���:�&n7a�u��nM��ҿ�S8�`��?�m��X�Kd��WovY�\��܌���k���y�p�H[FKc��A�3�1�g�%J�z�%.�3d����)Q�O���'@)��\���@?�/R�nɚ��|�*���x5��������-ucJm�4T�jS8=bU�>,����n�#y���K����f���࿱�;�+�Wc9���@��E�����,�qt�d(�h�1�.deo��H|N(�����M1��4����<�7b�p��Uv��WJ#X����������w'Ǆv�[W
��W����*ڂ;��mO�0>��@"�n�"�S�����%m̕�E�q��e��9��@��h�{W>��a��$�y�JH=I_���g���W�@6�/��V7�f8��;��a`LЛ\�iQ���@<+PP�M �[�&�
�o�	)�j�T�ʁ�f�s&i�/�v<	��|�6�������U*Rq6�B�yy����� �=�}�V�C����F���,I�I}�����f|�ͧy�I1&�u"f���Q"���],[&_DoF�7*R_]� W�/7��T���W�>�a垑�dGߕ��'��toU��gl��Cuv��Cנ|x��I��[.$p���[�?0�l��������$GUw��=���/Y�qo%S|���c��W=%"��8���K��u�C����NU	n���	���sKRe�1�vHr氎v�;��,}�Q�o�.�^��r!�C�����"Q�������Z�s�4'*��c��&C3ሯW}c$�	+���>�ˏ�� A^�B�;p
�0��O� ���/��n��jv��M��;C���j2����6�T�k���i���� ��)VL[nŀd;�Z�hBU��lϱ#���]ˆ߮�h���!���<	Pq>=PN�yQrELփ`Z��a����o��1��8Y%h�1%�S��C�G�v���@�j����e��a����J��'�Ɖ�&�A�,���8�F����jRe0D)�IW{	�}>P��!�6�R��N'��󁡙w�nn��oq@Se�]w�9%�-}NTgl@zO�Kjԣ�1�K�w(��W8ͪz3%�4�.��n���c��!����nǧ�4���d|��=��枯{&\u�by#�6��]y�:�zΡ��Le��;�	+�Yz5��]��G���*��wz�V���!S�[�����өZ���X��QA�N�����AN�BD����gμs̔�u�~��9�5�	�:`���1�!ن
��Aꭔ`���ʵ�l���q�0]�'"�*�],���՗�7�������QI��74���J\�)�D�<YR���M�`��C"Q$f��(��u�$�/P�q��21D�x����+�?3���_���
�9�����/ۘ噐����f���*��>Ŋ��a��J(q�ZH��J�ay2LJ֖�ll\/F3��rnԾ[�E���箛��S�D���X*T�Y�$X~4�/�9Q�/��Uv��y8��	�*�u-3���0�8��͞�2����ecQ���TTt����i�S}A��uȠ|n��IE���oY��r�-V���T�mS�E�r���[��f ����{U�T�4�-�/1�e�������7�����J��&�@�K.�3iA����᧿G�����2���U�O����<��G��8��hq���w�����a�Q	����7��_29�o�.��pa�n�ގ��,��}�np�G��'�%@���GՏ�vj������RŜ�O����[ЦU��2����9jJ��\qf,��'�����AU���Q�d�W��:��ӂ���2X���#���?
g�-�M�D�p����L= ��`�vW?R����cܠ�f�Z}*"��]x�J�>{�i��`5&����O�HZ��L�m���Id�\�{���0i1�C��w�[���S���Uy_a��dq8yS|��9H�)ٔ�kc-W+��:�L�&].��W���������+0�D�R�e�'f�v�A�?~(��\�� �*����[(>�|o����4����7�U&_~�Ȍq�*F٥��P�q��I����/ox��>B�l=Ю*C&�i�bd��mP?.$�2��g�1��ϒ���)��|~�e�}@������jx�nu�+9�u�/���'�5,�2�P7D���	<�Du��,��� �\��o��su<�j��e+��=8[�aM�,���~d�[B��C���uY�!�nO���Q*����'ȱ�d��!HT�iA��������$d,(�ì��Z1�6��#�߉��d`���G9fևT�#D�(����k�8�ZVY6��1��/�Ӟ3��A��p�^Xs�ZltT�W��ƚA�&���V�Pם�����ci�Tv�����N�ҭ��iЫ��IS�H�ƃ]�!�����ܣi��T$��-��EK 
��NBd}6��#m�"�-�w*0FLTKO�z�A#+�I�w0�*��|Li�Z��]���#�/_%"����*�[�V��)�`^I�u��y�J3G*���
╚�s��xvM�����+�\�0ܱ��}�kk��ɀ��߷-D��O�a�Ӈ�;Q��Z������Ʒ�0r�E��f��+G{Dz��
�����c�Scp��S*}����)�́ӂ$e��;F
��Rْ~����'!`����"[�OV:sg���V��}QfB�EW'`�g2����;��w~3��Kv9=F���M@��Ӷ$@�*4X���-8�#����t2����Ď��s��J|(���6�@���>���>K��E�ph���S���u��'O�ƴ_,t ����?�OE؏��e��la��F�
�]=�6%2����4BWs�l��i}b��Zq{Jz�I�?@	nۤ;ƕ��&_$|�7t������^�k�m�+�?��6dF8�kF]# F�����T���K<�,}���^����<C�����YU,�1�2J[,m�/��jǐ��W��i�=��|���3��8����#�:�4��rH�d��s�j��J/%��}|
��.K6�\�X���L��H���1�wp��<�X�!?Z/�o�Ʊ.�鵭��Z.���M��=�q�x)bp�j�y_��t0}�[�`�����-�\f�ư}Z�d�<�[z�o��oԮ�Ī@�KX���	Y����04�C����#�E�E<��� B{��X/�d�ױR�?�@��)k�go��R�;��9��Bn�����/��@G�'Or����k!������5#r���QgBu���7cSc3�W�=�k�M�)\52K���J��h�,�%��<*ޫ*��="�������7�� <z��<)��-�D�+z��$��>3�~!��@��j~N�0��`Os@������A� .�\�=P�p�<������m*b}��M/?�	�<�pE��M�YH��V�80�#~I��#O�хy�����7�B�
m��OJ��P�ש���[
0���X-Q���!����%�ޖ�I�J~�=藍0�$���ZϦ�V��*�PDS>0Fi�D�#D�@�$T#}��޼J��){�!�a�&�w
�a���Ж�Ё��":�-w��W5Ǔ0}�M�ψ�pe�y�����|��=ϡ�,z��Î4"{Gv��Q9DK٨��\�,&]pKWR��<y�ח-R��.��T�G��ue�������U��td����4�p�%��G��,��{ҒnN��t{]/8Xd�Qcf������uh�X���\�4:=1���Uߺ*��[��qrg�wz~�9|B��.6kx��R�.��x|�_I�g�b���Y�Ĺ�	�Wc��lC0[��>a�D��(��q��	�%�6��{k�f�/�!p��p�e��xj�p��ݡ�qѭɳ�S�BH.=UCRq0Lߊ�N�m�4I�/�h\���>��M����J���s&/[�A4�V���g��.i*0�>�8�4�O{촩+���>�5����kc����_܏�d��2����Z:��4�e�K8�
�3}̇�Wa����΍���KK!ZaQ<샢6��.H�%e�d��,a8�ܠ'Ϳs� ?'-Zn;��MN���֎��Ѱd��<Q��]�Y��R�����̳���v�L�IHV+�D�T'�1��iy���,���^�Bxv4[�Ќ����=�iΦ�������	a���Yq�}�Q%m���s�`�SLl[/�j4~ΕC��)�3�����wdQhk�A,����i�$�I���HjZ�AKUΏpIՌӋ&�5�hs�s��0����)�Ċ�K��Z���M��/�����	s)�����f]��C�5{A���by*�d�YR���}2���!�H�Y��'����ut�`ua���]�PFzw	��]���|�si��DFG2lŪ��u�)� �Ƚ��ڶVP%�C0܍f�����=�����q���K��ݬT4 <�:XZ�i
���?��ĺ� ��Z��=VRfC�;?�  �w��[@˵��k'�"�$<\]�?��Ql��--��O 6�OĞ���,��ߎ�~��M���`z]��E�!�1���5jF1��2 pfإ���k�`�z�V�E �C�G�1D��`�ϊ9Yc+	pi%v� �N�͛�{e�"�Z�y?��-ުɀP ��(�o06�+P˩h�j/3 Ě��(�&@����V2��NI.]�ٔ�ng%;n:YtU���n�a�U?�K���l���UO1�JJ�f��@W~O���-�e�&hE�*G%Y�{�Nm��|`��Q}N߁�7�߮,�RVK:`�qU_�y3Z�f9�Σ[A/y+��@�ti���ͮQW�=l?$�&��B�M+B����1qA6<�}����aa�����@DN;�C��	�,;�|r���H+L�����{�2�,�����|W#��!��Y����!C3k׀�c���Ts�pʃ	����Ĭޝ��s��)�3�7�u�
��h������U�iBԕD�!�!\aQ���P`���^���_^WA}�����E&]AvFRk��@����ۿ�1ǵ�<�v
��X.���`�L�Dr��f4��{���Z�q���k��%}Q"��(r~㰄s.Z ����;�$�ฑ2�Q��O��d�Z���((�aH���N0~�`(��J�+�%�D	0� ��O�������j������@iPl�m�G�rOg��������l}.̩�x9m%�N{x�,/`�4�83�x�ܛz���d��$	���4���6C"}��I�5UAj��0KS�)>��غ�:��k }ڍ�3n�'p7���9��6����|�&��_�Z"s�Px:�xY`�1�:��]F�WШ��	O�
������LC֬Qt-I��w;�g���L�[{ޯ_�`�~AЯ'�4�=��w�,P�B����f�d���y3~;25�	~D5ɓ�Γ���|M.4�l�O�z��{�݌�ۏ��w+�����3Q_��'D] ��%R�q�bL|�����t�Q����F��8�����y�1F�7g�Q�A�kW#�b�ִ� `]g������DvuNB�\<\q��}�D�m����;�	��b�o�$������m��3H�$Xybr��`���T(K�'�::��n�`����%��a �=ج�������Գz�
�I�q�+2�VWg��Dm���)gQy2�_( �D����0�"�v�
s��%Z�/���r2��Z�R�R�#8�����u"�q��>����+�})���|����1�>f�#Ճ?��#�nte����/i�/�5!�бX)8��|y����י*e@Efß���A����&�O2�>�'�릱�u���.��;y�� ��}��'\^Y8����M���)~�[R�������S�uH������P���R����[����0l�A.���5Ć��/L�&EyG43����3|���y8d�i��Ň�]
���q��l�KJ�=.ӑ��e �z7Q���Y�EȠXwʲ�����c�k�6�>ǉB�"^���Ӡ��xs�e[@� +���&R�fV.ľL��&�r�^5(��}|MͿ��w"�j�08'"s�|��e�L�&�<���r����H@�����w�q��6T�B�yϼel��̅��?�L��fr)t}�|��nǄ��	ܮ�i�B3&1��I9���W�Ѐ�&
�Hր�q<�x��$u�Z����[��6jQ>�����ABH�۳J�$���������\P��H�����%?�ev��|@��a��f ������Kq=�W��KZ�xX(^�i�����|VJ8�qfu���a���Zn4�q��j*г����=2(:A��0?� ��B�j�8$iz��D��oS��_�B��9#-�V�o��2�B� rh�w[ܖͩ�evӲA�ZFV�)�8sH�u���FLu�R���JG}�92�W�Jb�^�$1���~b��Y�8�bGbI�<'Ԝ�d(��\U��֪_^Q[k�N;c���@iK�����������şp/����\�N]w\�nZ�~yq��N��p- Q �������~���sDŬ�;h�-��8h@�|��j`��ي���ԉ�,"�3���X�f��}�(��NA����4���Z�H�^�68s=�l0C9ƥ�ց� gv0h�߫p;o�Jo��E?n���O�0H�~�B�$i����i�D́q�nh%�@�θ�稀'JѴZ��솋r����,Э�Rxq�n�]m�R	��_i)T��ϡ����Z� �C����
�P:��*�zq����Y�w��d��娯=���<�e�h^G�i
�ؘZ�*H��;?*� �J�%#'���taS���_�N�ä�I#��`�t���/�_t��&����.�
�)�����������3zCΫmD^�<Γ�5ĭ�"��m�̒f]�	���Q��+��@��<�m	�\R
v=\L�Գ/�򋻺78�#I݁�t��c`���̸R��� ����XR���
]���_�e��5&���`�_&=}ꋆ����E���&�X�u�?43g����(�����FjI$▤gHmDbf�)�z#�5B��R��p�Y3	��Gx�bs�� ,�9#5���.n9�᫁��頬*'r>�-
+��<2��2�N=��t.�U71���G��n�mu1P�NvmK��ӷa�kѿ_�h���4s?��b@�e�~��婢���}�"�a�,Ϡ���0@a��VhhY�v�FB���H"��?��~�+����vu��76*��^]S� �&�<�����+25ۀ��+��<����ZfI�q}� �u�v$HځS`�ϛ�]��갳�r6�^u;��t7����~�{"
X��!y���]'��ۆ�)�mР�����h�ϴD�Y,&@l.ݲ��脤uc概��s4y�5�� ��(x
S!�P5��[�����+�By�)�x��j�x�1�ߓy�v�6��s�-���J	g�W:��1~�C����wu�E�blX��5&����@'���y���2�y���s�;�iV�j�HC)��iin�3Ą�n�LL�@ɼ�J�&�D���!

e�����ږ�]�d��n�c����a?j��9s	�n�[@��/�s�7��`(����?�R���2��0���	y��I����(��!p��qf�J�1���1�Q8�O;!KG���_�f Ķ(i0��/���n�Y����o�X�ZJ�Բ��P��#:/��?)���Ӟ4�ތ�"�ܛ %�cDI��.Z��rqtH��N�Вi,�ŌX �sLU���/��-�}ܚq�@]z��3U��pǆV�(qc-��]�W)2���S���@�ˎ'S�C-2�9R8��@�������YK��p$A�D,31Z�H�*��\�vTV��k�.@����W0��X�'ʢ�
&n�=��h94������ �&��QY,фK��Y�ާ�YžA��� j�����Λ�g.�U�68JW�<xK>-C�.�`�����q���F��U*Ň�kdMy�Y��&�1�T������(j*���8��E5G��s�r
�'U
K���%�9oT�c�b �H�9��A�a�,�q���f�и8�oc�6o�员[�j ظ����2�ִ����P��cq#��2 ��2�4d#�;򐺩y y���a0kLټ���j	� �zہ�g���}�>���0pO�;�&�o�^�x��:���'��d�2B��n����W�S��vO�x5 !�ˡ��a񇍼7����#W>�ʤ�b ĀN���7�+�1bV#�a�_��2�엳� +h�]>2���V�i@���@ҏ�a;��W�}M�X�ٔ& ��5Y`���s���`�g�~4��<Y�u	����CJc�W�B�Eb���"
d2E�·d�lǉB����׎/+ǓY௿swy��e����:�
�wUA�F4B�T����)i����9�&�-���En,	i(�[�2�*��W��]"s2�hS�8�O}`��/ȧ|L�Ȋ�Ve��� ��F��W�V2ݙ�o4C�!�n�Qo�/�PQ���C*����)?A�4�썰eU����oc����˩��Ng�LkG`/wu}���������,�{�S�٧�ז�E���2�������D	������j­��@��z�&����P��-2�ڪE�I�S��N�ʨ{�Z��=�O���=-_)MJ�X�0v���$(ˠ��ο\a5�A`��%��v�������v�������B�V�X�q�	^��#CS۬kT�^��D����	 �Z����\ȥ��|@2�����+�C�	���R5�\.HDf���%$���}<�Ŗ�o�����͌��X��z�d��o�����*�M6���c�ǎ^:)a�>��8g+|X����rS��▻2�#��ΣC���(��JEp��$�s2+ ^�w�)��Z&����-�A��=�/�Y�M&i�J[V���o�ez�Ø��<�1`�o'�qk��$��li���A�ВKu����>��dUCT��������-�*g�)3�y���A�<��2�v*KYρ�R���[�Q�O��Q��L���,JR���m���U
�
�xP�g�Ơ�H���ng���=b/���gޤiw?!��)��#�g+��%Y�G[�i�Ax���G�~�9��!��E⇳$���;��"H;���ZF˜���+8�e
�W��n�=��P��U�#��8o8�!څ➚��+�	� ]!�C�)�i\=��̚<�����]W*w2�NG4�L�n̕g��U��P #�ڎ^���we�x0L�]�md���k@�YLB�G{۸�z\��� v��<�7#�g�_�W w�VNㄱ�)�F�QG�+��Agk���\���igt��R�,� �T��/�s�wEO�U_��7�]�����I�a }����Ќ� �,q���|ܧΚ��
<_�:���$���+�@�2�c�X�P���HQH��W�=oo�nғw�8HѶ��2�D6[�݃d$k�PO
�^��Qɿ�ٺ�j(Jl��4��Y�Puׄ������D�N������u���]`펍�A[��fo�3M@1V�N�8�n?}�G[�� �f8C[*#Ba���~i6 8��&zQe����G��>$C���f�,���ig���K�k�]�lQ=ac�U�A�����@ \9��&�)䉪���LI5
�G@9�1��&�G=U�ڳ�qx�3�"L�,d����w#�M�4�������Z3�z�7��#8�TJH��p�p�Mb�II;��[	%�$�k����qU_
�6�h�$�u�6�E��?M2|-Y�/3ۖ��b%�G����AK�̐�չ��`�� �!�޳UW+$gjZꂗ_B��z���/�`� ��[tBtM!���;Mg�H�|��c���W~����e2qa�����_�s�r,�X�Cd�H0���B�����5f`��Om)���^6�)�|�>�|Le�|��_�V	�M6%�ؗ�H�P�d��2C�c	5x��<q�u�##iGe��d���C��aO4CvDm���B0�iü{iOIw�`���<���#�_���Σ^��V���8��a�������҈��z��������Y?�^�ЊQ� �W�����+�-#P��Ҩ�Jz®��i��a�΂k����=$rZ���_��m���{[�{vO��I0<��c���KΘ\�����᧥*�#:x�ڰG#���@6.忞�	���@reSlvE�Pv+�9�?��/Қu2�.�U��������'d�'�W|u�t�b����8#���-t$��5̗���V��1l7_8�F��/+(|נ��x��E�b$�HW�q���Oݷ��/6��*��5��we~+�N�;����9��DPn�̈́
3�L���Д�Jq=��AP4z}���F�O�#�;�Q'��'y���5m�۪Th� ��^LlL�70��fﴽ�Ŗ�����d�,
��EU�A�CN}R[n����;k��Ka�B_�$���~���	~{u@+��pS>���VEȕ�Hajv0'%X/:�E]P_���|�^�2P�?�3�d����_���iK��ū��qg����-��'���w��|�Z�,A,;H #E��jR��RZ,m�7۹_Q�η��x)^�l��)߯�w4��Wuz:��5ݖ��I"S�;}��������iuU�7}zxZJz%�Q&קh���9�2�1y�y��p�C��8ڏc��Sx�ԩ����M�s�)�����k�;���kV5��(:R0M�d�;j5s�^+e����}��	�����^sb.G 1�>�gJ����V��l1Z�4��달�@���@$��J;M��)��'��`���ĳȪsո�_ȷ��t�ܾ�0{���]8�je�c�����[-fox!�ę�����e7W�&���Y�)��,<b��Z3�^YY�H���I�('i�jp�o�A3�P�M���ъ~JR5��ٙ�,�p�<o3�W��fHG���7<>�ۏ���b��ڏ�����p���^��Y~e[Xf[/���+ϲt�#�=l���0�(gZ�C�MR�ј(l���2/M���Q���_�T^�K��BSO������=�0��uui�����3Nb�ˢ�=�9���j={d!���:�瓒��7|t9����U�Y0xC�M~s�	�D����;�v��<%仆��pa9�����bq�F��>���魇�I�	ڎ�*�����
���mH��z�e��{N<�	��4��wu@ �C.��zo��_�)�\Ғ�
&u��>q�-+�H��&���j�f�t�u$[\�U���4�Ĭ�:���@Q��}���z���ʊ�~�L��Bx/0mgOs���KD���Ȗ7@�v��\��t8���kV� �Lp�u_-s!�β��[�Q�cYOଋ52���z٬Ql�A��K9>Ӡ�Pa�r�Y��FH������S�vWJ�<f����S|Iɑ.���)�>�����M� ��V�,^�{��Q��EI�+F/MD�nii�$n�VL4˜F}UP�:��� ���E+P���5��6��+2"�_a���N�&zx\�c��v��c�KS3��#�����2Xg��k��i��M��?���"s�
}�ڛ���Wַ�~�n�h�&
�P��uOՌ�a�10\�;.r��0	���ݜo�*4�-x[Q���+����I&��~̾4OO|ZIE�?X ����ʲ�<ph�����9/EV�x�2�[o�!��'����L����W ����]�"��t%����N�0b[:��&�����;������v�O԰ec:L�ּ���od,lɅ�����
���+����ױJ�wT��ߡ�uC|@xC�\�䒀�@
K�k�� �;� �ٮ^? �6Ä2E�ds�����.$��\�����w�d`���l��o�����6*���n�q�^��BC�%Kj�}���ګ.E� mZ^>�jO�g�����^�C��f�
}��a�;��}���-��J�yg/��%&l:C����XW j���g��������>�������C����%��I�Z�b�U���댛$L%Pù�Ń���빯�d7h�YŎ�=��:����aϺD���HG������^� ��C� qߚ����%�􋜤��oĬ��� 4�m@6�Oba��m��v��z�#.�_��T�~�f�싔S
 �NN����h��d���.�=#2�=<���O�m������G�q;�7;�b�~G�.��Lу@�X�F�N2,s��z��C�+;F�jI$H�9�
,Qhͽ��0�c&*��|�ы�tŁ��v�@G.���+e�LH��A1Є
�Rmud�m���")��%oo���[{��`���rw��:N[/�	��4*�P�,L1H�������H��\{6�hU����� �DUS�����S}U,/~Yj��įB�lI?���*[�Y�0N�\���XbpQP���K�����#eH<�ƨp�׵�~i��Y�QJ`ab=>� [�$"�Jwü"�X��_zL��q,4��-���-v*7d��h�����ڡ3�
K3��7�=e���C�2�\����˞š(Q#MN_�U��_�BA��;�ޱ;�-�M�&mg�wM� �%�.��	ȫS�,�3���d��ʭX7<^b���Qȥ�ڙ8G-�Q��rr�#W��)� X��,�Q��Ұ^��6�Ĳg�3��t���&+50��S�g䋵��Qf�}+��qs�#��_Fac�t�����f,lc&���c��N5�:K�xYm!���~���Z�.'2����p�M�����Ak1M�
Sp�]�	)1'� ��$B��/I�cF���\���v9�r�.a&[����g+��=��c��|ꒅ���3~�QQ�Y ��6T������/�;�:��ۘ�4/6<����:k�XЭ�F�a��Z(!>�m-w�w���Z9��4��#�njy������.��ߑH��]|i��7p����������n���[�?Z����������#IL��%3\�2:ˮ/�G� �C6
��J�ڪ�cVe$��j�E���&W�Gz<�5�"6�}�vn��d�BSt��5Y��O�T�2w�R�Ru�0�E�W���S�]�_��k0��r!k��+0Nz'�4�#�{�0\Gv�����,�m��~���� ����N]-MF��'�0�\FP��f����5��gEZQ&xtŖqq�^�*��4>���6@�n���Ӈփ	AP
W��W�W��
�b��v��'�W��Z�˿����\�Q����]Ē�G�Q�$1�f�/������6�գ�d��~��!a�=mza���hR���7喥x�t��8/��'����r��I&QM�"ӂ�/�g�~%N��<�\{��)��7���B�0��C.z�ˠ����ި1�a:�I2�ӓ��.};*��|ӽ��������]�i��ǵR�J���\>��̞E�e�7,3���d��'�O�Uq���)���z��!�H��UV��fq�`�B�u�/wM[�|�����x]���m�.�3l8�@M�S)�-<�7x,-��?� �z:~��rՐ�v(.	js9��#w���~;0�b_�rɟ2w�&��yA��'d^b�+
��t;x)�'�>��&t����N5E�;(V�O4e�U
'H����u�p&��sh�R�N��
�>=i=
K��*��e�D��6t�g� Q��m�J���L>/��~_�>�.Bۈ�C+g�Re`�VM�:���K�&SЊ$+h3���"�R�spN�����91]�C\�)��u�}�{'���S�*�I����g�2�
T�m�����f��x����
��0���ޖ1�B�+�����)UB���Q�ȣ��0g��q�b~�)LG�0{�ͪ��4(�ײ�[j6���}�4���k��#M���
�j��8�n����Xc:.����Ѥ�<�4��|J��Ȓ� �n�f�,���s����
�t�c�LXy�
�����P8�l#r"��"v�T'-��Q5K��iE��\��~r�I)S"E�U$N�����J�C��}�i����A��,�TӀ�T��W��%Q<��b`�>ڒ��<��?$M�a��&���s~������Q��d9L$�yί=��Y0M�;t�5�'S8�%4$��_ IK�]�tWʨr-�A��Yﳬ�V� r���4���-G1D.�i`��� �O�>��s�@|�v�;d�}l��R/lH��$	m��]�H���G�8�jZ���^���Fpp����+�R�kxx��+���?&�Yc���P�xvòǏj�k����{pU�fv��g��0�k��A�8�k����"3�6Q��F�d���wL>�֧a´Bh�c���Ų+4����:�NC[�j�*���"_�t��
�F�������-E���=�`�?M
��wY2r}P[tX�"3�׮#�����GF�����Os�`|���"�+�����ܢ��}~'�����[�aOE�i�tY7��N.7]�._v��;�X;>��^@�"�:,��3�^��W�װS� y�cY y�$$UX��O�^��n�֗d�9����d�\�*G5�25���H�o��� ���M�V`�Y�S����{�_{Q�"�R׊:�zP縸ʷ����}N&s�r��Vy�08 9Y�E���c�Q�֒��?�	}�)0�K-e{�1�y6��B�!߽ ��ɫ��6P�dT�X;V���:�˲��s��Y{Z#��(J ���B_5 Ô&�qg�����X�m: ���ꏏf�Aw0b�+��vp�G�S��$��xz�c��'V�hy%+)�YI߱�΋��-O'�M"ȸ���r�uL)���Y�eG1�$Ǜ�S�<um9���x��?L��=��[w,�����(�|��E, C� ��$ݠ���:�H���4�\��c*+U�1���LɾRqK�1�?E/���x>/�:�X��9ϖ¥�<�"�(�x���yS5 �7�=b�|Ý哴�S�!L�c1����%U~>?쪉ۗ:A��A�z�O��M�h�h��{��y�+Y9"g����? ��,��@���m���:C����N�*`}�7���(y}+vP��w:��$q<+����?k"����~��6��M-��H�Q���Ze��Ju�sj��;Kj��Jv'�N�qǿ� k:��겖�60�t�a�ڲb �n���I�Px:�l_B`Z^Lv��S@��ݜ|�q|g�{����B2ʺ#���`�	�ћr��?��rͲ��>�sp|���f�EV@ד�I�2�2mtKJ��ܝ�[�G�Z��s.C��<G�uເ����C�qvl����� �лoʕ_N�����2�1·�ߵ_�)R�d�o�Jܿҧc�������h��N�?P����IL�Jp�N$1�]�,އ�OF���2f���e7��5/bȝ��;�Dm�6�q�
<�`�oGSxD��S9�'��3 �X�L�*bU'��`�o�?�����v���D>�-��?�>��s��l�}J@�ъЪn�n�����W�N֦��fAP�&@�T�Kx����xt��PPd��,�"�t�����aX�lL\����6�ZC/5X�Y��(���B�a��R���[��B��d��'z�G�޿��Z����B��34�����7�Gz*LOT{�SO9Og��Aw��7=�} ç���W�"~��I���hrS�2RV2�"��4\����S=��Ѻ���zj�E@Ґ��w��#����@;�U�8C��Z�X^�}����ԓ�� �5n �~�n����Pg�J��?���r��B�7����{҆�_&uSh�Ǔ����w�sM���jq��߄� �wl*ut[fj_�@$���G�(���)�F�}��ӳKBڴ浤3�0�]�!����5�=*�_�?�s�`B,�A|��� ����p͓�.��7�"��$�p ��E��E ;�1��e�Z�I������[}v��@S~��w���G�!@+bu�0�)�k����CP��5�~~�Ք����^Љ]e�:y(�KI�ꝷ%|\��V��J�9H�y@��:���bS@^�yZ���� ~ /��z��ȋp<�k{�{���=A��=M�n�$���kF��1�y #����S���O�AZ��������ڵ �	Ѹ���	�?-�l���`�K���;��o��0����ˊ/A�E��1Хo�ޏ��E�j|*�<,a̍z�����Af0ĽF�����_�'�0H�K��)�ͱ[�+$|{�e�ut?�G>�]���'[>�Y�٩�kH����'���<0hе��������-uN�|�?��dI V���u��=?4n'LV)|7�_���OZ��\�K9IC�n߯�S6y"����Ӧ��!�4GJj˒�w�2e�nX��`6���]�LKt�287Xn����A����\Ä��h6}Q�$^�3Dɾ���\y�*������#�'j{�A�#�����-P��6�����)M9dE�ݐ�������1l �H0�s{ƀ��N^g�I����!7��V�NQ��*�^5�dϕ�D�Vȷݦк��"ٖN�K�Eä�¡s ���{���|Ǡ�ߘ �C�xo��lf_j��a2"_���o&���v�]%�9,^w/-�A�睦'O'�c������meC��˿�f�=�i�r�ԩ?�ڙ]��j�����</l_~wH��~�er<
^�l��R�����+l�]�L��j|��V��}�k����H�i��E�x��:e ��w�6<�K��X!���+\MM,Щ���þoK�Ġ,�2D��s�'E��Z�LR�X��E\����/�IJ�<ԅYW����qvo|Yԧu�������S0B�	���ҋ��<���͹Qϡ�����|��3}�S�	������JvLjr�}��;3Q�c)脖M*�ʚ��V&�i����k�{H�Z����9�[i�`�:w}���1�0��	n�
�W��쀂q������#���+�?�؃��Srj��$���)�4��Eٜ� ��W�D���lzr/xׇ}��l-���)���h
I�A����O(�s�����)ݖg����+<����L�I���Sp����	��r=fwuS�&9�Wg�-��x!�i[�[d�9��L�7�=�ۅ�(:����*���DS�QB�/���|b�%�[��K��&�f��#�[H��AH�VA:\�6�1"�h0Vͨ֘QZ��Սs�լ���X�5a��^[��IʕPd~9���a^�hG5�C.����ٝ���g�;��� t�7)�#�.-�C�K���N�3�FU@���*7���^e �:4���?jQ$����[��dܗ���Ƿ{�*7!�ֹ�T��?�7k췄�g枒�s�k?��}jS?���6�"~G���S��h�\K�	քje�$��1'J��!���Y�E;s�}W�(T�)����3�Es�^U}i�1`a��~YN��s�n���;��Ab�����z�Z݇63����K,���#YD�ߕ��[�g�d�t8�d,��i����+���#�!�U�O�	��Y)a���Θ ��w�ߘ����HBl�?M��x�� Al�	��ci��*�
;�x6�9��8 ��n��s�:��8V��o�3��U�2#���VD�$z��'��,��;ϧOO\�L޳�.͹g]�tԠ�gJPn��gi�R�"I/�s��F�\��N�&��D�Dcs�Kf����B���)�{�Ѣn� X����/^&U�˶-����^���U��.O��rX�8&�Л�/��x���Cbֿ�*pn���� �֘�~����V6v�ڋ2�t�n[q���*wm��b��_�X(/��h�>6w���?b��A������?m ���Ϝ>}��w����K }�QG�mr�'8�L	n�D|`��ug�#�k�)����S��
Ydyn=�d�2���c�j,Hy��R)5|8E�0C�q�-��D��+���qC���8t��9��T�@�`KW�N".�64�5���1\DO�51�	,��e|�}���8���Q�n���RB��vg-*}F�@z�}\�jz�XnZǚ;1��X�-�l]O�5��>J�&�������2����'��V9˯P�x�Vio�E�e�a�����f`�ԯ���h�w�1���`��Z���1�Q�os$)�")�QY��\G�Û�ͻOl�xO��v�G���D���	�R�A��m�re�h�Qu�3��%h�_�bxj����=�lC��؁8��}��{�^���f����fu�19�y�P[�=���������..V�/����J'O4��N'%'��a�\��1��_�,���}I(�*��a;�gU��a���:
=8��7�Իx�����H�9��q.��4z�Ȍ��)��BV��<hp��@Ft����LÄ锸��r�(�E?�Jߚ��G I%Ą;'M����S�����a���:r��A�k�m@�fO�/��#�ol��~у$S6��_�m\[�w8��y��F��-���1.�uѝ��}��{Cpxȗ�1H��ڈ��C��K@ Qg3 ���g9"��4X�93UW�a%�T���6hT�Aj��U>���YJ��x��+vS����)i(q���?чߊ���'�*�[;�K���D���Iξ��y����L\,�T	w�|�����U,�R��`��ȝVY��i��^�2P��0��u����t"�r��K�{����J���n�F�-�YA�� ć�d��@=Mg����?�@���<�v��n�?����%�dTV���M��b�n?�{�4O�7�$����N���«��HI���������Q�8�/(�k����S۪#l1��n�y�ob��h���i�--����4�vBӧxfb�P>/����l��of�	D�8W�y5u�bIl�b������(�S2ʮoW�H�6W�آZ}�ԜH�@��w|�M�q��z�I�{���?ĎuB@�-K�z�A$#���Q>��V�=P��UE&qH�3j�#���۽;J�|��08t��9���P�M���OM[��b��M�� �\�#�?��@�!�ՙ��CB��<��q���>���*ٲ�X�M=x�?麟=��q��6F���Ag�לa�9:1�������a#�ј�3��7���9��f�0p}�G	�Y_����p�� u��_�n;�sY�<�`�?�Ǌ��?{ǭHP���� D񉑞��K���L:�V00�o�V����gV�lC^*�H�l��e����Ԡ-�'�*� ?�����ŭ�?�elvU�?.��h�&g".���q���΃B\E�sl�uv�-��O ���ʿu����.�7�����T��?ߝ%�ͨ����^��Q�<[��/(��E3�4��u��(E��/	ZP��ߚ/i�1
<�c���w%X����� ����ژ�S��J��k��ݍ�B���`��8`�7{�E���,�V¢;e�9���T�I�.t�h
W�cҿHh<,���m��<[���q ��1�Gh�^\w�����O���)���	5/�m6W�&��1�������c�),;%m�g�J��~G`�<�?��*�Q��z����Q�4k��ц��/�쀯������pv��dǟZV���l�~�<fF��|�*�G��t+�6i�z�>��,rk=H�H����oP�Eۏމ��5/�9��Y��.�R��H���Շ�f��	"l�ӏ��K
���hm2��	�i*��C C�UDX�U�q쀱U�	��K�^>�.�� �Y_��#��&<n�!����?G4]n�&��-����쇽�q1���2�UL�-�.4I�t[Y����b�16�1_�ّ������{P����E���ju#�;�&:��&Aq�oN)��wW��� M�i^8���.8�����vw�u�*�����@g�� @b��mX}:%`��`��^����n"c"6ㆅ��:n�勵�-K��@9���i
ؕ�d�8N<�t���Y��$��n���;R,�2��?A!��8ɾ-�LvJ,�)h��1;���'��c{��00tEq�����w�C��;�?#�O{����S����P$�Y󞻭5�hB&�cp�-_�g��v$��F�?:j��{y��]�mL�`�W��Tg-<����Ó	�XwP&%ũ�
�g�㊛��,� ��Z�>�m#k$vM��xWeX���1�=�7�2.����zE��+N�,}�5�T XI�U�1�)>��W�Җ�V�.�6�����W?�R8X�S�rE��8��T��;[=Ƞ`PVs�c�.��8�-���\�碠�5�!�hlN�Q��m�S��0�n[�a���	��A[D`Q���v���Q�:�������B[d����zT�ɘ�~a1t�Ǆ��h��1��iTu�x^u�p)�%!4L��t�Z�8Eeg�@X�'Ʀ�Je��Q����S�
��']|��佧	���n9��n�c"�7��{��H	Ig�����U��l�	Re�"v\���`�ڵV�jI�	!wF
�%���2�j��Kq_�П�����h�*��!���k�`�:�2a~����Y����N��?�����jj�
���u  � s��q"n�|�,sU�ĴX���i�H��C���7�e�z�"o�h!�ߝ;����y�d�����������������ơ��0�T?���� �^�T��������x�X�u�T��rBI��w�����dRƔvC`v�`yR���RP��iۖ���ǀ�����|Q2}?
�bCc֮�R�1�/T��򷡢�lZJ�Lbk�����7�e���Um�j����E/���� .��Q����K�K�:tʛ��t�/��mrS1s$����I9�Gʾ����W�8����ϫ�<tnM��]ь=]�'d�+�=BNl#���>�ﰩ���:U�j�6K���͓�g�`�W�ō*>;sjG@Ź���Iy��mfۤ����״�<�D�ͫ��!����$K8%���Ѹ�Le�^�Z^5��m ��?�[�Y�@�X�= IBq��E!2�>�ǋ��2@_+�@�?K��vA$�֪�Io�*<8�O&����.�h����?_���H�㯈���{כ�\��g	�ؓ�(GP��2Aa�S+Y�23zaz}!�ܼ��(��(���-��-�=�r�r�x�g��l2m-�`!V��!�s�&���.ʏE�X����0��#bߦ���8�W�U��`2tOT�r�5���[� �h���GH�	I-Hx�3 9!ڨ���W�+b'����#�����CƦ�9�����33��w �y{��7R�S����0� dl����\"5�ς�XB]M���8�
���d���j���Z�5?��O��.1N���-݄��Y��'�֝�vsF!������gPHX��^�}厾e\�2�hK|�B��J���/
-�]c���K^�����ک��\�#p�����Y�?.�4���n��z�:�Cd��|�PCB8VQ��� ƙ��Q�2�v裏���2g�>yV�� ��G��')67�)dY����o��C�2��Éc޳�t^7�����َ�qR�H��#8��X|
��E�O�а�����,[�a�HAٻ�����v���K���p�hz�ϲ�{S�\g�q�U���g�u�q�;�A�n�8���˔�?� ��>��	s��9=[�$�6Ո�cV#r��F��mA�Nnb��ma�3����AmУ�vV���E.�2�����\����ef`���I�i���t����V�$�B�^�tC��{������@c��o<�_!>�Ţ�%A��;�	�)cS"��x�	<*Ѱ�I���^q�*U��]�-֖n���G��	Z�I��Uq��B�ݢE�
W���윺��/��#����������c�3ޓm�>(YR��ΉF��zI0_��K�����2~�N����@=r6��bǘ�[ci�,3mf�����߄ûsf�p��ړ���ԏ*e�FdI��~^�ɩ�Ij�/`�,��D�J��G��u�m-��j@��9�G�N=��5��o���	Zm2m��f}	�V�@N�T�)�� �hσ�nu��!��>��<���9��^���6��ǀvL�,�^tU����C��Ĥ�	Oq�`s���zL�;��XS@�r��#+aҧ^�&�8�g:Y�7�$�d�`���o�0�c��/�B=i�Ӣ�{����kS`�����֒H!
��]�M��=Ow��0�8���s`�3h1�=�4�P����W~�M��[*{b��7����.���E�NZ�dC%k�\�y��x�o;��w�{
@�=��T�K�U
���'	R���~Ɔ��xi`M/��skA3�ƟF�_#�bh^��v���9�"�@Yg$���5�=�7w�1�@>�D�����@��*�Q�Yy)��eP�����3���
�wx�H'�Z�i�������A�.2����>���E�c�l��q�6�֥f��kl�I]l�R�Ye�Ι(�%ٱ��T���Ȱ���o|����4`�R��_����n��{6X��s�0؅���pa�n��EUl˜^-�F�:��K��~���I0�'`�/b�A�K(���ăz�0���%��h�J9�
`=�H���8gL���Fl1����}���Ƃ�7ҘۮK��ȫ܌1��j`���]����ǿ����Tɑ�]�wB$�����z��4����`aB��8C��L��7���v5<"a/�B����xn2 �8�����I:%����9W.�d �Nv�eg*y/���<6���剗9��#ϥW�s�d`h�_�&��*R��g��,x`V�@�ۺ��1���G��
�K�У��m�al�y�1f�+e��o녛r����:�Òo���������+�b� B(�1��%�x��g {���e,*�ڝ'��Vv�OP�)���>���Q�_������N��-��mg+x��ƺ�B�R���Ū\�c%n#��䑣�h��i������@�1a�-���
�\W���;'uRi)5�0O�)>�6,�����=GG�N6�8��ofkE�x����Br�FP����km��_[����r2I�,����~�	�����w�A��'������{�uw׷q
u\�]<HH����y��9��Kcj���v���M\���^���JD��g �=8��z�	��^&�g*_/�@p��T3�m��C�h�������d�|9���kU��3��,̗+aLj�?���Qp�����7!�=��Bf@�߆�U�L���i�62��8���c�V~Մ�Op,Ԭ� �������~G������̂�ϗ��9�܋��!c~�w���(e��а��jҭ�X�'j�gT�˗ASV�Ӥu��{�B�S=>�#���5�F�'Q��>�Y��nq�>Шթh�
�������a�����#�V��R�o/��h�4\�Y?�D&3Hc>.�j
Z��_a��<dDe���qJ[�(�dgQna{n��E�R��L猻��<W=�7��CJ�r��r�Sͻ�7YyY��S��{�	<	P��T[/}w��S�/�� �sa1�g���~�
������ó �B[�1O�6�/T	���3~�K��3��*����%3�נE1؈2C����E7�z��F�$�����μj�_�wV����7��bL���3Q����Ct�p���3,U~�'&� ��k�&g}��b%�_�y`N��j��^��[T̰�";�u��+���/�՗�~�$�Qk��i�	��,�a=M��\y����IM�{��I�Žd��zmZN]��<R�n�#��Q�BTj�>�VӶ-����T-�C�<
*s�+u5oƮ��V����g��<����0�{��='�,o�	�������ۄ������J�Z g]\���\�paj ����͑PPS.'/k�����͓؀#���2���%;���(K�>)!۳J�Ʈ��y�h�A�o��?3��T��o&���%'�D=rS�L��Uw�N+8�A̓%�p��*��H�N%"����M�D��Z�z�药�i�0$�'�	&���~��joo	�9�n;���e����A{ʗbB�ɓ3/E��Z������H��w$�2�S��_�%�p�w��x�5W��>kz��|����hbؚ��F��߁ΘUq,�`D�߱��l5�3e}xJ�a����e�����?�Σf�F̈́�u�me���Zj��V��j�sߺ/fvab���p��ɭ��>��c��O�?����U�
�g|�� �f#�_�n�.��`��F[fԶ�Ҩ��H�- :8	��N�pzf8�
V���`=�����zǭ؟���d����W����!ʯr^���u|���F�����
^���ah.�l�D�`�0�`���%] �V�	r�J�_��!� ��oG?��a�FK~����,��T8w\��#i+���`_�|�묔μ_e4B�h�S8!ElW9m�ZS�:W>S�q�	�� �>;����@��� k{����Z��z]���Um���ݧ�<;>6\P�D]�S���\�] F�gJT�� ��k���Z�'�'������q
i��ܭ�7Q��%G����x��8��M�����{/p��c=��'�ht��y�������Oq��8�*����L�l�X�a{���|�IH��
���ʽC��
��\5���u��Uxb�7�'��9:��ar��se4�~�P� ��p~�c�G3x��-��e<>"�\�����P�}8TP/��%uJg@?��J���|}M�ȝ�V�k�Q�����܏qIt�[���t6����D>�1��n��Ɣ�7��h~ �����9�z��Z���<���Ȣ/�(9Z�c�NoA��X�^�;����y�r��^5Y�r��}���ZP�#���}�]�/F�*0xd�]�ܴ�E�|�
(��1��50�����3Ͳ0�e$(�ɷպMe�yP���3ԱJ5 9����)������:�%��71�O1RK�f	�hx�&�=FI�D��&d�'eIu�{ۦZ�m���?]B��oXt�D=:=�j�F�'R��2&�����̨Wѓ^�m؉� �62�O��ht�ucF�]x�1��̂	� �є�)�,�F)r��љ�ơ�6�?�*�$�9=��VХ鶷�:�J��*�˞��瓢~�0b���'$P�ˆ��\�t�;����&0(�^ݔ���iީ'�YA������)p����ec�=��%@_���~���SbfD�+�U�����2�2d�K��b��7�4�3�ع�6�F"U	3�{��.��÷/\ɠՁ�ަ7����	]��Ơ���7x(�HhXY?��u�/��t���4��G������ĝ<�������E�L�Olq�P���R}Jt���_�y���������y%D�C�x��9���	��������o�R.��!�Ω%s~y�O��6�C�B�r^�I�0h��r�a���H䟄C~��j��WFR��k�|
��|y���!>p0����!X�wΰ%��^ӓ���{'u�-���M�F���h% �w�����Su���4�Y����G鴩��t���b�^A-�=7)��~vu�]��$C�Ů�H��mln�:�`��۔9Q������G�]��O��%?L����k�_o��z���E4eD�N)����p�����}.�({0�u�)�E�8�S/ ��E�<&�ױH����,G��H *���JS��6�����<\�U�2��]2��K%�I<I�J�)w���^=�]1�Y�!�H�?L�'W0VC�xC�9�1Q��A����ga㖚e>�V������[ç�-��k�&��y/["S�Tw�bX�vÚ���>�z���z���B�EȌy96@!f�� �sOĉ/�;cT�&Z+C謁^[��ٴ꜄��F�U�ډ�@b0���S�f{W�q�h�J,HbW�n�Z���gu%Y�@0??f{-��V�i�*�jZix���>�SB��;f�M��RO��H;�����h���7X.F�v���+o��z�½74)�.�Z�p4�n��1����?�H^���2�|Y̖{� ��(��;��xԖ;���i�պ1桒��,�uW%��4��m-�e�����K �H�� �}��CO 	=Hs��H�@r⪝�ϒk�&�z Uvfß���~�spE�?.��Ü
�s9�!�)6��+׌^YE��ݷ��,���/�l�K�(J�f =Ũg�.d!�N
��m��@Ō�F�=�����j����b����?�F��&�n�Q7W�d�g9���2Ϲ��H#�N.*Dv���y����ueo��W( ��P��c��*l�y�Յ�J9y�������
?����a���b��Y���`�"g��:�ʐ����|��n[��F0,:e�I��@�^���j .�/�,Me�YU��� ��߈������GI�b;�H8�+�u3�����hr�
���μoP`��QϞ6�6W5)_�&e,�~�ʿ�{��j+w7��G��H
p��(qP<�<?H�XɥKȭ�=ЭIeQ&�s]�����C�������]�*�Eu,�Y�����9(�d~���w�X���=$�ZCN7�E��b��8M�"���N����6�V�|��pM��E�N)(AW��ǟLX���C���q���x �Q�����%'.�]�%=�@ɀ�$�&�%V���o�}��a~	2����{m��-�g&Y0q���O�v��=_J��QƬ>�܈�~��HA�ZBw)j!�[c�u���e[#2��љ�tG����Kä�N%[�����
��կi��X͏.����%W>^�4��n��4��D≼^�����k%�=�|�M'�\���9���CaA]�F�/1� 4A�oX���LC���?��Zd�\�*��zi<��X	�4�)<��B��!]O���γ���j=��^$��%�i��rP��?K`e�rg1Z|�f�X�Q� nZ2��B�L�8V���*�y�������=�P%w�9�sE�8�A��j�i�.�o!r�uY�i�ꈝ���
�nN��8�߃'ޯ�~[���*{�\�Q_L�h,�il���8��e�t��XK��f��L��>6��j�r,5�}9-�Q�L��G�:��=0������
Aփ�܀k�I�G�Pݥ�՗P���TI���ۢ�)}R���J���ͪ�ì�Bw\D��:�>Xc]��_�E��AS��5l1%����w�I�TY�o6ӷ��䗦L~�-�ML��5Uj�E=<������L�D��h9V��,�B��h�"'��帚����~Iҝ͉��	��@�}���� "I�|NАȰ���y�q�!�J7� -�~���n<uh/d�y�ז_1��i�3�{�k�yY&Im �x�����l���}j-_xo(W8ߛ��ц��y%��Eb�
�����ɔ�q�G�f�������검\�����_�_"�%��w"�U���ܢ�=��KiI� d��kY%/kZu������(�����(n<x'��L�CH^�֬�]&��9�5	�\^|��rR8t�����2�"�\��ӿ6�Z͜AV��f.�� �*LЁ6�I/l%�����%�~(6��īX�2y�k�9�[ẓI�����NzDym$g�����8��`�6������ڑ�`O7�1J.�FH���X`����~�<���\��F��@,i�p�UB�[�b G��_�Ce��@�_v��(��&����s�v��gEL/���`�B���)�ٕ�3��{�6�7?�}s�5<�v�y@}k�W�Ct��(�N�fD{RA��^O9KR�\��D>n�+���ʤ���Ƴ�X�~�9�a*^?:�i�G��N��c��QV�O�ڦ�K0Q���8ҀA�
;��xW��޹�:tcp��V���"�떂�U"�PNe�)Er�I��^�l�tSѾ��9��E��_�r���B�UE����#�Z�=�ݎ.���.ԟ�}��$ͅ�;�x]˘Q�FXWFa��Ș�&&�t��dz�/���<��\�"�(��g��X,T d�i>����Ϥc���֮�>h�c"�E���sз�L.b��lSMܱ�NO�{��C���^��$;5,�ay���f"0����k1�lʤ�}T�C|1���4�e��B��&�����fW��T�+q�J���?�M&�� 4�}oX&�n8���	��@]B�;�Uz�&LـP"���Ŗ6V�����"U��P�z�z�����O�eQI'@|~�ۚ\�f�;�ʀ�ý����
�
�S�,�d���͵�W��N�)���<ae󾾣9��k�Qgy�g�(]|7�
W���*�����F�U��0�1O��Y�7L?X2\�C����_�ev̛�1� �ȺA��kڵQ��+�yy��X3�1��Ck�8�YS�D$K3�+��-��	���ƽZ-�:���8uοۋ�%�E3cXUZ��!Q���RO���X(�jȗUBԨ�J	�Mw�����0�U��#2N�kr"i���K�K��(&H/=;�8���	��;jvO3IŋⲼGͭ�!��4#œ!�'h��0ⳝ�o�W���	g��7��g�l�S:h�iR��tp��]��5��Lg�R�pbN@����z!��(�������1�g�7�t���'�Q�\T�n���PSZPҳ��8b�t�X����]�k���F3-f[�"�~Y��4��+RF��a�sz�,SB��<'��׭�D��CC@���b�_�{ ��p&'zҰ�cQ<`�Q�cZ�;��Xh�s�6H�j����xrh��.$u�i���}*؍����V�,����3��>��=�@Ct��[Z)ȔY"<�GB���>�����45>ⷂ�퍋�5м�_��X�:��~D�,��,j��n!����1�d�� � �o�����B{;�(���E0oڠ{Y	���imҍ�/BR�g:'EQ�����_a/�uC���Ԗx��)_Y�n���R���l�p̨2fh%�F�� 0	_�;21�p�gw�z���L���͙&�)Ŗ�A
�H���cv�'ł�|�ܾ�v�W��lں��rL�Q�(��k��"Wh�W���ϡ{P��Zb���{�)��~E�?�!���������Q�4��%M�K�ƢW6��6'C2���֓�� a�k:��Fg�A۸�����.A���[��K'�
�,#��:	�ya�(|@$�M��p�Z��A�Ml�9��;� �i��1����ȴ��ݪ{���iD</Y��o�LB�H&�>�.�����u�||����{E��M���a�/�ξ��,3;�7���kb�����ð�y�.�w�Y��t��J%	����;�l�YśI��[�IC~��{)����t$-�X��{%�O�R�\=�<�t���Ȯ�N�v�EWN�o��/�ʡ����H_����#���>�f��&DTD����xS�t9��ǦT�Y���m0U�l�������kI��)3�r�����-��0�ǸQc�4�$�Z�ڃ�4�[�� }h&�`=�Ij�,��BX�JN������z���N�."�
��g�"��Mc;��>���D��I�.�g��T��1BƉ��z 6���Ä	�a��=<!VWq�ӿ/I_����+��7͍���Ls��5�"�l�ӷ��	T�1��(��E��������6O�_ue�
2j��(�E]A��=:? Sk��>ݎ����l�QG�����Rs#�e�E^ZN���'!ܑ��JR�CF��^��^� �B����P�v����?9Քzi--M��>f���W}�J�B�"�������#"�+��!w�F8��m�D�@%��I#��P��5r��#��f���]aA������J�'�Gk�Ȱ���c�G3�ð^^�֞)v񌚵|�mjv"u ���a���A�x��1�h��<4rM�t��'���R�_��>�����q0�l+]�\�i>� ��rR9�m�\=��W���0�� Λ��� ��Vw��ͷ�i;pF�t���8o��R���-Ʊ��6f6mE��K��"��GdkNNh�Z�:��!����:Ŷ�K�<����AI�Ŗ����E=4�QX9'A߁�Qi�P0T$v�M��X$�ӥ2���|��D�@�e<yvE�R�8~.+�?es�5�=��&ť��yL�#>+�[!�fe2{�M�D�M0=�9&a��c����a�����I���0�X���v�Q����	��Q�!�}F�m�e���rW������@B�(h��!2J��"�1E�~޸��nZ���l�j30�Ԙ��*,�$��� ;t���ْP��\��A%?	/ ����ח�ܧ��zG@j�l���ԅI?,=DP�W�t��� ��D���V����%q��a 3Ⱥ��!1s-BL��|�;���l���T�qO�����^
0!X`:�&�R�u���d���5$�wU^:�L-!�kVe�a��L�80�
� �q��|����h����|�Ş�ˊB
C8�bċ�n�مG+v��e�&���Σ��ϼ�6�N �~oQ]�K�"������(�%*��KH�k>����/�Y�K��_�vs�qH"���ߗ8?� ;TK*i��/J��~p�U�쿯�A���ɋb%&j�hu�)#1d�o3�ݣ6&K����O�:�G�:��~�<��m��2�X���	Z��A��;̹w���K��xֲz[��K��m��ImO�e���ߔؑ6�{"�=~�Ɯ�n�������?�1������z9�Dz�^�$��l����%����\��EQ乱[9o!��	����n]dNP�d��u��A��
F=�� ��}v~LN�����aҫ��8
K}�v�"��"=���b���$��<��x���P�\5�܍@(�kr�Ɩ��<9ͦh=��c���i����wQ(l�ҝX��
p��	(%�k.1�!�	�=���b�
ݚ���Mmbc'��������c�&�q0����Z��W���!���#vf6�ĺ�F�t0dB��)}0�<vypN||:��� ��c�i�&�����U3!��^�ђ����;�zȡ�g��X  �.)B6~J���:v�(�Z�6�TSؠw�N��4����U��M�=3�[���q���5n�T����O=M\�7 �nv�\)��̇��T�8�s2\�V���ʝ�xk����#�Cb�7�FI���t/c_$��T,sRh��6��/��wP�@|1�Fi�1m�`No_����H�b,,��_�K=����xS�:+F3}Xt�(kG?]<"H�8-nE$�V!�%������Hi�?�Zm��;z���9�tۂ3����W͋,ȯ7����GS �ſ�f�@*��b���GL�o��#�̀�3���6�N�Νaɸ�v+<s3�e�fYϭ0@GJ�B�\1�9��û�?$A.�e��m�S��d���s<�%�sX|	6�K�2{�Dy�Ip����s�7��wR�9?�x����
&{�V�|�χ��	2�Pb��Ƿ�P����HH��U�6�����$z#F���@��`��Þ����΃aFI�)�f)��:�ة~�L��Nr��N��[�[p��&� �k��۔S�������^��Չ��M��)#u+L�f�+�9�ѳز-y�.���n���N�t���p�?X(�d���t@h2{{Ÿ��QS���Z9k��M����*��<"�ƃ�F��ݣ0�D�A�nG=�j�h�P��	H�*��Hܶzc�~���%�Wɖ?T�qB-���0�~�3��� ۋd%*}���(�d}��M�) �(r�P�!��(В��B��O%�N�w���g��oäf	�W�S���%!�nۿ-!��S��o�k^������ݛ��y��OR�w�L��+-�[ ��s�,�$���'��I���͈�p���QT�ItZD�+�(N��g��L�xlV�M}8e����&V�����i�W��W]b^�&�Y���h�\&�G�̲e[�g�cf��d+�{+#+�-��m�������1B���3X�v�7��#��/�{�\�d����[���ݛ4+×l�l���딢�-��N�R)�)<%Z�w�^(�;؈��ҲE�wcvPO�s��P���/�%�䢜<�����0{�sp��R�m�K�3M���.�|$t�|5ɀ�$���qR	X꣣�,C�����n ���#���˜����R���M�����d�x{|�gͰd�w$E�a�p�d�MdG�W���4��Ivt%i�D'ζ���*P]�f	+u�l���N��q�&,�����(���<I��l�)<4�eQ�REB"ļ��
v��L�M��o�)
ee�*>z���9�ݎ��1�l0}3���¹�Nptc����&�=�pܜ챸��:a� �b���*�Dl�K���;/�Sν<,��.�*Ɖ�W���Q@����1F�r�0��y֖��غ�/sX�ryF|���� ��wv����}����po�L�8m΂�P,�3�=��;�s��䠵�F8�WDh@}*'[��O��o6��",c3D��%g���ؠ\�܉d��+լ�K"��&���+"�Jl̃�~<�H�O���o�d~�Ӵ'+VBL7����K��D =2Ɲ�����G��_����jF�+h@�����+����~F�xe���`Zޒ),� <�໣�[�)�D8���L[�Q��K�*�ό8ܬG����JQ���B�@=�Q�<P?�"��`˙� �}�����o�R��h䱶��Y�T���J$e�H�Y:��pa���e�^Д���9 84��gj�~����x �w��L!��`Ӎ��y�@ɔ�/Pl�B�?2<��L��3dW4l/��{���_B�9�L0/f�^�]��@W�U��T��d4�Vz�"BJ���Z���)<�!�
-Z>��ӋCJX�.Ť��Bf�|S��sMՖ�K��&����^�������	�~�x�*l�
d�gɴ)`a)U@w�yX6���N,� ���u.Vɱc3^T9P����W��EO��n|�[V͈f��/F�Km�ϔab�x�ҀE�}^4k$���6��|�e�Y2�o��N����m����ak�r'}��I kW��J�`ğ��嬘E�˭�d"p�<���Q�[��%�E�Lck���
�k���9H�����U�Y��l�ō����'�`��P��.��G-����M���Ħ���]�rh._3���-6�Y%�3�-�xW����У����plh7�1�=G+���HF�Tr�3��o�s 8�z<yE��M�Q��D���8�ʷ4����OZ��?_���̯}��)Y��s��Qb�&(�#�A�Qo/���Vs�Rw[��7&c�\T�*"�ũ��ƥ�8<��R��;�q\:Hg%��k�y�]V��}u1ס9� /l���U�������|-6�F�E�9x��K1�ɫ:#�2��>
r��h���z�Iڎ�C_}�F�!�u��se�|��W��ё�[^`d���i�R��̉Z��(h���� ����������Τ%��75��Y��b��a`���\n��"p{>�WTß~y�m�  �{��)t[z�����\9�W���ե3���
�h�H����(��O<yY�c��'Rxs�1� O���0��9p�݇���;!H�:f��
$�Ez����Q\󖧐 ������1U���f h�@+����y��g��P�5��xH8�{�\|X��%�f�jM����Uo:�(�q��ް���Iľ��ʅ�ǉ��[�W�{O�,Cd\����9㣶g�������#JclT]�|C
U�6�&@�8��ˍQ��P��Oˌ��&�>�
��s�=���)�[��۵�����WT�m'�__F�U�$=��`<eF���/�g�#����Au��c�]<&R�X�2K�D41�v��
��)�z��e�9@��].ڲu5�*���k���q��[�%4i��c��cU]�kO�ҁz���L�T�������y�{x�. �g�)٫���ej� v$���*���5��B
,a��JT��$��Ր<�=j�}o�ý�o^�$%�h��Sc�Zd˕�k~�"���\�?�z[n�XA�?WoV�tI9����~�Ƈ;ԌnQ�K�td�ϋ4-/xG��I�C5NހN42�䒭��`s��*��t�-����z���E"$�8A���C/��k��?U�y1�o�􋷷�'�U5����%
&�[���v��1�(�eś�V��+[:k���`�x�|9"�G��H��)}�K)����T���L��8��<��ؔ��=�����ܜ�5-�'bf.F��4�כ���JH�V_����E0��1��/�o�B��w@�Z���9h�6�=�AF�Ӄ*�w�2i���M�5�'3u��PJ^������e���X	�8�Aet�K�}^��/�4[�P{"�w��Q^ޗ���P��b	�/�<�ܔHuSg�aq	7�������ZQQ��A���j�*�w$h8@fr����:H�'��/JE��P�X���P�ohZ'B�������5��c�4�f�z��5k���֔sl>�SQ��7:2��H�i-�;%�Pn֘M&o�Յ[��TS�9�1T^2
=a���qV����c��1��J��0��ƍ���a`��/g��󀗄=�JZE5����-�M����������䠬�Qy��[A5�t�����J�r�q���k^+'��vHÊ���6b5wO�y�W��q�fZ�%�	�7�R�8h��v�3zu����;�����l0R�mp��8�ٱ6{�bN�K}�\��,n�b�6 -1�ٟ,���KR���/�����fy�w�q�A��qz^ ��n���L�^�E���&M�rK�U&Z��naKیM����i�s�d#ɜ����*�p���N%���eJ�H�/�<.�|���
A�>�(��Mň;�s��j���iI�\z�
��n2����m?}+�k���uU����<�v�q\���l��8��ȕ
�M��P�.��ǹ��ء>�1��B��٥"��J����Ap�X�V��t�V�.;d�_�ۼ�+�0�ę�p�t�G0�2V5��:뫺�*)���w.�*x�9����ŷ')�uҫ���~�����M�g�Š�uU�߹.n�_�d��L�?��h�|"�k�&�:M!.O��]��'�u-c�R~����UՓ�CD}v2YXak�M%�U�N<�+���G�CL1դ�g�Jˁ]��/i���"�ć��C}�:��"��F�<vܧL"tjH>+�a�~7Z�XKkB�01M:o�O�
�;�]��J>�u9>H�o]�k���@q�2t�5�T
0y�ݮͻ6S�Gus
}n!�H[�煯*`�h�6���u�$j�*6���_���.���2h�">�*���D�W�Ur�P�/n�P����y�tu�<8J��0�����E,fi\:�@��	���d	�׌7+F���|�X���ϫ�i+S3]���.E}�c�5	 �v����8,����[+,���;���u���/3�0��mx����tI(�a��dL�>x�~g���Ysq����	|�:1��߂_�;!9�eZ�S-�?J�o���X>�TfP��_�l�XPh6״y8y�l8�b<�����y�ǘ��	v�[1�ls��뇊
���.�C�_w&����ƈ&��r9l�Z�Z7�
!��7��I��r��n]���\ ��,�"o  й���O`[�������J�����i���J���('��R�q����nH�|���\R8��U���E���\�!����:kN$�����4�=HH<oHt��R�Ӑ+	҈�H�ۼ�E���wDo���s��A�SF=D��_vb�͢'���͎�Q���g�ڑ�(P�A/py���J8z�æ�D���p#E�� T��l��J�o�iݸ���p2A�U��?�\�#ξj-��z���C��#q¥�d	���h��Nk��ש�d	��Ť�e��0Q��{M��OE��������0�Be=e������лN���7��1����`���7�*�[�����sI�^:d �ZN�e���^XX��R6�A4p��ҁ�6E����"�KF*0Ec����\$c�k�b�[�!c��0��%4ⳙPܔ���>��}�|�݁SC7��oyUq�x��'�G��+4�ӓYhEw��x��vop�3s:hE��r�z�O�j=n0�zh"�J�ױ'���w�^���g5�Ч����#t�;m���QOL��i#��5/�|�͞�C��e�W�b vƚ>[�� �"��U�gl���%�g��`qXF��LFcfź��l��()N@��k�r5D\C�����M�5�n?$kP��JY���'�*�K�c����Ol#�b਻~l�_<|� �
���o�`�о���_�O�i9T�8��X�6y���B�5
�d�&�񎮞��i�G���.�zxa�(}�-t_YOP�?Ҧ����GC�����u �t~pи���ؚ�>.\��]����]���Ǔ�_5� f�(���t}%5T�}/5x�-�Eʤw�K��PB��mX�\Ǖw��}Ȟ��%��>	�U>�N���)X2)cY<�����&��	�(�GkS�"��M�I~s�����͋�Y)´���hd��K����x�,-��'HX
. �����E�dK�ڞ�^p0Y0r��39�:l{�ff։�/Rp#�,�ũ��P���������q�Ռ:*'�XsѿI��j@�&"�!�m�X)�; tz��pd@J6mH&�:� ÀQ>��
�n*��"q�Ꮍwg��^/*9�W'�V��B;���Zb��%����N;q����C\��C)��(REđ�H?,73WZ�U}t�*�t�-V�J��l�8��� �n�N㷉�����j��
Ӽ�tZ�'ԁH�I#o���DD��yE�Zp�ؓc�!�&���E��D� n�&h�axZX�5�q�#Ŀ ���s���.����N�q��o�sܰW�i&c���Y`��WʷD�P���
݁G�LI$�v��tj�P�T��OZYB��6KDd�a�	gXv�'���Yڎ�s���pa%�NK� ?j�T8�}��QWar�t?昃u2ǟ�CTl2S/!+�J�~�Y��\[��?�=�z=0�\꒔��W}�	� p��ml�}��� ���*��*�=��4*XT#k�*����Ո��LR��w�=XU�/�ep
�\[��&���>�\5�
z��&�7�Ź��e��L���.K���Y'����>:�:8yI@��2`<�P	Z�=o�|�w�5���5+~^`e;��fp�%*���T�F������o>p�ha.r����?]7\Ζ�&��(�lc!���cV����S��t�P�ҟ2ay��"��	�X���"�o���� ����&�`E�s\�.��׳�hٺ��<b�z҂�ȑ%bc�����]����f�3*0c�wV��-��]�7�!˝?�2c�3�:%g�#��T�P�y�?���]�&/;�\}t��= `ۡT�~�8 \�����	�S�!�dM'���s�+���A���S`�B:�Y��;�) Ը�1O��'7�B�܎Щ�HO�����_�� ���d3�m�7E&�Tޥ�:A!$����ud/-`�v_�AZ��U�����'q�4�Hg�o�1x`���� ��[}T�uJ)��ږ���ʋ��d�,#�u�aw���T�-��8�>R�XC RDv>޾�I�8��W�Gn��8��	�X_�!�Tp��0�2�_K�`�r�6��C���s����p�gKAtAt�+2b�����Im�o#qh}.#U�9{"�a���R���Ϳh�D����4�-V '4D8�@%�Z��eHRz����O}'�[����������TB� ��lo���]�t�-�Ѩ1tk�K�"�r��~]n�po>�V1M��H]�C~����oj
s�l���y+��0��`�2�*'Z�9��|�_˂�V��t��4�"�o�~´�p�	c���oG�̧)tO}�j��s�����H�xE])��\RBJ�H�r퇤z�����$��g����R3\O��d�Wl��4;f�7��3�&���iF���H��r�౨^l�6t����&eJ|o���1����E�qWܭ���1	t��Vl��Ԅ�[��j��_���#�=le6�@Ê^���V�Q�z�
��9��Վ�����X��Bl<���vi%8�A��]+��~ViA�ፅ%�P**�>+6�t���7&���a5"j��T�n���=�р�ۭ����N3���&�В�ɅN�$�yL���:ڟ!�1��VF�6����ꀛ/��C�4&���y�U�2j=�P����h��1����q��4��uC�g���C0�,I6f�ΊVDYq�-�l.���Yq�E`�[e���l'�`���$B�J���K�s���+t+)���`����:�s5�OdHk�@L2�
�5�qm��(��K5���u�0��՗zNZ�Y{����97�$�;�(pu��}B|,�]7^T��n`ƕ��C��b�WsM�0��Q�.�a>�z�G�fNǴ�2��./�s�	��eղ�Zq���~8��P7�Jͧsl���&��S~�fr ������>tc;��}�� <�P�Ƃ��ٟT�	0�,��G�&�Ǐ���Li��o�&���p�E�aE �m/ظ�6�����`������V���o��.q�7^FYz���m�;{�EntY�6�<�hB�.>��c�Ad�[��O�H��y���ջ����z���
��~6\�S�Zʩ��R�B�Ӫ����0��Wd]71���0F)w�(1 �6s��r��Z�?�)$e�p�u��Q7Ug%,L]�*>��iVt��u�M�ƌ�h.�(�Z�o�i�%u$�#�H��@Gl�G�U�H�z�+�WL�y��,e��&���99�U��&:$����F�1]p)�b4t���Ƈʀ`��#713�H#�q%�i g4k)]�t����V��ȵ�w:��
����E�hLz�����*�K��m+a��o~fu�V�'�E�8��#�֘�4AX�z���Y�a���Y=��_��p���b�3��fq}	��!��:,�'S��V�C�a[�+r!;w��%ee�1�yU�9��K�ijHs�qz��*�ӆ���ث�s?�ֽ�&���-��[�Ժx�^S_7$j�yk/�Ɔh5�z�}rR�i˲�o�M�(}1� I��}1Rk�;���u�����K݉���s���W8��!ۆĒ�H ���Fx�"��O'�I
鴛ov���N��N��&k��_D�V�\_?��*��C���m�I�ԑXH��"��*`q��m�&���;���.���.8�=�e>���X��଺��w�)ʛ�`f(XC�A��Т���!;?�@��<����ڇ"c��N�6?E��Tw���`�˻�l�5�1[�hTE�O��[�@�FO;jG2�l�s�.l<]�&Pa��Y���|#U5h4,�� Z���0e:�/a�.H��i�n�Wң��.u�e��;E!
x`�!v���|嵭g6|.�B�%Ǵ�I\�P�[���W.���L�G*0�"&.�)%�9J*���������
�Ư��H9b=���i�iZ����%A�SL۝#`�[ol݇-�'ؙ�[��l�ĝ�5����.죾����v�zX����~�4!�
vq|h����3;v��+[�4�����#دrb.��Ս��"��J+�Q�I�{)�2����\r.���O1�ن����6��lɵ�)ݣ����Kq�V�
_IG�/� ������{��CZ����<� J%�;Z��ܖ�p��e���\e����S�]��$�^|�G�+�D�/��l���c���x����L�p�n#k�����޷���ɿ�1��������M�?+�ͨ@�A�&#D�����S:D��%�G���8+&���'���V��H�*�s_d�c^`K��.u�L�TD�N��n{ЇT���-D�Ց����-\�E_�h�Ʃ�C�~+��xks��^U���w��lC^��#Y�d.�h�<�ũ�ٜ��Wm^�%�J��cv�Ƞ?f�$wX|۫S�=��	<����_1��2C)�h�[��2��� j�Pz81���U�\������)���T�{.�N����{9�l��,�Ur-�Ta�j�G��U�{�1������)g��P��䚟����	^�صK��Z*��d�'U�����t���p����BVӍ-�9�O�����7�"?S���z����+!H?�Lԉ;����!�J����;�Ӏ�MI*�P���x	�B0�:ld'�B��@������eM�ƚG��Q�D���ᵤ�<fn��Hsp�g�*쇝��[�U8@�Bƞ���4���n:W&�����\�l��@Vh�d��xbġ1���D4wb����6�{�A5É�y��69�N3p3��类�6���zU��qM��m�
Q�:5�^��Z��!̣�|7�s��I��A}�`����]�9%���R$%�s��9��I�v����39�m+��@6h	��G���Epʬ�T	�k&w���:�}"ښTX^�Zt��Hض-����s7��Ěz�u��C��3�>�a�=Е1	�
�.��Gۣ�L�C>�ZT&.�7ɡ��tp�F�/I���}u�ηqn4�2Qd�E'ߛ@�F�
�q��W�k�T-��j��zI�s.��������g]���I��?<S�9��X��j�sٷc���Ȏs�������,��t"��YR��Iè�/ߨT�K
�?�;��ZcS�a~�:�l�P�һQ�Ol�x�'.�@�~z����dޕ׀�aЂOn;iŃ�A�%��ʻ�`
��� }7bڇ��b��i�&F�F*JAӆPz�IS�4��5�� �j�]4��L�����%���:����<�Z��Ry���:��H·�nTV��C��0~=L˭X�7[r���N�bC���������.��3�S���)1�[m�@A�%�U;��'l�f�;t�`N�	W2�y��]��ۧs4�[�h7b#4Z=-�`�B�.���YS������L��R%s�B�'�����4tX�������f��EO���W�@��	.�����&ö�~ɉ�;��
��,o���p�SA��S\]������t��?���Kǽ���tׅ�Kw�\����g��qw��㾴b���D
���[�����!�=��XT�v���������P�C+
�^�����B����UB6Q'&�@�o	|�(��T��Aթ��fF��B�74qi�I�D�2�1�h����*j_f��d=߄���|S<?�<G!��x^K�2�S��ʰ��jF��푖e����zmR���"�2���q�O�6�e�~,��iN��j-0�it�]�;�+���[�U�|�����{�(��/ Ϙ�5���\>�,��2�UZ�_{A�Z��yj"�9��!��z*���UZ��iޕwS5�9d]�h�Vv��:��8��U�ԋA����/O��Ϧ��wn۰L� s@�� �0�/Y~O����I�Ǌ#��Y2T����u����C@;��>��m�^��3��h��wa|�'3��9��������)�� h�`��j��0�S9籢d�D�CeP���ot��b]��'E��)�����g�]�Ǟܚ�:��	��Eq����F�[�'���A+m�s$�*��wN���Z������x�L<~�		J
)�j�n�p��^9ry&䧕/��s��+�o�5\�A��=��#2�g�p�}"z�ɡ!�	R�eB��@�
��bC8:�	Q��K{^��+
L��_�+�	‬��7���y;ś gʄav�M�qլ�P��Ux?�w>��� !O�pm2��Q������v�Ɨ���n��﶑������.�@yFŐ~��K����ѹMG�u�k� �Y?��ykN&,,�*�����+���`9��Y-�a�BB(b�s������AHX��^�7ބ�c��a�ZPf΂�{�~ yC�edњ3`4-�+i�B�!��s�����,K��>�U1�-���*��a��|�F5E֭��Ӑe���٤����/~ SN�-cS}GJ��n�~�3�����k]�mM����ϻ�d�O�.�e۴q#iK�P����A�L�͝�iwf���b��Pb,���(����	(�`5�w���p���P�'~5#=�"-˘�xv��txd~�����*��DHkN���-�Yj�!�~����1e��;NY<�� �-ô��^x	Vd��q�0���*�q���p���9����p�6����)�ù~v"������b�B�����9���x��,�������\�@���p;�����ɘ�sQ�8ؐ�H6ӂ�6��}�%�w!��s*ߊ��D�]P�
���΋4�0k3���9�g<_�P�3'\�믝8:�e�d�\�K�:ĆZ�ޒ;LȾ��\����ѝΨK(H^��h%rz3�C{sIV��?2�q�hcƟo���RS$��Q���׃��b�����$ۨ�1,`����υ��دȂ>�)�-`a)�!2��缌�E�(ﳤS���W���tz8��
��kt�� �N,$?�_xa�'�)��	�����-yG�>�V�v;��Ab���ʘ>˄��$1�^�����ef����3�����t�+���qBʊ*��-�LB?@]�{��R����΄��*'L�/9O�Lx� �o 'w^0Fev���uJ���{_
�I�����f	Wt������diG���|��ۑ�O�L�@��ǵ*��(�����j�r8UO(�P�����Ar�U˭����4\���3�������>D�)<��ƗK�����n6���-fr���1�`�8�AY駽����2�,~G��2� Ϋ�M�3�k����M� p�u�~ꩤ�i�v�J�����i4Tķ�\ļ!�i�[�|�t��5�:������)�l�{"����D���cĎdtMT!8
�!Y�^O�0��,�C_�-)�L���C��M�M%w� ��U�[d�w��H��u��K������	��)��ubG��w݆k�����J4N,hJ2ˎ7�����ܟ�z{bܬ��w�gϽF�o(W�6�g,#f����E���PT�[c^U�
������U��OH�dRI�E\�ә������]��y�
uqzFj^�[�{hz��	����1jr�v����=*}��v�����
�҃ٸ��T�0�Zao]P�L����}lk�^�Q�渡��#�ag��T��evDK�;c��n��Mm�ć�21��2Ag�[>����G�)�*�Lw(�;�p� ��w&Q_J�[�O�8�Ȫ�!�h�8�p|L�7i2Y	7��ܘG�Hj�����[�n�m�o�rX;�Ag�0� M�5��x��s2�#kT9���ͫ����̶��4�&�K?�ͥ$�7�i n
��:������b�p��+�z����	>���$?&c��v���\p�*���V��4h�����6|5�6\z��c�b�.W^����S�����Q�����ۿ#w~�l��p!9����F��^���Ĳ�.�T�F�
��&���ی�T��R��>���-1�&F���gQ4p�ʌ ��{�2��g|T7�l槞,�;6�=�о����FF7$GM��9�W%���㽙`���˃�=���o�'Mb}��a޼2s�K�*d6���*J�ss�~.hx��B�%`��BYq汲�ygFP"F\aѓ��]���)ۣ�M�z��+���:(x�.�bn'��-�\l\h[�π\���T���BE��A��N��}������7���ư�O�¿��}f��9hɟ��WT��3N��0M r/{�Nq��'�8��Xu�)��R�r^����ޔui�&u�f���`��Z�"v�\�V9�l�J��C�����4}�H�(��B�UV[F�4�/�s��Xm�;O�6�Z���;�Sߨ�!"~`�B�*�OX�dt���ȸ�8��<M��Ԃ�5<~q��bԮ0���c<1��}֟�z�LL%�<r���ɔ���m�}���c)�V3F��MC�.�zXCml����K���������Ai��)P��1�L�\H���ٴ%�(Fb��7�Z��B������͔��e�����K뙋�*ϻ��f˽q{N���_�0{�����*�oo|�KHY�G,��]wa�i�����Q�w�1V^*_~xJwE��Iu���;`ӝ	�	��������I�Ha�Bj�¹!Z�e%��;
�i?��;�Q���3��Ͽ�ļ�ޜ�B�6�;�LF�8����\��W��Iv�T}�j�1�6���ßë��y;t
�VGF�<�M1,R���=�XV�I���(�Q@Q<!L2��)ULr,�V�NS���MQqe���w[���,yO���J޲�pRu��e��anh� l�U��u�ѯ����YUK{�) 
��n����}��;�t���3�.��+ (�h��:"� ��+F�e�� ڈ�V�9j���J��@֒�����|�}e� �3������Zz5OR���^��f��G֑�s�,z�\jAc.0�(�QR/����G쑶�>�v`�,�fI(�C�K��5���Y�d���������Qz`DC�T�\8�ws�A���['�y-@��pO������rC�����)�އ4H�ݎ�E��a���5���1�Hm��9&�T�TD�������6�I�X}Z_�����%0���l�څx/��V����a�Å�4	��q�#�-A�p�2��T�9=��y/�#�`\��@E�g��E8N�1�����V����/pj9��Z�6(�n �"ͪ�E��`�L=&MV'/��(V�V�+Oy�jc �����Bw,o��B9�Q��Cy�3%���<"~��vl|͘�a^�sc��l1z^��g�}�����h]�.AzQ1UdE���EI&�K�#�:lCj�Y���e.	�y�;��y/-*eǄ�B�6�VS%��Q�_�/�mj%*3b#^F�s@��v���M�Cn�N/`�,`�H�R��ܜ�}����?�Gi�e�A��r��䗲�u���<�0��2���η|<��x���ru�7������V�S 9�*dX&�_l@�z�k�6E�a��1�i�&�$7u���'�J�[�+�᳑e\��K1Ŧ;����������;e�*���\������T��e�����u[�]p��`+�����;�iJbf��c<*�����&Q��l��)фGTT.����˟���Av}����ˊ�M�N6�8��\�r3�JR�6uW�tq��ɋ֭+�B�FDĥH�[(o�X4�:,���2����+wM���'+8�j5������7&TW8����u]YOu��_@�u� �����ꯊ��Y&G��+*)l�7���2�N��� ZŗM�d����9Z�lW�z5	%��I�ְ<�M�Bi2�1Eٯwȣ�� Z���֨�z�9R5
�里�%S�êD�O9�uL��u7o��7��
�k��,J���y��_p�0�hǹzؚQ���������dJ�޳Q^ꐲ����Go: T�XmT R����m��_���m�}H[T���f�.�-X��(�>k)�2'_ۏ�(M��Q:�.�i�)if*E��>D��=�P��0|�y{�co֮pf��t��L��r�zp��f@�-���w�Ԅ��1�Lw��57�*�w���n&+��To�i�
��T}vf���d�m��TkA��D�e�,��ʨ��=|k�� ��/���^Y)R�?���
���X��g��$�$ЫU֫�� ΚSL��}�@�l�ه��ˤ�:bGS���jk�"?��"
]:�;�,Qj��2�{��Co�e4!��R�9���9Iƾ� �-�0=-��J4}�@T�[��W�ag�08j<��x����&֬%�����������RU+v�V�@&��گ�c�6[?�un�f������D�d�͗����E�r�y�Oe��'��i��8BO,� �	��aa2�4!G�/C2�jO���m��0��^����O��N����IZ
�mY��}S�<�C��T���6��	�K/���,��.��J�y�5|�� �=bh\�W;S���$�^�Wi�����6��2C�,`� -@�M�"����K�)O9�Nя%m˴l��TR@|��~*���dF�׃u���d�39�0Յ0�.���bZ���%��s���u��2��H�t3#I�XKA
hy�����������d�T�	�e�w4�{��ẁ����������P��P �}�l1Q\��"�sP@��匼�U��t�0�<C|)�Ç#�����Z�/��y�g=0���b+Gr�֋@���*+dj`Q��hͪY�A�7��,
n*��\I(B����v�dwj�:k23��^���SU�-m��qRǉ�".�Ҷ����d�ռ0����窠��V:�A��16b���"��U&*�)�G�-k9f:_�ch�Qt��v_1���#���&��(�X�QSI|�~��f�Li�Fb�J�r�]�3v��v��6�k���9�k�5�8��t��ػ������=s$�iی�ext�sI��rY..|��#S��yS��¢�j�Z���M2"��'��5d�3A���qr,]�)���vv��}Ǚǥނ�n�)�.�ռ�[}�� [�Rt&��K�VӐ⬤uA7G:�a?&����F8=��M?>~��m�8Ը��.������$@>��A�Z`�]�v��@�%ƉG�����7-R�l��bQ��v�xIfB系���~�By9�PZ
��t���XN�&���"7���>#�e'��1��iA�m��f�V�4#�ص�F�Hp6�c.��&&X����NG���S��`H*�+O���N��#�4eC��y��{���z�@�J �.�۲�>�ۺ���4��Α��P�8\n<�=>e��zܣ!׋�H��?�?��A3����$�b��EPY%F��p��_�t�ܺ� �׸.-�>ͬV��W����#�W+��K2��"e�a�>E���V�طr:����v_��gbG��	L�T��Z��c_��P�����.�`%$f�>1א�l�E��L� ��^A��̶؍�N�#A4��e�����PJ�Վӵ#xr��.t6��R.t�8������L�V�i]C��a#����4�
ߓ_U�=�ƻ�� ͓��i����|C�n���^���e��k6�"�ʔ�=kht�n~�RSj�^'��K�%�D�ʧq>��V6�m9��+1tÞ��mq>�)�V3S���s�`��n��!r{�Y��@��1�5�/�M����F�%!-N�qV��@�\����C��s�a��B�� ���eo4D������19Dt�������*���	L��3"h�T

�������Z��tk<{�X��츕7P]��>��Չ>Vm����ePL�a���k
��]���X����}Z�yNK��H#���D���!Z��N|�+KsO傿4���^��O��)|��!_��0��e�&Vh�:J��P^�bۜ�2_�Q��y�´�^Bʚ���k���)\��%?��>�����y�����4��
�֥�v����v�)�/��{��x�HJ�`1;�n��o��d�}RgG9�bò�CAo;I�ob� �z�!�����G��ĪC���	�5�\���P���	�2Y5�e�P�>?���r�+�E�'�7�?�����=p+��T���/�p\U����������N�Rڻ��k�+�ф���E���A�+r���>�U%C^��j&���MI���N�rs�7�b {O>_�0��LWm�E瘝O�t�Z�����/�N����@q3���rn]	����w�}X�_g��.}K=0����!x�e`C=B���ǌ��ag�Q��l��qB��\�8�a`4K�rGw�ɕ���@x�g퓱���>d4l]+����PH��fTZ���Gv.|2���#�7��EW����po�C��E~e��=2���j{-��Wp=���A��r@ ��<���9)qM�VP)��XO�S嘷d~%�o���x8WI�ԙ�-=I�Z!_�,3!Z;�87�*�V��T,7šy��J�X�f����8��(���X2�?ŤlJv����B��A.{"ᨑV�h�g�>�ީ�ݐ+�qy}�IE��O��I��Uح�8%��V�J�G��j���N���-pxa���s�3���qo��-n�S�R�r��"*�p��Lr>n��-��
.6�՛7�ƃI�q4���oR�I Q����CK0�}��J��ti��	 [�7.�g�_�)y'�4�u�ѷiL�hd��'��1�9ץ c��[��O"����N2�ӎ����C�1E\o�����[���8e$=����d���z��|���h���Kp�m�Z��rۀ���Q��v���/�$�C���v�*��ӂ��"x*���S�N�F����,����`Ѕ�-�z+$���Uc?5*��Ȩ�i\�OF��F��ϲ��]PC�E�A��^_1�Z8쫆��j�7� ��@u�Z�iƔjh��q7�4��dE�p9ݍ�mjS�u�Ă�h?��Rp�{ �툉J��So�7�G�G�e�@I��]8��`&Q@@�<�bV��xR�l��⁔��(g0/|�� ���B�D-��`?u�d��� �*�2� �u.q[���
�.Y%�KS�)j��������5���mc���/=�|��?��T=FOq�[Ov�i��6�2(��Lg�f�{�bή��( {_C�؝$&�+���q�XSƷ��`I�۩p�|�&���mφ�"� _��������zI��Aװ�'��(��'���.��9��������H���y�R��_G�����^��3j ��b]�d�-ύ��R:�"#��E�)����r�i@��mcVQ!'ށ��q;�~aT$�`W�ٺ�͕ƨZt���&�	�ӓ'�gG^������U����*{Fn��*�yjD������G�5t�h;K0�&$��U�[�����9�m�;� �B�ظ���E�����NV��I1�zә��וp��`c}���/�ï���/`w|sڟӲ�k�0Y��b�y$H@׉I�>�����3�÷�g��& *�Q�I$H�K�:�{gi��4�j��B8���UOn����B���e���R�S�%<��U0*�L�]�E!|�u_��N�|��I��M�9M1Ȁp�zy�Fݢ�>u.m��z�՛���:���(���<�[�ӈx��5&�'\��41支Mg^R�É x����C��=���O�Kce�z�h�����Y9��~0����E��M�I5�پf�$W��H�s=D&���� �<�`�M���FL؃��m��{V���k��N�p����F}n����߷R�ר�s�˦���r	!r߲N��R���5���[���9�/qB:U�i�j�#�_1���dzf����a�u@6�WH�/ 	�����%� ]$<e2@�߃��C��4Q��%�{K���'��P���j�&���B �h\[�T:M�W1����^��ָ���7�g�F�z0K?�~�l��OFQ
Ձ�Ƿl��ڟ���tq��S}O�jc�D6V����
IJ���
NyI�lس	c�y䐠��?p	sEȞ�������c>ha�()��|���I���(��)HKC����62���]��y;rꘙ�4�s�z��Q�vx��;s�j�����.������A�x�ϔ;���mE#;�^��+H*Gc$4�V�s�X�;o�)�~9>�oB��g�[_��LX�r�?Z9x�������RG�=zWU��u����3��K���ۚ"Va���[ ��`n��۪�������oPz\��ϑڦ�b�$k����v�Hh��#����MY-�p��>j�Q�`�S���� �x�1_9�0��z�X���y�g���~�����3�,u���!��"4v#�SW�¥�C�ϥ�Ⱥ� ��"/(p�NA0�T��_� ����:7��Q�;���.��3�Wg�P����^WQ^Ѳ���N�>�B}j���Z>�2to3�l��3�y1A�m�	V�"��u�͗])�I�[�E��NߒI�}����{�x��I��5�!_�4p�%��LbL�S3�Z�0dV뱩!9��D٨��ȉKY��L��z�!�E�w��GKʜ�@Lk�aDًw�G�fnht~w4�J��Ė�����"���ZoV|A)����Ka�g�kT�؆�&�'���A�G���O�6x+���6fȗ�M>�@��O0��2���"�Qy3`��R��qXfl�s}F�'޹�6�ɻ(`q��6�C�{,�{���&���e��/�]�]���} J�M�٩^β���p�DַŔ��ٙ4�����.�?�\�敋\�.pq{���#7��ڧ	�ʢ��eLM��(���w��:|	)X=n����~�<m�	J�rK����vX��EC�=���rGc!"�oz�3��6&䦜�~J�34��
5��.k��Oɕ�8�%�~M��~~Y \����G�ݶ�b�Zȭ� ,bq�w�}���s1�6�ߢ
�!���z�#Tp�o���f�����l#����IC�y���/RO�a�Y_��kW�|tvrö����ؙS��qV�wHZ���u�a�4���hW��!��as�B������`2�%��%1<�����a��Al�6bM2#>�/򂲙�eٝ����Y��Skq�켓��������u��?�B@�O��*�&�Lҭzӆ�o��m���9���u�R�e��*��i.��Q��!t�ךֈ�r�
�qI�����$w�y��8v6p�\��������;I��ӕz�G�g�����}�V��Ә�n�ne��ߴ'��#M7��P�M�Q>`���2���J]�G�$����zGE;&8k�~�3)e_]-�-3�H{��{�ז>q�NS�j�-ΜOR첦���\�2V�nE�F1&��C+�9b�0�XMcOi�c�qP�I��S�1p�Ōf�]v�%��xh@Ye�������R2/~�̤���p}����[��B���a��*)X�DNcV���f�� =�q��l;�F͆a뉲���=�&�OD�m��葧m�
�L�c���������=�7��ų0�S�J��oQ�����3��h4��F��U�r�Ot6�����S�;���TW��<k#(������<%�m��5�߆
�R3��n(�6���'�zP�w����'�{�	h^Y��?B��x(,���W�o�I_z�܁7��.q�,���)����+0��Gq�p��X#��hv�	���Fÿ��Ag���,�؜�=�DXZ�1X��_xȥ�	�{�uv)����=4L�W��D�-|H�9oor!d��@�E d��'�.:�h� �`l�*�:1ja���s{eyTz9�#S�w`��G�E���2�?B��
��3�6`\�{��`�T�����pd���'��pM*�`�
����_ħ*��
�촞>�M0a��F)^�IEd��Hj��MT^*��ͣV��ߤhxz�<������U�K�n5$�0��VoL���8�p��{�Wu�U�^Ij$`���@�j4@Yj�=
�:��J��HC��*��>g����Y��l"�ǗL����}����ς3!�����$�Ť����*���<�8�d����5`�$�t)l�}[N�q?Si���*���!]�1�Q�4X��ͻD$�'��'.�	l����f�)�-�㰗�Q�/�ݩ�G��f�3E�-^�#"d�70 ~~��4���c���wa�u��;oq���.w��b��۝V�w"uB��D����èK�/Ͷ� ���_M̑�����	��+��G����Y�󂺤
P5餕�$�/����u�KG(�Z8��@f���םl.k�4�ӛ�����#v��΋Y�59%��@���o�`	���8V�ݿ�	_^#+�%m�z}H�+����ҋ�U:�C��.���56i�V>����c8���������\��c�fDo$�V�<��qA�=tv�M5�[V�:���}�Pq��&D ���ε����P|�т&��7ɇq�����I*Zο�K��Z>P�`d�l�
xj�6��y�k@/�?6���ht k���b��;(��JE('2��7H�����F����ϋ�Ϫ���\��v,R (L��]Z<p$�0(�9�p*4��Ȍ�".%��G�).	���J$�q�e�4R_�̕r	|}e8�k��*�����ML@�l�΄�,��#�]MY3�Ϩ\]!�P����r�|u��#O%(���(�@�£:)0�#�a3PC�{�I#�K~�7�~&�=
ǎ�+�X��� �,�Ub�l��=���jFK󗵠�p�H���s����>���1��*���3��ye}� �du
7GO���W �x݊����j˚g��"�z���?�߽�.�U=}�����gŽ��b|�j�Ь�1�v�y��A��-zc;L2C�K���-�����d�:0li��S�s���8^#�#��Q{�a��|I֐\r)��������"�ᙥk������a$n�]
�̨��������lkd� _R�R��զW�a���5��\�~{L�o����V"�G�-D	4��`ɤ��Q��B�i\�/p28�[��rH��h,�o�Φ�&�]r$4��*:��%ul�����G�82{�Ɋ�����ƾ��,��g6�>�B��U|&S������2�FfNz%�A�$Հľ��Y�~�V��`���m���?��X�Jx�|Ip��?�Q�#Q(>H��O�xQfL���y�N�B�8��(���Lf�)�S/DDt؟J�`!aCp��b�}��tR���zyAɣ��S"�g���Пem��+����Һ(� �W�`+���Y+PF�4�\p�s�5�*v:E?���j��\{��r'�?�©}��Un����1v�ݵbX�0�.��vĪ)�CPe�{��y�6
�<��ud�̂1nR�5>ǂ��<9_���e�׎h�dZA��-*�k�r�|�HtQy��{L�G,w�N���U~7��AZ���c@#%de�����"	�L��X��rr
*[���rv͵����hp:p����
_i$wb8���6�fq2��p�.f��;n5�� S �].���֗m $u���ѡ&u�OVd�>⟣S����ϲ��ې��屷��\��O��i�:q�:Ω ���;�gٚ��+�����[-���

��ۖ�pu�e.��
\���ig��ףt�Ϣ��D���m���	��A��ª pG�?;���~�W$[D�BtY��A��Kd����g��&;�׬�C�j�Ҁ$�~���<��84ܲ���M@����5S#�����YP��+�Sa�)H�t��ƚ;v���fY�K�\coW�2��.�?\0���B�#Z�w{q<���)��'�Er���Fi��7m�1Cf���]�����ن�]�x)�BjX�t"�tI�?�T�������.���y��!^C�������eb>[��U�7&����_��˷J�z���K	�(�,Ӓ�'���7zϚ�MC7��~Z�A@$@�x�p� QK�%���m�R/B����#i�I��; !��!�[/�̫����W�+#�����3�@�EES)vȤ
�cu�V&��7}�
���ǐ�M7�b�%G�6�H�,�����h.AF�v�e`�Hc}�h�o����7����2_�D�Mt;2@0����Z?U`R ��nT�͉��%�������s�
�:Ԛh��@U�VzI�]`�mKbYuD2<���h�"��4����g^-�څQ����mc��ݬ���9��ۄ����2����g�VKd�&��h���w�1<d�as�t���|��:'��ӟ��2G��]w*x�֬!%�J�-��B�{�;v�ID$Cp�������[5A��Ħ����z#��1�L;�B~�M�+�����f�'� C�.cn��Y����+��p�3�=(d�C�4���g4�QH�c:zǨ������}���~�A���\�a�u�#���ebR߀1c/=̼��r%���õb\U9��y6��§���b�D�u�o�{���GYV8~A/�D©ڤU�B�R������3����&��|�b���o7$-�_e7��׷��o��n�q>cy���E�e�Ʋ�����᣹���/`�U�?'ڐg>�-�Qp,�"Sw����MJ�ٺ�4��B� �f��폞���K=��;����������	S�r�bh�1ڜd����{!pW�;� �^k
4
�f+�����f^ƽ�s�#R�T�9'�Ya�]W"R`允
�aظ*R�c��=}�|��I���s�5��ū#՗*>�f)�S$�~������P�43J�K�$����lm���5��;.��g~
'�| �H�Gȡ���M幽޷f27��O�1W�NPf��ݾtN�����>����,ݕަԡ��������H��j�(�S�ȕ>I�3_��3/7eMx8�]��'���u�X3M���T��FifY���B�J���7S�xE���(|�u)���N�;Nl>N�U��W��{��[���V��0хM��g	E�Sc�wH��@6�ٹ짗��;���o�Tx�A�FC��@K,�2�������ڿ�]��T1��@���&��z�d�������?�^�k��3���a��h�A�T�N}`כ�p����@-9�&���5���& _������l��Isͱ�oHk��z�5Vt!�:�[jEd�p�p$��ba�E�����^&�A�Ҁ��q*Q�������T�Z�I�?=�Ź�9vc(��KG���ͤ/
?�\	<GH���)��W�oz�Dri�q�񟌯O��]qpu��)��O����)6�+[�ԕ_��8��D�$�I��95+�n�y��~�C�4ᳮ��:�����ʽR�C�?����P2#<�d���\M��}�Wi�|v"x����0��C�!��R��Y�V<c�_sw���� }�@���6F��&�#��cu�?�f�>�{a�&4$��܆ɐ�ixkQ��3�e�5aO�$F�=����:�4D��_SKˡ�C�jdƀ�%��`&-F����fku�/����q8BNE���N�S�'"�h0���uA��h��}0!������OU��'�жֳ�\ϳ������Hu��W�HI�+5s�OF������<C�a����rc׳��M�M��Dt����;cY��Ui��eŰb�6�/�o�C�<��h�96F�l'�x�A���+Zj-e/+n�	�4#��a.6zO�1�:�MȔ��恗v�]��b��b:����#�Q��Rɖ��A�J�`-!�Y{E��K��Cޤ�^���AxD��`���!a⫏hd$b�;,~���������-��N�Ck�6�s-ݹpp���P�����&6(;g�VH�Q�4`�ŭU��0�
�y�/L=Nƀ��~9�Y�ͣk3�_��@ߢј�l̊��ҮXD+f^;?�d��[�k��Mc���e��+�D�BBƊ��$iC��{Sr�"�u��3�T�����=@�o��h��>�f=j'���#oR�#2�9��?�'�+R�W|PJK+ƿ�ғ�c;�����a��Ҳ@ɔp����vl�b+sO&I���B��mX�U��$I8��	Е� B���5k/�S��B߮���}��9����a��b�2�-��0H�4�,�#��\JS`�"\g�ƅM�(ZEp�&�N����6�G��\az�Vwo$4��V���$��5	�.S��(��&]��H��%�/j�愄"5"̐���q��cݥ��ˆ����O=�����aa_~pD� �Q�>��?�����g�CQ�1=(��m�MW���𽽅�A�\l��9H�3�M�l�|�[%o�6�@~�XL.�l�\��F��~-W"��B�hG�:uO�ɒ�M��V�����qc�b�����
��^`q�H4�t��B�ۥ\a�o��ip�AC ��}��v&���C��/: ����P]�����m�ԡjB�%p�M�^��I���`>X��3�����4.�X`8��Ł� Wďp��#�B%:&_</]Ȝ��i!�Y�'�M��Ke�h��}����O��@Wb�S�F4�N��+�3ڂ\o�v�q�3��?�)ʢ��A�6�X����x�3Sʞ%`G	K��Egf"9Ժ*(�6?�>h�2׽�}�z!��Cp�F�&J���O�M=�x!s{�y�vQOER�?�
��4��V�4\l���Pxo�iM��?�}�~Ɍ���cU��켸{\�$)�;��F�3�O8��v���[�Y��]&ʛ�'L�;]�T��$���%*u�q�!���jmm����w���|s篓>��2��n㦗UTP��*�؜��Q ��֗UP��%Ե���Y�{�����qR�aD��[_:#>�h��C P�D"�� ����\a�:5� 8���3���:�^�>m�űt!�dqR�ة����/��s>;y�����m����f�_��j�kR����:K���Lk�f�u2b��IXQUyY��{% g]����
���sJj�c&h�!s�f|FB��]�9��B�h��<K����E�zۀk?���g�#�2W�]�,�Ю��q�0;��Sy�6��Bk@��-Wa�i��;��^�Z������S)Ȓl6t��G�;o$�<�)֍mX��^q� ���Q�a�ԃ�k`�m�����J�j��
_li�5{'�]<�0�^��ql�n9���1�W�Գ�E!5E���+(Jٽ��%?"��'�1iL�F��{]v�Mb�zQ�P�����!|�q~��XxIn5���ۧ�������<l���K�Ջ�<��S���=]
E��ΟJ�d�
㾏���S�G�ę�E����dځFb�^�[���U���\R�e�Um�%dGl6f�-�O%ܿ��gy�l��Y�D�|����($�mP/!TPކw UC&��O�U�%�-�4E>ni�2��y�g�Ta�`v��� �=���a2��nߘ�v*��x�D�_m�np�	T�32���T�ZM�ȑ��ݱ6aI�Y�� �K�K�T>�c@���n���W�>��p�>�b�[��-�A�L.@��L�i����O����d�q���A%��R�����f�s���n�4骬݀Z�]`'�H�3I������\0o�kĐ6c�*O1��B2��&	���N�?��1E|y.Kt����	ײs��q�k�XS0_l��F���G��<��l�<oݘK������}��A���C�g�#�B��j�r$��ؠV���o�<����T���m_��㌟x2�Q
�Mw���6L�n\'���*zW�b8ӭ��1���`g9P�����+x%�9� u��\&�y�' �����Ӡ�ƓH�	��ȗac�K�M��ĠBs h}�F'�.F���G��O�8PՌo|��j�_I��W�YS8,��j���4�1�#B j_�t�m��J@T��s+��d�SI�j�ƐZ>�_���yI�J���B�����]R;f1�z�)��V�e@HM�Y��yC�d~�mS2��u�d�?���D�k���uo萉��Hj�2�<!Vy�
�R��p��nn�#K'#���%����@�e��Vu�JH0����t[9�dӯ�w��ri)��� b��'�n�]�t�b'�iR�c}h��Cr�C�vjuw!$���v�4�:��Џ΋)�D)^��vܑ��w8#7<}j�I,�+~ە�*2I7*�Xt@��
I����b>��I{�W�O8ж�տ��k[�������(�N�*���&'; Nc�^đP�"A�Lb�r��{G�K�v����~�6M��h�?2�	خ<�6#I�!�9�v�{ɘW�=3��ǋ͂���]� ����EBpN}����'N��x��o90�a�=����R��5�uH�QAZ���1ܥ�ic�'&ۜ,�e�����pNB�F`����9t�&�&HS��J�6�&����)�����r�M>7����7RX�!4wTW�$;K��Ht��N��uz���S:�g����ZP�,	��mr?]��l�N�z�w�F�����7�3��墰������<�J�0'�l��g`gp�M蹗h��H�9z:���+�����ibv�aݼ������"�����s�B�@w���~ZN��/l"d��欰����g����%��Bn����o���d�F�D���X��Z^�83��(�ߖ��a�6�n�h(�8qM�˫h��	b&�q�B�;��a�]鶣����8}a�)ű�y������s��ា�;F�������f�^���Uƒx�X����|ty�
x3����r�<X���^Z�/`)�==���Є�������2yn���:9��&c�B�=���m��CX����{邏�e�d�=Z4��/ƥ{�6b��b�߰3J��jI����.�b�nR�:&���%�6��Ƕ̧7�9b�z���qP�ox��u�u������&#���B L���vb!�Q"<�,�S?XB����~/d�Z�t��yvZ�Fk��+����q�����t��<^JNR���*��z���sֲۇe�PKǊj	��F��RےA]�����Yu+�V:n����J���[Dd�9�_��5N,X�a�y�b���~lw����� \�)��-���p��v�K�>I���eB�F��_d��c�=1T_es�z�Ə~�V����/���xb�y$޶ӡ:�Z����R)m�m]~
�z��G�c�t��y>Ȗ���l��e��X��l!��,1��VR�
4�ٹ*�`ɖ@��4jdΰ�}�.wXN�3��� 4��ⵋ��%�.�	��� ۶#�ԁ����Ы~3��g�d�S�_/�<�o��ҐZ�"��%v�4�wsR{e�["5�S�f���*C��q�]"� 3ք|�+�P������-�` 꽆W&���/	=�p�9���mF�0���j9����h�� 6G)+@(�fx2t�OJ�H�T�����"�lG#�*k2�Tj�����AӁ�W�C�.��v��;��>�D�`�;Z��[ü�Fp,P�b���~7��ͦ��m^^:�슄�k�aϙ��n��t:F͵&.�k���3 #bc#i˲A҉zÅ�>�U��UY�J3/k���c��4D�g����9��1�V�Ti&��9�9s�r�M��r�:MAp��K�Q\���z�����L�2��JU�����v�YQ/���]E��~�g����R\h9���TW���반h��쑇���9D`9�*gC��:Ӓ��$�?�>3"��9�3A�E�#���$��&h�0A&\���Mv6:w���SX�,���'J'c8�J�����$�Z��
N�D.)��?S�� �p��=b+p�V}����܌��<�ʂ��8,̻�)~<5���!%zol�^Y�bϣ���an�&�)f(���"����!�;��1��e߶qK��+2����R�쀒,�R�^��?���T�v�����$��U6u�Y��mbʰkkV��9:�2p��e� �u�/8�
�s�s�����߉��W��x�Q7�=�He��'�FJ׌��E��V�ΪI't!'e�Jb$(�
�P��V���\�[T���圷������Ĕ{��dܐ�-;���-��X�0�#���q_�z��b��A]��o|�\�%T���)B�>H�;I��B�̧�֕��v{́�)�P����=����O8��������w��=#d6�=t�߿��M����/H��"P�j���M1�~w��^B�O;E�%������r��	$��mY���.�lh���E�nf<�%�%^a�5o��'���������suȫp�����w �!~�<b2Qyn;;��{�^�N�kG��4��]n��`�h>��6~�%���<v�b�������q�4����[�Ђ���I��v���"xc�sr$1�ѶY������'q�`�u)kA� �L�є\�%�DT��!1�Q�W�f��*nz# �̋�߱��O�|4���U�e˰)"����W�+��A{�P`!��0;�� g�!z�w��$f���[_����\��b��sY8ⶽ�L�9R�k/P�x>>��d������t북_P��odu�A�'+sfibx)s���;���&5����;p��-�����w��uU��e\�Ë�?Q��LP0q����!�m_�i�M X���QP�O�<��g�7Tdb%�}=w��g��y}��ʒ��s��f�����N<SG���7%g�*寖A@Z�U�b�Rj$�yy�
fW
�_D�{!���C�: �3݃{}w����ק��V����𣺐̧������ ZCp_�
ON�Y�m�EIB���E�c�ψ�s��6�|��U��č������VE�� Gg�`��ݏl/}���o��M���1Vz'T��Ϟ�YKc�x�dR��-H=3m y�;
rSS+���vf=M�`��WN�����ϵ��Mܻ$1@'#b1�`C��@r���\$��4�x�"�fu������ox0=�L�AyOynG;�ʎ�����gB?�E�6zy����.i���7#s���:u�[���j��FuqZF
q�Y����||���,��ڤ���*�m��}�"6	�oxrbn�m/�USN1�)^�M���N`�Plp
���s2� ����@?("�_$�b��l)�����ZEPm�Kk�A���Ј�9� =��Y�
�L�����vR�"J�U<=H49K�a��H���M��R�堁�[
�B���P���
��Z�T�ӆI�b��M��+e[��ݝ�Uo�*���f	��[b0��Qֶo�Fjg�wF�'<c�{��}���A�GKL�L�4�-;�cW�A����>zg�Z�8��:4�3\ 礐�9K�b�e��<֗P��`g���o�V��Q����� g6�\aHj����)=������֗�����%�\��:�5�@���JH/�K��˶�&�U���@I$��N�����>��p��d�W_�[����w���5x�]t�l(�����PF���H��_@�> ��&�۟�D�Z�!W-�I�)"�5�J��������e�^uY�GI~�2�fWS�Ա �|e��ω�굂���/'�B3i�-َ�T:}+b,|L=1��9w�z�]�"7e��wSfi������־&�Ǧ�OÇ�nV}O`����O*��r�;qЇ�nkIٞ�+���T�g�����_�߲]��ج��ДL����^���C{pCJ�� ^��uŖ��O�M��x�m��9��Kr_���QT,��D�۵E���$8LLS�w��.���	N��6:euԷ,V�����p
d�_�@��FG����+=���J��6�����T½�e���L��7#��h�AIl�߬ ���b�c���RB�����G�!�!�E�*E\>�髠���ֿ�����*C�_�c��c/lU���a_L��x1 S8�-���ڏ5P�?-�2s%AYح iw�`���G��c�,���]��ʔ���y��ק.V�ߞ}���K�2�j�r��� ��J�{+���L��smLs��&��u�	
W�SD���Ji���ޱ��2)� |��R���2W��2���q@_HԖL�C���!>sf"�B�с!gy��,W�	�K9I���� ��}�P҉��9���ޔb܏��ˁ��	����>��� ��=�6�i��Y�P�[���`��c��nC����C��A�c�R
x�9��vɾ����l� ���=�,�|��(��=kNK�/��e�����-�$�ZB��6�@�_�j��A��:AG������(<�p�4��9���?��(�Jn��H*�1�����e����"Ѕ_��/�&�sO3���1�hT�-b`�������}n�W������jڊ���qҥ�������ޣ+n��wo�zj�]���9��8{+��y�]�;�	�d4,ʵ������nD��6��=��<Fqg��m���h���)?ԑ��m8>2UT���ܑG�0�s)��G��\5��v6Tq�j�0�x�"�^�k3�Q,|)��4�$���.�O
,��ǀ�*z�@'ཀྵ��L����+�T��1W���e��R�b�В>���ST�����8���˜����o���%%��,��A#��f��0��Y�|s�!��}[�촍=i��"(���<l�H���Z���G����R`�������	���g��J(�9�e��ऀ�c�*��+�_�`���G�a�|p7�?��eB,C��Y��{6�Q�p�Y;�)цf��l���VAc�ZCje�'=�v�d�������+U/��gZ��-Ġ���G*�ڿ�H��*�t�����Z�<3����W/Ũ�Y��Γ���P��G�"ڐ¨S��ARn��<��맳73�q��w0�H3(���_��z����&�Nd�wǔ+�&IB{��X7��ޖH�WbT��Wa_��k}�p�qu��B�Z�l��z�װ-�z��I��U���.-�4vp3P(*;�x��X.x��U��r#�mv���UZv+8��L70?F��*���o$�o���>0G�	,��t�a���3�׶��rP��U$�M��Ao.���V�Ag�
|�Cb�a.<S	�sB��2�ƶ���E�d������k�uT���?"�[�q���r?�P��uIk�wS7��$��)Jxd��?fص�|ׇ���-Ǻ���;�Ã�QH�:��Aj�|�q`H��dr�G�&�k0xG�-�1��k��}��?�\�}�ԇ6��XĔ,�br�]@����]_��*���6���*k[�E��$�t{sv���ZP�68�g{�;�5I��2N�6��
?V����FD��Ω6<��W|n��p���|�`���s��-�8��~Z���#<~ـD�Kw����
����,��69jϼ����_oJ�h��.���ͧ��-�x��$�J?��L0	0��Ԙ4�8�����Q4�����"�'A@��DK/@�Q�U�w�q
���`�~�o��SǏ�[�N#�p���
d�u��&K�^�-��״��;�>n��l�劜��������/��5Zx1��v�(n ��o����+�P�ng�.��"��� g�r���yۇZ^���F9�A����V#X�� �K�j��}9�M7��tte��%��;9E1IV�JH�?�ӊy��偯s#"ȗO�Yioö�*���>�X�w���j{����W�q+���*$\�|5�>r�$���g��	O����p�a=Ef�p�G�_������8�e9�/j��m֩Ms��Rd-�/�Xң�i)���ZG��q������D͂�*{([#L�P��DX�N���<|R����unu�&�'Z��j݄7�4 ҅	����4��O�����M ��Njn�;up�RS����������Mg%ݟ��b3��<���t�T[���ؚ�ϒ+����̊�6�����˿�Z��Q`)ә�,�j-@���s0Tэo��IPkv��r9l��
ϊ�a$$WB�	��#4�����Q���0��W1�9S^�"x����N�m��Q��P���1ȻP��J��%�O��X�B�u�t�]��7��9d%���z t�AGξ:���C�Լ5܇�r�ޝu<_�4���*�,Ư���I�VC�,��8!��) ,����cY���0['=^l)W{���c9����D����"�u��t���69�	1�}�%.R��ǚ�؇(
t6���ሹU�<����g�f�N�o$@�;2S�KP�b�Kq�w�����V��V�h.UB̘�PI�lx|�<a&<枙s��f��39�o��F��"!J..ճ�۳�\8�P�r�ɱJ��0A�P������M���Q�A�����ɾo��o6M�B~���
Jʯ��:q?�5���<Zan��F�L�~c?�a,��8���X�^����T�Ǉ��(Č��-��hh2A�� �5�XS�q�4��:�fQ̀:���zo"w�a��2�c�$���Ii"f43������! ��?����Nǩ�ּW���K����o	vF��##Q4��T+�|y�V�,r�0����6�^ӂ��֠��r�sL���WT�#��e�!��W�EE	�%��ˬ'Y�:�;(Q���S���- H���Lr;(�C�� �#D\�ÞxuO�]!���}���+�X�G{3�IhZ�:�c�r�]Re&v8��w����z��ZC=(J4�R���{�	��9��ˏ��ԩ�%W��$��#������mI�7�p�LO�;��U�=f�;h���8�.���	LW����{��5)�W>{玬IN/���^!���J���Ӆ4O�����@r�ڣ�u+�e���X,�s�J+�)��b�A�b5���7uwY��T����ᕾ�s��Ru��I���@�.��LH�C��9'�l@T_/��'5���H�b�Z��Z�
��%d�袜�-�.������,�J:�*�Y*���h�]�بb�:�
��C�������)�hc���
��2U��[�z�Y�N��[���7�F�,�}Yf{��y�7����*~��R��W�r: V6K˳�B��j��V����V9d��:�6.rT�ՙ��5{H�Tā���OD�����PS �|>q��?Ȋ��q؏ʲI��t���`!��?P n�� �o b��8H��؇i�>k�{�2���F2x�+��P]d�ދ��3�D"l����<�x�pҿ|Hy
u�4��2FL�߽ک�$�R�B��s_ۓ?-U.^���S��:G+%�B�=�K����Y�ğ��7�vǈ<5�q�u�J����UKjc&D�봭B4~�+x����LL4Q�~K��BQ0��o������o\zb�~u�$p�W=%R�m�Td�;q�*h��l�� ��[ ���1���
Y\љ���3rl�K%�h�e?�
�5���y�W�axCW\,�B�/�i|��������]ӰΉ���a�L���C#�J���];������O1o�~�)=���W�H�b=l$ǉs*�m�BY����q�@�V�t�乜e罙ł֧�[g�`����~?_ׂ��<� ����<~Η	������T�J�[!�)��Q`�PҘ�-A�l�u3��T{+N��ȟ3*�p�:��e�|׿.Ŀ�(���jSJ��[Itp�(�U�\�闋�����l��=�dN'��-#63�� ����h�`���^;�`�7[�j����+)����EiDJM(�8jo��Bn�ji��q�S�.��FG=/��~�y�6F���p[YG�y|J�Wi�(�DUr����5����y���g
�44���u�%��!O�!��z�N�1M�-Z�ln��XP')g���J����]:�ㆼK9���sܣ�-���G��$P��Z���m�ۆ]�����Q#��*Y��iR2�a�z��]a��z��?��]�9�率�I����4x�z��Rݜ9�U��Ç̂���c��\�a!�9^���j˔V�Oe�Tx�~v��d��Q��Y�d�Y�Nw,'Bl;3Z�Y�f@ta�+@��a3e\�;��<}Z������V���5A�'F����������ˊ��?|:~d�&m2�ga�{�x�ۯYL�۸��?~���TS������sINQ&:e�&�8�pax��`k����P�k_�>�-�-��W����M�y]��U��gj�=;�K\8��'���G�/˨+��9�9�2!X��wC�L1�ʕ5�h{9R(���G���!�ϑ�K�"Gb��Ϫ;Ő�3�",�"�w��	��џ��(=�6d^6��2�JyUo���l�ܑ<�
^��B1�Y>�5��L��3e��<��j�j�i ��.�&V�� �?89@Jdk����?fz���]�SM��z�3(!8�U�OP6a�\X5�>�Ӽøj-�O�2T��J�x�g7�ʹ�g�*�2�\A�ү�sPʑ�k�E��E���z�U�j@#�,���?��|k	4��F�(�pm�H����c9�����'�)�K��JXX��uC޸8^�<�ĉ��G~��U�U}e\��Ov���c	��,��*�����uF���
)��;G±,��'��ceڏ�z�1E�pw-��&ݓ)7
��Lo��
W�DϜ	G<���]fi3��wL��n�輞�L�us���y�ts۝Ϥ��ݶoU��i]��L�Y�]Y$�jG�n.�� �&w�R�R���#r|.�����÷\X�0��g�bE�������v����� O��0T��?�ca]>W&��Ͱ;�1x�V���ﮒ��/�13��*�ok;�c�>�H���	"9�����A��I���*c�O���|�e����caWű.���߱S�`�mщ��:{����w�C�'o��V<f��7����ϑC��$Aγ�[m��%Z��H����"�+��LQ�5����O�I̼�I"<E�u��0������>�+�ŵ�>u�v��(��<��D�!|�>MZ7
���B�S��ȗ:��Y�������ȉ�N�j�tDe�|�Ͳz1�|/"^��;��Ћ�gk���B9K�����8��,���0s6�t	>��|_A	�hV�¼���7�{�����7B��:�O��'���}��5�|>�P�O_F��x���I��&�-��n�6-�v���+Q�q�;~Xx���E�u��F�����5�
5�j�NY,Hq?S�@;B_� ��x��j���ؑ���`R�Ƌ���T
J��1ލ��8i�Ej+1Z�sY��H:~�;Յ��Mr�Vv����/hJ�n�+;
�e耽��ƭ��L�	�����_����8�Ŋ�P���Y�<��2�z��*
�qAU鑱C+��$�c��ʝ�b�?ky��ͱ��ѿ�x8�?�6����uy6��t%��1Hݖ����a�R���T�O�����!SXL��'�"�s�?��Ap'5D�iB��8��+&�Rl$�I���h��S�w��@�ߛ�AbL��� �(��{���^��R�}%P�n6�An����1�[���W��tN�`�%�r������i�PR�V�Uʎ�(�A� 6���q���:�-����L�V�Av�QrKsc]D��Ģ~o�1_�0��@Lj��C��0o����z�R@T�����R���}.��G�����~��&��(3���k�0;A_ =шM<���F��f#}F�8ۆ ;��,� �s��X�5�n1�H\u�R� ��o 	X9�H�f��3���`��8;��3�����?w����X�� ��v���(nu�M� �=�C|{��<; ��7�.v�͓0��������O��e2�6pKsZL4���ȣٔ1��:Q�l�o�:�����!�(5oK�d�~F����WJ�����bI=�,#%v3�F:E�e�������"О:W��a���l����%��
N$c�+��Te!Db8B�8jS"PDqF�y�;�������T�7g̘Ì_�HP�%+�L�`�x�1&��>�&A��F_R���yRX��B<�n��{�d	?!�d;Q4y�>y	��N�i�&W��WĹ�#8ͤ"�)u��,�w�ǝ�i���G�;�(gsƷ���o�|��1!
�"��s���o�ܑ��v�-hpj#hbk����Z�
���\m^~�nP�s�EHx2Fm��Բ���yR�� 2G��L���^zs�q;���V�Sj��cK��o��#��W�0YC�e�*��a,8���W��M�8��m�x��іX2ƑU�h��D����,4v���,�)�0qi���F�3���E��w��ƗDdP��'�U.�#����6O�Dq����_�P�QnӉ�>'q&���h�1�]*��,�X<T���Ht&�mK�Z�&E
�Ӑn_Q�7rcBS��`N^��.
�y������4N�$��28E6���MdW� q/s��®&F/i��Z�m`)�H ����R�P��t�b� ���A�}U�fGӳ�kʝ5
��c��ZlyJ� ��O'o�9���t� �n���L\NOjl)1p.� �n7ns�"i�d����k��lb�׬ţX���˥�4��9��W�\)9ƻ���a����l�߄}!�1��v�XƩ)\CK��1��Ę*��&=�d?�
Q���S&�q����.�Ÿ�)���j�@��T	:l-�G�ؾ�P4hkSχLj�7<x!�/#ĐR���-��D;��j�6��	�m���Z^�c���db7뿧�\rL��;���#�8@�!`̊�����������N�;� �`��]��B�$�q>��~�ZpAs�	�e
��u@P�<����U5䯾]�Vj���s��3�u��)z����[�]��5�`OW�틜7�"���k�c�� ��y=�[� S?���>߫��f��nõDL|1t������2�&;B¤��s���+HƒA���q�3�Y�P���(Q����Q�(ԛ_=d�_�k�{�/>�-���t�O�/����5yAH�T�q��U�1��R��Ȯ��i�^o�Τ(���UYI�~,��hz��ȾO��Id-�2~�9��Y|%�۸ʲ���u��7m$f�<)h�U�͔{��5DIV��s�7�z�(�~���D1�t7�e^1Cf)` ]�E�>��đzCEu=��j3a��^�-�,���r�k��G��MS�xC��i��9��8G��W���*I�X]��j�W9���B���O��Nr/E���ݾo�I;����R�9�&'�O���?-�?Qv�/T��!�T����JQ=���U�,&���eS)<^<��)D� ��6�bI݆�A}�� ������D�߳~���<r]��j�~cN�S��
u*s ��ՒT,Z�j�uď%�QpOĜ:�{�����|�~&bo�9RH@��@�@���g8�;��pQz���P�U�j��7��s05N;���8�����+��i	G��Gk
	Rڠ����Z?���V�8���b�f��$�ga�����^Zq��]<��BO���	�����L|�b0g�dx�k(]m/LC��e�J4rs�s�wE9"�B6��Vr��ei�F���]`׺���n��t���o{��r�ժ|t��ne� �+�y�nj �)�j�u���+{�Ch��P�FW\@�;y���2�j\�.]�XȠsk(�J���-p���&�D&�{�����戒A�Z�x��C��|iapR�(OW���d�S����\�z�K,"4,n��Ν�˹3����6�>-�rIV�/���0��A����������~���G�I��ы�h,�P�NZkR�r�䯫z��0%�!݆�o��*������=��_���eƽ�nG�&{���ʍ\�V?�^��ʻI�� ��n�q���JRƨ�U33)Lu�t, ���JcԴ��Z)�O@�C�cW)��=�����6�(��:���!�?��^�(O�2�U-�請vڢ��V�{��*�K]x����6��I��l?x;�����P��6V*;��!d����\��b�w/�\~�!���*e�l��|��W[+��Df��͵F�] �l�����0���� ��W�Ǡ�>����x�ڃ��_�*�+�?���deW���3��#�Uj�*����tvp�����^�8.�e�
����Д�*��:�C�Q���M.�ZϽ�����O���Ҿ.��iT����'�_�-���i#S�6R�)�����X�'S�f6�V�rүT�?����"����j-_�d��9m���M1����o�y׀� V�3NLi�,!t�"!�8q���i���%�c�}�$��]E�\z��ۘ�ChD�Ъz�������ú�3&\K�wD05�H�C�.�[�*�O��� }]�?�>��rQO45��Ip9�Jx�4�y�^H ��+�=�]�� ��@�!�d��^�Z��S_넆��=$�uD�g��2�Po��~"�7�՗���;U�}�A�#��s�ں�]�uc~�B��9�|��+rޡͲ�F�U����E.�l5Ss���/.N���ӄR-4Y�K��Ūxo�'�2���*h�g:Ē��D��+�9�T+~w���U5^Ad-Q�%�+��ψ+hʖ&T)���\E�_��h�x<�&UK~k����ʘyg��x����Z��Y����#�����n�Q׀�2-U�����!mquG S;���/r$φ��.K�mQ�QWS@w}a�R���-� �D�btA0��n �~��K@�x���E��O�.�{%�*�Rf����ip-���^S�=�E�Ѡ ��}5��n����b%b�]�����W�Xr���b�wh=��jWs�60W���!H9�����%��}���?��ޞʏt��������Q��_`�ǡ�0��a#�\ݰ'QC��x��um�#��f篈�<b���4tT1����}��qF�ʆ)��q��i�A���y@��u޹Ε�]�-I�0�j��1ߋ�'�	w�&j���D�p�赽�O�l���ץ��̶8f�Ax��1�v5z��Y5����=_�b+��F�%z��$��FgiwA�Ι2Q-�[�_�i��F�j��5uњ��nKk�[�N�M�z�����=B_P���pBŪpC�d��G���\b~g ��n�z�������U��I΂ͪV���'wdO�{�%dl6c�B|UR�]څ����M���ls�c�׹]m��κG�7�rq1Lbr�0�������v��T��~"Nu��,�OTr�%i�>尻w�+`]�:,�q.�C4��F��2���[��*��𑔄���6��H] �)B`�7H����M	 ����i~����:H�b{��Y,&��P�3YX�J��q�+d�2��_$�N]�0�W�7�h�%��c���G���l��t#�^[ޤ���8�KNVS���Qᤂ�#Z�m�z#���A1`6��Ԋ�	�\�;g���8�e����󦺙�Ko�v�h8{��e����k,E8��W�N3��[���܈*���`-Ǉ�D^�i9����.L����'������0�~$v��(��$��U�/+��St:S�9{�P�J7I6Vהv-,,�l��u䪃�L(����f���-��l���"U1��㆖e��,LJ�/��T����P^�N�W�|�)�q
�-�^� ��Ϣ)��ԇ�J����ٗ���i��z����ެ�c^�A��F������g�s<+A&4�?�~PY�����A�B�0�c�̩�z��(�`b�H50���U�~	g,+}�9E� ��֜TB��֭����ǎ���V�Y��uA"�!��<۩j���0�1O��A����z���g��������̳�-����(Rrr������ڧ���zm�`����z�).�z�8'�F*d!{�x�y�����/Y|�2P�hX�\]�v.rz;ޮ ���3疰�۰/6��~����gFH�K�[EW�\\B�7P��9���RN[�v�H��{��7�;O]��R�4`S5�̀�$J��	=\)i$�p��2�-s�0��?��VѼd�[�����AH�:r��L�ǯjt(�YH�C�'ۙ�TgJ.t90�l���=�&!��io�E~AN�o�5�� j>���� ���6�Qw���߹RK1�*���R��~#��e���vw��h�X�{�M����+眭� W��;g�����Oxw���o�&�i�c&	���c"�~��s���O�WCjŧ	O�e��i�K���ҧr�[�zQ�\ 1u��'b`��(����9k~j�'`[��� F>5�=x)��0��S�ui��*c���T�7*�k�(3)C��ٲS3�.�C8�<������f�f��O�U�;@,,5YY
F�Ո����%3"a�>�Vc����ھJ<u��X�='Ւ�@�.�~K�M��Q�c5B��f��u�<��/�j�W*K3�f"�b!8bQ��Մm��i�������>����[���# :��N0�b�"rs򂔑��=�2+B�o�P�	?U�����xHj5㯸��w��3y�֡8�3af��d��t�Xe����ͺ�� �k�(3e�J�V�	JЈXE�M"�(~���O�5j��=��jK/���;�F�W��Ѳ;��k