��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1���e}ʲ��cg�t�ϙ�a�:�KR�%���ݧw���ȼ�B��~Eв0A�>�F(n� *��dfn�>3� �Є28�k������ �y��P�M�7ܯRZim7i�����Ӈ�FY:&�>%�º�j�\=�1��L�>����dޟ/vΘ�K��BL9��;u�EP�bx	�uc�CU�2.V���+	(���}��H�&����7���{�iq��ͺ�iB�:e���4X��n�:���aH�/]q��DV:����fl�U�(J*���F�SG�xuJ�'H#���I��Q�()؋�,�/\e�)������E�hi�&/M�@�('i���� ,���JQ�)���T*�����*��P�0u�*�ė3�҉�:i^����_��8P-�K��iy��߄##T�ʪy�HE�[�8A�*�Yq3W��G�j��C����^a�ݏ�IT�Wxw)kK���kc{�KԞ�]����g\_6~
X��-5~c	e�L�b�}y�\�����Y��|��@��ӡR���w��d��w��Cۅ�*(s���z���H�:gD��3uu8��u�L��u��ݔ� ����`$9  ����zϸ+�.�3PG���,1O�)ڜ4|k���PD˜��LDd3��j��u
f�� ��
M��eM�&���Ɔ����F���Z!d��ތ���M�\~i
����,9��ݪ�b,=�xM2S���4�Y�y��-XK�9e�o�/����~�^ތ7l��h�r�z0��U<�ſ�����5��Y�t�"����iK�C�VbtVc�F��2H��da��D�GY&�.g�K"�шM7�~Or"�%�J!2f�#��
�R��v��Ȭq.�]��^4�:��>��E�"���?�asb�3)O�Q��x�S��`�B�+����&h�����Ժ�	Hl�j��{���m�S��5�Fk�����-=��1�y�j��m��B���/� ����gfŁ�aޠ��\��A�#�;��m͒�h�˫V.���&����C3OrΞ�?Q�Ը}yj�э���U�͍�aJ7 �p���O>�9]�^�S�ā�Cg�w�������Օ��H��<��=���#hP����:X�M�WUTF���7)�)�UBK8�5�ø�鹸U:��4���f|��6������ɍ��M��љ��>a���>��U��	6!�v㶜�U�.�^��>��(��.Ϡ۾�p����d�4�~��@YZ4�f�OV|�%�b3��P���ߌ�g���MW��?��P*�c?�ɭ �JE�_c�d��D��ՠ���%.�Q4���=#�"D��l� B��)��g��~����X��������|r$,C��h�b��3 �"̕4n��%;z���A�i����Wr��e'	�R������OxG�A���QЫ��D)˦_�K<��Bb���k�i�v�F�4��9PQQ���p��{��eӋ}e.����h?9�� ��!�����#��۔�Vx���u�6�v	ߙk"GhT.�[ok'̉6����ٱN��~4)$ϊ�`=�����b'�9߄֎�u�ԫ߃㮘JI��ʥ�V�r-H||�\8�b>!�ŏ��N���d���q��`��s�1vA;fT�Kp4���ҀT�Y��Kj:AM����K'�,8�0��?�z�!˿��͛�_2��Qs�a�ڦ�%���|��<��>�_7��1J�@lF���r�Gs�BM��$_���ڨUwf�$ɗ7R�bج?#�}�W�7�r#v���I���2�t�5�a۠���&���ƙ-�OrF��;/lEd|(d�(��J$)4G˺�[�Kʎ.)�>3s@�8@>�0ݏy'���B��E�Sw��vrG��G����Q}�Nh��D�x(�&U\�Ѷ��'G׏NM�r�ч��~�,�Ѵ {G�r���D=�Da?�����)i`��{�_�V��� ��=�`�N+H&]��P�8x�j���x���˺.T��2�Bņ�؊����3k쵠W�OxE7���j�#�(���:P�Q��(�w�=�~�Vpw�7�{)�Pb�>U�7��6��â��6�D.���-Ys��w�?Z��}�Oȍ��w��"�>O�W5�+%����f2��h���>1��վ�:��2,� �
�{�f�ׅȽ�i?q��r��qU�}�3;T�KyT(���m,"
1�	�d�A�X�]�_��-��Bd���m4�v
�*?j_�tk�(At4u�@W,��LK��'���=�M�`��n����P2��z�lk~>(�O����7�D-��p��4��h'񼾹����Þ&~���j����H�o#z�P�X�)`4mX��IH=4Z�o�z ���w,�I��V�NO�ǲ>��ɾʻ���%Sh�` 7 �̙�F��&��4l���L���S�
�\���49�iS��[����\=�R����64%1T�����2�my�;��
Q��/��b��*z�E7R�(�NƜ�#s0ߣ�]Y��� 	�H������L��:�ʒRԍx}���O7V�`�L�Xh+Q틉w��k�tP[M����qK�\��V��G��Hb?��Ot��sQ�䘧W�<e�?; ��ڬ��q9F�ë8{=pT�b�0%�=�BX|Ъ<^	�`$X��M?�"������
��?U!y`�/�ʟи^S�DS�;:+t�E�9���J��8��N�J\4�+��=B�#y#����H�ہ�J�b|��:������������_;����4N�j�G�d��D�by��,�m@s1XK�|�� ��ּ�C+>�>���Ԛװ�0ܩ���ҹ�A�� (BD�!��j<p\8��ѭ�n��޾�>F�`Z浐o,j��ve\��g+��A�R
���8�n�#�i�pu
���,��PW�s�B;��1��ӫG,J�����>0{�1�N�!����|��"ʬ[uL���-���W�Y��4��;粒J�+s]��iT�&8�J�=�&�^��d��C�G5�A�%�RUs.�X�f��4�3�&"�7�#]k����ۡ����ΑZDFޡ" � U�OZL�('�p�����B��/���	�۝�6��DJi�aV�N��ȩ�J�����9\�/Y�%����j��A%�uz�D����Kҡܟ���p��tVK*�6UF_-�!^�zu������(?x��ko�1X$���=T� !�^�k�n�%�K�i��
!,��~Xqn�6 ��溇���Ky?��|�n�^g��V�����#�����%��N*����C���Y��_��o	��dl����ɯJ\�!y��<=��ȍkfX^Q�Rhzn�,�u_��gîۖ�ug}<�;���=�a16��}ZA��0�tI��*Tj=�%��g	�:1����O�?�/݀�g�7pOn�s����ֲe��zq�,nGO%FғQ��G}���Sm��
B��p���S|�^s)���Ή�^s��F>��ڋ�.`��%�?��8f����(p�v	��	��G�a��cA�J���WlV�0.;�p��0�J�'�=CX������Qr��8�MzCo��Euq|C8��;i���uA:�y��}���*Gh4ẘ$��k��.����<j��G�-�v��� p�l� �A!�f���ƾ�M&����Zό��m%9[b�F0�=��M��qg�,@]��A����_,�8}�o2ӱ��V���tT{�R܂�i�dm��W�j/�"�)ҳc�5m'ݝd:ƁV)!p���:`��c�28r+��� ���u�P�|�r8�㼫�%��j�h
�%oUR�O�w��+��~[�m��ժ\mzG��D=��il�t�S����=*7����ޛ�.^�MY$]rVk#L���7�����"���!&���W��d�	jA�������@�vwc;��̚H����
�����˭\�5Zx�n���b��H��E����&�!C��\n��4��Tzn"�8��΍�	8Y�,� ϩ���19����q��7��w X�d�Wy��z���x����֒�Wp� *�r��(�Tj�QS��t=�#��Eڿ T6����! ٻs���_ 2��!�#=��(o�W�
 ��/ʸ�4q'��32�a|�(1�J��j��J��^e��4�Tvf��p��w���^�����E�����R�y�8�X�$�ރ��� <.G`�7��V���4��p8�r��H�f�k�Y��1ۜ��t|&�W�4r����%���O��>�I
�����*��c����ǧ�F�vp��1Vy�# h�16Id���0��i�60�,��Y!TO1J�]
��˂��\��8檮��Ƞ�\c�2������O�h�����01��Ū�|�\��ퟞi6Я������n� m��ډCeE[Ū@�R����uB�m!��K�K<��?a��� ����~2�/";I�c�'�Z�W"��b-"��<z8w�����]��bl}b�=˞�鉡z����[��O@�#���^�:6���ڲ��^�ř��Ӷ˯��	IQz��(#����E�D��&i����>ƿԯf䣖�O��� /��6��֟`c��������;�P�T� R3�H�P#�1!2��P�񓊱4�j�_/�ն������q�6��� DE��xѤ�R���a����AO>GU�<���6�n��VS�=�Yx����/��'ෲ�fg\�CU+����J{=h�� Q٬|i�׎ը/��ٜ���E�i��>'H�LgSW;�����RQ�)ĩҢT`��Ȼd[wc�8������w_G��1 �Z�G�!�l�T�_XwH=����*�S'r:А��x��ؖ�wJ��~Sn�.����g|�������.
�J�k��wlOO9�'�ѭ1�4QI�	� �n$rQBH�i���}��M���r����]Z�>Ϊ ��%94�$��y��t%�@��-E�Ƞ�S��S�kw��ѐi���c�?�j2�d1pT	D �8����h�`u��W�5i��u� �>&2�/����Y����T<D�u�lF����(��3_X��@�Vo�XXM)�W��N�sA.W�A)~+����Vw�52��kYHq���:(Ao�sg���[��y|v��m~$e�o�|�'"�A���0�?��nz1}��L��
��w|G�7���bёF<�OP��7�/>��rO�c߱#hU��P��ֲyRJg<���� ��[���Sn����0W� ��+kS��ݔ�P��ARv"}�������������E��y�]������GW��@�D���ds��"\���^�/U�W�'�I(,���Yg�VB���X��2�x��Ġ�kw7E�W��֮ڮ�
+>��/<g7]�x\H��F�C��n�/~�H���$��o�G�G��j���n0����T��%1}9׌�w�Y�<ͅ��Xf�����m���!RY��-S�Xx5������a����/I��<*���"�C�����]9wC �ٲb�'iw�1W7��9�����bK�tP�2p(���WUm�A �
I�N��>�A�V_a�bj���3 C��=lS�
�A�U��c'�}�A1���L���������n��{��S�>�C�C�M�$��3*��1u롃Z^����X�|��<�����e�/���f:��A$S�V��j�!qȳ�	�U�W��79���k^�rQL+��MS"z2ﻒЬ=��9��Z��[�l�c�/t�Wj����Ef��\2�ϙ̊iM����%7R���+�,�m��~o{�˞=�u)��#n!�g�k��(濚�PL��,h�r�$﹅���]��/
�;[�4�	��f�l������!��9r�Y��e��F5���0����4bƽL	�~�u�}8K�U��)@�z���`_|�V�"6��=y�NC�����taScQ���n?��U�=e&W�qf��\�@}��h�k�8/�I\1-&?9�*�DU�,E�r�Xp��#��kMٙ���-'>�u/��Mص�^���\W������$��&��M��=� �
�Ӫ�rPQ5�46��c��$)�
�@|���#9�+u�wDe�v���H��ĄG���jM�5�k%W&̥},��^�U��"z����x�������^����:7��H�)�����Vff��I,h�Y���Nh��S���f��ôlC�Q�+��Z���Bg�� ��E���.75��f��0�GW�o�(�0p��ϘŅ�<g=�'�@=����l���8�X���I�!q%�D��F���1 ��A>��Q|�;�bc��I!����w�jB��)�F��2���ڟ��v��Q���xc����uӻ��Λb&�{�(�Wܡ,���k�Gi���=2w�DcҷU`�)��ua��H��}�_ K���u�#��xS��3������܇f߲INK
�^�	�ն-�'�-���2[��P�l>�I�T�so�߂ՙ�)|�Ax.�����0�J�����v��� P:���s.(�s#� ��zzm�lnW�,���^�,91�_*)��#w�&(�.� �~�rGD���3�P6�	���8�oWЍ�_�e�)#�h�>\�L��m����ؒ��R�� Έ�k	�6Ϋy����d��Kv �Yt�rXr�.��(�� �y��c�V���9@nb.8b.�t�M�'Y��{��z���5a��cAy'��~M������ñ��Լ���	��_7�~���J9�15	s5�z7��^/$��@SK��8� �0K|��Xz�B�4��|�g�oCd)�#�gɞқz�y�~/.٩���..��@aƢ���vzS������a|��uz��C[&j��5"�-^T�����2���$�K��OT~5N�i�`]���>�ֺX��ָ��tL7�~"�H��E�oႵW�&�26$|�$,[����F��G����&Ҷґ�m3�� ��/J���e^��Q!����kЂ�@�@���!yoW"8�h[�eo���|#lxّ߽^̡Bm9ҸP�%M!B^w��A���A����_x��c>h�rz+Fޚ�w�`}SZ0 |�#j�G�Jw��o�O�wޣ!k���!�C�
5Od,��\�Wm&����0-�Ӥ;�-@?��.W䳙�\J�ʲc�^�ז�st?��?걆�K�P��*bh�����ʟ����(Εs6;o�?9���ё������pǠ5�#��B1�Q	&0�k2Ar�ХQ���<��@�A_C)lHƶq՗T��A��{��&�U8`.�v��F�)��@�i�'%�1s����}Qy��~�C,HU�jM8���W�O)��\ؾ���)�VOK�\�k%b�R�&� ����̯�N֝	6Q��;�?�������p�C����?���2�<~���C`A��n�<j΄#��� �X�XC�W�I:��_D6SL��m�♦�.�\�d�N�V�.d����˯3k(�o�X52�����hPr�]\5solc���ī��召����B��\^�$����_��Ԛa��:+�.*���T��༺˯��~$�S.n�x�V���T�Ƕ3���<�$ #<��Vz��b�Aj���W���W�L)�����^GƄ������X�zH��S�>��W���nۑh�x�!��w�&^��]��u~�r_p>�l�����	����c_s�p���@��Хh�����>��O�u]T�P�8����A�h�?�IN6;fR`��6��	�*�UP��]��z���?��^�L\ym�:#���������R���I��8Ŕ��B\�E�X���l���U!����#�P�Nv_���]lm�����&|4;)�!#Tp��K�	��,�֬���J!n���H��2��@�T�*(����7��=���m3[�� �� �8 �Q<!O7�x/*�.�V�Ј����"���U��G&|����_"���5�<4��F.\U�����]���C�cT¿���y��I6�
��`��U.C|W��أ�c��lƫ�T�,Xyw\�\2W�����+u���j"�����$E΀O�42R�&`��8�FO78�Y;�{߱�0�&}%20qZ���%
ˠ��g�P[�~�����X��z
�6c���2ym.�_�T���H�`�ޒg��ţ���A�<"K��T��(2*�I]C�=��2��hT��cQ>,M.�_�5�?�D�����"#��(N� |�'�1��,a�H����[��o��sH��@������+`]�z�8���PP=��`�N|�V(�z�w�Q��s{���Z)o�w���̶�Q��=�X���5�S�FKvf_֮�;��պ��Y��8�<7
z%��}��*
{���s��)��?�"V87�)N��Iy#4ǀ�Mv&�j~p`�"Uh��ڡ�3��{��q��a{��o�#f*޻t���gi3X��2�)jR���c8�+�ao���x����p�G�jV��࢝:R����m�_FO���y�_���ZG.\Z̓�W�I��XX\t��:��[/rw��\�H�>���;D�P	���V^S'�(:���"�~B�,�qZ�e�h��J�j�Ԋe�k&���ܾu���fҷ��|����Z)?���;��?H�	H�o��P��r0�����hKww�u;G@-�O��7J=�)r� ?���u�%�´�v\p���ɇ;��*��uٚ��s�[�������\ٿ�<޲h�۞A{�F�h�mc?�X�����ͅ�6����A8_M��w!���c}�b�{��B�@��ί]J"�����Gi��T�Ig���f:W-f�1s�Ne��-���`�� ��S=~���z\��]�Z�$>�un�a�w�͵=����J�#i�3��/r��\D�,�#%$�}�I:3>Ϥ:[��xa9�}�G�Y`��֮zx"d��ӭGbn^�!�+�pF��x�Da^�~��s�O�����m�x�#]���Ȟ,��|c����n��������)��>p�4�c!J����W�)l�4a�βS2�b#���>���D��ӳ���@t׌�8�%
��r�W#rXn��{�6O8|��Y�L�U�-Uvh�|Fg7o�N���N=*�+M$���dHr�-Q23�Pɞ�^��R��
��5��O��" 	s���l�cwTZ�ǘ��8��A�Ү+�A	������%�r��(��-��;m��ќ9�[e�.�M�~^U�� �v�7��4kG6�ݛ�B�YEL�:�cm�sE�h�SX^�j�M�%V҅�Z?�dz�9��z�e�H(���v�W��3��I�_i�q� �����*�ʒK��n4��4�Y������m �GV���<h3݆�.EW9�ʡ�]	[w�ٟ1���s�*z���5V���X�S�y����eQ�R��"-�����p��~�T�ڽ�%(�������/���{���q�>��m�Q(=u~��1��*f���t��b�=G$��Ey��Z=/�G�_��� ��b7�m�ʐ��7�G	�
����lޒ�`"/
�wA�끺�����AI�(�����B�Y�E#H�Zoc�d���b�J����x+��A8�A� xr����{!�=��_��{sV�Ŧ�ѽS��G�����Z��1��B3�z��(���w�l�z��v���bX��"3
(�/TL>�a�P�p-���z���u��}ͪt�T(��ܻ��Z}�Ҹv���RTEv*��h^��C2HW�F���G���ԍ�﹦��U��ii(.mqq�'����s9a��d��h�9����^�t�F� �������>Xa������Ld z��<��d���7�\�A��"H���^r��ʡ�i=�o����#n�k[?~�L�Fq�b&�OL���l-�ީ>xy�>7��p:��VK8��e]*�R%��L��T�q
�G��(�B��4,N�<�3a�a|ܙr���?���яA���?:;,��E�E��I����䌧���۬��g�>��z�yË�:u�^~�5)NYRb���2�޸�/�p�.��z��%��礃������_wp���m���T6��z'�2p�u9�����zԩ�������Cw4ʥ�fv[4��V���U�����,����[t� ��Qhd&��H����_ Op���O4;ŲT\WxPe��&�f��:Sq�ь+F�*������yE*/-.X���~Xv�杤����u?��.��١_#��g��1�5BC�j�O	5�W���&����#bW�Bz�d��ظ�O�'�d�j��j�VM^�R��ث��kd���ʣ��"��w�1�3	(*%��p��š3
�C��߇ر\��Ū�_�w`�(%a��'�|}��KHѲ-�s�z���[ޖB+�d�൬oMu_���UL��r?��_�E���2^�/�,C��/�u��:&�}���K����#�]�����o��1g\��i���^fq@q���~)��i1�B��+$�cY�~h	�� ��^xUߝs!~�q�xL	/�G�2U�QC���Z�I��OUO]��� ��(��C�jra\�
9VCƱq�ۣ��wp/�&m3}9��!�i탡4��%g�!6U�((��@��LG�5�� ����+l�H"�
<��+h�cƟ3X���:9��Z;\�q��O���
Bfs۞r'3�
Y�*j� B��p�c���h�'�mv%�~S��; ,ƅ�������Y��*qFiR��Z�ra҅�OP�ՈINh�3{�A����="su��������g�x���"X{�<�,�1�}�E��I|ئ�>�if=@���m�G�s�w;);]��������(,�F��{WY��lS�N��z�(�駭��i����=.�8OqT���`�)�+8�E ��D���]�	��j�D�<gE��gZ�L^��W���CZ�����3x��ؤ��_\��X93cgC�Qz�J�a���ۻr��)��e�/��V���m��S*I@l�A/���`�1ċ�ҥ���@�l���G��9ȉD<���'L��<�'��]|��>( X?*Y�g$�m��8���� bݿse�_�?w��7;d�fm�K�d��>GFO�ڧ��HF�4�? ��3�%ȁv�O+�!s���CS�����a,(��6����\�4bK�J�˲�I�*_n�%w��y�U�rj�}���w��b����Dx�e���p��ZS���Ih��!V8s��[�6�����~�����H �M�0���}앒L�T�<�Ĭ�_��bt��g#�� W�Ҏ�J�M�o��.�<K��ؤ����]{���5P��5���p�r$�wB���ዮ�M�awfx��蛹��1A���,"0��Q=,Y�m�r�g԰uJ8	B�����0 ��wIq^)�b(����������f_W�k�lSB�w�	��m��=t���N��
x��8#��:�{hs�t���t�8?�_{�QW-�F.?�JNb�]���"2~)樤�o�N8��y�A�j�0y�����FcF-z@�;y�_P�0r���bOh��WgŨB)X��C�����0 �U G\
�»����uMYy�B!�/�S���
���
ᦥq]f��@�];�c�����'��:i���))6�U�?�h�@.�\� ��by��apOY@�#;s�&����o�͐e�k�v�������w�\Z�rR���Q�� �o�P��Z2հ�P�F?�:���Urn��{���P�8�H�5����0���p�Z,��V򗱌�瑱'����މ������6��j�1	�+����/Xv�M��!q���Nl^��;z��nO"�󲱇&�z��d���ɊFW�2��������W{���x�n@3NUm/6����� ŀY����C|�Ġw������4C�,��g�G��r�@���ИO=⪑c��N�R���݇ꄳ��ۺ� �),b��O���&�s\2�����B�_�4�T3�dd�����5/�(�͵��/��)�Kd��a���E������k�)�ډ}E2�����Z�i6Ƴ��FU9��z�^/����o�ݧ�Ꞑ���d%�/��z�j�L`�k>�E�@�  �p����yӦ!��n�_�㣕��g��F;:�+7���ô)���⟺�{�g��d���O�l3t���N!����sC�CiCJ������-�2J��8_�g��@���3*^�J�����U����D�}6S�n@Q��/.����4�9��MPk�f�N��~����m���ʨ2
_�Gˆ��ǎ����=<��;'����8@"��)0�t�"��h\��|�#� o�⭡���x��LǸ�b3�Ǥ��x��=��0��8J��8f��l�k�\�G�i����R�t�
����=J���ÿF|��\�Ud<z�QV��XI0I��Z���'��R6��U�]ע�G����9|�+�������-u�B�.��Y �[�[��)��7�a���{�Bz��d�郞��Ā�u��Ua�k�KKݸù��?~O���Q��Z�7zx���<m�0�����|~�Z��`��c`%���Y�,?��V=�E��ګZ�ęi��}�)yY��f��  +��H�_J�<�3�nY'��&>>��4�ڈ��t�a88������B��PV�Fʹ]نE�[��ps�v�5���^&��C����6�	���6qDf��],S_u�r����G��ޭ��]���+)2y�М?j]�V�y�����`MԙS��o��6��c�j"Qg�BF��������?�Ė�ԗT��5�8�(D�bBϼ���[7nS�m=��]e�i��LH_�@��;{#��_t��_��aBy<L�1e`��B*o���p-j�DU� �!�*�N��D�-���͕�p}��Ab�^��H`'dzr��I���s4܊�vI~ סn���]��Z宨�fϧ��,*��!���ױR�/HUF�� NL���(h-䧜��6N���X�٭�)?��A�^�ѣ���L�Z��E(�P*Y�Y蹵7@3�p[��!It�Y��w�Z��MM97 �۵��>�Ͼ�J����&���FFU������i�%|�����z���h�_��U�2��'u(�Z[ů0̗��;�����㯴��[�9�eH��	����~��)f*����A�D�܇�]�0�u��"00d�P�-M|伱ԑkx}���`!�6��E7+���\� Pn�,��V7=k�\?w ���#J3�Ob.T~�i>j�{�D�����FBЈ(�_\�1��H�Y��k���Xx3�~;스�vP뤮�AqFx�i��$
s��E��CL�m.3��j�*�o�)t�w�G�]���p��V
TѸ�/��U"��x� ׽�x�1�U(���N|����K~\UJAl��p��x�4@�1ơk܎�i�N��>�E��^�9+�u �b�� #�d�ϓ�%�{�ME���8U��`����Kqi$لz�����,�W���yN�B��%~�Hj��m7 ��.�vى��/F�@	�~��tTv�Ƽ�����φcx����\���Dq�6�^-����(�=�j�]L�C@�˲�)��aՙVxL�l��S�-u�&�W\�Д�w�� _|���$/�E js�΋�ϭ,�4��4y�2����ϫ��z��b�&���>��A�qD7�� #T*��Acvk�,g Ѥ���e�%���Zd7�L�_}T���`�>!��]4C�QG&/j����#f���&�if5��,�����z�{G ��	��=�P�dp���L�z\��>8O
 ��su����}�*M����}v��w�N���!�G�	ǻ�*��y'�[�n�@9|A�����*�N��v��4���G�5����y�v��c����!��'���-�Q�4�Rc)����+C���F%��5�����eRԠ�D��������P��P����H�Y�틈)�+�턾���>�1~�4���4o�%�O�0��Κ��aX�Qt�[�)����B�������k��Zo�㐵�s7���i��ͻ���񨌴]�@I;r�%s�A���;X*֜��={�O"4@�G]0w+����BY�r�,��T�r�DJHmI��.���+>�r'P3v�	� �^
��l'<[����=����ۼS~�#ȨR2�o��� e��Ѓ
�S����ב��W�@\����~|
�P��`���BR~������Pv]���q���cJ��+���e�ZO���m��kѵ!R(�p�n��7E��3�O��:�>��xN,�f/��L���4P���k]2�bB/?��}D���/	=�Cw$f�^��C�FR�3��S>(�?i���Rg��}�;����A�ȇƣ" �}��J>�{?K6r��;
����h��޶��({��Z1N8�aK�����Maa��}V�j0T�囹L��ڽF��\�Fe�2�iĹ�N�]݈ ���������꼗��Io}Ԩ�����	��^��@��W�l�C�"�F+ ƞ�i�>�S ��|gW/�zV!K��n�Q���u��8D�;�5�xf5U0�A1�;�_�����`^�N��~���?uOݾjm�E ��*��W�n������4��Ŭ���=]fkw��~�Z������l\B�<,$:��+��`���cQ|?���w�����}s��  B�k	_en9�A�޻�G
���*�o�\a7f����T��i����I� �s}T���(�u�/�پzy�|h�w��]���5}���b N�{q�����(5g� ��P�Ʌ�N�,����p:�����bc��h
K�>�x�r��.\�&���ƍ��A�OX:���s7���s��3[ 2���_�&FH�g��YN ����ys$��' �T����e�?<!��W��4@I7AO�A$Q���[��&6�c�D:`�5hs�E�4�2g�/��21P�}��ZT*��l��:
{m?m0�
����e巼H˱�7���� �H�Ԑ&
b/Q�� �ǟ�,��B��X�jZ�ń��š~}�^��g���0������B��e9mߗ(!q��
�����6u.�8���i7ۮ�w�\��uu���&�N�p+�~��6�G�x��~�wvQ^a�̕~�떲�`� 4E+��=*d��VS�,D�-���#/��$��m��v��}Nd���Dłcw��5����zϦ�S�[Ml%}�6�~��Y �㔢V;�q⠅��K��싕��3sDl���8ڿ�n�ғ��o�ʬ�6AX��&�#
�,j����C����\a�`G#w�Y��Tϋ�o sP�!���Cw$�C|[h���Œ�tN\��H,1H�����_Uf����B25�c�J-��� �TQ�c��	�|إ�t*�P7���<{]vC\��̮6��0�,�@{�;)�=��8��q4�gT`�S8$:��֛�P! �V5�����fE�|����g���eB�$��mV�>#�'�$�Z[�ޟ旒��[����f�bqFD` �0�y�.H��m
~@�Z�#rp��̂�dd�t`H���,M��|(.���.�H�lx�`.����ģ�Pa��E �'Ϲ-P	�"�O3�C@ъ����H~i����\M�u������|�!��
�̅!�:��'τy`���7�bB�p����梁� W�b�>.���}_$���o���b'�����`��R�/�%�3��OxԿ�W�&�φ���񕗣�TrK�����:�1���deX-2�"v��jӎ��d�Ӯnf	��7"E�%Q��xW5*N@�W*^���C�� 2��UQ��}���~ź ��P�E#���N_�rNW���}�e��-2J�qP`S �]p0F'�xQ���Mv��&�([���%�¹�M��Ӌ��ɣ�	�k߯��!���U�^��t�a�S?��U������3��+K��;������^������z��9?`^�'I��"x���ng69/f餣��A]+v�Ǹc����#��H����X�着k��@��OU��!k�r�$�d�����P�l~�1��Ծt�D<@Z�_0�)U�X/z�bM�mJ�;�/婤�[���D_�� ��[x#H8q�_�γ��8��TK��Ĭ��tIȄ7��,�܁ �Ev�0:�b���34n@i��/[|bT����MбaC`�<��k�sw�¤�me�;�T�;���"�'�D2_��Yj�� <ʮ<b];Ո�f���ش����� ���C5]H*�HoA{@t4��y�wF)�T�\k��y�K/-�G0�ƞ&Dw4�oP���DPȘ�4H���)����V������{�@�x�,��Fp���N���f�C�A<��2ޔ����v��9mW`[q��f�܊w��dHB�R̋�A��R6dZ |h�2���̗MD�*��ܟ8��\��e�0rl�
�D��(����t�s(g>���Jm�.���I��mԶI�h�8�����o�N���b]��6g77L��N~�N��y6��w"�f�ў9LPt��)z2�\���x�,�1��l|�)��;����,p%�xaB�c�mI���1��u���u`5P�8�Z���7��x7�QC�l���\9�K�Y�ĽB��Ǧ����f�^�Y�����$�ot��kY#ke�ӊ����Z�v>@�r�b�P�<n�2���Q]�q�_����gy�y�z2��Ii�z��bl�b�L=Ϊ��ݖ�נ ���cH��@��;�8�������+W� D	;A���m?6���~�����q���m��&F 1I�C�]U�/1�"�`���Eq�q~~����<�t��6�^�V\�`m��w�m��bC6�ܬ����Q���I���{t(%IB��9Մ�a�����b�zoO`��1�(�n�����5:���8v1��b��U����4[Y�G`n���:k
����@9?�]?�S�%}�ͯ�����'L���!yS�;8%)+($��#����^��.sN7�ٵ���jV�G'
E����`��tU/����T�9�����җ�rCO�o���¹�읲I���/ ����ݮ�X�E�v�Դ�0��x4	���T�PwB 5O>˵��R�,�?N��	O�)���R�7�Z��eȈ��c�������[8����*�\:L6����t�` ��M��Lɴi/����I��B��3�n�$_|��I���X�i��͚N7�Y�6 &�H�'Ld�1���\Qt��^ɼ�g�=&�jxP8�n���<��Q>�0�`��xp�Բk�_91�H,1K���bjs�ʭ�"�Ld>�~ g�%�:"y/(q��k�nG�Y����*�4����K�0�7[��ȅ����r�����Yimi=�n��ğ��F�w���d����M��*�������p�!|�nՅtKTJ�A�P#z�>�7Ll�m��%K���UAa9&�Y�9ےD�?�v�������y]"9����k�F`@f��K�z5�KO.L��s�
��ҫ:������O���2UB��P��mm�1�A/�zѺK�.b'�{��U�
���2�����o�\�fUj/{~R�7��HLG<q=_j��q��4�������3�����[H����J��Q���:lu��~	�t�SB?h�C!l6�Np��+B�g��3�� /�X߆�Ns�;�gw�u腺��ъ5�~Q�0Tkӯ��M�ħ0e�g�*�<I��c��jV>4�rl�1dD&TA9Eb�HѾ��C���T�`�����-��h칶��uK(GO�yR�!1�#��a�kɅ���])[�Ř6���6%����y��b!dE9�:�����U��/Z�Gz�w۷ɦJڤ� ^"p����̿\J�J[����N�U���4���6� �=����C8��x�?��hYn�D;G/�c��G��E�6�o�*+���T�. �Ou?�[�dR�Jh��X��)�_�_J��7b��,�X�5<4�c}}����sI4YS-5w���T�M��ʳc��ڲ�����Tx�1��4��t�h�` %���7h��_��M
(���N���ݦ_˛����&N�-�.���P���'����7���vО�������G,X[����k�W�M����Dt��Y�����t[����*��\�����w����<<�'(qg����5~#�Lڞ��Ɂ�ЄF3��*���Qcj�MB�^rI|� 
�y��@6[D潔a�0���� 9%ȴE)X�(Լ4�
�N�<n�?ՌE�� ��&ynB�*�&G0�����`+b���%�<e��J�&T���0��p���������`�2d��f\��`���Q�y6��GȖK��C�xD���������P*�.���
��9����
����s�K�#ݛ7�=�C��-�ĵ2�H
��^V�#ka(E*�ξI���7�w�T�Q�]�fƥb��mυ�'�!��BT���zu�s��(;)�p]�Q�A�qw%!�,���q��-����ݒtJw�� �� �L�	��ۉ��1��� dQ�S=�A�5D� ���T�_tL�״�M�13R��r���,�;�e��GĂ��W���=�l.��WE4�^�lc
���.�b�d�sHNL6��������N��N'D9��E�-4UV�>�R�ɒ�L�e��?i�ɭ�.EMt�$nu�	�O�jR�/�<w�h��D���X-u>=	o^K�Y�+^�N��2l>8�z�,�A�A���c�TyN�YU֣�S7�Џr��L(�>^KϞ�o�;q r�|'��`�������㋋��I�p�9Q�smDnYg�?R+{0��8i��?j��i��j�{�R>� �|$`�%Mܘ4����l�g��z��z�zӋ�d��hC�M{�~]�:Ϗ��p`���hdC�T��mG�]o���C�9�_�r�V�o���Zl��ד���?>��!�^@"�r�ӗh�e����Jv�A�T�"��ܚ`}�	�|q�4Uݰ:�:0�<���g��LA��ؖ~�U��wԲ2�8����^c�P��^4��J6u$�.��(q_��X˄��4iHE�d\��S�E��i2F������2k����!%����ľ8m�3��!n���v7�E�H^��c�}y���&ȵ�x��\�U����C�_��<�:���@m��a�_�W��	H��h�&VV�PY�c�f����� �TO��k+������7����w��nA���v]3��B`�Nl���BQ �3[^v
��F|�\�[8?���Ek�w�P���m��ߖ�Zp�`�DO+� O	�U\78�=$4�/�>����{y{�R��=5s'��A$\ܒdNGҎz�ef!�T�A�љ՟7�f=M�ӵ��'��jrtc�4��I�(=¼�f:����ߴ2�5y�V��iٽ�\��~�mǢ@���p�]⤾�O�g�>"9M��ey$'þ�j��B��"�����nh/�Es]�$b�{���C���V�,�Zk��`*�mi�l�;~�����nV�K5B���K���~�@a�"͊�A�V��2�HV%Ly �.8��c���D� �Bg㣮��``��@3���P��h٧CE�>�@@�1�(���W��^f�|�����$+�9�~0�+J�:�D�K�)ˆ@�ʴ�~��/�p�e��͠0�F���~��U=:R`�[v��'iS��D˃.���˄��Y@�v���T��zK������@ ��o*V2Ҝ���C�=8��ny˹vCƛH�$5�;�;3�^�ک��waqg)�Ā��&������.�����%b(0��}��ɉ��:����Ψ�y��A�]���b�3�b�u���o��.*O7�IRB [��)����
�GY��jhZi�\7Uo	��B�M�\[�פ�?g(*��ٍ��9 �i�,���0��u��FR�����A�Y<Fc��.�m+��}L��(�P`��5�mD���3h�����-�u�~��x�19Sr8zhy���Ou����Oʁ�`nM���n�^�9@��`��2\��E[�G� �2��>��/8�䧮��ĳ���U}6E�7y��/_wP���b�tV�����LJ~C�>��D���� z�p'�
ԍVQ�Yۚ�����>ٵ�����x�O]��n{�<a�U:���}P"�Bdw�>K������j�ԝo�܀���و��]7��p#�;���_���hf���
�v�dԘC�P$~��/^,K�Sn�Ȓ��=wx�ފ�(6��}�8�T_ �Di�����7����K<��]G�DǢ�-���>8j6B8f�L2�����s::�8a�^3��U��={Vr��CT�	o^��,�<�`l ��6��R��D��n�N;��j�ی��1�����7�ʴ�6r���!Cd�<*Ӱ�G�+����6!�t�zR�������|�ܙ�,�l��M?r��^��k����j��$?�u69������FC��S���w�	{�}�h�*�@�oc��,Љ����U��ѓLPf�v�Q�P���<�R��[6%~m"��Ā`x�+VOc1�X���Mv͈B�H�i����(�B���?W��-L������h�k<�ӂ�f���w%�]:ʟF�Z�|S��y0�h��
��k�Qv~V��Le�[-�"I�6�`� 0M\�\�P�À�>\�y�P��6yW��i"⁨ްJH3o	��I���j��C�+K�^���߁���t���qp���}e�p�<	�2���K
��J{'�F�b2RW<^�|�j�7�"�QKMg1�������H.��zʳ0���ؐ����9�`��2�o�'P;�x
B{���פd0�1�?k�4Tx�[YPG�\es*��u�3s�!Ք׳0�R�4�b�0���<\no��qD)ֺ������5�];����a��ʃ�U)s�	`�%�J2�wFjd>�S�#�V�靃u�(J�>=��+����1�̣{y�e VpS�$>�dx�Oe��+j�5����o�(���Y;��rO�H��j�;��1�����F�E�	�h�3To�s���_
<`}��N�C�1<��Odcɛ�ҿwhn}
jf1��V��F��Kb� ���wAvQ��Jv9܋�1�N�n���Q���yV��F�[T/:�����/+A9���,MD����� �M� ��Lm-�1����)UNЪqU�H�Y^c��������\@��C���!��ZF�b��(��gߐPZ���T��Q";CG0��{��o�����fXsk��?ө������=9VB��Q4��IVZ~�{i\j%�Ò��ɶ<դKFm\��'����.�Kc^����~+2�O����B�>ȁ4��V���
de�imY�i���}��B��Y�,胑��x)�����n���+��H���ӹҧ�M�__���hͣF	gh�n\��F�Zi��lgO���L}O��(Hx���9ן��I��VZ��X��)Jw i� ��|�V,��s�Ӈe�}��{fC2�39R�����r�o��i������@Y���F7&L���������N�Ƴ��Y�&FfH)ƅ1����I#c�G�Z��K���%��\4!�8QF�����M������bP����f���A�{'bҗˑ3�D��v�Ȓ�ʖ}o��Ȭ�yd�-"����#�f��&�3{��\�t�0���H&���aփv�ԝ�T!w傕3we-��q+.6WO8xipZ )Kr�y�-[�zϔB�h-׉�̙
Ky 1����?|�z�a*�4�R���~�c���v�e�	#A��4��c.�r�[Yl���W�M`��F ��q�*_�s4��C}?1#����� w���TR�r~E{�Z�@K�x�N%�L���I)T��-K_��� ��3T���l-�!�6]dM��X�j4Z����E�k��G�C%��V���M\Y��5�X7D5吽�Q��uϳ��v����<-zݔ?�R�KҰ�?���,rdog޷Ugj clU_߁6�>��>8c���%i� j��;j�<T����j�c�B��E��cQ��J~�칡*'�����8D�l����?��Nl֥��ul�����\"}��ԡ�����{@q�ù��$玊[@��NPP�y�&`��Xl�hv����c�w��/�:ڞt�Ɔ�}r򈄅�*��1�H����G�e�J\EH�hjC��%c.e��s�нmK�U�(K�p"����f����9��� �P\8���h�kvh��^�����J����������lH'�N#�����hWB�5���6�v�,�����4�7cK-��g=�w|5����k3��Fۉ���Qn��J���N~ݫ��{t��%�m�^�.2�4���Vum2(����"�f{b}jkb�JiT�U�5v����<�D�z�Z ��X�jK>恨�e�|�M�R�x0�',x�k�v����1ѷm=�c��c�tsTG���x�LH8�GK0�)��a��SG/���1�$�.��#��Ѓ�� iPY٠��b���q%�����$L�Zǒ��� ������[xL�-��Vo�I��9�ַ�4!�%��ʡN��Ox�3s�(͠��66�k(6t�P���WX��b��J�"�Y}�p.�ڧ�-�H��s�M��p�]����sv�U���Ύ�1�G��"(�4��B��E��iw�)�Bw+-�+ϵ�^M��i����L`X�XDg�j�~�e������-�hW�݁U���sŋ����1����^�n�( g���� I��Lׁ�|4�=���X����]�o#4� ��{��r��x��ރ�Lq���5ƞ��^�}��mn!�uP���[�S�o'��'Uc%�\��ā�"����{��΄���q@K�7�8��p�:��a�M娮v��u�N�H�U�-�`t 3%����gX/3��a�'s����������v;v�)(`4�gA<T����|*�{��䔂I�	�G�[��x�V �	�����t����+�:')�u&dA�Zh��h�-ub��bֿ�ל\0���,��.��]��/x���ݘP�ߡkY]�ˠ����Bɀ��էEF��_�����:��m�����&xbؐys2�U�G�=~f;x�=�A:^��1��E�d>�`$ ���C���m���ߣ�1�5ղqw�޲C겘O�J�bYj�Z3��',=uF%f�=tY� µ�Q�	��4um�� ��NV2 wp��;_�x�]�&��|���OT�
��ղ�M�%r�ƶ#������W
&��Q��}����6�MP�x�	�Zr��݂�U+U`��нB�!9�5�/"uwnN.�:
���1�W�T(xt�]|#��,y-�/��=����]���O*R�jJL)=��fC�B�c�0H��=�{�q�V��Yz�R�J��8\��\���]<j��4��zlMy��V��[���:M�xv���gD�\*�<��� dJPZ���>���o{Ҧ�h�U��#2����^���FT�N`�c
nY7� �N��N<̀j�t-	�ug񫕻���8?۽7H����QL
Iw����znS@� K���i-'����z�� ���P!�	fe��7��Az�[��Xx�f�m;�F��n$�tS��(�MB�	78g�0��!�T�)j���6������-dy&mު�i�� �0�0�W��QeAA/�5{=5էqǟ�ee�FT�ЌX )5O��伖^��G�.��-���6�6�2��I���)VJ�������!��2����%d��:O�.���?Ă����_�)*`ƚ�h�<CdO��w�9( �n1�L�N�^^���m�j��!���~��!x���٨�Vc	�Q��mېx�zeE}��)!�{\�uL��S�"DW7Xs
zP
E�"
+��j*��ܵc�'�V�b��-��D�K<$/��ᖩ����q�S���b����H kXNG�(�ƥ��j_�ʻ6���֕h��iJ+��{��],[����:T}����c��u5�f�i��b���:�-��n��g��-81���sk����Da6zLHO���?J� `a��9���Js	��������)O"�"�Wp_u���L���6t�	&J�xWJ�^� .��s~�c��Dџ�-U��5���#m|Kc����Шu��H͸�K��&f�;{����P����x �n$#x%u:�M],?I~~����� m����O�O��Gb�� `}���Ox���l�'Hz/'h���k�[�9a��iN��{雌>��O��}� �&6*KWX� nJ!�f��:d�l�C���F���ʹb{��J0�V���yr�=wыX�����:�;-Yإ�]�24�
1sc�,�T���9����k�N��M�Z�wS5V��vry}^����4����	�ĉ�_5:5�^ś�b�Mh���2�f��$�����v�����ǀh��'<(`؇j�t��E^��\��0�k2�x)z���L��P�~�.��y��6M��&�c��j���	�?��|�T�ؘ �
URTUo�!�=f��b��b���ڸD*ҍ��NN]�#��눂�Õ*��j��Q��$(���2����q{���ϝqS�9�:Ո���V�#rg�o���Y��~n �
?j���n�hү����<�\!�d���)�p�����3x��twM�"ł6�T� �j6tɸ_W�^�w?��V>J�����9��YVD�QA��]�##;[��Y	c�Ă��É��q���Qw�F�M���Æ8鵴t�W'zꡓ����,)[n���+��о�R����)�s��k搈īE*�2��uc �y8��.)JޠY�c��2��rR��e-���3��Ҳ�r��PW��t�O��d߷�f�*�F�LB.rŸ����H O�.P,�l9��U����t1ܽ�����e� ͕�Z4���
�I�V�@g�0���z�׵�֌��%��p0�RD�Κ�v���:�CJ��ɻ^�j��l�OV-!=���H�S
MXK1ϼ)h8i��h��x/0���AO�[!.!� O���U,��;1�'���k@��4y�Gw8�a�d��JjSHH�2��$��������K&a>�:4�%���ПY�[�}��IHf�B�}��m�Ӭ �lH}��ܰ���~:������6P�w]���&TG�z��s8>1�;� [��M�{�)L
Q�U�Bo�T��O�9~֋zrǚ�yH6�N�+f�g���192����>Z�O����"#��z��#V�6����f�r�i�g��<�F{��_�D�x���%f	��=ER�5�P���$�d���P>&��o�M]_�e�.v�
_k�I�؈7`�(U���4���=~�����������T�7���e�V�x��Ȣ��y�foF�R�S�#V1#c���g��s~ �`�����Nߖ֎u���$��B��tB�������$T'8\��/eMK}.z�!�}�3pi)��ǧ	p5�� qЧ� �.�>����t��;����<��M���W��Ƌ�hf?q6��b���|O�xHb>���N�.��[���ރ�p��D_hx��u	�����T3%�yt"ğ%�2:��y����WE�\�(�bq�[U���,Z31]Z��]<���ѫ9��0�8�S�Ϳ\2�����mXhlLO���d5��]h��_�J����;NѴ���=��;@:���HdhX��U'�1��,v���Q����ĝ�
^:~���F���1o�<f&�׬>Ru %�Ƴ���e:2�F�{�;f�o@����ZV��B�U{Tn��`�(0�����u�p��0� d�S�;�� X��y�N�Ԩaa���D�X�z|�0"`D����hͤ�1\T�m��9p��#AVQl�ͫ�O�h>��*/e��FL3���'�ļ�[D�i�d�	���w�!�_#?+��gm��o 2���uw��Q��&5�>Kh�Nm����Ps�Y�T���-
����iR���)B8�_�Č w(q��^�e����CP+p/���oJ�rH�fِ�pM��2� N�G��4���m@��I ��o����ڛ�с�_/�^Mb88�g�or	n�ha�_��!��`���,�q�mw��� wX��Ə�,Dj3��P�.Um���b���cyaNO�˲%���O7�U]�..]�䙍(�&�;q�a��D��LF?L�:�\롡�6�>M���avC�o����LW�.�K��f�
�0�ĳI�H��ڨ
ź	J��*̋8��V���`r�(�[\c���4�2���T	�m�o���,{�Yi��ޯ^��*L�k�F�Dz�x�Bv��/qh7���9�A`���:2�H�s���<�IwE��M*h����8v����@����Us���'��B�(Ў��r�3eN9�ޒ��c�}ZW�|i%��/S����m��$�l=�DD��|o OI�r��S���6/ᷛ;�Y��.d����=�3>��` �'e��_��L��z�h#�fz���a~rMa�5�=������V@AdH_R�,��} S>����Q���L����:�_����C�e~�*���<�M����I�C)x�'&1�L�����"��g�ut<��}ē�g����"�߰��Yxn�A��G�5����]M0��fˬ�z%����t4(�UEqK��j$����e@9���Í��VE�ߏ��=A(��#	�4�[�ON���ۮ��"�G��n�J��21`��O�hcU�;���	�,����8S��S�x]���kBdh_d���6�5U� s��i�^_�5_� ��q��clW�%s�Dyйf�mx�}j#i��|X����Slt��{�0=���H�����w�ɣ�V�;��F����x�y��!�\�)��T�Φ҄�����5&Ҙ߈�VNc�%�U���TE����Dƌ0+�Q+F���O�}4���'=,�S��e�;$�#'�9���Zw�E����]�%]��^#���2�%�jEA�qb�m�b����]@ó�M������3]M�]���GCh@ƥ�#�mU���I���ni%���%qx%��H���Ҡ��Q%.�, 	bcb�Ψ8�����L!uӁI���o��l�5m�S+���77��3UTc���/���3�9(��}"㡵��ߪ�a8>C�>`d��)�c~���rP�?��+ �JoF���y�sǁ�0B_kt�1��׋ǆ?�t0�a)��X������FA<�����G��kuHUӶ7�����c�γ��\�Hrd����x�7�R hW���be%q2����\�ʶ�|�x�2��®��J+*$$T�/`�(���دD*leb����ȇ��_;���Â7��Wϯީ��9��C���b1o5�9a�0������#���(y�T�d�)8��)�~�8G_rۡ����J�$-���|����`�c��h㕌a,�D�o\�MNeX�n>Y��$Hׁ�d��UV`�H��az}C0�6�6>�����w������ʂ�q=��#g�󔍏�\��c�����g)�0�����fLL`&G�Q-TH� �ڈ#F�ޘ5���{i��\|��A!N����ʖr��!��}�N7՘��TС��
��L��X� ]�w��Fi���,�gV4b�3�?�T%c�.��2@�� �-WY؟���9�y^"�;����um:q*��n�i���Ku�u�W\�0pYˑd������f('�w P�>ew��ļ�9�?n%	P�J�{��W�1�!g,)@�z~�������q�"�B�d����V��?@���y�����m��'�Woc�U�_�a��H�П(���}�����	~��=���g�� �X�Z��d�"�ox�%����9]�p�.'���ɍ�蕎�-�6'V�|ؚ�e���ai�F���F�8ً' a�XgL�x�d��Ȧ�^���+��G�s9M���~��F����j)M ���׫X�f����z���0�q�4�=/�PE���ZB>Aq�+�@�a��K����>��w�;�<���ږ�����> ڼ#	��� IUX��cjO�J!���λ7��$ೆ������uB;��A��e
E��_CjW�ل⊃-�װo^Y��ყ79�0��5� � �i�e}0�Vx���1co�7�?���(d�c��4���,S�L�?�j�:78�30S�$�"N���?���f N&O!����gt\U�4N�������P�0���)%�z�T�rP�1)NĦM02�J'y��N��R����1Q����@�P������B-QUb�����+)�E"��q�F~�[!�Bل����y�\ ��F	���Wfx�,$�l���Z�� '"L�5��q���R���"F�',�Ɍ]�Y����|Ec������P�3���R���c�
d^+�Z>B�$R0Bi�.��ZxiY���Bh2�K<����bM2>��Mi@[� ��.��w�%�{���%�?����_�Ҧv��/�A��o�	�ʻI_�&�D�vr�d���&t͙���b��;n�N�e=�'��>B }��+��)��l��@ ܅�"m��n������	����듊C���f ?'�&o�^w�lʛ����Rq��7���K�����jW�rt:sB���I��/�I}y�e�ی�C; ��Y�?	3'���ѥ��H��.D�;�HW�w�V���9��˘��쟬<obc�/S�b��&�'�W���n5?rɺU�8���ܽ'P�&���u[�=Ti;�6N^�k�qWz�u��6�wd	�0��J]�V�6qH$�a����H�F|r�Q�9���~���?�M 2���%�QR�`���[�P�t�rԩ?��@�2`��$������j.�I���%4m� �j��Vb0���l��B��d+��-�Q��s�/t�W�"�N%o��8+͘}z~�Q��@^�g*rWff���Pa`��n^��.r�׮G�c� ~H�빂'6'�n�� qLb�#�TE����t��/U�΢8�+�`$� K ��d�&D��5���"�<�;aQ8q)zD��w��8&݅�c�4o���]���������\�"�8{�L>Qʍ�h����`2�AӧM>2�ֻ�iK�"KʕHb��Ч#�	�d�\�U�YM�U�T��R��Q���u6�|�-c�G��R��2Ƨ0��ASE'ao����g���s��a
'Q.oT�Og��#��Z9���ѡ��)��ӜX����8L��� <�ӧ J����#�I�c����$�'���K���	Z�I��#F��'�6�|Y�Du*(�~[T�n��J�F�� ��,l�CIjJ�s�b��g:s��ܲ��L�ti��ژ4�Yh���O=MU�ݾ.��D�q�HFF�]85�©�6A�~�"Y���j�l���㰭n��5��k�A��CK�BB�X�9��M�Z9���bT�5tق���\0������8���q���#���ѝ�ª���|��sC�?@EQGDoYY��1�-�7�8����2��S4�yS���X�y~�l�:��=��J��r��X�)���%�[GR|�
Xī�UX|n�U&9P��t��DA�;�(�!{G���x/�2m�nPF��y�Q7 sŻ�,��fb����/ߒ�݃�(�uh�[Ԯ��4jr���r��xs}�
��a��2H��4�>��E���t ����3pr���77�d���0�q�6��W����sځ_\r�T&hӚ��������:`��s<�A�S:���Ȋ�>���(a}�I}[	��Eנ߼�u��}q�Q!�j&lJ��R �]�4'�[��H܌���:����cT�O��l��i�W�,r�w��-��eL��1 7��q�Q��I�l;��7�h\f�堲n��'���^'v���V�ŧ�IK��ǁCwlL �_�V��L�W�^�nz/����e���������&�p7O��ɴ�Paq�;Fȵ�a�o]��֮��2�@�,�8cۜ&���y�~�
����ؼ��<D[Yʉ��<Jh<9�&������]Ԡ�ZR.�l�V�u)U]<�g�$cŉ�{{����Гw������
R2!�BȒ�|��TԽL�<%p�b�Ž��l��+۲N��ZJ�}�`�V��Za�+TC��:�*�8؀&{��{
6��\��v�W䲖'�y6��|a���v�/@q��H��B*̯�c��9G6S�?/1��6ŝ<2pA�iA�2!�7.9ݼ���@���x� �@���#��vr�_�J+��Ӳ=�Z9ȹx��.F�_,գ��oa��7����8�>�Z��ؓZ�B0*���%`���Y�T{V��uY�q��r'%A��rv�@8��� �/ ��v����WGl����h��?hk�0W>�{�q�C�(���[%���#��t�X���	�_���TQ���?���E�N���c�ȥ��Yn����ֲ��*�w,p�gV�V���&�n����,�s��ۚL9=Ooq�	���C1N�|�D�׬�労A"��i�������](�^�|&�IecpoR2�-��F��P�y
X%e��8�}@�rƫ9>�{��[�2��t��;��G�4�/�����6����x�sg�Z/o��\� ��$}"���M���&GS���l���
U�Ҿp��<
<SGv~������=2z��J�F�+�27�=���o/)#AI����Ώ�I��(�N�(2�RA�zT':ӈMf��b}�`�����J
��o]t�j+��=���*@br\����k�!���_�}w���['u��j�>/sSj�X����yI}��1����z^CW�qnIG�,�H�q0M�ҙN�֗�Ũ�T�GZ��=� ��b"6�^�T�F0N�k����HM����X��!a�.�c���،L-����</9u6�k��G ��a���rV%���֭�U�ڰ,��=�����TH9)�f��e�$
�v�rq)�(�B.���N?� F��ؾ�f�%`�ڞ���g0+s��D�{ŉ����>U�M�6�Ǧ��l��Ս9�	��Si�ɍy��|�qM���+߹�|�Rк���$=e!V����"T~��4w�.Y&S}�	i�{l	��ֵ�)��y�:����q/�@#�]Nn{`���ɷ;�I9�>��"����X��u�����|A�=�*��z|�r�$A�<�/�������SN� �}��A��SJ(J���xUyy�\�q�ca$G���V�*A����� E�Ff(�Ώ�P�����8�w�Bաż!��Ә8��]�4YQ�3��Π�A�"OwY8,nڭ�V����ͅ�����l0��X����a�s�+1N/c�`�Ud�V��<���w��1�"���G��N`\{@y�T�R;*@{' �\�#z���S��ľ���H/B&�����k�c�/c�܈�����D��w�9�rQ!:0Ȳ �k��.?h��$|�uL^'>eyW��0['�K�:�������~������R�F�Ř�y��s�ľaw�G�͇˕�/HM�](��Iܟ�NrT��P���5�繂B��nl��R�*��o�v0�q�
k@-7d�͋{c6����(u�����5�$:ϵ˄��9�f�L���h��c�ɜ΃�$r��B5(�|�F��#!L}��JY��n]Ok����]�����i�Ԥ��C�)ـ�w�}�|�	���#�47�h�-��~E:_�g���:U~������Z��#'��ڈz`.��K��W��0u��T�t"��{�˟�x�Ӂ��[�3\��}�k�o������m���K>�h�	��`��~�P��]ԓAܱ�h~�3&�,�����`9���.�?��ц��yE^�BJ��>>�i[ぱ���qn��2�EVJ2��k����)/�4)bf2�Hh�u�@R�m}����jgm�a\�,^uId�j�#s��`T�u���WR;���I� �{2����
o���5�:�8#`o�DA��'���#�+(�6Ǿ�	ʪl�O�'[����Q`D���>���v�(�n�LTwv:�2�4���'��^����\gA����k��G�RW|�.4�'�b,�8,���&�{J��u S��EZXB��)9�#�e3���A�[Yi���� �*��k=�GO�s�f�Ů���c�wPЩ�&�7dT�w�W��	��6����M�})�1V`[cj�[���R�Va瞕��J�[Q�l�\�������?�B��G�c�ёb)�Y���:�����@��
@�#�Ď�I�D�H�q	V�)E��I�Vșv*������o)ߕ'��%k�;$a���0�k}�?�W#P���EO-܄���Żp���?_�B}�)��i��T��@5�uT��?�W��a;"�B�r���3��~Aq�a�m��jj��S�$Q^w��� 0E�f"������q&`�W�ZҔ?`�y̋ʝ��5��F��֟?:��3jK�2̈́��0�]N,��ym��h��z�	���0�L�xEs�*|7*$�C�Z��W����N�� ��³��#���0|���9�M��B +fյi�,��S�	��
4�N�Q&�����LJ3���h	��|�|0i$�"���ї>��
LJM��A���C�V�������)I��r�k�̖t���z=���?�V�0�Ŀ��k�J��~��2QK����n|����~z2P�b�@C ���0
�.�%�ۖ7,Zk$J���:N����O�S� �WBv�]v�a�q �j�j�Gi�
u���c��Oo�6�����2�?fKC�"��V�w���2�1G������-T���
p�Fg��)w▬��l8|(9�-y@8"ͽ�f�78��.��Y���w�%�'��$�Պx*U4ۈ���%��c�5�+5�C'PИőG&���M���bI��c�I�S�qT��c\�tߗ���I۝/X�1�'�څB�*Cqv�g���)N�GW� W�S4�7��a��U2k�U�.DEW\�k�,W-��,�^+b/b��L��O/P�j��3_1臋;�Sd Iηzy%5=�4���u//�f�+���f�V/�������)��L�9\�OEW�a�z�Χ��^g�0�z�+�6�)�Y
e�M��[w�`�a�"���A/� �
�h���>�4�>o�7�/I-�vh�N��4'�\�"�j� H�~�+�B���D�2A�J��jߪu�-�0D�x��� �W�P�u��F��5�l��U+�_����]�gW�J����%g�|C��;�z��M��ޫ���Gq�<�۵�%��zP�y��S���9�-�Ky��������/�w��8��~_!m�u�z�Y�K���:R�x��G�1MV��� �Qr]�y	��K��`l�h�F4���	!p�3��n|!/a�+��m�$G
��v�m���|mfP?�1�U��~0����9X&4q�ݛ�e��?�Di-��R�St��k`�g1���*?���:�+��J�0�6~m�
��eۊ�V$�[�N~~�u�%bQ��y�R���2P�#Y�:��a��k'���Ѥ||u�H<�H�㷳s+q��ӳ�ܓ�:Q�"]�<N��	Y���>Tv�>A.��d�sڄ0 hP�fFE$Eg.桚�/�ڞ���]�Ls�����7��n6����IOs��*���^O�gģ�Y������['F�1Ma�)���tn؄�_<w�������Gt�Q�"L�y{��`'�Fƾ��<~g�f���䛲��djN��.w4LK������Ws�E���g�a�&�YW������8^��s��Zp�2nN��|؍��V��ߍ�ְ'>o�d��9���A�e¦�������Y����kw�H�_�w<H�瘔N��e_�DH�5+mV�ua��y���`_�pxG�������w��;�m;��ՊO:�Ł��:PBL�"��՟� \Vd�ՙ$l%�}�G`v�a>kƦ�K��q�����.��\�[7��i����:)�����W:���1�E�4Y������d��Ҕ�ۈ������M�Rr>n����es'�'� ��-�����|�z¿ώ��。 k<�-PH%X[��N���g�hp�cZ7��h���]9�G����7id %%�І#x��2v�Q�f��06�x��w���L�{�	��s4��G?��ƈ!�{H咒tթ#����F�C
֏�����mV����� Q�� z"���k9b�ȍ��v�ן�=$�Ah"`��S�U�6�Q�E�9Ny�i���Ti;t�/���ר6��S��,��M��
��{�;TMK=��s��%��M�-���ɽoræ�[~����X1"��V�	y�����i	��W�r�.���̓���(bഄL׸R��쩅̔^ �D v�� r����w�Kʫk@ץ S8�oF�	 /����K�7��c�̕�t�A�Pz�) cR��Zc���"��r�Ƞ���7�?��C��`�xӾ�~�C���t����=*I�om��ެE��+�k<��/�98�Q��/;�)��3�3��ؚioڌI�v�%'[*�F� J����C�e���#e��p�	�]��e!9C�w+3�'�z���ư����Q�׏F��9����r���˄@�����3[�����"C�t�l��@�T���X��G K��0�f���j� Q�����W(��z���k��"%&v����6'��qŁivSQ=9謵k
W�77\>x��fs���O�c��_EV4G��P�Q��������k�M�\[|4��0��Cb�
�6=����Qg_Yk���t�D$����8Dk����;�������& }0�}�t�h4��F���+:ncr��mϲ`�0���Ra7��+�؄mY����"�Σ�Q��^�C(w4�׍�Уdr�5Wz��{ �Fb_����%�C]!N�B�0�AF=s$��	O�5�ʾSeOr�E`=��^�@��&	�<KHl*��"�T5�M1�Z��}����
9;��l���h
��i���:Y��Cʭ�Ü�N.<���d�{��*0J�,k�R��=�l�\��>�4�{����'�C����e�"?����{��w8d����C��F�S�ð��w�\X+�Νv_��:�e�]
��B0Ĭ 
��M:E�TJ�#�o�*�wuX�o��mC,�����^<�Ԧ[=9����C��;=]����S�m_ AC�	�%��v��D
�϶/߻�T|_WT|GńW�P�&��TLa�
�lZ�/m�ٗv:g
Y	�1�H�s�`�s��È]��?���ZDfxՄ��Y�4<?�� �!R�������>��+]K��-xW�W����b�p$����r[��_��h���e� �8�E�H6�Ȏ˒���Q8�+�i6�ZS̟a����4꣉A�gg=o�v��Q'���`T\�0��Ɋ�|O9����
��2��C�*��׋�zs	l��"�˴�n�1"���v���g`�|��7ݕ�?X@�3��>:^���ϳ;� CfV�B���R�+��̃��$X6-�x�b���h�Ś�iC�R=�僩�%]���H� �=�l3|3��q�þ�SWq���Kb[	���M��uG=��|�L��>0�#	�4��=
�:]��}L��&gM�dRӘ�T��[�{�en��#F��TK�xھ��г���fB��8�<��Vj"uǶ(*�d�a���ą�ڷK[�B��� �D�]���Z��;�sP�+.�6ߧ�؈N0tEvF�b,�8'��0�{�vk��Wء��jV�x�M&��T�È�t��oq}�\5��������m*î0ɒB�7k��4�D�L�m�������ئ	-,���h�FC�9b��sFPF�0��?�~u(���f�_�DjӾ�V10o��]�$O2�x,�������ڮ��l�8�6�fͪ�ˑ����!�H攣�G����?�Vt\����@%���~�S$���p��h�/����r]�`��)r�^bI���y|c�Ι��=��tp��հZq���yS�o2��%	��#��ͧ�7�!���*�^�2Yi�l�;І]LC���4/󄫡be�0�8�!z�ܶ� �1nWu�m����iG��@�ߠY���:���;��=�E����%��1m��O-�a�*�w����b\V��: ��������|i��F��$��b%V���*p��Y�I�!Ω]�v*v�V�*r4j�Ά'�7ؿ���Q�A<��l�x�n�t���%�J��]�}+��M��x���{�YP�}6B1�{�`$��^e?��׸ڣD�W�AJC�Q7�x/��c4~�W��t�w.`�p:���N�)�-}�A2�kd^q9Z@�p�a�N�$x���;u���L2��ќ.k# _)^�{�\��u�n:J�c��\ALJ@������kk�A{�����$֧�Iq���6V��w4��[��Gow�/��UTzX��-�7��袤��� ���O��R���E->k�5#+�USք#=�{FE�I=o�Nk�Ѣ���F�5�6�Ed���ܿ˩��b̫�X��n!�l���i���x;x2ۭm:��
%��($���r?�@J4�:ƻQ��ԂA�+�h���fl���߳����T�{�wO����p#*=Vr<�Op\��Crv��+�v���)I�=,w�FuI_]M `$a�kt�/ۈ�
��̅��;�I��R����[���$�b�H� �X�BMwP��"� �����Q�@����8I+����2�E"9���S�g#J���`�n-�ѨЮV���<��6��N!m3�]DYf
��g"�~�D�!���* ��xuh�~-6U�ɳ b�d��\ֳ�R��6*�X�G?L�#1��T�������?'������x�DgONo�"��.�m���0&������z�W7;3�mԥ�z��K׏~S�6B���P�O_�%p}�����rb~���'7(6(B�i���S����#A�Υ0�����Y���X9�'"V�����`��X8�m�f���6�v����lGְ��n�H��Ƭ;v��|�@��j�}�ɿ��90
oc	�|bl�eS=9�~#�溁\���D>!� �?-�8gz�Q�W�_-��k���� ����}8�=}^����V��r��/�$�G}��#�&���P�n�1z�cI[
u'�:]sPD��g��I���"�`�k�Yﳰ����<�a��C#[?�����񟊋`z�j4��ZW�]���y����u
�������z�;K���7�)g��3<r""��3G*,���$t��á��8�&b0�)�P�ۗj�M
e��0Mih�+"A1�|:W�p���nJ�@��:ު������Hf(7ç�)kY���`b1u%��@i��X#Co
{�2��\��
IN:-���ՠ�{�����$Ց0Woٱ������
!�<����� �g�^�>����/�(�nz��y'T�P�5^h���f�[�:�^����o�>��YHv��OKc�Ȉ��w{;���駹��-���W��J)�\��af`�R�ћ�_l�eQ?�*g�B���������Ɨ:\օ'���%3!��Q�V���m�|�wI�҆�u�T �����
�RX "���"�%��?��32x�3�`*����m<HZj5�~A��I3�-7�x�U.٣�'O݉��3U�=m_G��L*�bΤ4e*KQ�,9�)�������鸻[���!N�q Vз`#R�	�-ӝ�kA([H~�*2����d�x"��'V���P�T��ˊTalt�O�è��G�F)��S��IȰ?��vt�������΢^�{ߙ�-!�A*�Kj6v��h�L��>a.���g�����p�X<<ZB��	�7K�aB}D�05)��+Ϥ��!L�-_}��m))�_��������{c� )�E
Ӑ�_��;���\��oF������jFqcҍ�x.MZ�9�B��	ov>���oe,*nI��Qc�\toy��#>�PQ�qp�J$���"���E�?�c�^͟T0c�����⇖g8���r}�~��˅�%b�JH�L��R�p'�vj�z��/��fP�g���aې����a���!��{��y���H1]��r*��>W=M����<=�K80)��8U([��ɒ�g:^ݲEa���U��(��,Ƈ�tZՉ凾��t���ݪΒ`/��~@W�Ǔ�(�Ř�1N߫E��f�5f�����0�q벀7���g�/��3��U��؟5bB�y�7 �Hzw��W��⳴w֐&5=�P!i��t@_܅��#���wd��Qf��GU�0ģ��Û�n�G"�P�Ei�x���<�#��[�7�h>DoaMvl�y^?���=	.Uh�����u��olo�i������~�4K��^�6�C+�#���;}�{4����<�j�<�m�ʢS��r�=�������������2n�-���Gq��)m�L����{.�&�V��� �8��p�`��(O�ن"�:��n�4��50�2˩$}��K���U�[�<p�5���sU&�Md�y�M�ED��x��[B�v����)�e}ȗ�56�ˎ&:�	�L��&�������!#+U��"�d�-����e�QW�'I1�=���X2pK��oŰ���=�T�V�^Ǭ_�`���P������**���H���JO=��� `ӱ�F]�q"4,�9.���K'��[ĊKFm�әfD,�N�.�Q��$�_���i&��R����ԣD7�Џ_���Q`�4�D�
��4R��&�P�<��@`�HJ���HP�������8�4�@傭~s��n�^��:ж�}T:]ˮՉj[I)oh�W�2-������t�N�"�[�$;��6�����,s���m�����hu0�q(ȓ�7ݰ�2k��gF���{����1��'��L N��~� ��լ�Zf á%��I��np)�����D��>��[5�PWB���N4���9�����_�B=\m���)���ů(uˁ��������G�l6��A����Kh
�@�L��R�p)d�K0*�#�z�K>���r�Қ-�iG�C�q^�ѶG�گ��R�*�D�8��S-�vڣ�E��xl]���XCϭ�CUs����8����ʡ��@jJ�ѽ�c;\��� ~yd�CE`20���Tl�xl$�7��́@��th�Ou�t�~9���^W�������o�dSmT�R��45��-a ��,�k���T�������c�P���D�x����'�Z���A��ߋE%	H�C���r&m$�ҳx��ؿd�%�V�f~��&_����� �v��V1ZsBt���Qĸ�(�5��	��ei�)E0�-
�@��3�d|0gu������@�kJ\�t_]ڞ�`e���q#��Kz7��+Ģ<MT�ޞǷ�מ��\�F��t���z��6�6���1.e��8�4��������$̱������O�g�pk��$�T_f��?.�����al��YT�CU�+y�B|yx��fa
E��GW~P!7��^��Q۫̈XVH�������2�Yɮ8rP�����	X�w��B@��r��QFSuȼ��qe�=�k��9�%�*bf�Y|�i�����;�Pȃ~$��Ӵ#�'���#M��#ѦJ�+�L��vPBb��<���m�J}�C�Vs軘V��t$����DR`�f���ӵ�FsB���||�ͱő��x�����6�a��yc>t����-9e� ��U̼��
^.���tn�:�w�K,�1m� ɩs�t@^g�,Cl��o�2����1��O������?R�N�N$��ch/���@���\�M�A�%AOg��{`��&�4�l�-~�ܕ$��Y�|�"�-M�q�/�ޤv����t��0R-��w��)��"�,Zw2ہ�������Y���	�Ș��t����Qߪ���+q
�S?�-���I��ܞ�|�E Nm�7ԏ�]ډ#�HU�z��X�v�������f��sR�9b�́��ԥ������}H1�o��_g���{:�K��Y���P���a�`��^L?�8�J�H!��gB�3�O���]>r�<��@�mb�q�k��t��ZINW����gH����o�[��9�/����l�}�!�C�X���z�o�~{8���Щ&h�N�A�e�R���"{�SY �,K�.f�:~BL��:C��:���V���N�"��#L5�)=�ĕ�i��T���P��j>]�0�Z�p�'������j:T;���+��A�]�P�2�dГ3U���I�F�kK�=[[A�&�u���AT���Rnh��07�^Ž	k����/��&�Ԃ[;G�m�ƓA{��4K�UB$�e��;�����eBӌ�� n/o ���%��
oK�{y`66h��q���N��f��G
�����
_+�W��]���pAEQb��<���Q0��x�2b�ɣv:`e�՘�X�<�DUBw��d�J�)�?��67L��"8E4��Y�D�G�{�C+�v[��d�T/&W��?o������v�	� ��b��G����3(P�������3E�fn��i��~�,uƚ���p@�7�~��'[Y���62�yEN�;1?����W�w�b�Y:c�t�y�lZ�~ �zKΪ\�cSq������}KpI�	Ax�V��N-;�|�`|3�;jb��,�4HX��t8O�1KX���g��������0�8���T(o6��=���l�F�
K�S.QE�K X�˳�{i�}��r���:����)�*E[���Ns�{D���!Ļ�<e��(d�,C��ʶS*�P/y��%`��G`>�����X;��Mj~��U>O�1���'���?�=�R��w���!$��Ƿ�^���)��~W��)(��qVT�[{:=Y{�G�(�D��P�	�!Z7L�v�\�������l�Vꣽ������W84�R��(оpJX��<�G+_osa|h�~��4�Q�۪&�O�S U�r�ES?F�pC!:�*.�����H�Xp���CRb
l��*��\i/�7�逑1qD�3�/Z�j�� M����q���zNs��B���b�f����&�襑���}��A*�J$V�,��k�z!��Tn�L����=~��Z�����I#H�L:�{bI͘�c�Uv}����n@N�V�)_ Byx��������/>`��8��HL�m�QM�Klr{D���+� 6�X�;���
�.�a}�˃�Y�J��"�n*>P���\��6�!k�6�",��S�a��K4����P�$i�G�WI��+l�J5���B+�~��-�gٿ�
��:b���Ѕ[5����PN4Jxn�v�v1��r�ê-]������`�8����?\{���D�F��/r9u��OIܷ˵���+�d	��4�'�7��4,���Ҙ��r��u2��PQ�B�Xڕ�P�W����!cފvM�V�{S�w�����-�ד�+�y�����f��竬��l�� [��6��w�E��vǠ#b��p
X@�k#�v#��\�i��cAټ�,Z+���X�:��c������K>���"%���}�8�(?�����?o��yjϽ�(�ѣ����U{��+R���� �q��@!���1,䥭s4D�/�e ZED;�A$(���F��,&�K!4
��I�;&�*z�d�נ��f7�$�Ɠ��e��Wy��!^��og�:�\��h��뢩R�=���:��ISENv���0;z�PZ�l|*�Le�}�s���H1	�ms��6P:~�<�h2{�֦���s����nU��]���E��u �	�)�B(G���^��C��J���͞f�����+����b�+f����l������v��)Þ!1�T��hF�f�s��o���(�s���f��>E�6�0��]cH2�u�;j-]�������ʖR,��#�!�[��r�x�^p�qs�)q�'��f��^5�;��#��0&a���lʢl��yDq��Q�;ԣ���~b�Z ^<]�sUv��r�mDYs��u�	��c0A)<� L]����~}�m4e���h���x\4(�T�j!SB�#�Z�ir�F|}6u�n�W��z��4��g:�������|�P�WG�m�.�ed���)����i�g�2�-6��'�ؠ����M%H�g	߻���"��S�i�9j�6��tX���m&�q�^Q76ԥ��������=gQ��՞/*Ip�[�g<��l��$l�]w���\v�9�I{��6��kT⊗�ś�e�%�M��4���=����#LK��.���Y�6�f$�^���k��in�,QM���N�	�k}\��&�1K�2�s�*79��7�)��JU㖥���&1�e��T����x��Qg]W�������ã�-�D���DZ����&�\|y�It�T���vfr9���G[�t�C
�(��gr0�����Ҝ�\,^�͑��փ����a�9����m#�����(�&�ȩ�X"u���6��]S~P�|4�S>�x�RE��g��\�O�!�`�z�;lwQ���SS�e�[Ѐ������e�W�ij�����Kzqn�PJ@d%��n��<II6��&���+Rرr.�;';�r�����W�� �[:��o6���a��!�sDǵ%-�ްy�~pzǖD��C&�����<�0���:+��<�#l����/��σ��-]ʻ���)�N�X��?�!�$.:j��q��]��N<S0D��\Zz�ϳ�ֆ�\���*�O�_c���-\Yp�	�E����:��ʾv@��`��b�a��kpn>��z��F?�ɘ=�檡��S����7�R���4������1�y�ȑ�i4�M1c*��F?0G-Q&���,��Z����m�A����Q��~���sIF�Lg�<��c-�).	���Q�o1a�Sy����nϡ�^��s��.z#?0��O�=�'��!��d��Z���b@����<�k0䙋�h��N5{x%9p{X-b��o�����8v8���ۅ��^��q��c�}l^BE*jf+����,+$�NX��s��8a|ᖣ��c!�܁�cW�n�����	�yg���&���f����42 �#w"�R|Ȃ<]�i���C��A��H��ik��p�/l9E����ި���H�_p�ܻB?}�܅X�P���P����hW3��s�d���1����8���g��Tځ�A��I�q�z�OI.C�\�w?E~�~���#�3g��5�Q;�z�������/%��'�k�Sৗ��|S�j��j�_�H�iL���"p�i# ��1-L�^�~�IP�E������������8!���7��c���һ4�n�L�%H.Ѕ�H(�mTrFE��,�zK��t�~'|q/��?B]G���К�'�3R^R���Oe&uFͼL|����;�j2���h�'��k0�:��x�Y���;O}
v�j,�*��u�0=A�.O\�kƶ6��?�ii<����p�X=�%	;�BU��_����
n��a��¥�/%�����4�
n������m�ߞ��+��$�2��O$攅����4ř��rQ���_fp�+��,�Ա��Nlߓ?wZ犵�a��k$?j�M�
R��T\��Q`n�T��A�0�dQ�C�5T��q��@W�=[p�I3�
�D>����	-`gz�篙���������������P�W���v��W�w	����G�����o�p�r���\UEJ�7�������}���qKl�XGM�fo݁0���ն��Xvl{�����;��lXbѣ�09l��?�;v�2L~�+�
�-���>�����{���{%G���<_i)���
��?J�4kϔ�\ d�H����.���A�Y��^R*�y
Ʀk����<�3$8��rG�M�G�p�|�������y�l�;[�7\P���DmBY�S7�v�,�I�i���:�w����(�X��F�}�<i�7��쀴��pn;�lJQ5�5U F�D�^�ָ�ԍ��821�幌�%��wNS��!=����^�DV�+�*��X�/��'~�d�>-�~��~�\HV�I�;���>Z:��!؏Wa=�FT�8o"�A��8���P���!W�$x��A>�?6!{�]ʿG8����P��ê��
M|j�U�*�:��h�e�w\��=�_���B��I?���4�����j�L��6�x.���<<�P'Ҹ#"}����ݣ+���3��⪢>aS�A�E��B2�s�:I�E5�搞B�\�F�g�j�G��Lb\��`�}d�آe[F���5Tn�A�H{��I)ȽdB<@~T��~17�oR@�Ŗ��]�PX��.˗܃����e�G��� ��'^U���aݹ4ꗫ���s���:Sz�m�n��(؄�8{�	�0ևX&Cd&��w���9�4��@�b���JĵM�����8d�@$H@#���#��4�d���H+�� �#TN���9����k�ƓC�Q�N�f�iM~2f�w.�F���*嚑�������¦4�-󉺇"��Y�t��LK�����s*�Ry��f��c֢��ߩ�/�X�"��}��>R���_/oуT�V��|K� `@�Zt���/C�ꎍjџ�㵸g�/��e5�b�a��cַѵi���MF'�D�5���J�4���_L�_sG;:J
�UF�4cOf+���٨Pt�Zt�(�(�Q$Z+=!<�g_P�9,�d���2��C���b��z�~*�xPW�H[�(��xs��6�;x��쯯.c���>2E��B��� ��N� 5����|���{�"9
���0���Q[��g��Ӊl�5c��k��AO#Sz-jU�� �1���Y1�}�e�SEQ����^���?��H�p�i��p��ƥ�c^h��H�z`�<��A�����b�_���r���6� �Fwz=p"de���O��]�u!���T�j���H"��>�]/��P�{��M�o�<|F=I+�D�	&]�:���o��f�Gyx�ZZU�Z"՜Xܻ�O��<�E�m"Ȭ�א���k]l�\�9����	���4<ʢ�oK�rC�xL���AaE^t �/t�4?I%p'j�\i8�����[/WsVᢳȭ1���j'{���]���4u֮�f��״��td���%�[^�]�oX��3�@��I뮙||�b�ɟ�
Ϡ�ڑ�^yVZJ��H�9 �t��7�'���Q~�p����XD:u�N��wx�_p,���wՍuW�������L�m�{k�?mr?CUr�/m�t�MbǠɘ^��+oXI��~�`��X�v��C���/}?:�zƤP����p�}4,?��ɷ�o�VJ�}O>���^d&��"���������|^G/D�ʭ�~�O��:a,��:�g�̰\]%�sWcG��%�R7�"n[�%f��.T'��~}�!��;2��U~gy�3�y ���Uş��&�
C�yW<�7h�I��_���B����|��!����Q(���0�g�&
h�߂�4|5=C�����Z�C�*�+����	y�=wzأg�v�]�����19���	��6rJq�qf"��f?I�����F���lV"&Ȃ���^�
i�j�]�;���;:�♖�4q����+�{���x�nC0{}��}	��K��0�;.��:e*���N��r[�o�;[1�Y�v��f��S6}ޖ�������(�Zn��͌bLM�"E����S�����q)	{�6�w;5Z�8��]H���U�f�V>V����̾w^�����f��g�;�F��j�)��1~�T�L��
�*Ս�#Wъ*9B%	��O��i$l
���Ǟ�;���я���\�k�0j
�����U�E߲F��I�R���ElL?����2 QG�o/f�����$^��p��)>�z�#��.G��5�`;�Kڥ,b��l�W4�Ps��b1j�d��qQ�0(E�^ ���[춚���eB��4Ӗ�v�z�����V��Uݐ�QQ��*��/���ĥs��G��FuIƤa\[�+��v�i@U��Y)}�Z�[��:�7�{�Z��*��*���v�>:)�ɂX�蘹���~1j_(��gb�� �Ɋy�|�Y'K�%�r~�D(�v$|����Ƞg-KmG8Ň~P =���$']�����̶o�0���x驪	���Ki�¦�GP%PKP�B\��SR�{:�S�����JV�+�h��4��|�XwV�F�d����O�^��=��Q"g�X����DC�[`E��őod(́ԓ�r��x������1j��оa��j=��"�dPF�M^��������ԉo#H��U��vJq���ֵ�,>��:����Z��
�8S��o�_(M5G�5ͤ�G�9��(K�����^��d��P�>�q�Z+�ŋ���)���֟�aK�����+5ә�aK�0训���J��f!7>Eu?XF�?;��Z�,�~�zל�`&��m0��b��}w�]�Ź�e~(�Fs�k��U���E��伦��G�7:��;�����]�`��d�-T�p�M�"�y���P�32����s�ϕ=!O93x��0�	cg_�]��;�ϫcm4Eq'�A��q$�������̿��+���-��XG΄���ub�hT4��'Z�TI#Z��E,����E�38H_j��嘈�3�d����w��/����
���^l�=�}��m{��IL�lf���{P�x�AJ��"�	Ń����0z�?���8��#
uC�hE:����R���N�ߙR��$Gc�!
c�_��i���:�/o���	Ƕ`���S����ɣq�5�ZIEF�y��O:�q�;�(�a�d��#ڼ܉t�9H?����^$cd�Az�p@_�[�.���/Ƀ�ׇ��Zɰh��K�Q����W����uc<9�X<9
:��m�ܔ9d�|��i�DI �����uS�%�6���L�ʁV�W�G-��;��'A�Yo�7�{�TЂ�PY��D�1r�8c9�Y�B�z�jW]"�0N�������ʃ��Fۯs��ץ4��Xf���r*c��W�)������)��-B����0!,"6�D!��+JzR2O�Ӷ���hH�t��t��l�\a^$(#�I%wV�:l::�dm��)��8��g�>0���Q��a��.�F��M���^{ VЫ3x��側�kv�%puߚ��q$��1��@�8;����K���A�0<�>{f�S���4�7�����Ⱥ����{�����;���`���
f��&�4܆��������Y����%yj����r<��T@�bw�D��7��Q����HF;�ABh4���Ȗ�tPV{�,�E1ٺ�̒n��K {w�iEn;�9��lw�(�H)�F��׿��v32C?M){�3pxK�7gi7K�5
Q(�h��e���%�{�+�fǋNsF��$�N�c�5��� .h�=gV�M�,
������&��i�T�7�;�S��Ѽ��Gj���*���������Z���%S��|�1(ʞ&	��@M�M�d�6� R9�de#�xٜ�W������Jk�C��%���cz����C�vWO�E>P����+�� �E읚�Jh��>��ۛ���w�?����ë����WB���c���a*]���p#��]�,�2����*��< |Ȍ��/_�LCɘ�)�Ȏ�irP�W���L��Y0?�1Y�`�	�1ah���"��'�Q�Ȇa'�!�%\ȍ�GG=:�ׅU&�U�?�pOH\
��&���q�b���9֒[7)�#Q�d\��3(w�'��|�Ek-��m�j8�w�y��0~#.��7��cN8`�M!<ޠ*�{_6D� �6��/gw��?
� ZAͼ�b���
�	F*�?_F�JW,��(Q��/vʁ���,��.ҥ�F|@�W���R�d@��kc��ɍ*0֭��޲�Ks4X�Nw�r���U�i��Q�k�y
X	2[���Xڢ��
oFy��R��8��E���%���#0dG��9Q�A�iN��?1^���qU=֊�����fQ��C�n���y*K,o,7�ǑC��.�T�y<�֟B���D���� k2��;\�aj����[���E�3���xî��O�����.px'�mй���	�x$���s����s�0�$�� ��:Vf�ܷ��y�v;Hk�S��q�R3��������4�Qy��x�� ǒ"t5��Fh��.�^��G,��;)2��
����>6���oiL��
fv+�`�`F��qzq��!^��&e?��~ֈ���v���S3�\��:��|.s!H�'t�W���� SY��	}�b���f}���~&Te�:uz������):��ʷ��d�/�с�qnsV���{�����o�_ŨI��4>�
�+M ���78��k�H�c�i2g���'j�wu��:�8Jߥ�.�A��4�x�LQ�2FО.�i�O������;�2' &WW�~����0-��8�����i�Na#rWH�	��Ia����Ӎ7�5��~�<�&�m5�<I�_�@2f��ӎ["T�w��^	c�F�!�'&"Z��3΃�`�)���W����O�����Fo���m0S�:�E�īN̈́��  �KX��F�|�"$��Nu/�|�\��]����#g��%G�#j%��d����{r�$$:��.�Q%�[��m��a>�kQ7��4�=�6E�[Pަ�"GCH��� D�f�NF/
��qu���Bk�F�44i4���J����XcV������5������Ik�>��T��.9�Fp;~k��E�j�&�?��bX�d�߽�WYz��R]����GP��_�������ƖL����Gοt@S��y2	�׉�|O�XIVOH�ؐ6��s��7 cV@7��FM������cj<�Xb�Z`���*�ǭ���5����3B��ϓ�"�L�4�z␭��{�h3��-��aj��Đ}�� x�
O��n�,�j$m�f���?㖢��j*�g��b��!��Q�4b֗��ٺqʉ7���2����p�M��;��5��O�!L���x�67��l�W0 �Kh�as]�D�D��kWgH�#�ڬ�x��͑�(Z&�&!;���g�Q;�m���w�!�f���㹹g�la}���B�i��_�08��$i	�,`� ��H��?Ad���C�!s�Ր~iNC5��_n��C����D*k�2OH�-��yH��!�ܬ 5y�:6�a���C⫾)�1��l3wIU9����C��Ϥ��h�;���ˑnq�[�t\
�<1��d�1 �ϒ�`��*������%���達hfaF�5M���Dw+�f��o���q%�e�c��?�z���Lq)��� �]U	�n��w惰�ϡ��
rT_{����l�S�~^�#	���Tz"N,qN��f��%^{����V4�%�|��W�B�`|m�?��hG�y�*�B@��vR��کJ6ĽA��^�%\{5\�` ���-)a�u�R��x޶K`�1[�h�p~M�MRǒ��"��E�u��X������ͼo@�	MJ���5:#�Su/�!'Yq�����Lz��]ٖ��y�z�_Y�����o��)�bt�Xp��wO�����ݔ�x�k�"�> $aGBXٲ�<���9hL_yس�ˍ�m̛��Tq6B������=��f��� ������6
7ׅ)md�
{��a󍒗�V�P�*U#��j���n���HyWA9ڹ^e�}5or^����ќ��s;��vPt7}%=3�5���7�~�ZeR��w�*�y��ݣ�M�~���x�.Q�9�P��ĵ�b^���ư� �Z���n��j�����$���4��|����Ė=�|m%S!nS��z����v�9M�;�'�P��`�B��p�Uq|8e�u�'h�zTV:�/{�����`u���S�	|F��>�W���U�果C7Z{4ZJ7G��O�s[��< ���)�M�g��!qC�g}����+�\!�r��f"�n�*G�ҡR����̒YO�#�U'|T�UZӼ0��a�У���?�S��V:y\�Cɞ��`��B�����k��;����z�r���T�y������ݐ���B{ϼ`S4lr���T_-�~���"��	l����w_��"|?!��Y�:&)�⩜i���7�� ��xZvC�LOB7=|x@��+�������BP+�pNl@���i�m�l��J�G�*����>g�e�Ӝ�9�Z�֕����h��e2g���h
>�Qb��`I�If��+�j�Z7&K�ޘ�p��b��?aN�)����q+-�>#]�^��:?����J��6<C��
ۤ��
KT���h���ӡ(����N�R��D{�,f!�Ʋ��SN��(Q��R��N� Y2S��QD�������	h{��ĸ����6���'߀b����/2u�^��dq^�i垿�W�-�<��|N������G���L3"-�kc�\"U�[���c��:��o7�v���G�d�
oB��ՊV��Х�b2۽b'�B��~۶�x��`F
��l��G��>/,��Uu�4X �����PfI-����ӔPı�B��.�'E�x�֖v��� pV�^��� �����r-Gy]���ˣ�`�@��p-W��K�4���9|-cJ�ܹ�2�&�H�ж����"�4,����y������7L<t�5�L���-B뾅��f��+W�JD.�J�Լ/X�_9ʅ"�p��cM��z?�+�\TBZa����_H�VA���u�(��� �u5I���`�-�C��4�C�$��ۘ���s�z���;�f�)ڥj�z}���F}Dl�?68�q��W~�ƒ�@��AN;�'��c����v
w��ǩTv$T� �a}4��m苫:�P�|�q�p/���v�������;i9���V�!Wf�Q�QӰ�m��1���Og�oJ�:�����h�sᔲ��t�H��7��ߟoD°^eoڿ�3�xǠv+W
$�a;vy�[�$5`��&�(��@0(`�H��V=�|ݤ�[�pvR�T���k[��:�%Z� ��|�j�غ�d�	�@�q��
z]��{,��O���_fk�/be3���'�\w3_�pOgn�������v�,UQ�P���$����L�Wx�Z�L8�Z\���cSX��?W�W�K�HT�8���n��G�B��b�?���^U��4�r��K�"=�r�Z��S�(��ӊAڧ_'}����T:��9̑���H}YM�鱅�复�d�|�G��n�7S�l�	H����wؠ!�N�0z��U�;�����(jh�k��0b�� �O9�/i3rN-*8)�>�b�Ⱥ
,���ٌ� ˟ǴL;��}<R��H�wr�`s܆��1���x}GOU�ܘ֯�S����g�|��K"aCz�����'��C�>'7��X����#ny:V����O��j�A7~q����I���K3~Ż������!X�ȏo��z��x����z��ԎƴϏ����>���G؊�c��(�e�_�ʸeGj_���c�{��Wt
wh59�&q�����O��J���X|"#Y@*�OD��N�@ZB�#�-�L8ػ�V�2k��T��z��-0��|׬ ����r	e����^	$~]���3ݿ5��Zۈ�洞�M\�a���˴��EF�SQ���Q�e��фC��z�{�;*��W\3�*(ىS��rh�zi_���Ūʪ��_/�t���>0ͫ��>!��ѻCQ��|��w�7� �mc>SJ}Nȸܭ3�	�� Ϯ�c�2q�p�!�g^�^�D6.oQ� F fQ��u�<]��NT����I�2��z����G�A{'����F�D��B��_7W�R��)8�X��W������W���=�d���KO�A����~�X�r{!�.��.�@=���z
��@ˌd)r���[���ZYQ�I��Y��%�7#N,1���}�O����17��&v���������=u�-���C�2.�6>�}�`h�z��sz��\�#ƧX�$N�+���LE����k�VE�b�2�R��C�Mx�I�i��}�,ѰM?�x}�� 3RT gU�#�\Q�䬹Uyx��qB���x�MH��5�q]�G�D��fMR�^�������Y*��fP�Q1x��L��"ü1�R_(�k���x<�A�ב���Fc�(�T�lA̤,�����˵��q�ˊAi�KZf�Ӛ���sE0:�#7�G^��S�Y����@7�[�C'���d�~|]t���a	�C�
�2�%�Nn��!�d��l32�����i
6m ���
��K]��B;����Z ��~zW7��$Z�+ʬ��9A�똝9o�EG��p�V
�M�����C{�bx(�b	�70wf�H��p�(��Ĥ�;U?����o���P�(K���9��H�1�1�&��r�!�����Os���R;}�g	��db!�b�0�<VV<M�9N����h	C7�Ѝnwc�Q��r�Α!���շ5_������r{�	0��bh��ue:�px�36�.�HG"(*B�~#�l��s�	�^@)w��_7��vM�9pJ 7BEx-���Y؋2�[4�kRJf�$�f��`�>����(9
����[>��e: :,g�^������*�(
~3��j׵���2���F��iW3@"��cy$�����`�k��mȊ�C�0�i(�\��x���PZ/���M�`�W�)ȼF?�˥s�4���ÇT��wy�Tv����*ΐm֟�G�;qc׊ݝw�u8X�<�����?LV������ً)�F���|ƒ���k���"O�ȿ�[�"�i9i��/�/�d�s�����f5�
U�}�ix���' x��֩��p
��}(�l��LO{]:���7-Յ >l,�>�'IrEi�\�,bn��ocم2��!]�$��������, >�U��k�h�O���c���nw$�j����Ҟg����շ&�!	�9�z�����8>߽Y�JD�WEr:@|�k��rL���L'B��ۀ�1iׁ�#��5�GGdz�v�"��`(Eme ������zeio����b����]�/���Nz���GQ��<��Q��+	Z�v��K�c�Zo�7��f*t�����黏�(�d��N��`zJy���Z�Y_ `u�|�͏���i:��!�����0��ޔ��2������)�Z_�i;�d5���V�qdX�PjZ��~�'��G�Nt��a����r�E�d=5�>����h��WAflAP�޸]Qp6��̊Lu.d��0XB�4��X�!�5,���g�Q��z��8'��O�
Y�"�qf�=�o�h��o���w�@]E*�ɷ�=��_�]	]П+�$J�Ǵ�)�3�����C@t��}\q��(LԎ�h���i 1���V�ӦB?�k��'Q��	-��@%��G���nI����׾L�ot.�d�4M�{� ����.�L`�Q+�Z�v��� B�ٮ�!��A*��vE鹁��Ŕ���
ˮ#�C�F�30޵S���!�\�J���]�Tx��1�FR����)/yZ�"���F��`�Q��ҷ�O;KW?�8&]mBKLŤ\2�+��Z���6�I/ׯ��5�c��r�Vp�M���䋃ݷV�`����Ȅ�|����b���c��v*Tpd���[ǔ��E�a+���E5˄�~�����*��A��N��.*PN�/P�TQ ���;���Z�T�E̵��D����9��O��bEAS5�5�p�m|m��,���Ҡ�+r�+��fh��>��C�kw��V�K�^t��
���τ�>l��#�J��!,;MLcW+b����z����D�ļ\�ά}:b��o���3붉ݥÇ�ܠ����=�$zXѲ��;R��`e�~�yGJ>�"�"�Fe����E@�RZ�ӂ��E(��@A����Qòʚ?aWk9L���*\��5�К��K���!u�P�����9�̺�mX=,�����Bt3�bW�����S~�j!uy�%��������ڜ:�zz�� $o�v���BI�a �@b�|��m�@�i��V�P��L�-V��6O{�&����YN�^x	#8O/�횴�/�g�qk`)+`�M�4��KZ�勄�;�jຨ*\ECk�4�o,�k�bR���^^ⴊ^`��*�"Z����5���"U��8��$�<��� 0�w���O��õb܃��ro�^�,��Td�lU1ٓ�-2�Ѷ姛b�T*�t)��>=�iI�fy �K$<�X�L6�����."���-.x1w,�N�>mD��ԅ���æ_A�h��i��~<��U�}h�5�ԣ�N�W���3�^:������ 	�G�"�4��9&KR�;�Q������;�̚�w���q���V�
;cb!�qH3�J�OI���>�����ygU3Nk����)E*S�/'6V.��;i�`o��`9P�3�?�L�bT���h�}.�=�*,3?�V�7޸��x��;[䂒K/vl\�Q�c?  �jp�����ʹ�)�
dH���� ��OĕYM���)2T^CB�;*���#�����@m�I�� imE�V���X���5x�I����Qp3��8�pjdR���ԇ��L��P+��j3`ΝT,IN�hi��U�)���Hݢy���GR��9�C� +gs6o��=��t˳G����}��%*m�L�I���s���+���<To�"�p�^�h��+�y[?}�]�JY!{R�ԭ���8�P2w�g�y�����B�{�����<}=U���ju�.�lŃ�j���AZ��
��\Ex���4	#87Zʴ�dw�KH/�Jr��h�KY�G����N�]W{�-�B��h�x2�I:S���z��ı���OW�8�b�3"��)&TG�(O6Z�9G���,_;L�P�fp� p����[����������~]9G5YyUi^��G�a/�P�b�ڴ������W��G�b��"�=��s��뚩����o�(g�±X�0��W�4�����q�T������V��fZbS%?9�y��iU�h�x�%t����TV�����u)����o��̝�Sd�4�sA�����i����_מ�Q��k�lO���vt1��j�� �+p�<����S|f�OQ����$�+e~At��k��X	A&[�$cΰkıg5�K�ń�!������ϙ��p)Og#S�`[�㜴��ʤ��h���2��$���_L�ӥ1��J��D���k�%{��F v ��J�E%"�ր;��k�;�k��#Kӿ��p6c��}2�&�ꎨύ�R���F$����\/���
�Co�uK�H׏t=K+[�A����ָӅ��h��)��N��xӁ(�1���a�VH���s.��Iț5��X�a�$�c	�h��bk)5�g�͸�f5�����H��F�Ҍi�F��=*2����enB�.���R+H��=l=o�o�hS�>��U,�)gͬ+OX�ѱᣐ\�d��4;��φ��O�
���+����dwW�sY�]F�Z���� �����1�k<���1ԕG�����n@(��w�;�%�����)+\AJ�`dM�zT��de~�^�'f�QcCQ8U�p�y cp�����G0z`)I�4��'��֊�^�b6�Tʭ_�?uXv�z� ��f�K�֝P{�I�,T	������r+1�������fAjћR�<��g��!���Ҥ��'�W�T7��r��Zń�������(�F�N�I�%ߙs����\��(fuq3d�]�Wx��^V���$NC��9�-+�s)4P�wR[��'�.8����'5��X�^ }��@c�/�#S���/s����Ҵ)��ZL3$��wr.��s\M�_�2>�ƢK��=8`�7^�^鸅�E��vߍ����X��ޫ����H���p
�_7��Ѧ�� ~��	��p��r��w[\��O��1��9�C��-ذ:�$��2[p�`��`_=\e� ��Z�Q&�l:ʰ�Ԧ���B%ʃ&��J�p��yC�S�kCJ��γ���`��zm���?m�l���O�lҝOs鎠V�"�B<j�n�d��_j1?��;�&s�g����aF]���B�m��5ɱ��Ù�	��+"���W+Q�7yW顃f�D	�0/w��%�;�+.�LMU�O���6�7��YC�Y�, �W�1���Kx�s���3ub�����M{�o����P'G�)����0�Q�h��${J>��|R��M���q	l��' $D����fb��\��o	~,:z���!�v��h����Y.I"*�>��ACz�t_	%�R˳'��� o[�A�3��d$#���T� ���S�����|;���؅�m�X^���MJDZf���$��ED�nq�>ejv s���b��	�"��",�{;*�;����W~S��
��o|п���������9E*rS̩�i�;���g@Ӷ�N�����+�bx��K�
���<�0�ߌ@n6��6,�Wt}���ONVZV����Eon��\�%��fA�dꍴ�]�ESO��s} �0�%��*���-&  QA(�Q�6���G�L���� ��\��nI��
�~W���Շ���3��jj�7s���3T�&��ѝ_�,�E���U0�x�g�q�Ұ���#U����5�{Z��LH���
"�5�D�׼��%�l��o�\"Q��Z��/��z%8�#��צEg��;u�k֍�~� g8&b����N��>y�)�iB��@�4�6V���BK)QJA�*�J�'�F�c
D�Qgu���!�*�j�C��=��hc�Q���(l�)Z�dq���������ZW��WdX�5^�0�ćm�Q	�N7����ad�� Bx�&ف^���q']�B|xb?p���-�è�� �s����]�TA=�6��
BJ�R���}Z�F:0�ɔi�JcF���%,^�
���,.�`���+�3��|�wFeWG�]�lp��1����S)��j^��^^ގ��!n�
��P�l���đ���4���>1�2/�ǫ� ��g��N~uD��<�����(�]���3B��F�v���$��#�R51yt��$���ɻ�se�]�O�s7��&���8�%�̚g(����C`O��@P��={���)�D�������j�z9�3�a&y��2zC�\���b�Xx�/��مӅPj�q)�w��9u�F8a��?����s������\~���mxe�	�S3F�.����'\���[��4X��ө7�B���y���xq�0@5I��*�]���y�����^�Z��zŴ�}�� zg���8�m9z����oĮ��9Ey>Xw	��W��߷Kf�GoS�ڻ�˲�߃�*������n��Z����zn]�k�V�`=�M����	X�햡�2AIP����[� ��Ⱥq_����q`k�����P�Y��K������^l���p`�#F�y�<�`O�yQ�����#�h�s��2k�u��B0|�m�-l7T�J]UD����@'��΁ٔ�k?�C�<#�k��T�O҇��1fR+��,�y����T�JȂ(���ƚC2�B��y���6�B�+o���Ε§/���d=Xn{��J%��&�P����H]ķ���F�+��H?�|B`?�XUo�ҠH�4��΄��C����"�ۑ�	���4qZ�hC[�SN��.��uƋ �A|X���3Q��3���f��}��#IE�Z�lV���m�媜]�3H�8�3�O���6v'2����:x�0w]��h�Q��7]�g*/0�z����va�j'���n����S'�vqY��<�l�zO����g��2<Tm��!����C�$t5X�/T�6}73+C�bl+a��[�ǫ�QFВ@CG���&`x���jNÂZ��8�sMeK�{�n��H`���������S9h
�I)�4!����K�V�fqĴpخ���(�?�U��$Ȋ��>��ُ*��~R�<�~W�ZH�R�>(�"�0���ht�Zy47�ɐ���@^���G:M�/�,P ~@E,Qx��3�.W����v�� ؠ�t�SO/yyp��2�w���$����/�֊/����䓞�$z���H��&)V5��<�S9d�/�@��i.��{[�����8~ج��l�A�����ND;���~|��Q|rUb$�y9'ԣ$����f���'�?H���t���X�UU�\^�G�c�#n�8�ϕ�4wL<��#�)��9�G;�i�w��3�C�à�ܹ��oS�xF�R-�&Z�n�L-1�0����Y �/u��.�倥������i{ʜk�6�X�lm��K�ͺ�~�8׮nǼ%����9m�eoU����n|9dJ��a�N��G���N���ǨfT��dؾQفݳ���K3�B$�)K&Xq\�Gk�y���l�!��N����[��ES�*�2ɣ;��}�0�~��W�JN�v���'���Ȩ�J�$�'.46fD��C<,T��-�c�c՗O��Oۇ%́g��}4�w�e>��C>�dwвT.ʚ�ӟ#L�цl���S�a��SWc��7܈N���X��S-�+U]�T�
�-E����_�;9�_�Zŀ��%s�3_���$qh�FiW6�uE&W����!���m�J�����R���b��9j��f��vpɷ$iF����$>��0Y i�pm�;{��.���U#B��J��� Yt�4�y�f��/^uoAJdl�3���瞌�Չ.��W�#���zQN���>�-MT2��)��T����G��7�¡Q�2���p,�z�Qx�Rw�ޜ}�:�S�Z�b�����}j%±;��gC��*%)	�)�X����D���_~7.������]�a�!L�=�\�&"��H�`�(�/۔����mKN�ܳ�wQ�Br뺴㹴<;С1���H�iw�y�H29�r$)|���YU�:�#5��SȾ�k�I����ԇ��+��%�?	�L�WE�& a���.��<�!G;&aE��Ҕ�(L�=0��>.����7\��y�86�r�ʷ߽1�)�����Q@���?`���>E�+'6DR�"(�H"����:$S�<c&��HSs�v���
����2@+A��8ٝ���>�D��pfEOM�d���$j��
ߚ�BSAJ�a�Ք�+��G�/u�z�VɌ\�����ۣ�+���b�UV���*i#>(�ڰ�@�?����i����Ӽ0��0{F�qGye�b�P|��I��jPV��I^#��������e>,���H�?�<�Զ�.�N�q��p?_��>Y��bv����4�8^cuim
�7%o�~L/�c�*7Y���L���J8E��}��/��7�S�O�&���� �K�
�_���܁!���	�e1S{�R�Sb.2�72�9��蘆u�B�.�&y!X�q<�r�#Z�[X�`���tr7�mK��o]!lh�F���)�]j��{G(l�:�S(�(���,�:�0­:�)Ē���D�XT=շ��r�ąJM�����5�mwGHQ��� =�u	2�H��'<w(��<�6� "�����knP|�7��݅��jv��h���<?�"�zE��@P��ZjH��W��~�-��IN݋eF��S��؏���CE��\В�=��<6�7��nï��п\)�1Q�;Y�QK��sā_l-�w��\��57�,Z�_�P�=���m�p��ȭ�FG�� x3�D|�Շ��1.��k���\e��}��w�ӹ�����1���� �
�l�V��8KlХ
]�ځ�`L2���Ytԗ9��58�m.X��3#p>6A�|����貈���������fs�Q	��ҵqKև9��]D��9���@��d�Lത3�)268S��VGb��\!���`����f�!\������ţ���0{�dX3`�-
~|˃ -̮2g��~r.�5���Q~�Jk-� ���L��%�8֐�L\���6��l�(���-kUq~�4.�U27)�)u�Khۅ��ɿm��(�_�ӂ�ۑë�JLo��k������d��s�N(��&��50�Ύ���horS�����gHb�/��T�?|�u�X|�k�=�T��pU��9�D��>�6)�zd���8]�E?��{nUa];g��)1j*��W�J;Z?1�S�+S�(Dy)o�M�E��y:�����l�D���h\D|��x���s1�W��boBy����:-���V{��C�����x���tB�H3g�6�9�2��T�D��!)��,Hʍ3�~]�A�z�o��ň %�q������Q&���^NLF�KP�I�g�$V�{����r`�b������<����?��Ҵ����)[l\#Z�a�$a�&ᗕ �P����cY�����=/XBK��}n!���'�z(�ߨ����[9cZ���T\�(��UF��������:�e���sk���Ԝ��2Y�(�yՁO"d�w��_����F��uB�\��o��?@�*����}6�KXh�&q<�R��^]��]�`��ջ������g��B7kz��24��X#|B��2g�)p�f�Gg��jW|j->��	#�I�_ނ7�!�JLʇ�χ�s~o�h�LX�9�*wRȲܐ"��;Ѵ�DQ��/V�PSiv�*���<+���L{�s��Y����A%�=�&&��)�$�fֽ��,:���)��~�b5ކ�E�Ĝ6D�<�0U���S���0��dK��P8q�|�,׷f�r�j��L��n�H�}�pWXo��raS���qk� ��0e��_����NUO1�`{'U�p_�<�!eN���a�
fq0�LɄy[%�︂���4�[u�,-�r0�Q�K���b���ǯQ|}#�r`�n���k<�����E��+%�� '6�^�[P��.=ʜ��uN~�B�o�����\Æ�)z�#K�>�nP�sz�'-ip��e!�eUI�V�"KI��R����C�T�ؑ��c79�H=�O�6��Q���/��EE)l>p��P��uY���I�Q�o��J;`㦔dQƈjr�JY����n��b�萎��`~6��v����Y� ����J�:t�����Q�_�Rj�W%����1���nۖG�P&�����K�X��T{2�=H��X��ְq�ҽ���A'�XF�2�, � ��f1����֬?��_v4��2�͹��c$�+��ZD;9��Q}���oc���5��|� !���#�����L�ш�2V+��,�M���U2R�yv�XRbp�XǑs����_	|��
�]�fQ�n�[(d��FU�u�*Ä���nU����%s�(,��2>�TM)�J��~�	#�.X�a�rߩa�Q��Jb�q��e�h̙�1[G��@Vr��>�8�2�@� ���.�@�L�(X|t�V WB����\���p5X�~y��0��y���o����M����*PX�l �KA1���O�W IP��װ�A6	̫v��w���4$pێ�}@mM�^6E�`�9[�� �����9-w�#��@�'YbM�����R�,����#�,Ei4hq{���t�]�k#^W>g�n���a��%$.[�*���J:���8g'Kv4�D�pf�{�f�ic�#'[C�����r���'ޘ0�~u@�  T&kV�E���G�OD�4"��Į9�'�Ἢ���Y��n\��8&�d�U�9�%��}o��⬣�C�g+s�t�T���x4�&�g7ޖv�9�����],�#��ګGS�L���m̃��Se��wեB��)x9���b��b���8��_|�	�o��	g��;6�?�M����lbgT�Z��b��e��mw4cb����x��GM�D�.��8[g�"ZSK��/�pKD�����;b��G�U��O�^�D�1+�cz�+���^�N�l��S�'��i�!o�Ip'�����/1QaJT~��
l~���3+�p�!ڮ��3@��[1 	���'���}Հ���0e��0�t�$4��M��$@j/q�Ƒ%X�~��ϴ�v�����������{�Q�|;P�/� �}��c��������x��a���N�he��6	��8*�Ӽ? 'v(O�(u���2��:������q�̨��KOo��-�Z�7�d�.�8����aP�AV��*�k�ba+!Ł�N����O8	��Թ~��ؔ`{��Sr�W#$�̡(�6�G�FM�@U���ޯķͦy�&������X�ˈL'm�V��r�	@��+WǞ����4X_�X^{ev�ь��H�࡜�t:�#�:&H#uʬ�oB!����	�la�}�0W^���Rhʧ���9�(�|AG�H�s���� �3�n��S;�8@|U�_�1u��UJ+aɑ���R)ce-�T]��	�+ԥ���iNbH��)?t#`�T�X��H+8�$���+���zއ�sy��}f�= ��`�}�0	��Ě͑���w��3���z��u+��HUL��(�2cPH<Z�L�df�k�#�h����c�b��?8;�gTuHI�)eZ��+6��o�#CQϮ�R5M�-Rm>�+E�����G3���#ܥ���I��PDF���4i8�z2�*��Z�;{�J{�_�WDd��,^�봇�\1m�N0�n+��}���[*�;�7*Z������vc'�_��A.��63k_������`����,�Bo�����Y�^jagg5.�ͩ5rm�z/�Zu3��ͻ���c1u�R�)-9�)���!k����=�*�:'}]Y�4a_]G�Yd1��Lʱ_ԫPVB�L{�W�T�=�ga��c��H����&���w`i�8[<w�{xKv:D0�'�����j��B��c�V�5\I{���xn��g���sx�īh����d���H�c��/:�+F,ԊZ���mw#��&��~%v!I�wAL�$����(��D�҅�ߪ�]�C�&d�,9���!9��(K���z�@Q_�.�ޤ˷~v,��
P�z���8�X�|h{E�43�����߶Bԡ���TOV�Ώ_�t�j��]&��UqET��hO]C�|�f�� �8Dd�މ�#�K���5���~v�8OrR�ʬw���m��v[d'os��I$l�'���e�v�3._䐛���]�s�e����b�� |�`h?��o[s{
U�G�i�0�����7I�z�I/�d�Y�AV���#��ݔI?�V�U�Ao��W�u�:#\	��Yh/yڼ(�䝴���)>��DkA���d�#a���)���-���Lܷ�h�=�ֳ��{��� �ᄛ\Rw�χ�e8@�Θ��8z��]��֮^���aﱉ�IM���L�wh��t��?�qixZ�";��
����Q�d���r�赊�:lC�� �p��pa�U��|?C$C�^��pRr�Fl@ɧ2��֊��2 ����yx_$�����mL�٨6Ƅ�V2��l���2	�F�'7��z�T/��eD�W��t7�ua�Q��I�y�
� �^jFO;�R��5�&W��*�L�Gk�?���!|��#����6j��#���J=�0��l��_0ː�Z�v�uoӇ��	��$<a#�=`�q$���Nw 3� A�����31�r�Jk̮W $+�	�3�X��[�>�Ԇ�Eq%_}rS�c�z��
�ۛ��Xv��o��_�;�lM�'s�B�n ���f��kj{���3(C�V�l7�Mv�>��N^�>k��ȶ�d�ZO}��?t�Ҁ����|TUw�
gQ]ft�j|�.�&�P7i�����Q�!)i&�%$��~3eڦ�"��L��}�)��Iܞ�1���4M�{"��f��~$����,L�����>mmϐ˩��pX�f�g��2Q�� ��\Ѳ�|����z�[����`�i]�7�y�y��ݍA�1���=���H}C�(�|8&��dt^��|�v�_�V?��*����]�e�W����=��d�G4F)�����pڙ��=W�gi��^(�M�Y�:�a��/]<�
�;���������=W�50͛t�?G�cC_��i��+�-���;��*N(s��th�QUؒ�:��2�,�~"�.p<E�I�]K�p��~�Ӣ�aخO'0�T�h����N	Nj[m.]�$�C�EQ��x�eKƍ 1���G��Mn8�����ӡ֥�T@UD�9Ӣ�Őj��S��P�"�������X:Hܧ�hv�����m������5r�T�:���I2�}�]�eچ��� $FP�ґUt3RR^��m��a��$�cQ�����{Ǉ<(6&�k�qm�e8�P ),1&�&19D^��\x��7�TM�����G\�@�����qPc�K�%�P������f�_T\�U-6_C�rA�u55�c�	#Y���BD=�śD`�n+4+P�.ט���{NT�^sKC�Q���9�Į�v�~�����7�,i �cxo�9v`^
�O$��6ǉ��]���]Þ�`�"Ah��J庤6�g��R,5��mwp�	�u_/��������������7��{�x��!�h�M�E~Cz`/��k�3����-��F�E	E��K��r���"�(�0{ڳ`��p,.0� þ5�����L�Z*v�`@���˼�!�m$f c]qi�?����8C;A��M�uJG��6i]�.��2�l���	%���pE��;�p�\r�I��|�-AF,qGQ3�z9��
7�v�P�͌�,C,\�j��;V$���<	�U�
f�e��˜��α�i�v~@8��Q+�b��O�z:t�y�:W�����H��U�إ�y��ŮG;�J)�$�y��.
��Zy�9"v5tu������|^�#��OƔ�����[����jl�|v�O�\�f��_�Ӷ�ꦩ�B1�B!JJS^�u�h�xd"��.��\���[�C�:�I���`��uS�hk���z�s��+��2�hݝ���
��lm�)��u�M�dG���{ٜ�����_}7Z�%Y��F�����=˽�2P��b��1�n��Wz������Փ�Y�|�O���xɈ����r.V��dM�6��
Z�C"JmT�S

���@�yFz�i7*.��G։~(NL6y
ͧ9�A���l�9���������H��C��G��0/P/�iu��+B��ӂ8��3��]�l�x��CI�A$lu�_��d�G�����Z�m���ō�������z+m!��	���F��ɝ_���3$#;��O�6c�|��1����\�Ca}_,�wE�k<�ɀ�( ��^ ����6���Cꛣ�?@���/Ǟ�������?����\�GW�����q�F\�= ���\\��M�d�D!� ��V�@XP��Ӕ�;���g��ҵ�k��0͓�6�}�$���HZ�5پ��PU=�F-.c�s*�,p�{x�A�O��<gd��J�w�<�6aO [���ŵJ���B��R#
X0xh�m
�	����,�����dF%~XF[Ǿ�i���� ��SD��t9+�BFC�X0�� �h��މ�n��H�O��&����n-���-���\EM���5����������2��J��yI,B!�����[(h�-�RW6qh��Ga�me7�c�t22؄9u2Or�1d�u*H��a�҇�e��e��򣖙�!9�,ƹ�
J� ��.�=c>�#L΋n������	����?�q�0��d�/gaW ky> X��ϻ	�&�r�}?�ky�K���S��u�E7�PH�[�U�꺝:�9>�<'۸�� $��j��Mԛ�4�{�����j)h��!�E�+6�x�Cݶ
L���g9��F|��b��Z�V���P����##�|��������Ї�����}u9��L�X
Df4=�`�� �j����Q�IRsYX��W\=�_^�2Ħc�$��4�����y�hʚ0�����u��3(�u&�V���\4����mIC�F+�p_�ʏhW2���v���ܜf���S�,�!2y��)�4�/h���]池��g(�W�U4������.*Wv2XI0,����!E)�*t(9 �JzmL�p��N6}����ë�u
w�@h���U�~�:��FyBs�d�>�9�����"ŹXH�@�(�v->���ݰ A�}�����eE��VP�^
�������I	H")Vp�t↸-k��-����#> �pè�z�1�y�;�Xfn�K���$xU���H�=[��#	˽�EZh�
���ɔH��?iTE�n/���PM��D�����K�
ֵ@��՟��Je"�]�{xBe��I������8%���ѓ��f'��X��E�������\��+,~�8$]�
�?��ڎ*\����NmCm���wu�/t�K)]�7��M�X��`�VwX�O�-�s���w��#~�@��p��������G��
/YS�3�Y]��Q��N�z�ǌ�<�K����eM0���u�������^m!C�C#��>�'��7(Ir}�{�R�8�[�K���D�����(�v򤺒»��NM�o�d�6�zKK���xEb��ey�"�K�&��L���eq�X䋀�sQ�Bͩ��0���
VP| r5r�7�����5�Mr��Zۊ���*��׬!^������?ͫs��5��^0g��`�+�7t�x��{֙�L/�ti$g�����}B�|���%��85ؔOC���࢖�+�?2ď0��c���;�}�� �]\������������5�GrV"M5Š����y?��{�;Q#.\��1`�U,�RZ,��uR�*rjB���,�'�a��y�*�*M�n0��L�z�ҩk��-��\��N���$Rs:;5�JX�\�N�X=1��T�vY->���,�Ӱ�A^.�_{�)K��E$�!{8M�yV��pa�����G4�fS,?�1aZ�ۘ".�L��Neb%R�,�<&�2v�����N�zh�D�-��:�q��C�`��|G�ү�*������'RV����:`@�%�V���UL���B�͠bk���<��iMS�t��P���`���,���h�M`���͆O�����3�І�\\��悝��G�)���W�(���3�?H�{-��l0$VO����*v"0S�����ct�BV�Q-;|���'V����V6�w���2l|�]J<
-��d��9܂K��FufrF&V��]����SȵU��x�=�?C�D��s�Ǿ(��J�0�R�.7Ͻ#qgx��w>u��y �����<�:�\����b��ep�����[�Ρ��W^	lz�̍�D^l�*�6�dG �*o5<�
��2֦���k�E�7��N��>.Z�������B	ɻ�~N���/m��$@������?���t�K�N8J���n�Ca;yf/�Zq�A�%J'����k����a�sS+ϽX�q4����o��#8�h��Dx��:%������gr��p��iꯋ0+W��V���>��I�I�P:�����+[�\�0�ϙ��7@<<�T�Ү� 0w]�N�����X	�>��ui���y�Q	4��UT���B=�	\�bOiPڰcb����a��M�=�?�B ��4i�<:��w����U4M�3���K\�*��W����6x%��mVdc/��y��Z/���)_k�jw�X!��o�x���{�,��!�{�{}�b�T%�avx��ژk�fG���e��E�J�$�.m}g�t���.����qSU~�����Z�̗�D���p�v��JQ�<��qJwLAړ�_�������!o���n���	�"q��Q!��Ә�PS/ѽ�":]kGY�(�'i��
>�`��c��(�^�t��H5K���@��N�?�n=�9M�s�P���! _�+��`{�C2�����q�����?L�r�bTnM�vxu{SP/(7��vG���1&�6���3d7�����֩���+cUu��]]�����"i޾8�h��o�.��j§�����ޝ�aw�=\Մ�@!�{8�7����.������V���*��a%܃��a�e<�����V�h�|H*�Dj���	B�ΦxCoU�A��Sw�}��~P�7�8*XZtz����8[��$��7����ŧC.�焟\���S"��=�۳HP��b/�J�d�Yo�qZJ���Q�#�2O�8V�Ԓ>�	���r�<@2N6'[�G/���+KQ��|����!��MNH�i�#����~%]������6;%�	�c��am�%kA>V�1�j�}A�@oy5��A2�A{���R��|,埭s�}�`�\�_��4R6��d�RX��M���Bw�)u43�1�o�Q�����bi��ׄ���xW��Px��~�Bo9K$��7go��*@�Ԍ�tY~�t˄0������%�k>�2Éq����7$!a����,8���!�{��rHaZ����M>]��I*e����]4Ĝ9e##��DVh��jۧ�?\�@$�CS�Z��3,�CJ�H_Zj�mV�,[���1�̂"���2ވG���8^��"�ql��r2u�t4�`/Ծ�*x3_gM�-Jz�J]uizIi3��W+����,|�)��VK6�\�{+d"g�|�q���)�RH�r��C�����O��%ʕI`.�����r��ĎSӪ3�uwCy��jW�oE�8��l)�!� Y�ow%�K,�m��]��s� 7��~j�P���.�j�ڦ�lr1�bw"��|� �j
x����۸�ԛk1�-���	�u������$�l�"�`�7��x㙤�Ǜ��H3C��N7f�%a0k��z�!�Q��~Ѐ�v�p�Wd@�V�	�����!����a?����ƺ�i��r�|kn��m	��),�oZ��s3�3��'
��_���)���,��EVt\�&�]��ޅ>d��`�)�?ԡOox��y�ө&�k�u�t��s\� ?w+mb�VqV�Wl,m�:h���&��.�C(��L	����N�<���32�S��_�"&�z�>���v���4��=��S�&�p����+�0c���ޕ+���Q�Q3�<��Z��_kw� �T��Z�'��T¿�D�,�z�P'�H��]�ޯ[��ʫ��
��`��xK]�/�HXV�lǸ���ǰ�/O�.�k��U�2�'�����y��o
�υ��Fw��W��Vz�i@����	�e��"8����oa$���"��G倚�5o4���h�vQ��O��D%�ؤ��0}V�rK}wZ�-U#�	��M�
@�io��G��2���j�á|��q�7�2CM�2�Q<�*�թ6��Ը'~�E��#e�6X�Ջ5[h�*Ǧm�p�?��������M�}�z�(35�Jo�n�#�&�S�M�Ţ��v��LV�woE�Z�����\{�P`�z�GjQG�UR�r�jȆ{m:�2L�+=���Ί[�lԍF[���:�BP�nTܯ�2W�`Woд��LF9j)�l�� ���UV	o��J�,�M"y���/$�p��m��;J�l��Â�c�e��,
C^�d����q�5'�����4T�XX�� ��l������h�1��Bi�C���(C8	���M�B~��UB�#Чl4���R��!�>r����Q
%,��{�RZ�qH��OA3�'�G�&��*R��<ʮk��	��c��6����_�K�-�[��>�N:U���gн1TІ����J��t�,�骰F��Q�)
�w6���O6�����^{��Ln�,	1��6�cf��Q5����
�i������Ѧ��
)�����X�Ք�;������F|[�``�ϠͅXF��=B�-6�s�f���6�?��bIr�J�L��2�,�
z�l���������[������k�R/r��P8�����;3̇C-A]�(�[C�q��_0�^�S��Kݪ���D~�5�.1D��4�fe�B��"�"��ȅ�+��Xϵ����B�`R�j~��c�W���H<[ǯV�D����mg����pw1>ꂰ��0z��P�?~r��1ݺ�@�;�9���4L�Mc�o1�B�gR���	�ߨD�yy(\ٰi;5]<!�T�}>̥a�~�f��+�K�p���P�X�R�Zu1��G�C�����*=���E��,J��W	o��@�n'�������A2WL��=�j��[�ޕ�L���)����;m���E�ٮ��+PR�b�W��%8c�����V�F�O��!;`)Qy���V�=G�Q�~��B	���F��BP?�Z谈��
C�b2�*�G���Ηm�C��\�(/Vד�
�h)���\��P梥� b�-������ЫM�'$�ƙʴ'�;���KD�F4/)g_�<�-Gx"�jak\{ϴ�|q�f^@7�����R�}����D��Ф�AZ7� ߗ-�Z�1r�9)6A+VY���M�;F䬊�i>�Et\��Eu�^�����+��ݍ�rt���!S�����Aȴ]�m��3�5���@#�+[�qXŌ�|�Ԥ&��N�f�F�ԋ�;r��L���_��={Ґ�~�W	�wZǀ(Pըj-�x���t���h�_G�-IH��B��Q��+���p��Ϭ��^y��cM��]0�$b�Mp���nhޞ��0WO� �\�E:50��Q�4�	�e9Q9W��K�9�'n���K��WM��W"ź^s�\�~�F�B)������=0KX��I+2=SSe [LxK{j�#S0��0�F��h�R}ԥ�Q�M�EV ]�����,�vv �K�E>lŰ7,IB��}D�j�ghp���B��O�N�Ru'��6Z=}o�(�e6P>��KiyX�?��b�����NҢ螥Web�^m�+�%0��	=
��$�n�6��w{5M����H"r~��a>|9�ᔄ�Z
�c�7G��G��"����8F$`>F�Bm$��V\]b�"���tӾ���~�^�hr{,����x.Dh�/�����r=��D�Fޢ8!�˔\��lƣ�+ј���!�g��!�f��4i���$?�a�@�$�x����jv��n �1�G�������Ѧ���kz�ݟ-�R$w��nA��L6��3��uяA�b�G�C<�s��ة�4�	lò@�t��FG_јBx!�`,0��=���;X��U�r3x`o�V�$���˄4w��Y�q7k�><�i\�;*3(A`�4��ԣ����@�>��wO��'���I�w{��Ɯ�\y�=���P-:�� 56B������L�X��M}]q�Cq���/"ER�lzrw�p8�x�b�O~�7�N��W|����bţ��`k�}�]���M�I����=+�u�L:�		_È��b7�>�N����(�~B�b+���������L�j?���V�Ozi��㚓xY3B��8Ю��/ea���F���%�)��a��@�r�G(Q;d�}����J�4�1�o2�8Ƙ̀�A�q�晝�ɔ����h����,��MBW�ؕ-&��͙��ۍCj[`���9˪?��G�%M��t.$-�7N��F������t4z?Ƭ���j�1IP5�U*��T����'�``.� [$�l�GU�#�e�D�Nc^T ,~���&A3�^Y9�c�'|U=W�r��ܷ��*�lfu���=��$�$�vǞ�x�< ��| �`��ĳ������Xk��&�dbM.g�QI�T�R��ޑ���9���Ň (���_r�g�����Ɂ��ɝ�d3|��U����&�!̧��YA&����hw<�F�(� �>�6���;�)P�}��(��n�+���n����/��x�-�5�W�&���:�xd۴]�����b8�����`nr뙧���ދ����G�2 8��n0����޷��R8ک�5��i��[�hǬkcϭC�l5$�=�k�A���f�����DU�duC���3_�J�A��^[}1�7]�s�d�yCѮ	+�H���E])�'Ǳ�rpzB�s�����tA���,MR��W��,�J÷zg�
&˛L�|Y����|BO�z������^E_j���=��ޠ��W�4�܏�[1N��'t���w7T�v�Vz���T����m�݆��#G�dfV?#.i�V��;O~��DCd�B#V=|�?Զ�T�e�R�`K���}����m��JO7�b�%GI��Hq���reK��5P`.��/c�=�R_�<��Ӫe�i��
h�W-���s�:'"���U/���áw[��Y����Y�d(ʯ�p�<��͎pRX�T�;�o��-`��B�n�4B/����sqa7�[�ci�Gc�ha�iՊ��y��/p��>���oh2��J����zfX�./~�TC��`Q���<�=Q��^��h.]F֑]�f~@kCW>'5��-G?��;Q 3�/n������Y�s �)m�\����zX�ׅ�y�UDE�3��3M�A�ک_P���(��b7�R�V���'\�!a<�q�cg`�2)pw)��U}Z�*U��R5��{i�C{�m'vr�B���� ��[ 7�Ω&��8d	<�l M�ԧ�1fO�&*���*ٸ�>@Tj� `��g��Wfx��?� ��������B�kT�Z�/�8m@7�|I�ȭs�d�p�F9:`����U�|^&zt����Z�-8�I�����c��Q��$pA:��(X�q�a�&�r �e�E�N��T� �;wDS��6�	Rr�ˁ��k�)�/�D�;D�nk-b�N\'�8�*�=�N�6�5����|<��h[b��)�e�g�X&���x�?�v��bp��Z�.��?`n��Ƃ�I�x��rɚn�;�c"��?.y����DbO����u��qvڱ�3�;�!��T;&�p�{�_��H�d�̀8�.M�oN�Jzʚ|8����y| ���>���UڈΦt�'6oz"jI�	:��3�Q(
��4��?w�O�fE����z��H�� CU�"(E(Q�rѡ�K�޴�~�[v�g� �$+�ɂ[���sI�l�����:��6� Kw�#���F<�)�+�ˡ�a���X��z��C��C���&�Y)�XS��=�s"wӳe����\k�ƣ62?��:�
̋}�P�h���$0��$,����^`�XYfD�(�yX���gOwOŴ��l�Ag9E�b#�{ b�m \���KmH�'��ԯŧ��~e��F�n[K'����Oǂզ�y&�g����v�싛��#��[�	3`]����'4%*S$	�i2�H�<��T�NYh&˒���oԢ��9�K'��=�de�����vH&���J��Ak��%h�T�w�B���Ȭ�U�A��v�N�%��F��<�	2�.I_�[{�	�E��4(}d�2/x�g��I"K�����5iB�Q[{�
Ѷ�:��L^L�]� %��.��=P�j#S����_vL�܃���:z�|-/�#�w*I"��@䶊�WE����uXyõ�enNod�1\t�qVu�9�4�ҙf|YQ:vŞ��L�ଇ�J�s��1�?oA�VQ��YuXv�3�iwLH�Ʌ�����.�w���y8�����|��R�qR��;+Q*0��Z�R�n�5lˎo�E >p;�z�5MR�s�>�&��0��Wb��?�W�,����<��/f���4U��k��ۜ��.P�EEe��Z�]Z��#���S�[&!�f�Ŏ_u�����ᦪb�C�-�˛���>�,��E�hm�㷋���\��br��ɑ8���F$��ҝ�$$����<���E~I���> �i%� ^�?��G�f�����Թ뻙3I�?����ս�hh����<�푋w�����z��F�t��� ��߮I��7� �DGS(����׷f3���	x	nM ׃];���\�u�ćkq��+1�]�U@'8���
VF�����$��t<�ㅽ'�Ad�s�A=��*Zp`����%�j��$�B�-�2�T'N$��{���T�h����_u���bB�ԛ����sn����*�a��(W�8��S�dL�A��+�0�@�gQ� j��q�� u!���~?��!�	'�������+�^��t����Ńo����-�G�en�n1d&;�,�2��6o�ȅ��ͺ(m����׳���?�b�ر�G����B�6����s*�}�����6�4���s�b3��/F�x�mY^S׀�G�b͢
z/-�"��E�6:a�~@c}h����"��}�P�G��"���!�c$6��u,�m�#<36��z����Y4�у��V�#�1Un�t�!j	�q����3,��J�����y��d�-����i�uh�e������v�a^[:瑠��2�����]�فG���7t\�H��X�� {���ڷK�V>D��U�cw,�?���jvd����9��Z��#�/S�������� r�/���i�~�*��;�����o  jF��*�~I�# ����G�����JA����"r� �k���~����k���l��;�2��P��	�@ z�o�Lz�	�NZf�`k&�øj{9Y�����d	�w�W��F��K�\	���i���\Mi�]5o�#	_�1�0b%G?�EӞ|����˷nv�V;��%��$��� �[�_�T(+g_�0�� ����_���Cdy��E��R�����2@,�`#��h�P��0%��S��8�9�[�KI���"a���8-I�!��4ì�ӯք2g� �G��i^��9n��È�fqT�$B X�����_%P�Q��%������Vn m\�+ƿ��ן �y�L����#:L��T����42��7��.��Y�1]+x���ĭGo�x�S�y�t�S^�"���*�t���&�6�CU`5�B��H�W�G��d��'�g����#E4{���~-�,�{p�,���O�@�`{�j��*���0O�6���@i�7�I��܂%��b�n
�9� �I�@����G� (n����I�9�P�	�iAX�,��7�*\�c���/��Ǜ>� /�>N �'�|e�|�b�;/|0Cl5�>�@�	����{r�S3/y���^?�x�v�wBJ�2�7���?0bC0-}�bK�� UD6i�Ӏ�񿎗a���̿�ћ�K��H�^�>,=��#m�p�[�γ(ƪW���H2�-����\4�	�$
D������&y�v�U�p�%�������t�h��`���Sn9�~}�ȃ�11@B�m�L�u��"E(��J�DxNJ�0���Q}��ī�K�em�X�dX'����Uv~Թ��?���RA�h�ir��0:�N�f����7\�7ꅋ��.�YH����+�wf�C�V�W�@\:�҆��n~/����dF�{�v�0|Ť����y\X"<]���~*^!Š�����uk�������Q�A6���y��!�~�1̈��"��
�\� �܇#d̿�䡓�
`2��<��,����ل��ϼ�_RXٲ�#���}�nT�WUM�Lb�*鈈����'!�9c�:�y���b�g^�/JzH^�PS������P��"���Ye}'^#=@Ss�	@���sX�<�0~��ԍ8�Ид���w��H�E"�F
�Y ������2"�@s8������TV�������LW�$��x���{x�h���R���G��t��5��T5��}�P�7�8;�� 
�¥��Cg�B����/��շ&�|E�a�p���#V�6&�1�;sJ��V+��M�~�͠ش��}�(�k�݃�-C1ϡѠ)���K�p���d��/�R���5 �C��"��h����y�t�0�(:8�mR��&x�a#�#�0"#*X��x[x�g�OC��X�k��'����d����QG�(V�{�Y�� ��<�.?��*���[�2˝�k�V���ʌx돺G{� ���2���ho�t��擝�����O�e��s�n�s�%C�(�sI��#s.���FJƢ}.��F'F�����ʽ1����'�1)a��[�G,(�pl�F$�'O�׃h���Ys��v�ȨՂ����pi�=ux��CeJ�y?�d��)sj�?���I�	8�=�����@��������콦��Cw���@��jj�ߚ�NH�)�G1M�Z���!�Q�HCg$bӽ���Aa �nҚ�/�W}O_��$�̋��zJс�,~� 67�$�7А��{�K�+�͋Ǐ^�;�-,���rtf��ҡo� ����S��O^��A��yG�@<�5��w�\���-vSH���˧~��Y9a�x���.�j�� ��f;释��c���B�J��ߐ��u�7܇.�JĠ�k=�`,=�y�P�(YV7�Q#�^S^fD�����r�
������#6�˭�����N�����3D��a�T� ���Ǘ���H��a/�;�����t�]ڈ8T���[��tC#�6ss�9��Y9������0�I1I��h�m��et�p^)�����,1t�@��(0�.(LҸ�g����_���{��/�(�0��nS���;�u� Hq����E�P������nu�����a��*�O՜��&�c�L��Z{"�+ù�~�m?�M������8��Ƣ"�5�㍒���q��'O��Z�� ��U����u�]���]h��\�wQt�k���j覍~e�CiC)��n5� E|��� _�O�3���4��5����U~[����
u�eQk����h�56����S/��=a\l*�����:�מf��=�ֽr
yyչKt�bs��?�}uF�,>�uL�\Mݼe&%Y�d���-�C��[�'}�u^h��zT-6\k��6��8H�S�	x/�`��A�a�ᾣ ?VL���1Zr��4H�������r���ނ� U�&��:}f�jPn�SM����FE��sŴ<��	wL�y� 񕅝C���&��z�Q�P�y�9L#��|2t�l/	%y���A<#����E� Ҏ0�}�gP��х�A�=N��d�t�Jٕ��e�G�x-�C!�9����p\�J5P'�zL��f��@�%D�Ѻ'����#�udF�Iϟ�3�pr��[l��(����M�z0�de6z��*�Zc�-'Gw�':�gjFa����'?�jק����s��Gn�!�@S<8�8'N ��3����ʗ��O�s�H���6�XYm=�� �c`G>�W��-ذU�J`����LB�|�I�$�Ot����7�"�6c�g6Y$h[6(;�:�����b���M:�ɉ8s""�`��Ⱥ&^�ԝP�.��O9ޕv�ڳe'����Ot��8k�.g�s���>;��D�g��n� �H�v��+N�s���`���Q�(6�&�XW1�j�R&Ri�uf%��~e�L'����_Ӏ���W^5)�n��D�XW��(�6�����}�����i�W%+��r�X�q��`�M��RǾl8W��Gl���YX�n^#*�F��eǪ�[???��dT��_�� %�-n�r�0��WPǵM�R4��5��(�6_�߷V�N�����ĩD}�'��A�Ɖ!���(A9�&1��jܑ/~k�X�sX��&��L3�{JC E�Yk�<�>��J�|��,\E�#Hva�Z�Ǯ�F���XTS�-ˁ�e�@"vd.��K	M':_=m��g�ײ!I
�q��� ��
ң����
��PtՊ��׽<Y�`מD�	p�1I�� ���,Ug�Ky�wp�|�qb��,+�Wղ��
�S��Oqg9(���o���g�w�Y�;���J��X���:��0w�U.Q�U��(T�;&�wlGX��ܢ$�.�R��xAHuI4ָ��O;}�ˈQ�;�s����ʀ��v�'�<�z�z�(�*ƶ�� [~�L�O)�Z�܌��?`� ./�Bj|��mYD��ڰ����4B�JG��B���?!U78���9��3���j��	t�3��ĚP�53Q��H�h�����(��O#�v�'ԈO��X�CI[�I�W��*,���3�[��e|�L#�m�̵9���=��H߽��*�?<�ϑ���B�����K��<��OK9�)�	LV�"u�VL��.�nw6�D%ql[���ܫ�O�����:�?н=po���B��5.�S@(c}��S~�.��Z�����xN[�
�:��)O�"Il���&�,o�W��7]���gS��G��f������rm.��oE��\��U7^!^0D�4�B�:2U�?F�ě�T3jɕIs!�8���P~�$�N�Q�ȝ�I��݁�̮r)��>�����H�qY��-����9��z�"a-�rlJ���c#��=��/�Y�����Cy��Sk��!��*�ԣ?�IPAU�ΓƧy������������J����2�*�� {7��ҥ�d'^ J6��[�$�W�/���h�>s���4��]���WVid��T4��nِ�8>���P`cĢ�������"��a�m�5��%�"�F�+f���������q��]L�[�dR��/_�_R�)�N���wLDP�(��Ltp�|��p��*Ln'uj~͍/1{.�A-�T`2(��0w�U:���oNJ98�RE[�z�<�M�%٫Z`p���Ԍ���&�1q5�%G��
i�g�d�a�T*~o��J4�lJq&���^�?N�$$\D�{��gzO	����M߿�-���7^u�������@�	:�`���z���?���n5�Ye�ˮAF
/!��I=�����ӄAJ�*`���G-�b�0�s�k�﹠�I?�ϩ暴�V:��N�W����X��a�/�\*�gJ�|z��:��kXqII�e�Ĩ�3�\=����' f�E��0�+q������O��y���aRNƙӁ4�xV��3�܎l��mμ��k�_ZY#��KO�6�g�)0�/�=����+�\!1\96?�g
����*)���\[b�,�(����1��1_[�k0!�.�W?�N&�@!��¦I�N;�k���mYRT��:]�T��yc��-��Rh�P��-���лa���	`�A��+��^4bid+��X���|�ז�/U���N
`�$�Iܖ`��ctS$þ�Q�tD���Ѽw��	��,Nn{����=X�A恧^
+��v:>��о�6?�o��A?��iD�q�@^��t�� +o�uz�Wk_�Q��Ʈ�j�uo �,���#R7��k����������֋|t+�痡�u}ZH}1����LH�����#�!����g�Q���S�0_�����
�$c�=�	�z�������I0|��WJV��V��g"$��^�᫧�9��&L�@Ё[�:# J�ʲ�CIB�%�߬���E�L��5"�t���Ea��=�R۷ꛐ��*���D�wn{���zO1�p�v&���ꫮI��^���v
H9�,1QO��A#���,J����l�b��"B���$b�QbQm�b���O,�9�^/�#�T���[܆����>���\��k��[��G���`�|^�fĂ�N�;���Z��j���ژϭ*���Ƙ-�bα~E����eu�I�%/��Cb �=�����j�Þ�H\�tBD���$����z��=�_O��rBV��6g���R�[�c��N�n�Je��ҫ�h��5�Xe�'bD��	�i�i��0�S�Y:�3T�<Dq��C��o��c!�����qX�;L��a�&h5�&����,#M5��ޤ��y���o3���Ů18s���:K��(���S�KA���3|K���5] HW��
8C8��TYR���K'z�u������t�'e�R�:bF�mPc ��.��r��S5B������&#�Y����25}7���@x�"�@��ڤ<��t�77��"���1��^ͅjӟ@d1ي�S�!&o �$���˸Y�ۥ<S��)����єE����6'�⣦�٭������kKu|肌�hR�>�c���~䶻����tE��-�HB
ǅW�o�i���Fv]V���g�$�Ʋ��-M`^�݈����˝q���Q7}7")���*9�z�b�ќE�챗Ƿ,"�<e�eTp�7>>E�m#��Kzb�7��ؠ�,�U�UD�l��Q5���v[�}�+��-*������d{�#��sr^Tu�]�r�ר�^�n�T�0��4�_o�Ԯ�l�:����Y,^���w���D��xCf�s�o��9�6��T��X�W!\��l��v`u5?a]��3z�h�ݠ��uT���\q������i�Ұ�H�*)
�hKr�'/ f��ܗ��#>�ӮރW$f��̾��K*�dE�>�"�4�z��uɑ��GV��
���PH���@��b�=�|�ˠ��а \'��m�NL���W�Q��$��װ�#I.��p��H�O��~]HMf���;���=9�3t��i@�W�Mn5��_Â�ٸ'�+��i�+SA6<ekj��FK�y��Qr9Y7�ˢ�4
��.]�}gU�CP�+
���Z��A�"��dؔ�FN�s���*�rx'��X�`2��U� ��4�h���k�IL]�d�և��{�Bg�,I������
�ͬ}��� ��|��J����-
�r�15���v���a�f=�5a+~�2��D��{�fQR��c�oR}��$���\�"��O��
�6ꅆ��8t8����1oƱ�l�w�'\���Q�z���vu��� &�N�5F�:��!�/=�-���Ʈ����[w��9����Ή�n��)�qFS�0�쐟��