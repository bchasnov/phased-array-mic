��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ��)sZtYzѦ�#����������^{���f����@,�B���ul@k�"T�z-��0��{�oQU�<cM i��CV��Ǣ���j*��>3���B��1����ݿGi�b�2g��8��H�2m��@�}
�G%�p���.�x�T$X�v
��;�b$C����f$����D�j����+���DM�#��k/��|�S��p�k�ҘMw�����t���3��	�ΆLww���LG�\��*B/qR�n�d�"O��
���<�[�ٮ<��?^�+�#�����\`2Y�Ϗ�cR�W�G���	@oU�z%�� �˗�#�fŪx��>��1=��&��mErc��ϿY>g#d����WQ��Q��h�.�8� {J��=}�17=E-�挴ە&0�3HFq���F�W]E:ń�{�B:�(��=Y��َ�o5qxE�~�4 %te���s�6cܮu_�b+�K�s�_H��м����-�]�Ô9s���f�Y�5@�(�:Fl���t�����"���s,*�D|�ޝ�'/J���v5�������n���4��>� W����� ��驣�֢�7]�DÚ�\�y-DӢr�X��5����}'�E3c�j��6�۫�����0D>��Tf�G3�>�~�0e� ��d'ɔl�GP�j0d�S�T@|�;�'���t�C����K�j������E��n1�$b9��z��!��o��1V��%��xh�Xy�����B"�u����hk-)���7�b�ψ�V�*�㿓M�}0K���.��"����6�4�yjᔌ �a�o��������6�1s���S��.��j9��;�;��|K��Z�n�>�W�?ʝN����+��l6Z�+�?Thd���Z��w�RbԲm���B�����]���3f��r�H��!`��B��[`�A�k����ZU(1�>�ğ�,�ˠ`%��o��"�)ţo��[q�3�*R.(�K�g�(��@���"f��ql���h�~(2WP�	#��[q��S�u����9ۘ����|^m��8>�N�hЄ�-�F���\��6��&W}�M�2����/�/��^SzkuW�c�[��[�D���e�Ifk]\�
Z[h����P�^ún��^rU���$l��.�w	P����.DPqU�?3|�zN��|�<�e�_$��B<M~�-$�2"�����߃d�JAo?����K�M'��D������������td��>=�&�^r����~�+�	 ���&w���q���@6��y�5�kZX��dd}<��d����ៃG��	وh�.ؙ�n��F�eV��ܻ�=�0-p-�abo���0NG};�vn�?���{��!�]��D�!8��?.<L��q��%��R���%{w����{�C�{!ɸ,"�<�̧�w��Q?���p�_�\
u*.�CsI.��� ����&�%��Xx�;#����՜�&ab�1�����hL��<��;�A�A#>߿�B����@�`ő�%@*7���(�ԭVJ�H��
D$��w�q���S�˨C 
Z6���^H�p�j8����b���m�K����;^��k�e^��{r�ǟ*;���>Y빃T*�p���,^EE7���b����Z��\�F�S4ՠ'�`%�K,�Q�:�U\g0�v�O�<�t�1�eAl�]����da^�T���>H�S�y�`8�� `��
)��є!��Z���Sͪ� �᪸�E2\��C6r��+���_/j�hf(��6��ꌏx~1x�A�<	��q�y�mP�3���2"D\�RT(�l�G`���c>��ꌥO! O\x$e�}sB��t�ڤ"1T/<�����(~3'	Y��8ڑ/�>8L�$�M��=�g>q�5���G:��.NQkh|��j]�Z;Өwv�/X��e�^@�p�͢_�yv5HIԨ��^�*X�9[-�%>nX��-X׵ƛ�eW��L#��M���U~Gҫ�^%��h6��Nnf��-�6\�#�bD��,�whiSgW,'��$�3�A��u���>@�i?B"��8��Q���ט��^�ܯ�T�� 9P�AS��������N3p��f��w�^r�ûJ�N��͙��L�w�
��*qOW�6��dX} '�5} ?e\�I&���RL�`&�5ʗ�K��aIòN���6`Kwe^M⏩꜠�X�?��y����i �'���ҫm`�۶'߽������Sk����Hz��L��.�>R/�I�����Gn��I�'�qē�@o�Ɠ�9r�u�BIu�N���L�џ���.���7Ȏ�1�;�2����Ĵ��q��3%f��ѽ��н�:'BA�i>ӽ9x)�p�/\�C�fU}�Csx%��W2���i��1�q���|��z�C��r��UG�`b'�[�4ή��؎N 
��S^��
.�:�i�`/�4�\�-�"�Ո5e-���I�.�־��+��4��K"(�y� �<�~����5��GῩi��Lt6�-u���991�_g��6֛f5��rr�P�u����$i[I�E�r�#E$	�����{d�88��W�B��w}�<�ug�tl����1���������5>����ܰP�U1	�5����6�����C�?��a�w/9N>�h�e��N�qB��-Q���k�����@��o�",+�����s�[�#�r_h/��$7����N?'�\�y�Or�v��8QI̶�]�9�4r���Vv9�5P{����xe��W\{�!WK���T��J%��:5�bm��������m��x��эW��><*�����5����]!)�<���~ڞ�MR��X�[�H��e~UK�z7�qV
'e��o����-�ϥ8��z�24���KiH��}\-R�U�����ce
��佉�y�`e����Q�wW�����H5V�[wN�zC���-�hQ<q�m��C�j��W���ϵ�dmA�53C:x8ݒ��MW)5�bEU_r����k�m@ˤ)��|=�0���/�+P�4�q�����w�5�EO$��"�xϨ���]���v���9s�9�J�a�Q>���b�>���R�<ho�tX�_9�T�����5MN�/@uF�4���G�j��UG��� |��6{6>Y���tk������L��M��c<L�ڝ����G����$��B��I��s��_	d���2U���/FQpx�?o�3����5�� >,}����h�.@��s��6W���1�ZFՠ�
y1��w�|����+�;����<�J�vm�ɷyg��z�?.�����B�R�� �5`o�ܦ�e�Kp�*�<Ї4	:ry���t߁r�q����O��ܭ�� 5�z�r ��>[CWy�u��}{��2��Z �$���ף#[�Ae�U��a�M��:�9JJx�ɥ��B���-�&��?ߌ���`ʾ�Ok�;Ɍ�,��bI��1ls�go��IȄ�O�# ܠ�ty�Fu(�������ė"b�����"娎��I��ȗ����;	����3u�4�Q]�+����XN)����6�mȮ����|l�����+-u�����9���1��C����� fm�%��ԅ,�E�m�&	z�Xv�H�+[�Ÿ���<	�j�X�0�