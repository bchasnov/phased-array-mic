��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\����q�?��e�I8�b�Ǽ$��"����ׯ1�V0���ϱ ���u/;�a=�r�PZ
�]�d���$���4"@n��#����Ӟ�D�`�)R���=�"��5�8���00o*A���BDj��#�[�q_���.~Z$�Z>#洃��^�:�?cy��M�p2��%���W�a��:���ȆtB��^��Bgһ��a�SN�9S�dk��麢���{�XDx��[nc��#r�w7�<�Z�!�Xǚ;�YU�ײs���h������,p�b���ך�=!XѾ�^�v���S��z�#W���W�-}�|�5��j�iw#ٸÚ*^�mO"����*��,4 {T�Ѵp�4�K�0�f"�����(��O�0���,]��T+���qK?��?��2P��֢�7��s��0�ۣ}0 c1����΂9���3�/v��E�\Sz,�l;@`g&�?h���,�-��4p�wg��C�j��������y�؊��)�\o���ȉ�/m���ɲ�t����"��p;M���r��47�5����tS�	��q�o�]�'m��y�%Z�|�y"��Xb}~OJo�=������Z2��Щqz�X�F��E����%� �uMJ,nzI����Y7*п�'�? ��*DB>aT�	��!Y��_r�r����Ȕt��_�6d�B�d��^ָO��2ҍB1_q5��v��o�a�&�qW���� #0�"I+݈���y��p���(��R9�!I�$������А) �]v����V��>�݀�G��]��L�N&��hbZ�s��cO j��}q�_^��ݡ�y�l��`�%� !�
O��m�_u�?�������w8��Bi%	���)1�r��ij�]����-��Y�JT���/l_R&�C��N:������Y�#��HM�*��蛹���[)$�?c֑w�]�U��-���<~���	(��<9_ؿ��U������,^Y>8~ƑK�.���Б����\r"|\oc��n�-\�����	��d���Ȱ9�4�Ԩ�"�>D�&m�2a`Rc�9}��S5�2'A'�����ob[�cD\y�^��v�7� ���`:�<n��4��n���dY��w�P,bAe/�@����̛̏w�.�7U�X1�u����A�H���z��%((l��]r
z���$���sJ��eϑ�@�'������ `�4���\G��'ܟe-�'x5��2���8�vS�Ъ��ׇ� ^*�&�F�^a�-:Z �������j�j��g�?�����8㖂�������)��ǥ ���W������]�ҵ3�S:�A�vumb�+�4�-s�|�{��1G����q*��pd����!��r|La�f��	��ZVn��v�=M��ľB��j�d�q����� @���;�d���8S��P��z�o9bb�?='���6*��ݧ��f���ݚdI]��Uz؉��]��L4�b]K6�ް�`�Qsϥ��'�ʹ�% ��?^�!���G�n�4!ǗQ�O_kqע7�S�bp*5��gj~l��Wj-du���t��C��ܟ�u?�G<���=�aE��נ²��G��YA㙒�z�D���H,��g��'�z<��\ď�Z�A	-�R��V�B������3����pt��t�k<��y��R��(iv�u��<&&-N�F{�T̀�P��P������xb�l@�M���\�V4R�PUy��;Äp��{�C�F���.�j������A�`�B�f_�6�K��h���� ��X�W'dS�l���,��%��\�#��LunS�FU�2� )��u����U[�%#��b�"Jt�02
C��z�4@��tu��MP%!�Jq*d:b�+���J�X�N�Ry�g�<&ׂ,-߼;KE��S3@���Gq:?�h���Kh� B�(!@^�p^XM%�!ƈ�	���$!fR���";��~{,��-�_��V��Y=O��-+N���X�����k�P��G�����(kxP�v��j'pHA-��94RrOr��4�dZ��p�^��m���w�(|NZ�������n�ʗtcH3��tV������8$�"ęH�)�P9�* �Mܭ�G�3��d�7V5��Ww�F��gs�c՟.o�T�ʍ�����04��ϱc�B�+�!P�z�[�bn�j�վ��h!�\�th��6r�f��^����C�+u�(N���2鰪Pt���U�'�J=ॵ���`�PE$�I��A�cw�ѵ�b�a|1m��Ӽ�������"�5�HVSN���#�|d�5C��%t#��� 6x��]I�S���@a�&6�5��
C��oSErf��U�l�ֳjQ�t�j��h�kM-;�8j�;{Q��57�D_�xT��I�T$�T�' �L�g�!�ߵ.Al��i���l�xw1��<1w�,~H��K/�B���:.ˏp���vG	%�����j<�<�����ղ%o)�#7��*p:��\W#O��d��g���������s�6H{����;�L퐊��0�B7�͋3k�JG���O5rn��7��>����b]hxu�����j<c��
�`��
1Ecڏ�U�59�݂������M5U�G����ڼ���%/!�� �:�12�����,T���q+3-����Z�����ɺ&����V�Z���3# �A�[9��s��/�{w�L�f}^B�ǋ���gm9��LK�``!?#?����(e�Kb,T����_&�:�ʏp�'���|*����\D
�N.r_�W��Zc�����Fɲ�b�y��!s�>V�����;�,�zw������EF���J�r�������-<��Qtu�|^��,�9��^<5�$�`�QlrU^L\��ψ�\`!����Y����3��m�İ�1#�Ap�����#r��It�<�k(t�-�PV!���8KBֳ��\}�	6���>-Q,Eq����{�:NԲ4���֧_�&�Wfo�o�0p���Ne�o?��|/��l�W�씡�E�"��Ǐ_�9��6Y�'~�Mꫳ�b��ݺɷ��`�"�,$m%�&͓_�R;���&2�7V"/�@��6�O*�wu����%maQ]*u��WDS|�7�Vo�[�3x�v.ʒ��1�1r���i���q=�Qb��'�dr��T�m@`ۅ��B�h�DZ�_�R4��)}1i�����y�|^��'��6��Ȑ?�&��x-u�,��e6b����k������)�e�|���5DG�k��n�G�P��|<(�U�5�PM��GL�(p:���ɷ�Y���E��Vd6��;��6�߁�{VԔ���S�7��[aiip4�\�#��O���:�V�v*j�N��8�ōy�׃HiL��+H5J�n�DM<U��C�<��1!G����;Â*b��~O#���� ������H������v�� ��a�4����X@�KçüLD�7�.)߀�	AnK��џN!k�u]���A��"B]���,%������=l���2�r�r�b�*t,��?5-8�8��Q� �ĶdL�+��M�1~��������d�2	:�F�xR��(� ��Z�\:�q2���F��'�t<���|e���=�y�6�P��s����ܒ�H�.��� '�B}�`�{3F�1��-�x��@p%6�(��GnY���Sw�\H"�[)�w��<���{$��A�� ��(0��Y�u��*�.�݉�����z9 �Q�U!�}�*�@�{�"Y,"��m #�տguR�ݻ�Vos��J/���hc��S3�>W6��V[ab��Co�g\ *u��2�E5_�6A�(�}�����E�_"]��x���>��tO�+���*F�cuB��i��2�T��>\)�ou�.��a��k��c�q��i�߮��AEFt��;��̭2�
�@K`ۈ�	�Ȏ��t���1}ϏcH���}jA��珘(`�EK���sb�y���よ�0VW/�����t��p���i�K+��p:-=�(�HT�*�zA�1PG	�)
u�n�zк�>1]0)�W=!	;}�@�9�p�e&����1w���&=sd^s)�ok����b֬�[4s�#7*5�V�ac���N�&0��K��?�e�2]_qՂ�~:v8���p���(������6?�=�������=�0�{�f��sgUa���|6���J�E~�8�ɥ+M�b�'�D�1�e��i���4IC�,��Q����5'���%���L ���H�������� ƕ�|lU b��z0�����m���^0��*!]��F�|<�W�`�����d��&K�\���W�Oά`��Q�n	�\\<�u�2�6?�1�ռ�!���*p���v�#�U�[�)��}�A8E�6����ǣ��_��z�o��j9J��zazs-7Iq�]�*��=�7��4�-��V��f��/�P��Sxh�Z��K��dS���bm
���˅E�7�9
MZn���Z��@���F�fwHH�̽fʰ�|<�H�}�eؠ�	 �",g���=����v����)�����
����
0����v\{!�ؗ�(gPl�S�|Ꮲy@%���E���SI6#�}Hŉ���8�F �4�*J^$��Ι0̰J_��+ľt�R�Z9���Ɩ���)�t��՘@�a
��hn8 �byt�E�1���q'1�1m7��]U�9�|4�Jԁ�!���j9��c@!ڀ�����h��Q��l���R5�����35K��$����:Y��P�����b�E=;a�	�_�6��bu.Y�G=�Cn����U��M�z��$�>�I�Y��o��W�u =Nˊ��N�8&}�'V�djzW����7����q�|�Q2L�8ә��Lt�$o:�!���m�ֵ;w�Kь��y��Y�m_�s�Zs\�[,�A�	7cL�x�x�ƽ��~l��3�{J���o��x:��ߦݚ|�f�d��Q�,�ml��K�����	�¨/:����ulD,P霮��t�4Mr�V�u�����CYA�wM���@2�fs�)ڨ���>ʉ%�༵�:�e�P�,5�H�1j}l�N;@Ӫ2���*U0�������ǭ]��-"�wۉ-���U+�`���js�|�
?*&_��O���e��'�����ۤ��a����ý����/O�e��>�#�Y���>!p�|�SH���d�~/ki ���-�%Hu0,�$�?���1Y%�����A��G��J1�:U%|��ư�QM�+T���M)l�]�2�ݰ$`z�t�Q�y��8�L�E��4�J:�MK�O�eV�$IUlv��?xɘc�Ś�;���ک��AO����M[<y�<���mJ'��jpi�y�x���Zb�~��\GG��f�R��{o�
5��jw�S�x~�@�`�(o~`��bAeZ�0\���{���\{d��Z�u5�MK�=�7��&!�Xֻ�����//B�[|C���ݦ�.���R��|S6�͡J5_��p}NHݜ�E���ƹ|�:���$g�*����Luf^�ӭ���B�H�Sy>_3椰r��'���8�_��t���]v���{�[�v����*�:s��$}h���ءW�ʉb�	�N���Ɯ6"Towb����R��n���O�p�"u��V�3|<�dv����M`bn�:��67jlic��̍�^����R"����[����o{U	�,�Uf���2��Ib���{h«)�+��F��dZ��h3g!�����j���
�Ff&�����c�椓�/��_��(	������)�M&+�����7m��O	�^����ai�"E���&���9�}�m��ԯ97Xل���ɀU͠Y�Pg��/��Sn�Q���l�R5@,�G���.Z}�n�!�%l���>7&��:�;�H�U�ނI;B��4I��~=�,g���|�E��%�Fl��/]�V��E6gU�->����89;�{�}��\"����<�v������Sy��~л�9�PQR������)~ޠ�D7��N?
����[y�=9��yi�J�o�Z��	��s2 Ϧo��>�l3T~�����L�YCB��,}+)�~�ύ���UtIƎ-q����L�5�0�l�9��	�a�B͌H)�d�W�	�]�ᒷ��e�N��C������������kRp^��V�y:^�d��D�ԥo��R�M�hUc�x���y��4�g�}�Ɵ��w���}!z�B����t���n/%ƢCz�Ko���6H
�[9SoR��`��0gJ�,�LO�y�Z�/�[w��(z=�,�c#T��Zm�W"��(��(-�> )w�A����vtJ~ht�a�&KF�Ĭ�؇���kl�|d/	|\�=�aRr��␤3��֩�Z��,��ic�f��R���賱���s"��)g_�Lvqؚ�^�_y}�_����\�>�\�[w��<\���r���t�ո:�|��,���<�J����z�8S�pө�!kz��Q�����g��Q������l�c��:�On��=�,a��#�����v7��ʏ�vL��z�.ٿ�6����C�|�������F+�pY��yꛪ���8�5��
Ў��U��y�c\}�n`��׸�i�V'�@+�S���3�Bvq��aR���tJ�)#�'`PōӨD�HQ�,�ϓˈd����2@�pZ�.G�ɰ���p�ω�tB��b��ο
��c8���<T�UV"�U"%� �y��F�L])W��	s��N��*D�9�I��]*9�8�`�&���J<�P�)�0c�A�*$��o.ĵ.-陈�����ܷ�¢�:��Y���ՓY1�ũ�m�(ޢ	�}�to����D������W�(���Ao�S8�1|P�b6�{r������R���+e�I�M����*\+wC�Դx}���`ZB��~���_���e�6W���z�j���v�c�K���j��HۺCs	`#�<*��|)���S7�I����m���N������5&�jy���xv7B���������5� gG����ui��
�c����-�A�)h,[���~͞�'�h�W���n�k�#\�,�T�ۣn͠�p�n�6��aD��SYw��|��7wq ��0��1��`"9��&�C���̴8��1����!��	[��ƸCs�5 �A�o�?�y�5��&;k��A(R�"��_نA�Zp���L$�E��Sz�m���c|�x�V����k�?�oGF{.�g���K�\��,���M�Җ���l����^�Q�jD)יƢ�'�/�M��~)
CE_?H_O�Ф0aBW��P_�<GL��4n?z^ܷI.��H�T.�ǎ[�g��O+S���1v�W�Y���u�V�dX2������ۜ,@��5�ֺ�"�������^]��F��y6�V�)�2��6hG\���#i�4+'��ٔ
�H�5u;\H'�T�&��� �xހE��?�&�z����kb�ԋT����@���~�u{�5��l�^~BѽA���Hm:yUŋ_M�11s��g���!�C\��ʍr���{��1�BD�~;<"�_���� Ox7��~|�6�Dp����֡�������a��M��E/�/����$h����0�b�k޾�wֹC�ƀ�a�Rr�()�)W��3%9��Y5I�x��Q� `���n^ե�#����Q|B�s�H=�a��ɱ�{��ۇ��~>�b$�i?�P�*����YǊ�*W(��s+�	 �@\���T��#�un�`,n���/��Q�s�Z:�vk3a#�1ؤ�u:�l�a'�}��Z�O�	C
ѫe_)�j9-rh�X�&���"K�)��xb����]��}��e#'�u_eEJ�rf
W���]������fXk���%�L�-��d	Jґ]ROM��3Gi%�p)�q�&>n~MF�O��
>2�+��~{X�8���\��3$Y8�;��-w�24��H{Q��&J��n�1�t_�ǲ1
!�#9F�xdV�^=l�.J��+�t���:'��-��4����7j%�4N�&�8%�U�i�y�����B�*���0Rt�&�ɷЏ�����͋[X��U������QPZ�)�K�h`<�ˍ0��|[��]o,��u�(E�+�T���P�_@�����l$?��[.�Wf��fg�%Б�R�+���81��q���\�#�VϨ6z~�����z�2[u�&�=lR�Wr�ϖ��"�mE�G���nZ�@���Iڭ�.(�ڥKޚ�Y`�q��'�����$Hќ��-XW��v�v��{(O�.ɇ��N*�U�r������:�͒F˿��f~���J�q���#U;�@�[�)�ge�T�-�zMP���̅x��zH�^�����m����Ut���2�e���d^�+A��B�U�V�t'��tW4
Pz�ŕ�L�Nv�����ʴ9:{#.�~Gʶa��t˼6 ��s��(ɔbBh�i��=�e��~�[!��A�d�=k��iU�£�;L�,.��`۪I���
0�d��N0#Z�	�֋�A�>�g�Y����2+*�jZ4x_]��k�|���O��q������L�6�O��n�����w���?���*�����+Hݨ������/��"�[�ѻ^`��KC"ֈY�����t�-"���u..�8�'w�U�ۨ�����]`_�T~��^�X<tji��]-S[G����$tv��W�G����f���r�X����j��-���;�3�.�7��v#�c��	�W�d�F��7������yJ/����Ƒ/r ��(3O