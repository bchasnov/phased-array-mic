��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�]��Xȭ��p�oȡ�;u0ީ�^�)�>vys���2{�L�~|c_Iy�K����-��9!��\�Bi�D��{�Ԣ��r'T��NjH��ဣ]��9��|p���4d�#尭�ǕmpC��՘���z����m�0��X�fծ�+oa���}˗!i�v�:¢#�������B�JCv��=�g��
̟��I�Ɠ�9���!l�A�C��č�������kC.�t(�yZzN:�8��mݰ>��z���I���JD(Gg�6Ә]���I����"bv_�z �@�}'�b���!�j+XfIt �堡��;:Z ���fTĿ����6��NM;5Km��������T�`�Bп��S!+�����M�o�O��bf�S��,����%���4�`_'���d���ۮ�ďD"N��	�f]��@��54m.��c��5%I�d3�>��JZEz��Bz���ѫ��N�M��S�](,ݿ�!h�QQ}���n����9������s�tw��J����5=_��aȷ\����蠵\�,������K�������IT�C����$�P.kB�8���r]i*�*��K���"��,��}��(��v6��S���l~z���"-ɤkK��Np��T��3��.���;oZ��w�:PSh�+	2��y|m`�q0����Ħ��ř���� ��]jcV
�D%�}W��G�C{��==�A�R�h�,�:��D=�';�K����s%$�G�ّ�2
�,�`� �QkzȬ�Y�m�ŪS�^�pd��͋�E��v�X�U،��V���0׵�Iꧨ�$"8��z�l��2�,��H\y���#D�؛%�G����$3K1�����T;/V�L姭(0uC��\Л�3��[��@�qR��D���s�;}��� �#�輏���v���^�0���S�<����w<��L�[��E:c����֣��dm��gR����K>^��na�~�:��c7��!n����ی�㣖1��.��k?�/Y�"�֟/��󪐖��@����l��W  �`p�.�����_N7w�~��:�n�$`G1���-0�`�r�m�4bgGR�_T���'���.u���-u�)��k5�à������(����0������tE=�z��UjU�Nv�/Q��WcV��`5�83�4e~H�Ż;�d���1�=�c��$��p0[ք���x�2q��`��Z�ﯸ�k:�T�9��y����T�N�Y��	�g����<d漹��m��|/��΍C¸�����a�K7f�-���;Cx��}�<��p����Ew@��r�GH�k�h�{`!�hp-�[��=%]e��[`�}vCJ�Qg�Ԁ�<�~�w���6=��SK�Û�;���L�eV1�P�Nb����-z]$Xr<c4���)�����2�+{F|�R�d����	0�cP��s��b/�]T���*�:RI�>�uv�R��*W��2���e�)t�Uޞ)��s)��`��,*c K%�;0}p�$��n=�Da��']:i�B�#���8����N0T�<,l��H~��J���K�ԉ���<�o.�}h8��� >�
d�����[�䍩�Z@�K�-[�?(5BУ?�eR*#a):�Mjz�Z�� $עi/+�)6٩w�	�M��)��򘏂J�\�"7�M������N�e�H]4�ևu��� u[e��mv,�W �j��i!�}����A9�<����ԛ�ʾ��=�΂y�.Xa�VV4�jd�,��8�iw����Qzp7
oEƧ�����$9��x$uQ}	@Ik��F�.�tDb�Ԫ�߾ l���>��� �~CBU{�WFI�J]��g�fU}���ֻj$� ޵V3�z2YX��t��-�#h�ِ(�58xʳ�F�j�4x�c#f�z{z̋:�ކ�}�!�1Z	���/��� �tM�N���.'̠3���PN��y��ܫ�s�>l��.����r�'��O &t��Bx��y[QD�,*�ZSC��	=�yT��9��b������Ԋ��.���:�^sQ
#e�7�VM��퍷*��]	�	2��~�]6��cL���H�<	JQ1'��?��e��x6	k�R�S�5��<�܆��EJ�O�5գΠ?uw���0�X��3��t �dbG�u6�z u�^;�n��Ts�
>j,h�ew^��I��'{ޜ(�
h՗("���,?CphùvS�z^$���ö�A�d�^$��qÑ?����ݢ���;\PQO�|{��f�m���v��;
��]z_�X����c�2�Yf0J)��4��W���EΝ����j�ǇJA��G57�6�=8ۑ�9��ؐ6 i��%�k����Ҳ�5�_}�:���~�G&� ��?z�g'��sx�����P���=�� ���3���evs�d�E��A8ӈ}��<�&��u��7�l[AP��?�=�L%�Ht/��*��T;[홠���W?%�N&�hbh�!.��d�;�~����'�.y�/��<�y��`F�8Oz�_�a$���*���𥔿\���@zL�Nz6;�j�V����Im͹P<�x�J�ޑI��^��2�=�OB�R��$1/=�MτM.���L�tS?�mk��� �C-ӐD �-Mwj��Mao��,~QJ����pA�d�y��(4MZ��隦����j�C�Υ	*���]�*N	B�+v[�V�	������̏ߦ!z�WL� ՠ�I��:��5�0��;���"m:c��Y_u�H*�V�6�V�#�?Է�)�.]yZI�r%K L9b5���A�ꂐVK�:O ��[V'+j0��2���@T�(� \����͎D2�3m?;�I�]4&��({?�.���i"h ����wH�e�$v��jsU�Uӷ��,>����p�eP��(�q�k5�F]����?�S�aNL52�H�0����}$�ft7�瓘k��w�y5@���G�s��[�{n����c�@���^���"64�X&{�����3���QD�YZu��=6�s�zn�$hW�^�7���Q�ݎ�j�e���$�k.3�>�J�a~���:C��-���ə�(1�*�4YO 1����,�16^�b�I�/vz%�6�Y7��ݦ-��(�u�]QXgS��B+<�+�ª���2nR��H�Os[����@9Tч'�����c�v�����D���y�C�Ͱ��i�[`�}�c��2�J���t*�"^+��_�J�-B��yʶ	�A_lF�U:ߦ��w��I��$3=Q�� �X��1j8"��� a-�&���3઄�np��f{P��F��ar4	[-K�]��Lz���Z�6��o ���a�y����ൟ�:y��Q�ܚ�e+�f
9�065)�}:�
Zɼ��M�r{�)��ׯ�p������n�m�{]7L.Kx��;�2D�pt~]�vX�r7i.��9<_�	L�B��$���<�&T:�~x|�Jg�k�*'�9� 7W�ĥ��<&�A���`.�ïf�hr1C[�#�:��YEj#���%�L�;�����=��iZq�)�E�pm7((�˪5��WV��~j��OP��͓�?ɑH(����~MÜr�e�ƣ�@�l�<�d��*_� B���]x���p�]L#��3e�B�i���IW�V�ޡ����4����|)��QMâ�{Jj��y�pxu��l]���1���Gٛ���"�%����G�zyU}V��7�jA�|�n}R@���L{��gմ���D�C헳�m�*]HH���j(l(͇�� �UO�P�=ƪ�r9&79$_N��~�>F�j�g�U:��6tI,N���B5�%�y|8gQ/�&�Dsu������6�	hߙ�yH85�Dso������vG�>S{]�1���K�9�<������e���d�������u..��9��|�r��H/
�\�(<�Zl�T�+@�2���Q`h�.�ֻ�vyO�E����x��]��5�R�c!���e�g o(Xf�	�"��{�i �uO���!�I���P�t2�T#��Racj���:��}K���QsO��Gi6�\�Q�n�>�x@p5���Sʀ!�W������V�?��!�߲��Y�3 yI+���c���Ǔ<Rf@V��FUŕ#YG��DX�Q�{"��k+w-ն������lX�5%¾sBe<��!�!�.�  �"R�EY�:K5Ji���M�xfQ]I���X������jQ�w���Z"�Ç��;}m�X�;�k��������ɞ���E[�|:*q���^�-�
}����~�'��L���a����"N�&H��k���Ca�s,���S���ʘ#.q!kW|q�6��˭.&��n�-��.�]�Y�N+������~B47ʒu�i)���`�	A�m��}U�Hw@$�_�4:O\ҝ�(�@i<If����ޭ�ӪY
jT�G��@��/{?��N����V��6�eÂ�pտ��zo��4��{N��bЯ_�h��`��C������WT~5���'���$���h��$��9K�[#���â���A�ͦ�D�?�@�uU��"j�[,k�j�U�R��{�O2͸��K;�q���*pY����9��~�5������|&a\����=�"|�b�<�qT�tZWЖ�'5sB=�%�l�.\cz�J��Z9�^����/��n]�x�
�:��	���GЭ��a$�� -�����(��F�K3�?�\*�1���K˅3�����.�W�P���?u�
�p��ϫ*ύ1��Dٝ���x:\�^�rK2��S������/@�u�YS�奷�l4�T=�C7�pHf��zҖy�B��F�a�iJ�#�$E
-v}eP�Ww� V�}���������gF/G��BT"��Q���U���lzSH=�GCK�%fS�>��^��ߺ���؛F�.	�#7`y�7o��J_�1�Q^�ŗA&\�=��W�i^��l�ت�X�x� ��Y�����-�F���P	�8�{�K��-�����hWx�������S�s �2�I�:ވZXw���G����۰�jV�^��3�`v��M�v宦���/��=�-�>��[�0o'*���h������5���V�����*z�����m)\�[5�Ii�r�a�Vq���c�%������kWP������H���\�
���:�Fn�$ɛ�k�lm���i�wuH,�'��
�J=�TAo!_(�Г!�mz��"='K+�$D��$en�E�4!V��G��-��$v��%H��8Ͱ<�I�H��x�C!�N�j�i^�l��ź2��J$����v�l�+)�^XNT0��+�g����c2�����5$֡!T�X�����ym.��>ǆG!����:�ؑN��3�k�d$0����a]�L��-�0j'�P�<xu�fj�gS � �ϳ�)�T��2�߹�|��6�1d`{`����QԀ���:����Q,9�d�G�N.�L4J�XP�T����P����r���φ!t�@�����=9Z�&̮!35U��C�yj�k���C3��2)�ׂӳ��v;�Vn��u�׀s����Y�ƾ��l���
�� ~/�$��,8�J����tQ(��d��6SP&�dݢ��n��=U�f�f {A�p�gV����$/ԙ�Ӂ���4�]��+�X�g����-|2�a�e��i�<��٣Nh�L?��H��.M���j�ɾ{U�m�Q	�����z�r�����Y�,҅��:�E�m�h2�|���+���x'g��`������'얫����O104��4�F��J$	\CJۗS<]t"�0�T��Z��r�˟����&��ñ��[H6�Mt@\eU���EV7K���� 0� ����dϔ�������Vb��j� t>�.��
å���d���MOY%c�o��4pW�V�э������2O$��'��c��|�0�|�M��tA�VP�=HH��ռ��D�-�yMʋ�#B��dq=�äu[)@�ݤ@��3�y�VM�1m����fB]*肱� �`Q�} �>m���f^4��^�������r���c��� P�uh�������똗�4��ǖ*�i��z��nm:[�eO4+/���t�,�y1$9�B�@	ˣ��é���X/��@3>r��ÿ��i�*!6]:�����?����i�T*�ʲ��T����!�ۄ��Xg��N,���Z�?��x��Vn�k�OB���l�C�Z�}Bx U?�2Pۢ�מeC���3�9��%F՗	��H���'��������[Ab�JWI��-{[�d�9�w��;��z�.ԓh{���@s/�y̢2����7�g5ɣ�˯^��60mG�Z��7���?�႙��\��R�xo�c�Z
�K�C����>��A,�jY63BBBP��V�W���\���� �ڍ"2]��:�R矚���a��yO���%��=���?������~w�qbk�A����f/���|~[�@��3l�j{I�|E)��ibG�[�������J��a��`���
��=�BS��r�p�WEE�`b-cE�c&��n^���ǂ5>�l����Z[�F��C�2]R���LQ'����{�6�f櫒j}A�o�,*�9�̂�!�`�wJc�G� w���'r�7���lh�½��y��Km dl��A�����|�H؈1�:|�q{�!�&Ty&\�Fk��B,�zNOu)����8�Q�Y��N,Y[q[v[tǠ��mw�}�@qH`�Z�Í'Bx4�\� �P
�4�*�ɔ��+f��p7���,qu�������؜��>���#�t2���{?���"v�S�J: ΋��F�.t[��]�����Ej�,��8�w�#^hŮ�� ��еZ��t~A2�����=h�����<�F/�~
����[��1�hw�iU	Nǿ~mc*3���ULČ��_3�wk5òN7b���PPD�c�C]ܱ��@RbūZ9\��H�z����St?�<��v�T�����.:�q���'����&j�O��2,����͂^���I|��uWݴb������ �dh��?Z7�=��P��TڪuTB�u"ܥ\��G�͆c�F���di�h��#�	����ގd�{�I)��M0��������a�l�H��|�ƅ�v������/��p��G�ĭi���`�6���Wp�i-���4|Eӛ�7�F��{�:����,�t4��J��Rc#B��\����QY�$fy9p���E��Ě��W�AXdnw�,��-�~�.��׺�1���������%aPWv6=�s%m�5&P� R=�f�8�}`��;���Ts�πC������>�e��8�"��,{:�,v~�W�1�"/-_gr�t���D��E�.���t���n��QM�����vM��ָ�NoabW38����$���e���b43S2��a^�o���*+���Y���@L6�wrb�&!��6��v/���W�e;��I�ZK_kM�)@XI�l��{.�Z�c{Q=�����/�j��%"� �%;7����wX(�������J-#��s�b����}BZᩥ�o�H:ꢖ3���$REKEo?:�5\�ŮhB6��q鯲跿B�be��� Wj&��;gD���-���	7ɍG�0h9>1b�(��=��>�ԓ��~�}��t/o�:=+��̭�'�J��/�}��iL��)�w������L.�&C���[=��ܹ+C���v�/d),�5uLj6�h,��F�B��Q.��5���ޮ�ݯ���G�%�2 �����'.o�L��L�S�%��$�A�OM�tX
�!� J����L^���Q$��bz����~� ��I9���me:���Ԧ.�@�9������9Y�s���2A���'�6�&C�<A���t�7�n�S�!(���(�����)��/�+n	~FE�z2Ί�[�U1�̌��ǎݜ���	lx}2�L����l�;�&oܔsx+(�o:�ĵ7�����Tyv'��h�8���ӡ��K�4�f_۷�����Y�p��^;�Ap��z��6�eQǸ##�kj$ˈ��P2�5m/<̈́z	gA���&߷��<�Ɉ��9�kןu+�aK \@�4eI�����QԦ�O��X7���X4\ Ҥ48�%�A�K�Z������Y'1�?����l[�_f���=Ty/������~�UG���5�ľ"�!`�_m�7J���c��zՁ2�PB�;^������KC�؝=ܔ�I֌+1j�]�v��0���S9� 	��0�Ag�B吲�V���*A�o�r���p���}kW��52�\�R��n؛Ǳ�4���9�P�K�H��9P��I�l�"������T��}��(�mo.��]RB����8(hgRV��k5�̑	Ӈ}cu�+����� ��	�%,�;��AO:�v��O �g��3geU��m�<[��#�C`��B��JTT�������^/�u�E�?��s�o�Y��9�k�4���c��we2�f�	���by�0������8f4��