��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|>�qT��>����f!�r�iQG^Ѥea	�p��;$l鿬$�����ϻ��J/K��2��DJ�b� �d�$r؟�(������-�����R8��Y'm��#��:���
�jw�Ey���m��\��1<�P X�B"h�pe%�Y��˘m������^��lH��E�ؖ�&��m�
1|)j;IX�V��Ti�rC�� r��J���Y�}��Sx՘�O<�3K�"�Qei.�Xl�ݗ�y��]���իr�O?�Q��iΪ}�q�S@�P��{΁��&^h�~�K��ZG`�H�("�$j ���ͣ8�b���Drd�b�'i `�.�7�5�Ë�����-�3"D�'�&�ۘ&6(ۋ��Q�� �\!k�
w��̛J��Zn׶���;�H^vGF\�T�=��P}�n�.��5q�f=K@�����s���oi�	�2
�B��G�4���H��Տ\|5T����a	o�x�_�G6rh��0'�u�RM�Hx- �%�╉Mc~��y�}2́�S��\�.���kxP�ʧ���ϵx�iG��=����9>'k���ӑ]gF�yk5ɠ�L~]���Ν�fJ�o��������޴E�e��)��
��{���v!F�'Ik��ڛw�'�k�wϙƀ��kF�!A��#��/嵮�o���`����s.�'L�dH��:�!79R�ޯ�R�g��zT)#!'�5K�MCL%�6��x�m�?<��G��O�8�/�5��Q���9��/��I�%R�ڥ��B�u=�0J��U$T���Hnl��˨i�V]T��;6���_��Z����-l���2�d�]'�$΍N�l��A�@���i(��գS����\����G읮���)2���p�8&P�e��,3�!�k�}�3�s����>�w�-B-\�\��~rqrc��{nқ4T����f#�o�J�Mx��<nl1&�6{+�ɵ1;�C���~f?�⦁]E"�7G<��,�s%��rblx�Q9|"!�_�ipp�z�V��"m����y�0ZID�"B���D�J?�D�I��q�{����uq���+s��7������ȋ�M���ym�]��gW~Nˠ����o��lK��hd1�!p�	z� �ΧG��z�RZ��$�R�<�
��?�"���BgE�?:r�	������ɣ�2p#.�?Ա����<��T��c8�����8�w�S|��#,E�Fp�mi�+,��&(��0>L��(ol=�RR�'m�� V�^��?/8s1�,��l=��8b�ZǊQ���F���KZ���h� ���b�aW��0T¥�AҊ^*ٔCQ����#�pV	�N�'n�=��q5���"�x��m��o����m��!9�-\�0�f,��,����0���q���	��s�mpJ�5P�6�5�-A��(�O�@���L�}i�>�/DMc�'*9;o$Ɩ<���^���᷂d�6��h�5�d��G��a:DώMx<!]��?I1��<\�Crt�A��8����-қ�i$�L�Q'�R�-��΅ֆbC��y��Ѫ{���sB�"��q-�B����!�����q�z� �x�wL�yȦ�<�RB��-�Et��.i�ו\�EDk��b��e �	�����	*|�� ���W5�����=���~Ҧ5�m��rs�D*q�a71�s3�ڟ�-���=��6�$�7AGR����(B��sS?����D����1���w3-���i�~w���<0�aސ�F�2����+�7��c0��o���A�4\�r�ڌ�6i�;�7�+�i3��������?�RXl�/s-�$�K��f��S��*_�(E��;�#�3�!�+w��ΧH�.��=�D�E\�����u4mZ.�\z}��[�&ٕ�W���;( 7ḩ���.H��G{�i�4<q���8��P;�yt���
l�M9��$�ZI�uem�F�T��j���~f0I��o��ʍ�D�(��:XU���Vy��u�x6�ᤋVB������o�~��y����%r��� `��I�^��Y_�������%�qܫݻ\�֏]~�Q��&F��	�؈���R��M�aC��v��6�����k�pë����P!�#����+}��,F׭��2����Yl�SSp�VR��k)�q���&��F7�H�&%�2|�M��p�&�h�<�R�$�F����܋2.�zM0%/B����L��%��6MA�+PF i�OgtL�ɾY�/ﯵ��h�k˷h�

�u��.�5�8�������w("�J]9�#����bc��?:0��k��S6N����!:��AT�h�R�S7�ᜈ�z��wW�"ˣc�F�/b6s~��V�.�fvǤ�t�`!�1��zr���� j�}A�&���s�Cgn`�>5ԏK6�V��#��9�m;u����8g�r�|���OG�����|��$������ڣ��G�WA�1n�b�?�4 .�<=�c:/ ?��H��f��� ��:nH����*��ȋ��أo8�}�&�ξ\�>(��̺+��_�O�KC�R�!��ʈ��|�4��5�ޕ]��6D�N��e����Q�B�Q���3A�ʌ���dwD/S�f���Jн|��R֞N�C�NP"�K
D��m�Z
�d1{���d��B\��\��Jy�^[yeVI�X-��e���Z]�B"�L W��\�z����G��-�5�H�y����y+�~��SDk7Ky�T`�|J%Y�H,�ٽ@yA�R�7U�z�W%}+�ޟ��1֋B�AB/I�C��Y�|���*T�
?��q�H�4㢂��i(��2���դ�^����f@���;j��i���!�ʴ�dRi�!2�md���g�m���x����;|b���g�H'2<������|�VK/������Wt�C[�0_ѯl��[���:\S��-�s�Bﲐ��~��?�~G釨Rŵ��/���~�>��u�Ը�%�TC]EÛ��xXK��r�m)�D�@�|��DZ��u�s�F�zL+2����p�1L�Yp���2�q���^X���%���~�k�Ƶ���h���̦�����(�W	qU�A�(�,w9��U�=}������C��;g��DP�R�] ��t��˒,�?�iE��M_:2��(�B<��u�$�U�e͊i���)_#U@;�v^W�>D����y8Z��	嚮4��G�N����Xd�Sע�׼.4��N	fԍւhv�V��b��TP�hB(�*�$��c|fҙ�
�X\������720��N@ӛfNb�c�D��нܷFa"���,�d�,���{v�w�Ln���-s��`!<�N--�=�	��eH�F#�HW�h�
S���OQ�ʏD�'p�Z�/[L��=P���r��A����o�M
�t�ҐU�k�~tj/�\�p�U�?"���ͷ+����*�h���(��$װ9�ĝ��!t }��}.��$?����L�GO�\�^��R�E����dj����Ù
�hd��x_�3*;���mIK~j�U��	w8�-�`�@Bc��~�s&8fy:���1��1B�?��ud/ʘ�Qf�?�&����ؐ�VV �I���!y:U���v���fܹ�5 �*�m�_|�Ϯ�X��+T|�dE.
�.>�m�ޕ�J��X�F�`���~�IE&�DJ�:�B'Erh���U5�$����Tm��
�Yg�i%��-t��d
ko^�*�J�cH�2}rš��Й��+�k�i%v�"=bڨ�C��DhEDز?��Ah��VFtP��9�]�^��,����