��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ���L����ѳJ���ף�6I	��7�"�D�}ے-��KpV��s�h�n]��[��;,��*��_�H1mTu�<'�M� ����Z�H�H�#����*ծ���p����*�R@�>���Vx�Cl/_G�b)�z)���e5��=")D9d��R�d0�� x��Ġ	\�{���> �Ueڼ{�g�_ˡ����T�x�\mB��޿8x][������v�	1)�X}� E�� �_ð[#�b�$Xt��C�
w��bGe���ʹ����UG٣�ɹ�~V��e"ѦΙo�ɱ���0�-�y�v��CPܼ�Fڀ�2@�E\1l�GN��Ϣ l�iRP'�ϙ����Y������ T�*�g���DO��� f1v�\�w������Z�2���8.�QV,���W��K��� *�,�J�6��jH�;�B�n]��CKxv���R�i-IJK�vC�?K$�Q�Ai�L�����I��L1�Cɂ��[�������x�9ئF��ty/Y��Tdto�	�^�S���/C'iy��^�,��)�:��K,϶>�e4��D��#��#�a��ÉB��� m2���pv �Ah���q�ݩ#��?-����A�1	�)W"�"Q�T�y��]�,�V��~���zZtˑE�qv��C������+	�i�����Kc����|���F���o�|B5Q�L�ν�!������q�"��?����z���AL8����B��<�x4|��<I�*��m�}��E�r{���K�B
�8� ��p�P�ĥ��X���@;;%lcKrʓE���Xȉ+A�|�7q���vI+@���dK�K���.B!xW�����4��P\�T"�8O��y��_�e�d�S�7��+W�B+��ZBf��Zb6�u��8{�~ڔx���p�c�b�i$�u ���/�x�S�56"�Je��Q¸������Ces�(�u��'�<B�:+= �Z�*����_�I\�IAwb{�Bg�:�����6���v^���E�L(�C�y9�Ǹ������8:$DKFNa�᧩�׹	�O����yrӃcu�9��t���tKc�����׆��D[n�Ĕ5��֖�6O[�<����*Kzڝ�<�N��"ժ��HO�R�ɮB��(l�K���� #��'T'#��o�3�7�bT����?B�Ȯ@�:2_��L�����-0�Tb�A7�fl�sn)�6����]od�<4k(�����:S��e���_�>l�.�Y��@P���8@���K�^���j{�+j�|�K�^��L̇�|����N��P�7�B�}ǻ�J�6�7����ρ}���s|�!A�[
�īB� ��Q�g(�5�a�&?�55��q&�Fg��%�x�B��܌N�\�J��>�. R���@W��	�Ơ}Hu_�
���*�h�7����Z��ك`�XR�q����'�/����F9P��b�D��ÑT/�3�%�R����o���?��� H�VC�v�nĵ���Т��M��G��T6��Pb6�>�
Ű^(y]F�W�<�6X�~�eM�i��OO��{w�@��76�x(�݁�a�;�Cvb�+��e��ELOZ���R�?�R
�I�)X�����f����4rx49H���kf͒=�����$�ħ�[*���T�7��ɢ!0Ԙ��S����dƜ�,�|KX-}��P��4]�""�; E��A,u�R�U74�oyH�:�&;@�!�{�� �W����U!�6��(#����_�{'L
�+qYG;	�f���N�"��@N���:�k����.�Od���2p�9��l�r�
�}*�j03$�y��I�8��>$�����eŗ��7�h�_�f�ӳ��ml���`��8�"¬�SI#�A~��{K�S�	�Եm��ĭ�x��|���plL�U�UC�W�(l~�YǗy9�+e�z)c����qy���������E���ƉT��֞��LnG��U+�G����,��@3�+�#�����pz�,�&^|�����I���� ��R(n��ø�f����?���-]6�pϘ99&�i�|��}e�-Spܹ��"�L�O����Nh���Żvd_#T嶒$��.�P�c?�����k��5�����x�8쨌�� ���6�<��j7����S��}��l��ј��'V��_ğO�49}HC�`���r9��)[�Ը�a>V��p��N���:�!����~
�|
����q�&��F�w6�nGHi�Hm)L��~D)�ՀJ�+%-�E��ῥQ�߰���V��^�Y�~��G	4�����p�<i#)�wXWf���D����G����z<%��t�m�\� W�.��5 �4	�D#�$[�U�B��r��Y�brÑ��te��/�Ka�69���(⫒*�Ԟϸ�Cq ~�G�Z{b?�҃�fɠn�v!�*&g͔ح1��|�{��M1�#�.G�{
B����p֣3�4*%�mOT�3�Ӗ~F�o���l�ޢ�<�l������Ka�K�
�w�G�$��XL��������?
�)$7�slqPU��U�:�˕�Y��R'"�5\�4�ǌ��C9�>T:�D�g8:T@n�lb���<i�[O�{BMXI$��mha�oY�S�����{�@kz��Lt��!�U��꾕zE]���SV��-��7�[~O�_w��[�a��[,�Ѝm���X�Ʊ�v��v]��M�@�$�4X\���\g����<<}�|@2Gׂ�z���jGp�\̅⧶�?>�#x� l��.+�Ho��y�r�X����\s���,Q��Q����I�r���9�q�x[�	^C��4��&φ$�v�	4ݥ���l�Ǣ<Ϸ��I��#�	�]����Hy~�n��0�j��I�$j�Q>пJ�7�m��ӄ���,*Z&m.�z"�M����=<:)%��t]'0�*����8B���:�˗ծ~�kqw�v��Ff�jG ET�����D��Bݎ�3A)�CXs٬;F/c���ϫ*A���yT&���h��!��&Y�h�4�|�����#vTd_���k%��*�Q���h0i#����	�٣�\cY)��)��<lӏ2�rd����{ֹ�ƿ;Zγ@�#ab�c�������� E��b���p��Z�iE��	�G��(}��}�H�x�e�v�UC���&��|�b�'��v2��?�`���R���^�Y�F��\�&�+�#r���8sq=H]��`:� ���2�/Һy;�	S��ئ��߈����F@��gA��]�lOTș`��Ҽ% v&_�E$�6/����n�Pn�&A���8H�P�c2u��ȋ |Tu��a�[�!�[�����0M��,�OY$��f�>d�ǘ��SV�3�)�}ʐ���4zq��E,���5j��o����l�S?� ��K�zI*��A�K�Of��l�"��x�����l����W��?�����WmQSNl`=f��MP����vې:޺Q�	`�����Mbr+���9KC �/n*q,ۀ���S�M�^��/��꺁�G���	\/�SDs��["�:}���{�ӓ�R+0v�"!�����/��P��Q��{>��ٟ|M訟�IG�KӰ`�7���I�al@ ��� �<U,|L� ��� x?zt�u{\@v4�&'��硰��vN�����9�˖��1�:D�0	�k�M^�K��	�Z7�=����ژru�&���|
Cv���v�m�A��;cв�煽�z{���� �߂����3��{a ���\\�|�=:��r���ٴ��;���@7�;���U��X���ܚ}&Ā6gn
 ��c��ȫ[v��P�o{H�/a�37�����ڸ측G]z-0��a<�]��"��^�A-��[A��8���p�frʋ��#u=S.�y��q�ō�*��m-7����{�����1M7��G\�9�cz_�.\��Q[$���HW��[�d3����c};������"Ĳ+�)�)h9B�D+UFn��i�0�ҝ��N�}�Olw�Ӵ`�g�B�P:qb|�����0�ϛ��n�Ko��4�<�7Ϟ~ P{C��Ҏn�Jϑ���o�Z�5c^P3�R��4��%�.r"�������ٻ�f��e�e�#AW�9���s#�w�(6Gw����5H؃Z���*T�g� c*�K�+��{��A�ȗ�1JŕVV-}6o��{S0 ��yIu��P��D�M )���9m!}�f��YR�ҝ���%�o�N��b���]񆸢�Rd,�	��=�4u{�a��ǒ����A���M4�~L��Y�-�}���o~�}ە�`rm�b�2y�gq{!�XA�U^4jE)4��z$�������"!��u�i^���jhjP�zy�~r�y�,��EP@Wk$�O�8poDB�ҸV��� �|l?����ϊ�c<�:ʈ~���N���;4�Z~�֖8��)ѐ���?�Ѹ�>�b���͔6�[�����-��Ry	ћ��Ν ���g��F*{�n��Lb���CU��%Q�	oѧ�z|A����>�����(,�ŏ����~gd�	�r}���K;�/ή���8�P!�|���P?|��J�e��R��9��G����c#'������qK ����ŇQ�b!(?!�9��4%�ֶ�br�gwn*+a|�{eJ!'����G�J\$0�s�ZD/�d����v�q��!��KT^�:RU"U�i'���k��b�-��SF.����/w�P�49�U]�F��xG��u1��o����aF!�iѩw ���1h;O�Ɗ�>_��.!��[g_�,~����S�vŢ}�z�ޙN�Q����s�����w&cm�qJ,@F'k�S�k�h�w�zq1�H��Y��c�5P��~�D�I�7:��9�'��Z�'�>��!Ed�>lf�S�y�̻��=��l�}�+пߋ��zx�N�
)��U�$��'������B'�	N���ﶪ�`�Q�Ո`���#�߳w�n���j�D)\\U��3���#�C���׺f8O�~��x���I&j?u�ﻶb�$��P(8[հ(I���>3wbY�0���u��P9�cN�� �8q���!{�+�6815����]�/��8|�5�,��a�z���5����	�i���ڜkjn��"���"	N���|ޞ3���s��>��J�^��|�<c�V����}�y��O���Z�L�/y5�vz��Xm�����+m`��F�*��+a�%�
>���3?�����rs�?�������cr���8��@�$���9�ku+�	>&pk歹4�NO�>B|�h�_��*m���dN&\�\���1h��w|��MEa��d�f�羿�.��E�%�7�t�������z�F�3Ў�������zE��9��`���Ⱥ2��6��r���S���T�xy/��k^�G]x���� G�r#	d�<<�]	�Y���R�\Qx@s��/�/`Eo!ۆ�_�"��e�c*[y�}@y+���x��e����J)(�fv��	N+n�³Clkᾴ�*B�dOῂ͝Rư�$a��V����Dt~��~06��rm�al���53��Cl�L� g�� ��?$ݥ-��V��r���"a�����Ѽ��:f�+:ut���imD:��Ӥ�!��]�w/�2��~%���X�=s��t�au@r�r��T��,A�>���\t��
��4ɵ����bf�e��o!�]R2�?�$x����+YA/Pq��6�7���}��˗�O������H^�Jp�� �e��O?Wӽ^��Rq�><�Q���,���a���A�i���d�.N0�����;�Cps�Le�N��_{k��J.�UϤL�`�e9 t���m$�OEm}�Gt/s�'��%5�'��V�n0�A�}�������(�W}mLEd�d�Jۘb�ڣ�f$	��%��I�Z�'<Dbht�)������3��9=���id����j�YgY&�}�2kI����7J�E�����w�1�V@���@��žg�)A�v� t^m�@|��hٳ2Fv7Y�����A���|Ew�$��P�G��F*=�^�g˥��Mf��}$V���ō���D)�[]��2���A����Y�/�#d"�eX�
.��H���_�J*/'`��lP;�cB-�� D��4�.���!|�x���	�d�ط{���+��	Qes��~/!X���F@����e+&o_)2�����5�x���=��g�
���C�n�3*L��{�f2�nt����\#�ɘ�xM�b#QW_��2��^�wU�,���Lrv�<1ϧ \�	;끀�?N�qB�>��jә!M�-E��N#�ҴcDO5yʙ��n��#0������E?�q��Y3�$G�� ��6U����������w��xP �ﳢ:��3�qp�Wn{�݋��"�Mg~�/�X�E������%^Lځ���!�z�w�'GQe���ӳ��*�Ȃ��i��]x�^b(�'D>�.�r]�u������9ϸ$q�%�`Q}aT_�A-U�m��B�x����L��]XNb�.>cf=��]neQnȲ������YޮGe+K&�\w��r�����_�F�ô|�ϓO�Xͫե��I�������<�;?�0���֌ٵ���%8J�N�m���/j�XЈ�N�h� ���"b�$�ݐ�tw�����hv�Q)���3�e�+���K���!kR5X^���G(DX!-|��,��Ɉ]��e�'0���x����$lvK[�{�+�����	߯W�f4z��pa!8v�c�q�8�#�������w]�bI���#j����t-@�aY�5o��ե�*|#����ᶿY�_����g�<�����L]�n���-�(�.�s�6�@��eğ�`�2sV�ŵ��Ɔȧz�,��L���Zi��M�����lu�z�RA���Q��;%9~�K�N����o�փ���P��G(v�Ս�HG'3�!�p뼏��WWA=�v����Ҷ���'��=MM����ď6����;�O�(1C3�ޝ�r5�c��n_����h��Lc܍EU�̢��6��$ۗ`�\�0]� �ddr�o|~&v��X��ׄ1.�J�����=������ϡƞ���,��t�_�!�wL~��BX�G8���lg�"����}{�I&�����K=��:B����Ś+>����-�Z�.�����D��k�N�>�mob4�]�>�$���\�_7M)�ݝ����/ȫ�-4�$��r1{a��kC�']Fa���0�eLr�&�_0�0���/����K���D��9�A��n��;6ay�h��
�|[,�4B��pyc�s�q)b�˸�à5\��8��݂K �Ea�_)
K��k�F �=�,��L�c��K������(��˿�)���s[�|a���tĭ���(�rs��r10�}���c��A(B���(��a� [�@%={�LV
T$������٠"n[x���}X�\jԈ+F&�.#��Jb��_=� �p��=���G;�	�:(�??�/X��Ys��LhWۊ�:�Md��F��>vLb�;&T�FoG��)��9�nV�����sV���	(X�h�C)��LM��9=�ސ��(h��L��t�7���m� �f$�4�u1���,b��"����.Pv�L��
|��(ʤ�#e�w��k�cؖx{�z�g�x[�~m9��!Gp������a�c�T���λџ��*�j�*��,��@YA�t����c�
��Y)�#��"�4�F�s������G(�aaӜ�(�{,�5A��T���*����ҨAn`�F�Y�M�呄��mR��Ә�TB A�f������,ܞ�^�����_ӵ+�Sf]m�o�NNV��:�Ɍx�c��m� (e:��g�� ��Z�X�EX4���AR^�X�.��n�|��&�糋���H�s+Y���oS�L;��1���$��,���t�����P�6�CC<�p�BZZ��Y[9�@������̅>�Bk��U��&�������!�J�i>�o[�!d�������-)2|XQyi���E��1�+%��m��������-Hz���*6Q�ygk�0^�e���ȩK���-Ö���(d���M�.�����лԐ׽�YB��r���<����؍M�Tn�w�%*�Ŭ���+t��r��ғxG�����\%+3�A˖A�xB��e����V��휂>X;�q�q��Pf�i�g*S���<;�G��au��N�X(-z��Kk˞:�YK&_D�:�#�չ��5e���$���Q���J}����1h��l�1ή����w�
��og�\J�����1��M׌�l��R�b,��w����l�t�Nl~�$y���<�(_*W�t�F�n_�g��o�f��Q���*,�S��� %3�b0��*��O����N��eLG��bU��A��O��(�C����Wq�E�;*�¸䵒q*��ZF��"�����]����G�Ldn�^�2J���(Zn#ϑC=/	B��xw��j(xgJ�)�qfIwv�}���O�8������'!�.\�_��^ͷ�t�>=��ל���cvD�c�a��<��q��1�'��bRk}4���r���9;Y�| '�:$oCH*�F��$����қkr2�������XL~�/!�v�Xnz@<�Fs�Kx�~���ML��y�2�����8pYɽ��1�':��8~跒�>�vOMFI*�kƽ��F!���Oa ��9���������U��އ�|�l���Ǚ)����l@EEEo��Hy���p׮���19 �T/="?d�s����v�|	���.��J�9��Z�Z�+���i�4,�}�qas��S��
����ˮ:���g%	��l��e�aki�%@;��$����N8��o�6k��t1��n���=�����k]q)�F�.n�?_��3�'8��.@(�����{�0#E_��bi☶oi��Z ����°!��(���&�fF��e!��q������hU�p�QJ��O��j����{��&8��Ùr���x��#�y)kْgL�^|\����#�������.��b�Z��������qP�V��Ƭoo�6{�x��S�d'��U��vTB�Ԕ��Ъ��i6M'MJ�~ɹ����]4;=�!�A�����4�V�d��}�Ќ�~Y��d�>�N��<k^��V�~��s����I�#K��(����\_��4N|
�+g[9�����c����Կ���5R�I��-�2Ю�>X�Z�����> NQ�=v1Ϥ�W�бbC�����;��J&��^�'���6�+�;�����>�ށ��B��^{��pc�2MH�Y�f�^D �yt�!�[������:ԮM�r=��fK�_L�Y+��䊊?��݀))O�
�|� ��w��A��0��Eևzϼ���i�}ϝ#�W�b�9��[�\�-��YZ*�pɿ� �ǙR��J��T���]�<���ʀo�s���ڸ�jhǌ+1[ĝ�k�(�� ��K�*Y�v�q}�˕�;B���|Pk�0�Mh׽���1x�Y`�nς�S���e�f@g;m����s0˹Kw�F��.��b�.�4��4ϣ6��y�}s,\/�1�VsNH/��e�������5)ҹ��,OP3���c�۩��g�n�AB��d:�x0ϜѝV��}Gt��t l�aY�^�wo�Q��t˩��Ⱥ�ãg�q|o����.��\t՛c%n'���E>����]Ț�ѰkYY'��:�Bk��)����+$��}�K�љ��r������N%�q/^�ӎ�����=%Ti�
�I�z�to�]|4���!��t>��4��^�Tl��F����P���*�Zw�]>�'��o~��JY��.���׻��+�������(��=G�9's������u�9(�X�By�A/����J~iP�XM���/7'�yZ:ϩ:!�.Hjv|~�c��i/��d���6��J>�*~)��[9h#0���N�|u�僱l5WNx��|���c|��HU8Jճ��"�cU��bF{��,9�~�=���Y�E���R8Am����j�����,^�5d
xS��A%=�ר�˹�����s�9�"�j�kY3�]��3�V���:���S;�
��q?Tqm��Y�x3U���_�	I���:�5��S�07��X���-P$P�WC���4������*��O%-�B�Tc(ǫ�|(V�����ɹsݹ�(\��܏�)k���ْ�.��Zf/`����~���3��N�� �C�q��Ҷ���*�+���h&��I�\F�.�)y�B��Y�u��w_�[;pJMn[��sbsHg��n�ϻ��ь]|Bg�1��YT�Si�զ_��b��}����N��C���"�M���� ��f�����X��טּZNj]&�O�ۮT�e��.�=q��q�e �[1a~��'�EL?�����.�ܴN@�#HdUUW~����Z�?�	Q�>FZ)���a��&���/,Sx<ɘ�5�RU��az_B*:P����o���'��L7]{l�?��QEC�g��zFF���~�]~�'���6D!�v��7j�Ϝ��I�͊A'7�t`8��Ō?}-�M[�hL��*���]>��,��M˦Lnˑ�\��k"�Y �RK�|qqR�����T��ְU�g_���R���1��oQ�p�˻A�'.]O��! >�cι;@�G\���Z�_�5@l�^�Y�p��I�v�� �H/�1NAF�cQ�L 	aj0�2{��\�<��b��X�p2��	�;�m�Izz$��Q׍�������!S�f��HC�{f|�z�PԀQ[��Ri����P0��w��kK%qֻ=4<ہ����U&��T��F,Y����=C���Kb��7�\$cE�Pm�&�u����2����1&�7���J��R��&�Ԧ9���r7b������l�.×G�%��S�Q;���W�rt�\���9ZUW��#���̽��=o�]��3oh2���f����P�9�(��'��I���D����C�������d�i(M��� ��R�yM!l�s3|�y���:�m{�qc)	o.vKY#�G��3�Qw(�����i�k{/�^b�3m�.:.�bԨ�c��*�'+R�S��I4�A���ҀPҶ����Mo'���p�����l�1��s�I�Rw�~HY���L$������6hyO��1!��}P�<�rՌ%��� �熜T�v$F�N�����e������g�uD.e���5�{;���,1�9t��?������m{�ϖ�� QK��4�<X���s�������ZN�L�E3?_��Xu��ms�����[HGm����;`̄���+i�8![�@$	�p�'��6�WM�]�U��#w�v�.ޡr��d�x[��>v�@e��� ��}�)y���'NX4�X�%�
�7e:�a㢇Ԫ쇽z{�֒�� w�.e��HjVT��3��o��y�dK�E��Z.x-x�1�F@"�ƦS m�Y��*?���X�౹���\��<�^��QI�q��&���爺�m��0��6�^Θju�h-K���i��rv����lԘ�fF��5�˶:���ʴn\̩��LapQ՜u��`���V�"���/��2KؾE:R���:�'Eq�N�����_�'�!su�*��V��s�]�RZ����=��[�L�[�vg[H䘲�1�1��^�����t�E�6[��#E�z/���Fx�8'B�͈͡3�p]?��8�D/���|���_=4zo�S.C]9�6ƴ��Y9��R�EuZ4Ѹz���j5�o��Hb�(���X��s�.�� r�	;�[<��T&���92�Ӯv��U���ݙ���p��䬢"4Ga�B��Єj��(0��C%�
��oS8H�OU_��d8�F6�/�-�v��x
vQ������ǵ�^�����+/��IW�9}��mB�@$�N�x`�ё�����
�	���B�u\��F��Gm	�r���B����yH�VG�zKY&A�ZǂhE
$O=�s�6G���j`\���F�#W�\�����Jf{m_yz&�>=�Bސ����� Մ���T�^*.X4�����o����t�־�/~S�Z{.2ԉF��V+����Wt������!#�\��J�9��-�m�9Z���40슗B�j�p��fG:Lza��2M�'Ӂ�?�iZ���#)2�-㲣oR�}>�ve�SS�#���^Xh#Q�]cfn�]��oI�6aisF��ɥ�c۽M�~gq]5f*��/U&ᷭ��;��rqC�9��%�b�3��%T���u��Fk�q����� ����}%���� �C���.,4��U���l��8>{ ��c��n��1kO=�_i�����wŅ�1�k�3x�䨀��F��uՠ�L̎�(��` ���y�w��:~5�5v�;���N��[��?l��Hy��"��Ӗ�n�	��G���$���=��״"
�k�=��Е��v��� ��V���uC�I%���D�Y>+�RO�|�_��p<_�"��mtiP�V��{��$�����[0[ֈ��;Y�3��/a^���� ���/�[)~�)�(����)��Şj��؊����]�_�H�b�2�(��5�H�]@ڸ�ȰAxu�%L���` )ޥ\���5��T��{��tI�UG묱0��� ��t�K<Pȍ('���k�_5ղV��-��|C�C�kӰ��Kj��7g��c�8z�V�\oX�9�랸�:Ko��f�;�>�ژ,re���'�aD�YK8��$?�����05s�ɉp&��U�?�X�2�;<�K���#]�z�)���$H�t�	�@��A��a��i>27@��_;��5��p�ܒ�g��@��qJ"Z���zh���dɤ�f����Z(��iU��;\x��2�rA���ߒN���m�\��>q{bz��j�Ui(~�)��mOr���*�4��s��b�%���r5��s '��eU�dҺ��7RJj����_�B*XB�!\�q�h���3�iDe������1l�u��h���d�x+��y��}~9�03������� ��������θ@�� @$�L��W+�֧�<���Lj4Y+B����lL��`P��:G����߅������g�O�*���^cf+��^n����tK�@���пs8vm�X���q0v~�Н�N,[�Ez�ك,�z�f�1/@���S�Q���]�q*���eA߲-n�ׂ�RNX�D���;�͉� q�J�x\��lo�uU �	����d�H/���x��u ����!����o���ir��>� ���E�D�7t����g4���ʀ��8�P#������*�
����XƦ�g	V�'�9?7� ��(��ʧS�N�ꪄ��VGx+C����� �=Sb������9��#�Cصv>�ӷ�K�fݔ}Φ�pٳ���'��a�V��p|VYy��Wlf�!�R�)Ս\�lNO���x������ڽ��<S )�<ZI <�^&ql�����ʡr�)cB��� 
�'�y�/��Lڢ���k�=c}!,�Kx]9?����`�G�#��q�<V'������!�c���� �q���5�0�z9-"��s�ڲT��o�^Q�����������-��ÕӲ7��ÏY�>W�^����6L�@�톌�Q�����M��{聙r�g�qꢺ�ز�g�IQnX���Eִs=�0A�/�yЙ}��<�k�Tј2q��Ւ�7�}Q�rÕ�c�O��$U�;�Х{�n�F�8M1���x8Z�1��W׶�JT*����z`=�Zg�@�6>1���B:�4�[/iA�8�B���##��Ĳ�h jt�e�쟎dI��	�ˍ�-���Z�Q{�f����F���J���F�d4��4;%)�V[�"c}��x���fr�,CR���ClS� p[+:	W��Y��,�3�t��i��9�6
���f� w�ve��FH�W?C�_yM�&�b��B�l�3M���*n�0�thɞ�����`��b^��Cص����D��V�=p�|�	t��rJ�}z�i�Q��g�� �F��qn	�ޢ����=����u�"j�y,y��q$�:^�l�/>2'�9�zm�xK_LWE J	��q�2�"���c��<O���.�ј(@|���2���ݓ�1L��+7��>���YW:đ�v�!��������2��͉~�e�\PM��w�)Tbe�~��?Z��'�2�G[e�sB��X~_��&<���ڡI�ʘ�s�J������7����)Q@���=�W�&j9}��h�+1������9Z�j�f�(׶¾���T8u�֦�bFΘc~�t��9:��tϫ��:HUDۊ�@�G��2Р��1W l���/J��|��⌢��g�������Iz�ލx�0�&p*u�1��[%(X�I8MC�<�%R���[(4)_�q�#�g�Ǯ�Q�ZZ��f�Q�����کYӂxG������$���31	����UHo.�����us}@~��4�v�l��l�Sv,Q��D��7�H�)E�2C�Rc�c�^�mY
�0k��mS�d�#�\�q��.�� i8�BHS�/wґ�[�3�!/�4H��2�� �����\O|�������	%OG�}��@�S�ެ���D!���x�\>ҬR��I��0E�_ܠ蘱S �}��p������D �,F��O�G�S$���r4�.������-Dh�����ek����b�.�_��)���Ͱ_�q�S���-��O��}@�h*q��V�O�[W5D�"�J�$�2v,JUQڸp��R�1�����Kdɖ�P4�r�鄖XF��? �q/+
뀧K��/��q�t��3�ɘ�R���7���oF7e�m�_����<�;��皾C	 ���2��eC_��A���r)dBe�ǣ��;J��|�򛄶���� 2ӗ��/��ű�����F����y��$������d�W�KO��zI�Vv��������!�@0����G�x	�)#���$İ��p[���2dTI�vjU�����<��
�ݹvK����a0�'&퓼n\Ci�.\35��%,��P]8����(���X$�?#���S�͸���]x��B+��کl�����?G��pZ�&X���nLE���K�Y�чP	�B�J������Q�G�e7e�A�%9uюd�s�`ȣ��r�v� �qi���Z3�Yb>\�
j-���r'�V�f(��Ԇc]Il+~���<������{�E=P.cʆ���l���&H_�ݽ�t���m�݈����fbH���-�t�ğ�}`��������M��M�ar�t�5�dE��7���Lb�Q�F)l�q 3~e3	�*2DY�3��;�s��������� y�i(����.���&�������bY��ȉ���z��o���؝����"wo����P�L�=g[I�PQ4��p��Xx��9��8J��ʰ�#u��c��ӫ�qa��Ƃ� ��r�b��୪/3Ÿ�Zr�J���S4�1]jZ��[a��/���q+�-,8�����(lņ{�H�T��8��A �bb���R���uW���tU�z��Ks�D�(����WR�fZ!�9-�F�۴(;��j�P�!�"�s}�Rk��q���o.\�|˪���3`J�`�?@i!�|��]=����i+{�H )��@
����T9����=a�\֭���4s+vl�C�d%���e}�~ze��U(�PG���=��mK�n�``�+wH�Vj��r���Ep{ݛ��@�R)���py�Wז������t!����n(��ه���&���^ D���g�ȋ���-�Fe����Y��_��Y����u�k�jYQ��{nf�|I\ӱ�!�9J{	�.�&$B�����&�L��"�F��K�[�Y���"^;���B�kt_Ҷ���/?����� ��<�v�4-H�x�'��ͻ�^�әb��l��<�&�E#�R��~��ЩB�2�S(���.�������檔./�b�goxn�B���䓘�<oTN���o$ٟ����$G�K4��!Bi��M�f����
�G���fr3�H�W�'�>9�oV�=�`ӳӫa�7�MN���y����i�@�S�}v*��*�Z�-��9GR�d���{R��&`mI�:	���y9��"#�J1:H�[���
������c��[�?��d��op�[��MHQ���'S�w���D��lē�_������|���JeuP�mdLFڽ�Z �͘\#�W\)/�a�p��*JF��9�i�ίye�Ywo*.|@SkFh2��m9�r��VxXע�6Su8����^0� ��%�kse����cv���VEl��f�ű>�����DH�N�n/�L���Eh��Ew�?κ�k}8z!}la�5�9�cw���d2'A�|��d��`VtxZ�O���E� G	mt�+���9m�T2��n�z��t�*:GK�_$|B�)W��w%�xn�i�&���gL�y*�>���{���C�:l�1.D�T��� t�q�����e,�7�CyҒ�kҠ>��_0�QSs�R8i+PQT^[�LC*����1�l7�/�9C��Z��y93�:)���b���ΙAf���o(�,)'ۨs���=;�Q��5��Q4�tQ����_~�P:�2��ѣ!�o��wF��*�EzE#�
�[�ȭ��RL�@�'L�ߜNpxa1��zGM��ka�JƯ�d>Љ'��.��us�c�X_���9���Д�޲=�}��흟8З�K[cQ~rz:�7�����Z�E^����C�Oθ�����R^��y�9�_�K4���|A�蚓�'۳��Q�''�ڡz�]j����Sm��u� ���f��~5�]%W���Zf@ʂ��g�R��k��Ldm��m�;Gㅱ���;��iU<���i����A[n�� ��֏��������jN��$Ln仁��O���T{)�&��u�S̄9��ň&{���n����i�c�ﵤ)��t���N��''/u{q��&�����T(4d/�;v/��f=�#R�@�5KsX�v�%��Ev�M+�&|-yK6r���M6��3��֭%���<w��M�~��_�I�� }�_ã)���	Ʉ�=kAy��r;7�6X l!֍�)jq�����*�Z�В,��jo�plʐ�ϽE!�&ژ<i���6���e:�;w��M`��_�R].	�� e���!�o�}�QTeD�zHl��EmJb�:&��k�������-���l��6�E��{E��a�vtb\p�+���N�&�*� �Wd@��$�hd'TP���\�t��[��D����=��E�6�mz_~0������b��bO1in[j0��1���{�S�'�9>���~#�x�5d�S�%k��4�W*wGA�����QwSƩ8�~��_t�uPr�E�X��%O~B�X�3�#*hı㎬��[�W������N��6�#G��ęV~�v�)���e-��$`��݌<��#+��R8`tZ�6?=b&6�'��}�	J$�G��Uܐ�
O��Ѥ��x���V�\$&Y�:_��N �M-��>Ί�c _NV{<Z�����.~D��u<�p�Ѐ�����a�$��[$���?_n��6�8�&b8{����pu��b��3���2� O�j����M��
sX�R磑]~��1���\���}�Y���fL��V1�'�]�?�
"%:�����7��k��m��-�����5Mb]��TS� 2��jq?��&��� �ѡ00�7؟R��y[k��,���<����4ط�����C�e �_H>���R6TX;��k��je�Xʻ�V�E��Z{��-��s TMMXx]�%��wA���Q��i�=��"�A*5��>W�C��Իz!.b��ץ����sx��D���K7��	$�l!>�5�O,g��̕������Z<�m$!�0ت>�9n�)`jXDu�`�ز�.r��s�y,�U���[�4��G[T�^�J�1�� ���=��R�r�fE��v�3������/k�((��[�.�J����E�].hx߻~�ӭ/���sصc��M��Xm�)D�I:j��`�es/g?��G{�z9	Ol���e4�d0�x��O��6 ��CK�s1$*y�Cz�Sf��#!�/�*�#}�ñ�}h��Γ�s��f2��z꠵O����*����U��hK��R�,׸Q���a�;�W/M��5�bσK(���c��Id�`M��hv�LB�w��]�|�����
-\�ⓣ�?Z��
G�����d)�]�Y����A����H<=�M�۠&] �
�N��ͧp��H�EP{�)�����Ⲵ2ɲ��Y�yW1q(��u��C��g������GS[p�ì63I�ML��qϊ�gsK��A3-�~��1�n�p��8{�A�i�)�~d�	_�#�r{h�ި��V�7��'�>�h�G�������r�ΖGDB�urCԛ����X�__�;�XթEy�����f�b-"{�Բ��Ic_���S�
¨x;:(P��j쁛.�J�J)]�"i�}���������T���C��T ��Z�T;i[���ޓ��K�w;n}	"`0�{�#�H��tq32�����3m�:�|"��ZǞ�m�3����tІX�4Ş�w�� n. `t.�{3�u�|R�no�Ҧu?ID�����~�Y���9�ʖ'�9��M��(<O����08m�d� qg��J�gO�=����7��ӹ+V��ގ�C(c���D��O�!����o���.�&��ڂ�J ڪ �P��uXt(�|�}�G3��pg�1��a�+�-�bA�ӂ�.y��p��6M4Yg�v�ҫ�gU�ə@P����p�K�;�iǻ'��\���Y������ �<)���=U���m����c2�l��&�*C���+)�FM�ɣΫm�*K�eA�MQ����d�Q��m��&G��~@8�9�.v�d/�`1J~�1c9	7��Z�pU�GbEL�|9�9�;����6N��h(B�,1�R��ꂋ�}��w�m�Bn�}H�bj3KN�K���̴I��[A���x���T�����R����{Q��v`��4і#��o�B��?��o4��(��C�pى��i�B{X5ĝ��u��������P&���NѸ�!�^��EP�.�X՛9��m�%�6�^Qz�N~EλF����w.(�fn���X�\��j�i��H��ݢ������`r�ޑ���:�Ѧ���S�J�[��N�?C���k�V����v���B�й9Z��>}��|~��ʅ��ř�j���j�'��s����I��1R)�f����1���������o�?ԋ{�����Y���/�Bq�A]�/��X���h+,�8��%�+V����a���L����j�5ӟ�����qc
.��M��K�W��p�6|���
/f�S�و�L1x��Ƒ��j�� 4!��h,��0��*�0؊4f��%۪0eE-a�iE]ę0�����@X��<�j��U��"S!m-_ ~Ճ��<�~�t9څ>B+���[��lP%��aoBƍ��2���0��Nj����*��^R����cK�����
�qy�q �	��n~fP�EJL˯:yRK��N��zK�4k���u����ϵ#��L?>&�m��{�y�2�*�4�]�/)�b��������+)�zfv�X72F�����*��ar����kf��`ͯ>F�Կ�Q}^��
i?�K9�F"&�e�Bz���i"^�.M7`�>��[x9�-�i�;Of��s$ױ���F(,hʏ����K� w
�T�kY� �����D�9��h���Ҽ�-���t:V�f���IT��s���A_�>p��T���H,�JWQ�t%��.3A��� �-i;b�����[���?}z�� vֽ ����w���򩦵�n~޺�	~��.j��!���^Vo����8���K@�t����3k �Ѝ�4�����w�+/x�
*ٛ~��-����S6�q��'��z��)h"Lm�N��&1�VLB��� ���Ɓ�
��	4���f伹��:��yYB�y�Q+����B�D:.����Sp�����4N'u���x)c��m�t����H�k̼wA\�%Y��G�	�
tρ��`d�v��#�6Y��1�ų�'{�}���3���]�5}z����=�������7��*���g�ؙ�����^ڄ����w
�1��rm'[ࣹ�J�Q�G�6Gp�������[���s�����5!4�u� Kqo�e���ͯ��8u�Y�Ws���"^俠�>u����v��^{���Ɯ6bn�{?`��X�s����F���l(Q��ϧ�dIe����<�}F*50-����q��7�㲈Ȧ����]��If���|��{��~G(���������i������N!� g��
:jw��=_1c�n�(���7�4�ag���(K��|ᄒ&O�k�\&�o*J���T����A�/U�,=�ݸG�RҊM{*�pC��_������阥Ƀ���#�;o:d^��ᮚ�I���^)��:_�L1RV��K���*dnt��3�I�}�B_��2(3	T���w�N��ܸ[�덏������5	c��y2Н�C���8���d��X���ԋ�E�͋�|��7/�a�⸌�|�� �� 0�]C��&��Qwⵌ= (��}�ڕ'/�\	~�+S�TAQ�pe�S�uE9�j n�@�X��/B�|P���ު�p�]��>�,y2�K�V�4��-ťhS�Ia��ކ��"�r�e�Q/K~��S�ٛ����8�L؜�>�n�𦭷1Rhs:f##�� �K�O 5��1�3�ӌq%��?�xNF����{6�;?ר�'�B�ɴ:ꇣ��_Œ̐��?�2���q�d�B�ʯ�!��4�eİ�1A�
A�Vø{Ӯ�+�1|����6�G�T�3R����0l����Ң�X����)���}��h��G_fq�q��'�}aϱ�Cw��J |��%G�p!�	V
a*ve?�^)(�l��>R��zU���oYR�28U=��綨�`p� �t��疿$B-_P >�x��(г�bwkBǯ"�.eP���Y���I��
�'(�.������7jGEN����l=�VFP�ݒ�q5���VA���䪾�n'��
\�(*)��O �`����p��[B�M٠�HL�ٍ�!}�	����&K��sv�{i�u�x��o���N���bg*����N4�i�ΰ��18�=�S���hZaI+Iإ>����W;k6��Ze�4(:�-��#�9�%���G`��!т,�i|:*0��^^�tmC�z�Lr �V2��	o:��z�}.�]����pQT�}j�@��c����;(�viYtLhx��vK@����Mo��{�,-���PF�iQ�n&ʼf1=�+��u2��b�#(->"��r�q!������n�����y��&}@���D�f=�Ly�|�l0��Y����H��g�؈���(�2�����3�<شc(�j:f�݁���CK��
7!�+t������|t�
��n�s�YU����<h'�J��
?܆U�����Į��}p�!A��#G$&姢#����K��g?NA�N�,:>'��]*+"��Bk�[�����#�n}G(8ˣ컊���O�c�����,��YrԤg0;��a8t���eV�����I'�֤����⛨����XW+/��Ϛc翣'_:��G�El$h�P�>��B
�[����R֛#��,H��k��^�u<R
��:2���T��p�&؞9f��׻�*�-�Y0��7����ڦli���v+!�(�3Mh� q�S~�%QB�עP�ڰ!�o"ю�h������:��Xb;�
�#@���SؐZ����
O�r�.+�ͭ�+��)NY���'�6vd�)�ﹺ�ƭ P��xbĉ�q!;�`�H���@�C�����P�ݩ��F�b,��g�^i��ﺤG�\�K��Q�Q��od�i�%�F{����X"J��N�}�"!�Aotv	(Q�Ʃ�y���!���:i'�����Y��[-�e�;k��o�Z�� *�����	���.��(��P�����Z����m9mт��Q{ 9}"���Z͊"��w��_Ce��-��/�M�D\k�ѿT�C�٧yzd�T�}p%��˕�ob��oX��Ľ�1���۠������H5Z�brI��tC#�E�n�݃|^�%����������t� �T�>�
�k���I�:��X�a�ʿ?�S�D0�a���okj�O~�*��,y���6����NQh���r�ǥ�<&�x�䈯�c���h�R�d��%��_�f;�-�,Np�+#��X�:]$�E_Zg�2��u�&�m&`w?�P����/���ݾ��H؄�~�(�N�g �0�j���)~N6A�]x�tV�=��{3�o4�է����gA����!�����f�PQ�R�����mn@&�R�o��4��&���N�E����������Iڕ���k=�>�n�5�O`�%�⾈����Z��ʕ|��&i*.���x7�8�a�Q��Vi�4��;�k��-� r���4�逻F;>���!�pBa���<����ȼ�:3@-���s�9�e�O��Jp�������� ������\~��D-��L)����2�㗗6�At��b_��UD��O��|�L�چn��㲠���+�,^� �E}"|~1!O���#b��������˲�R���R+s�͊�����6%�rl����"}���@2�&1�.������Vc��.��WQF�d��L�F�8���2>��m������vț��y07/��僚w��'$�ο�m|�
]ٰ�u� �=Sv��A�=�@�%ӳ@�0`��TC}�������O���!�H��nH�~�â�N 
��0#	{\_���=V+(��CuIu^A��2cb+�gf<F�o���ce��	��y�7��g�$v҉v�������Ν&:H��z�DX`��5KA���#g�,���]i�Ԟ�?�.�}~�%��T��Lr6е��ĭ�4��8/�����Ϸ��8��h��>%5�~���OE��g��@�0C��KNVb��	*ιWQ���+���?�����0!�d�<�O�#�K�(��~h�g��>�[nF��k��M�ܓZ�m�{�F�w"�4�b�^�R��%��]��	��$�7�u��n)���ye�CY�MK��K>ǏY�B%�}^6�R
�^?K���{��$�d���)S֍��G3
�����ї� P��X��R��|���+�;Y��IQ@��L$�]�r�/؇c���U���`�� -�;�uǶ��
�m$�ӉN��j�[ /.��}z\��V��_���KL�bIݖ�!���	7TslR8�/����n���+���bZ�VS+�rK�E�y. ��:T�"w�����ӖU�����|�w�	�������y�M�1iT��m?-%eѿ*懤��]�J2'4Z��Z.s� ��2S�·�@��p�B�h<ƻl�!���~�o�0XL�2� R7�]��E�qZ��3���ёȱ��V"pw��\h�"��'y�z��������|�o1ީ��å�]�������X
+}�o�/�bg����ׇ|���dK���ve���^��*���٣���B�J5@�$9��u
�}Tݷ�_Is������!Ζ�Ry��l�,��q]~�P[���ģK���+%��K�{��@wd�ͧW��ڡ|4�Gy"tn-*�!�:>Ǧ4�;6y��0�G���a��[�ѕ��W��jr��B�X*��O��̓�𙓭1���+�����-U��;{�P��8O2A@�w����iGN�R����J
�f�;�),�R8R��F��PS+jzWsmuj��ދ��)��RT��,���,R,��P�>];U+Fz�c��*��ΧK���-�"@��7�@9�h7D�[1-[W�C�(l��={k^|6�f��?�Ü0D�@��ۙ���$k�jߏ�U�gT�<���*�f��[ G��Jm`�6������:��0l{C]t��H/G�|��
�+��_����8^�RG�C"tt�1a�ͯ+�&��є�~;`��Z�����Y��i�{��ڻ週���yʅ�i�T������h�	�˞"��ǵ�%tQr��V����iI=��e��K.`���.,�.��5�*�G	X�SW�ۋ�=c<x𔽄��V���{��D�:�V�X_� <���/���1Y��ؖ}dv��(հ�3��$�
28�y�՛���a��C��!s�i�f]���H�6�a<K��,@��&�3�Yxj�.��B%�Y�,�j��m���j����N�m(�&� �K���O�� ��#��9��
����j4�ؘPc֎2�����ED��)���3�݉���O�'U$X�6�˼��.e�gȲ���Q��ݦkChV��g�y��b<P�5<ʦ�u�T���.�F�����L'3ϓy�X�]���y\�b��q4���Hp��}�p���9|�����kLi[��r-cܵ�"�����4	��~��%�X�!�^[��R��,᮵t��t�o�%����1��<F�҇�徒�K'#���T�g��;���B�������J��k$'%��{s*���^��̋�)F������m%%RHw�M�z=k�`�7Q��&� �n:Ɛ�*b�\��Ār�oBLp���{���Gx�S_,rz}K �딴�O�V���0�x S� V��4�#�ap����n�%lݙ"?�$[�X�Cg˱�
o�,R����S,n[�C��i�Z�Λ<:�bڞ\&��ߘ���nEe��S@�S��p�gkt����qd�(���e[-=�t3�V0劜Ȋs\��������,�.��U�MR��$H
�<�Pe��0�e�M��dC$�U�j9�R���8uM����3�Ҥ��x�s��ٶӥ�#��\^a�W 
��Y�6��z�������a(����H����S���U����j7��:�v�򏶉�V[P��}������z=m��։����q�]N�I�G������Wq�1t����$E2p;qf��ګ�w��S���T����.6U�y�5�-tO����;�3�-Y�^!��Ƭ+���*�&�WBm��j��b��ңK81�+Ux�i�'�X5�g}1��:̧Uw�,J�4G�#�S(�XlHB�=���~����I+EϪ5��P�WЋ͸0 I/h}5�N�DM�V�g$�Uo�H�??W�v���#{��>S��1�r䓆l�Z/�\���=�S�y�^����J�����=p-as��7ͷ?��y>�+�Ӈ|
�&8nxg�*^�o-�I�z!�$�J,]C<ߩ�OV�������D9���bh�T�v
��� L�=a2�XG�F���s��v��K\	!���I+׫Ʊk͊9�xft?�*N���7�i�F�V� �BEڅ�J�:+xdI�@�Uw�-e�+[�S�m븏�@}S��YRF�k��bk,�]���Zs�B��6.s�'��\���5�7-�t�� ����T�J,e4�F�1ྜྷ���0s��Ӡ����xwX�k��i���mk��܈k`�s�O�#��J�y��u9iu���v�5ޅ�__�~aH�/vY����HF���oߗ�pvU?�<�[3@ &]GY��zXݓ����ӌ��U��3�Y��,�[,*�?ݤd���Sm�T9��O����R���ʃ]�܇��3 t䷵��X7z��Q�3�펽����k2��>=�P�߂\ �(!� �?֪�)�~LI�Z���zWP��2e�]H��[k��YS�>�(A�]��|�:�n��Y�q2zoG�$~�����6vVL�e�)Y�V�ι���9�����AY�������'���M^�9�����^$��|[��H�w"	)fs{�r��a	�*b�	��)�X�u`�	!3��v����\��9��8��q[�ĐS'"黐A�l�k�)�G�4��u��zj��<����t��l�<ܳ}��MI�B,.�\���w��4|���$��u��ʜ��\C*����}��d2�@ �����-Þ�z_[((�;
55��rk�E����~T�Θf�jT%�����W�|.[�����X�68��Hx?W��[̭�QI�Z1��|N�AS�l��,�z��q�o�hxˬb:��h���W{�C��ee1#���7��3{��C{I��%�к�Z��r�(7��x"�m%��;Ϯ@>]0���>�p���Fc�Tyر�	���ӎ��|s�����=�v|�Q�;��؊�n8X��j�z��-3ﯸߞ8HJ/�M��Q5���~�tT@��
(:�c���
3����٭�	�2�|�98����U��'�Y��&B��@<.��k���/*Ǆ�E{/�Uu��CG~�:pw�O�;R�o�u� 5�S� �|� �~I�=x�kM��sG|�g���;��U��k���%j��B���5Lt�,����y�u�Nq W�>\�9��A�ɕ���0<^���u��tYx��Ű��b�������)�+�*A�͏�J8��ڼ<o�rO��4����V���n��MEz��3�d���U��+�[j��p�r%Jֿ�U�L�㈌��G�f�>�i|q����:��fC�{��5~�Ei��0{]U)a�W�i����'b�`FP��ڙ�>�+���#g�v�49���	Qׁ�M���A[��g��滖��G}������*z�]�G�[T���9���Cc�Z�@ ��P��8�+��]L">��ͤ�T�I�=��<c�����E�LsD��Q%En�[/����s0��8|�=S|N!!����*K�pn
��~�%T����Qc^t\�������m�֬�S�O�%l�=K])�=R$�	
��N�͚&.����"�MV~C��N�*DLTR|:���n��O8��|�!꽰���<7�����I�y��XM+�8�J|%�~�Q_�R���m�CnY��;6�j�3I��g ��A��d�Ql`���73h�yy���=��G;^�Ӫ/2�F�AZ�.�Ǎ�	^OK�Vfo�I�[a)|䳬�f^��n,�� �(�v8��a�J?�)��w�w���ʚ[n��aܢ�%����������>��\ւ����v����P��v�PVe��A�l�~�zˎ�Ϲufť%ux�+�h\ip�<���Vj;�_&�M�0�r�!� R;��~#����Q��j��5O9E���*�"m @��6�o?����W���R��!K��#nG>)fR�AT��K��x����`D��j� f�,_hrK�& ]�x˄&��٭	k���=��z^�:���W�y-$/Y���Ǝl���7�?Ƃ? �}&fǌI`�}0�=H�%�yNT�u�=)���;��1�_Z�Z��cRCW���Z�!1����;���pL��N��.�<5�����O(c����K��y�_DXd�3"�_����QU�s�w<���/��JwAV����X)�W�J�(��Z"��0��G9���1]ɩ( �������HVj~��`$_�8�D�̭�|*�>[�����0�/�����S�;[,`y��r�~��L4ls�#�x)2K��(��I�>��td<]9{g�.�ȐA�畳�4x�Vr�>;N��q�)Oǜ�5�C¡��<�'�gX��n{q/����k
�L����RK=*�yLK�疮#�LCPy��we��&�J�����GzO g'j��ߴ��)�C��ت�Ő������Q$W�LT
	 ]�f֡�GR�`���	�_i7�u\��c���I����ꋿRݶ��LQrcs����N���JB���Ύ���кN�y�Ԑ����3ǁyI����L�&��j '�����F=�i����{��ql��\W��ݍ1q���p)�k�\@��Z_��CTr�B��J���w]��RS���e|po}5Q[����j�Jıv1�����r��0C9 l	)q���T+mt�/��2.�j|IY��]���c� 	C�n�lHޫ'�B����_eb�wAu)m5L0�`�P�qW|d��^ֲ?��<z�����~����g�4	���,.��%���z>����[,�"3�ߘ"��u�`��e|^o����3�����:���]I�Lp�=rLo�̈i3��A$��
\������^��k�A{�)��cw�����S�;.ф���=$\ԴJx2x+�v���o#�8�)]
�{�^6�[L,�z���gQ��5�.�wc|�B"��@�����h�
� ĺ��&}�Q���8$�4Y�=)[T�c;uG{��X	�s�~�c��+�>�晨�C�q�u�M��N�7ۉ���D���&� *�7��G����Ӛӹ�ߧ�s߶^	$UB��͑�0@~I�t�Ye (Yw?[���C�2�%��|��x�+Z"�P7mq6I��<G�>߽���d�{)B{bP���.�vi��9frvd�aQ0����ǲ�����n�C#��=��b��oT[����Ʃ[��F���rՍ��˒��Y�o�*xz?Y#�X4"���P�ʴvE�q�Sy�JӀ[�.�|�;���d��F�xx^>z�sT����c[����[<�L��-������������.��:��.3
YX'�vµ7�p�șN�Qq�
t,���Ĝ0I��L�WJL�f���Rp�:�V���������$���๋�M0l�F讌t���8���?���Me����|������ۗ��BU���i���P �NM�n���{� ٞ ����kzN+��Q�恬��8� pd\.Z<맵ݜ(���V#���-�a�8Cm
BI�I��W���y�N%��"-F��9p���T̆	��CX����["��a
8�,��4��W6���I��Hs5bL{QcH�����ȥ�O��4��r�
�DW��s@2�'0��AM\<��cH�UЬ�,�����'���/� ��ރyD�r����u�a;�h2^�-2>A�N�#%�/vT�?��d������S�1�� o��=�1�oB�Y�z���[�cv�Ph��EU��.m�����rWp�Y�ͨh�~����bI_˜r|,F+�cG��M!�R%҇PQ�w	���ߢ���ט��w��R�ZA 3|��ٮEd��n�{)���N�������4�9���<o@:q�;��AX�།9�e>����
�8�%���T��Ē�N<w��wS�
������J��Fxn�������Y|�֣���Ad�ujڶ��G��c�(�s�sJ��H�K�J�����_ �F�AB��o��(�s|W	7�P�?��H����t�ƹ���vtH~kG����;���i��-C
稚ȳpT��S\�ɮ�gK�Y��.(���O+ͮ�����6=�2�II�>����O�+�a�f���e0�M�)[I��^ۯ-3��wE��XG��Hgn ���#&�Խ��G�(�uk�ҏT�۠�7IH�q7��v$���.����/0�_7��a���n��U0�������\1aC���7�J�����Z�=�I�"�"�����������
q(��ꡊ{����=Ȉ�Fb�@������h�h��nHu�����@%0p�$�ș�����g��.���������p�K�'�z�v�l�QV����g��>"!�j;��c.�[	�V�୫�������u��A��A�;2���2��a$��d��&�����@o�x�!��DX^w�x�Ta���:^an4��|K(��2�A�q��ń�G�Lzf����u����#����|.R�D��[��-`O�/����9�']�?#��1�k+�w��#.������?�$�<��G��\Ha�⦉@�u���~�y��䇉��'DO8\%G#�≊"����	��������,��Ḧ�hƛ�ZAG�ygj�%�x���z	�`���$!��c�f{��s6M�4Uֱ8�G�"�-�\�4�,�;��i�ӸH���P�pSQ�*�@�7>ۙ�Ty"1e����p��Y�:T?'�X�t����Ւ�Y�����M�����*mmDi!�űc�K,���̓��Y�� �����Y�i�i:."�����5!����g%��Z@8k�v	�_:8�=�&؆g9P�� B���"���������UI�'2��Z
�7�|�y�����'w���4�O���7�v�4z+½.�+�����j�I����̖�n5AQ�sP'���
5s���.�*�:�ZB��������h]��^��R�BT.C����?۝
�t�ϗ~��݆m˓[��[�E�y�ᜨ/�*�,)�p�:@�(�P&���p;����a!-X�%��s~��@L%�v�\�(��*���N�7�MiS�x�����.�w��	s�o��ͣo�@�*=�5׀�,�ՙ_���L��Tn�v~�uNZ�����Q[ր[��zR��c��4� �Y�hJ�i�mL�76�TJ�r�V��[&�1w�Qp�Ȑq܌0JY�)�#��?[�7],�Zt��\Q�ܜeC+;ӳ���Y{���e��:�Wr�se�����H@=:ɳ<���]*k����H��ǣ�>�鏏���<��m/I4�Sa��
(
~�%)�>h�(���`�0�/GZ�Pd��ii�|�>��q� ����U�����JJ^B'�LK	�u�R�0�U�'��@X*��%���.Ή�����Y�n� ����aެo��}6���N�x���NL,s�ɛ����:˸~V����d���� =�s��U�郝������wrpT�B ��#O�5���%��F�T^��z���F)���"iR�W�ϭ[ �����&�spHx-d��fkk�17�����+�y.�k�Gn���e�Ons$g{�-�%M���^��\][��U8v���`t��W�ш_M�Đ[i��w�@�Z2���? ��hӃk�k^	�`�A�i)uR���z,heG��j�`8�v9: ��B��(˷���)3�l�#���n���זK�V��n��R��=�Xz��>���\��L�_�>�ńS{�����2�y���۩�,Q+g�hDh��a��y�H��:�������yh��(���v�3����	��+�<�0�@.�	-�'��Rb�����f���Y�h�K~�����'K|q;�/��[�N�&&��ܚ�a���;�V��0���d����R���L17���S�1G&|��T���i��84��n�qe/Rōp�HI,h��dAڒ���o�˖�-��\��t{5�9N�KL. �'[FGns^���Y.���|(S�qD��u����5�^�L�)FPc�\�U��lsCBa�4f]���C�b�]��mIu26A����z~��2x���'r�2F�pC�/3�|�Jy[b�� ���6�E-W�Β�ZϺk=f�L�*�#D;,�Ϭ�"Ԣ��ć^��:���1^�Z��ͅ���%�n�Zc8�T��3M̨*��GD]��*�D�7%�:Yg̃���NFT)u0��}�U"�J�=`d����B�3�?[^V?܄�����?�c��+/ZPhpl#�\�W*Y�1��s��g��=%������ޫ�7��y��;�8J�K��|.JZ�t���tX�v�V�U��9���}�eTUcuz��2i�D<�7tc�c�R�g1 &v(��E	K�gg���9.Q˩. ��'͔o��BT Vg�$�%����Y�h��
�ړ�*|l��S껩Kӟn��J=�W<�
Ajg��ɠ�0fx��A�����:�U_!~��mߦǅ�P��+����wH�#�f%lH���r��f����_vlc�������E;���L��P���qL>�*{�,��_n�5C���qĐy4_�,�(
�Ꮑ\�3b2�1L�x�9bG�D�+��rx,l��郒� �`V0d�]sZ5��^�h��Zb��#����gЇ28�(�&6�A��I2�_��c%��:�v�ٌ��J�WΝ�鉜`d���Φd�=��|B�T��F�����d	��ZW`A|x��IY�c<�vs7_.Ł�F�1Z�
49N>Q�\`ȝdl�T�\J���*���;��x�L�����Nry
of���Kf\��-l<'<>���ߘd�p��ĢW�h~NZ�%-4�x�*��׎Z���O0q���+J/��H��_8E.O<�T^���,�t����|�^�h��v&KX�He��0ٓB-�4/����v���[��nR��Y�p@
�_�-�dau�5��P���xf����d�ĳ$ �wx����t�����~�
�Oi�b����y�Så�.��y�\|p0��>bƞ&Ų�����Y���1"
��fȱ]C���,���ҩ����&8+2��xtZ����,�H�%E0},)���5�$G�f_��Fp�͆
��W��SH��{����O^a��A�;3��<�_��)�����P�Q�N=�}�k-�T�nt��:Cb���ZN���?������#l����}"th�I��L�n��APPz�Fe�+��a����Η�1�6j'+H�P���B�3ϙ����B0��C3+�A�᬴�k�r����/����Gj��� �DVVIT�����=5�x���'@�3�5Q�쏼rmD
��2����W���!���u��hd2�=�+9��;:�щc����pcW.�7��������({��i�3�NsnLtXBc{(�,�Y%N:�e4$����/Zz�|*������M�;�C��E+%1��Su-�{�͈X��w+XLx��7��4��`��M�sK��Ҭx-u0��R�珍=}l�N��- hM�I��u�����c[����i8eUb�h��KARx�*�Ǹ��"5����(�ظ�qtt�9��@�o��{���XK�a�[l�-<�
/�����}�v�F��QUge.�z;-�T9r-Pw�K}�@�,u�M�K��|׼`N�S���N>�$�̊���)�YSj����*��Q����m&�5V2�-��g��e�\.�as��ФN(�°�"�d皗��ȵ����a[�< �X���%7 �.m���h��&�Y#�K�����ӧ)%�@�{?~�Q�v!t�m���8�E�����} �;*}�ް���v���^/�y����I`@.l}�����`}.�Ţm�}ά�+:.���D���S�B'A˽�"6�IƉ4�ZA+�ʆ�1}*����.����m���c�(�Z��!	�'����t�����nʆgn�^:(~|�a�p��H��4�G��D��"���w�#��u<�i�k�ʑ���QH=�}�Fÿ��>�(���H�!O��Ӊ|��5l��C���-�QfqJ%]QJ�D�#P$��5��Ly���Z������*��r�q)�[�����54�NQ�Υ�t�k��"}�\�^O$~�%:B_HҘ��8�����9^>\��&~��r���x�R�g�ܩ�<��i߉���R�U����~�ل�����5�Rpǥ̶ S!�̱��i����X �X�g%Fn��g�1C_��wZ�-���#��45}��0�Vt����̵���-�
H�DD���u�~�#/"1SV�j�*Yr�z��p +�ƿ f���,���g0)��]\
���jhN���Um��|����P,��` E��$3�nH��x�ޡ���:������axu���%�2��B���(n��l�M1���	G��΅��0�y�Î
���&xS�[)���o�p˯7L�!��D�Y��|�t�&mj�P�2�Y�9���,D^������fGF��r��a=�l9P�}��[��֨٢5����Y��;�"�2PFT ÊNs�㞜�SR79¸�*�_���/��7�D��|E;�}�h�4���A��HIĎ�b�[�mm��h �p&i��.���@q�p�Br�*��ܴ��a\u��3���W4?��z�~�0�y`��"�2Ssh�{(a��{P�Z�V�h��}���4W%$���~�pq�����r���K�}�%ځ�Z��",��}�}~�Ara��.kK�
K,0�ǘ�pW�ķ���~��A��׆��u��&L���{T�?}��^�V��2��ؤ��2J�������ʨ�p3ј��rV-�Hm����#)�t�G~	�����C�bBd�P�Z9�Ǘ��֤o���V��9i��ׯ����l@������P9_��H�����
�������\ٚIW0�k�o�븣%��,>�����d$��'=C����4�����Q2՝4��P��1Z�b,s�j޶�U29˥$���������6�g�/t�|@�%?���b��&��;y$�8�l@Z}3�|�QujSO"�i����a8�.������_��oç��T�-S�Y��!�H���H���:�p���b����!�w���Lɋ"-�&B�BFɺ�*���j�j �&c��f�2#���u?ꕵ�ۖQ:9�O~�dbhaa�]>��MnS�H�V7��hH߅;P���럋lV9��Gn����1?��[+9@sY�je��bŷ�[����L�闑D�=�q/����/��F 5�`��wrt&�L�v2j=�FPd(��c��Z�w;#�~�#�p#���F GǶ�p}ө�D�ҍ����(m�n�Wfb�a�"LL{q�c�KJ����+��F+�����OvV�N�C��Ky��j�W0j<]�H��������)pȃ�"�av�w��E5ći�#N���r��*��re�
?��W{Js�h��H�b��Sc�+�=��##דs"( �
����G]X��p�|b��ܐ�-����9iM`�"���m1c�E�O�M��E\�J�|�V���pp=���D�c� �mC!*�MxM�Q<E[�!��g�X�Οg᜺�h�8g�^pwa6
KyԒWpg������}|�łJ�At<���= k ��f~���)�Z���Rޡ��{������"�ԗM�Y@�j�(�(���#��l����\��ή@�ǤՁ�#)���ۗ�6�}j\O琢 ��K�`'�L���7Ǆ	aibM��$��fC�F_%�������SU�Dr�qVp	o�=.�4�}[���B*,�E!��ʼ�)�H�Jv8ssw��BB��� N��_�=��g�����r�	B�^�
��#� ����8�Ty��+�Y��� G�_]�"S�V��W��O'��[i�����^/�ե�(���ǃ&�C��)T��We-� �5�72S�`�\��g���9���&ez�E�֔���:��u�Zj-L�����L4򇮡��(z��UG��sMy��{�'B��
��0���hrf�P 2\�OH��(��k�ׄ�-�m����0�2"Q*q��K�-�uFL�L� ��-�Ԡӏ�N����u���R�*S.��7��~O9C~w�D�ئ����J��⶿f�`�`�0�60����5�Q���(*	�m
d�Cu'�j˘����g� �9�K�w-|>�=t�`��b�Y���c��e��?l�݁� ����ML�F�뷾+M�Wy�S�;[|4��n����N�/U��SBzh��ht�zKs�����Ge�Ix�>�x�2ʪ��KO
�T�����q����O0��^n��u�����<޷w��:��0C�
�Q�g��1���*f��o�Z�Mݻe��a�����s2m^������n/o�۫<>#@nCV�K�[<��<�=`�Z���^�������j��v:�v�0����I����ڞ�UϽ����|���������^"�Α;Tu��/x �y�u
Q�覩?�4��,�j�� �e����SU�i}%�w�k2�ds�g�E��8��H�/FXA�ZH%
V��=�+%�)�ߐ M��]0V����+
���|������Z,�&��Vc����r�9z�� ��p��gV��/��Ý��m��! $ �R�����l���C"(��Uj9ߗD��N�KN��2����wG�c��V�
�M���ƶ���ڏ�/�Z��H���!^�-�b/"��n`=�kG@��� ��q� ز<��ٺ�_f33}���YG��ÐJT��R��IV+�)�ﶖ�3��42�|���L���f�J�>�¨���T�р��������8`�}�����k]o۱'p;Y;��41�ұ�c;�V�>��Y[�7�$ݔ��/����j&�1l	n�H�oL_����ݠ�7�0�A�L����Oo��44bݸ�p6�P)mV�It��՟����0UJ�Hi�og�伪��;t�;���BO�X߃\�$�a�q	�BG�.ͶQ��Ӭ� tL�`���|!Y�X���Jj��kd�'	)��
��_�0��?Y��yR�`���p��K�I�j��W���e��>4�G�c���#�L	�ϫ��s�g6@�Bt6;��ғ�N��ŧ�yƭ�y�t���)8�>f��|=��m*0y��
�����~|<#��#	gm�x@�	����_W�d��9��[�.�:����>�QPy�E�:yD�����O��~c\O�D4!Y�Ų���ƉB�)�]��)r��]�懲���d�BO���L3�m\/Dr��3���T�-:����>�Q1�NΩӆ����}HU�s�J�t�G�R�y��G۶X���P�]�G��j^[?�A��<�F2��%&�j��(2�w�dY���Hw�C�`��&i�2��GFg��t��el��dCS�x�=�q`������s�Ü�U��U��u��(#>u��Q�R��6-}κ��y���`u'á�ptܴ��M!�$g�7��9��F�u+��/Je�C	�9���� �l���y= ��We�I4�R�=�TV���-����η��d� ���4�yD�O ]�����h���U�E��[!Vf�r�|c�({�TJy��UC7��,�:�~M�X*N��K�T�hz�k}2���"��س�e�:�Y+�3����Q��Z%v�F�&8��̞8��3�/#��6_a��D�bC�]��t��'B�qn�ְ�;�sf��_���.�L�E�֝R�h��ys]OC�5����oß���
�'dW�Zʁ�����N���GVC��ڳ�O�$nn�M��K1�zd��RQjQ���S�;�	�H��
�R9�̘c{�6�$��7R����J,�� �%	�v�t�����r�N2�Jn��F0dw�寣�C�A���I>M�lqD��E�epGM:fs��T��eZgyW���p��J���p}'��A��B(�Y�p�b���5\�7�G�AP�*�k>$���f~(�:e6�J	O�hE�b����J+�0�ҕK����,�	�E���t�3jf�S_
�M��J����H����fޯlw�槎��),բS��`t����#7M�Xfzjs�1T�F��̝�i,_r�5=^���ڂ �L�WTan��Wj���f ��"?)����ӟ*}�ٜ�%Ѫ2
^�0�@sͳ�0����5]J<�\?�Vр+�ܚP�
�̟"V�\V/�,*z;�퇎��W��إ�Z�4��3V �tH7�X��AxqҬ������'<��?���)>OY��f/N�����v��J�p�"E�/6���EB�g�-���{
�"�bs���.V�q���e,��i�_�gz��������Ӕ�32����L�X�|Ε8���O�*�t�S�̲�LսɅ��b[�ҮDYL˱�k>���{����X	�=�~�L�ܸZ���{�RW�f?H�5��UE�{��#�Mi����2BJ(�s�n��P���,]i����UTk�H���k���;ߣ�3�xu6���n� � �J�i)�Ue�n�/��6���'׾�/렣�^��Br��.U�Zn!���NƐ�w8��Z�o����s%����S|�!�#�?,�1!�ot��MH1���z��H�I�c�O%Օ�������s��eܞ���|y�U�ypҥ?s �ʟ@�SJl]���A������@�� �sv[6�q�j(ʟ�Z�s�WR\Eu��o����� �%�}������[�6��L�ۚQ��ͤ�AB6���pY��e���d����V�A��y4rv�9� �-3������j�TL|��p�`#/iy`ع����ʡюP��K�{5.���8�T6��y)�߆7�B�����ބ�L�"a.�i�֪kaF�;T��Wx�����5�R���%��l��������vR��3��Աo;��+z0�A���(�觋=	�L�Q�,����[o�%9x�an �yu��45B`��D仲e�lDI�u�o�$+���H+������z92�ۡ!V��#Ԓ{f��%A�ߍ!.]v��&>�U@]�Y��+]��U���!�;I��ڎ��� \d��e�͊&ى�)�#�Xz�Ҟ_��>~���"�d��$��f�FgH�-X1/��m��TlrCEV��*E.�nr�H ���pZH�<�0/�
�~{��WcW���G��Mcf��T�֯g���y���o��Q�(#K��VC_P 2���U���!'����Y՗��>	:D�5Jd��>�٥X�L ��>�}-�P]h#<P��H��f�pn�Q���||���7�T�p�L��PٟR�~X;�M����k9[�y]p��=d%�ӑ��:�Sx�j�χ�7��b��@`2�J��yf�T;t��`z�����k5 !�f���_u+�Ȋ�n/B#�9�&���9���8�E�HH�DKŭN���U�����䚲�G�P�W6}bN�s���]{�qwi�������Գ��ȗm��j�b�|������������>���:��Z:�f'}]l]�C��^tL?���zB��.��ta)_"�B�B��U^F�T�������U/�o�L�I|�[O��|z�h2��>�oIJ��	��ie@��4�V��=𬂭W��s@�ft\��4%�T4��W�o�Jʨt*Xw�6 �[���d1�MD~�a� K�-�6P�:`x���G��wv.��T������s�
J��;h`�ů�D6V���9Te��c��`��盏�h0~Ja���2IGٲd�un�3O�V��p$7�4������~�]��
�ٺ��7�@E4�$W0З��w��pF]��7}�}e1A�a�Y��d~���k���r4�47k�!y�&�ߦ��	��}�3�z�d�Zo��h��Ol%�-���=� b=Yա��ðլv�t�6����k��Y�ƧO���TDe������e���oU��*���9�o��6��t�y��٭�e�V3�)���]�g�pg�V����K��<�Pr�V�aY�R4H(B�([S�􆋔��l��\ٞ 
��Vy�t��=�|5IW�i(\�iT]�i��؈]o��]_� O��yt�x�"�l����aCP�jp]̖M�vI �$(�_~Z�y�����a�m�IZ�W�m{�� �w ƫ�=�J�)S�H�q'�Q�2��{���Ή ��Zϣ��&���g�8�暨���膣$��#p�Bh((0�U�P>�v�\$[���o�w�M�(�ͯJ}��d?Bh9��)_���|nZ�b/�|��r$rCI�w��q��o�c:-*�����a�NQm��������8�^����%��㮀nx�q�q��h�n���&�W�8f����]W���N�z&��oJb��uA�/�Ь�Aq��>Ray[��Ek�
�;�U@wQ��hFnNj&�إ<��ns��B���(Ō�x���nؚ�k'��f���w�p����K|2�C*�+��c;xSpD�5�ډ���\�§��jDS�^n� �4~��lF�g�-���b�b������
۔ �rGJR�e�]6ݭ��7 ����G��dD1�)�ԏ��	R�(���qi���z�蔥��$��nYa��D�=m�z@�o5��u��MN�~�F�;b�|eFX�NPt�Z����/z�jU�k��(!��:l�cԑ����lK2D�L���|�y�}�-��QZ�t����S� b\ey\�P� ���Vօ����E���u�y���f�<'���"yig�#���n�.5�>}xM��z��1�鑡�S�h��+`n@8�iK���'L�[�/��l*֫Œ����)\.:Y ���h�D�����\zMp�A�I�;a���� ��@�;���Ѥ&|�o�;+���X,	i8���~�K�����U��/��i ک�'�����I�L�<�{�ŷ��Q�Zj��pFtzDk߅W��!�[� lQ�����0�(ܮ�&9��_���`��;>C[Gd�OЂ�է���Xd��,XE�&��O��|Sn�k�%t���2.��We۝a7.k�;��i��VW�뢱k6�8�Dè���d�['�EQ�h��ϣ�tc9�Ed�be�J�m��{+v71�o��e����ґ$!�n��,Xn1��H�;Q��q&�1���O��EV3"�[�W�+4J?�jw��1s�"^�ApJC_f5��NV7�\��ն�e,���2�*D��L2�� �h�����ӊ��Sf��@�B���~�F݉���q�i����1��~TN���Ad�6|���>nd�|�X���b�Zn����5A�^�&v�*}t�|�v��HW��Yۿ���^ÎSN��J���J
X����H{m��;��K=�� �[I������+�$�8M��7����$�?��y�*]�����r�Qt������>��
J�/��͔���@j�<-�m��mwUQ/�X�X6��c�}�W�.�6�d�jp�04$֘1a�S5o������!,mts��P�o�4U�x=�r���6P�&l�gy��-���՚�X��!,��f�j��n)�V�,��H�.�����fN�����ۈ�i����J�°�D�~X�T��DgS��0%QD��u2�A�"i�W&��>9t��������k�J�'��Q��s�0g*�٘���]f�]���/�[��j�[Y��؂�Nx���V�o���o���篋#f�2�5I�[:]�zI�*���o���4���P4q�Ŀ�#e�9�;K�,f�=o�)��5�*2<m ~!N��{�5��#���(!q%`��^~tv�oW���:����O�ɑ��/]UGF��%�T7�W�ݪ�`�H&�zhϿn�d~�r�n���NɅ�StG`�Q}dm��-�i��ʓ���m su,A+m,	�Q3#�Y*�*<��B��J1���[��W'�$��'�b:�I~pM�5n�+T���N[%�u�jL+&t�U���@��Wu/�p"̪��_�>��/�5�ض�n�j���N�~��9�Oe�@�{/}�S�8���y"�n�c��	�K�oՋZ�W@�u�RktS�!�M�y΃��6:�.i~F؍	dh�62�>����]r������k�P����X#�j˝-�2��e;Cl�K� @�<�2h�"EI�ޙ�� ���6�\��" _�8	ܪ����6�:�⋨�C��y%ش2'��e-����]q�:��E��m*�A�r�iwI���5^JrT�*��Y6v{U�u�Ȏ�/��Fơ��)��3m�.�lv!������`�p��`�	���O����Ԏ�\��!�\3�z\bs���ʸ!��eF�骾b#�|�?��Bj������6۞�d�x��뛣3�xYj�x��OA,ӏC��.���:��H%�@��m�W�>Q�q؍���h�y���M������Y0{��F�{`�x�᭲(�������eD� �Qӓ	��b쌵�
('ZX.P��?J�@�G��ΕY�rx��_6]*���z��PS�_თ���6P��$"GE`�I�_��{Z��on��] ����q�Z�-����FHf:�Gٟ�ڋ{k��D�zG�!u�~'��i`��~D������^��F�Ϊ��/_���B6�z�������-s�Hn�{�+��]�x��/��ө��0�$H�b
|��F]"o���r
�����U�ot��:��$W�W�[o\�"n�D�M���?����Q�%��.��*��C�ujD���n�S*�VI92 �_�
������F ��]�빵�l�EH-�%A���2�"���*��TB}�e�a��v�[��0��D�F%��v⪫-�յ�Ƨ �ɮG[�a��U�:<%}�}=�����¦D2S�S�9h�&
�k&����\�a���S���o��Z�X1^�:�-6'	/o2 ]]�Ӆ���jɇ�\��:��{|��+$�ϋ{;>���?Qk�{k|�*ܡ�\�w�vq(Q��������{�&���{:l?.�r=td��k���yK�z�_�W[��0��&������~K��R����J�U)�fHan�N<��B�$�����o�#�T:�IGg�E�!���I�T1D�7/���?�e�=Ҧ�7>�qV:�?S�C)�Ϲ����R��C��[�<3�Q��1m�P0gb������2fZ"�9��6�z4V[#�#c7��!���?�����n��9xB������&s悐���o�i7-KF�+��q�X�0[�E�Q�1�%p�[�|�a�,��;_j�D�U�BnfU��s9	ַZ�#_^�}���ߟ���49|u� ���O��	Q,`[0(p�Z2NȲp�A��׀�(�k��dl�3Ξ�1U��n�|���S�	|�s֣� ��'M*�3�+�f��"���w� ���Ѣ�,*W�h._�W\[��zG7�;�kT�=@��(�0��N$v=��K�	U��e��M�q(�z�	�[D��3c@�I���.拿g{%�rfV~��Kh��qg����С��u�E�5F�'��4�;�?��ս6�spOnX��@z�1!��;U#		j�u(}
<i�X�<�sŽ6y�b��?X��uf7җ9_F�d�ɍň��*� �>7�!�� �V��(!4�N����!+^��f��:�F~�OX��Ưߵ{��@P55���{	8�."D�����Y��f�a-�X�NM�ˎ72z���FB�п-�g�tE�_&�_�}��'e3�����_~����4�p!m8F���N���A� >z�k�����J]X�w ��ؾ83m���))�4#�\�	.Ӫ"�F�n�܂�TD��S���>�?�nZ,�yK*YN2��4:�T	%/�6��>?�+?��y�nU� ��$Y���9%/oA��B�����Ŭ˥��׎�v�Ak�Dsp~����l4�/O�q��J`�|��k�;��K��_�N�&,q�K�Zb�����w��1'S�|��������b%̓e�g�P�b�S�?�G/cx=�'�~{f���3�Pz��g%��A��V�'I�0�EB�0�X�0-�2y�bTk�@�W(�65�*���s��ByY�r�8�-l����R���r s���5���K��8n��q �� �8�r�h�ɦq7����O���57E��������2�>m;i����5�K ��94�����w1��顳�r�s�����M]`�\�x IZN�،�+L�=,'t�$Y����W��TཱིC�p�-���V��M���$Kl[�l]'RxJ�����ݣ�����W��+��a*^ j���*�OauoL50os� R�+f�(v�"`�fo�Hsuӌ�DZ��;��I�d�� k�xv����q�b�q�U�y���.����
�����>@2(�>���$���ё,ŵÿ��Z�ީ�L��=�Z�nk5�2�JDv�j��5B��Fd4���{�sJ�̭�V��}�/kt)wߎ~�������q1֘t@��K�wA�-��r����<OgedhL��玱p��l�D�P`��Ƴ��}��K�y� �!���>�$U7��)���eYk^��+p{�"} ���5��7���액�����N�?v=���r�>����QǸi��d;mQCYS�����DͶ�uN�V�/��}6ݪ��=���v]�����,*���+��va˞���j�yׇ�j1�Jޞ��oo�c26$��?~<�ȣ��	F �X� s��5�7�c���m7QY#�o+nKD%�w�$n*c���b837���Qs@���<t?�:l����S��:$�Η> `Ϩb��e*2�����ZC���u]����f3K��(��w�Q{�J�61����|Ѵ` P��Zore�6�Xu��/|8R;8�q�����(��on�n%8j��Q>)��u/�c��Ԭ�MFr(����NM\{s��vp-�=��@���k	3a.k���	n�d���@	,��H�J\<wcK�HG!�?����n+4!W��.���a�5&�}I�cJ��*&�&f��4u72WTMY�
��Ë6���HjG;���7tn�\	q�C�s���-������o�ʂQ����D��;h�ɜPU�_"����Z���!�@�'��(��1̈�a�1�Q��[JFnA�W�he w��a�)[�ڷL�L,n%;r��O��L���Թ��t�j[D��p{�$~��A|&�s"u]��]�.��#��Z6#��ϛ�F�-|�X8PD��a�e2�^yZ3�a��I��
/�
��P�>5�]��̟B�&���J�h��7�YK75�MPa�ؔ[�`�{Gs�u1,L�����J�N��
xR$�[IDD�]�����;�Ƹ���C(�4���[!gfX���$C.�b�ш����?�n����V�a�D"%��&�����,ޭ�@���ڏ�Ŕ��#�A�Q/4
���[p�uC�Q�k�YWJ��J��������<�
�֖��7N	�]Xl{��%�`9�|kb�Ȇ-"IQ�Ua�DI�/�3�6�ր� ^���'̌^y���^Z\hŴ6.H�9���@X] ��*n�\.Ľ����
	u�x�|�<g*��4	���w�v���D��ݙ�]i�Z�IV��b�D����V�+.&���G��?Ȟ:����Z�/��z ����	N�*U�+0��H�@8��T�?su�}��`��cO�O��=5�z�_���]������������s�s"?�E��<��kca~1����C��;m�^M�����瑪�@![ϨSV,/f�k@��͟x��*�u]�����٦&jf5�vbH�8�2�A!�`��@v;=-ւ����]'�r�H_�(��]��*ڴB��$%2 BJ5�K�{<�
��y��d����-�=��� �;L	���~#jh�N�,�(n�����D�Ɓ]^;lFt!�o��Nw�)�HQc�Dp�Xs~�u��ȚzNcF�4��U{�}�IT�B�^$����~�eucr��I?�h�I=T��o(�R+���1ɡ�(|D�\$O'P������GB;�`��2	�{C�_m�)4�2���O���'L1��Ϥ��f�F|- ��p2û�U���5�^:�|��3n�e��'��V��Qf�1`��R˒Е��7���/X¨(�ePI��F����Z�<���)���7q�X�
��������#����A>��� �I�Sq�>)���1�yX<-��A�Oe��T�6gz2���H��D�`=+j���n`H�P !`�7�} B��+ٺ�Beë�u�N�CV�AW��vY���B�wy(2���+R���,	�`yS����m�ۛh�@m�C˗�Hk�!��`�r���eg���u������3��~��:+�e0XR�������Fy��4dTĜ�tKx�y���x6_�2���7��\�H	���Cy�l�Ť�O�"���_�m�a���,X��>��#%Dx����0g�� �'嫩WI��^r8�Z��/�B�PP�?f!-b���H٬H��J�ß~�^�{���	�:�U�����cu��27̽� ��^��ӊ�۹d�>� ���SH`�lJ��,'L<�%9�����ej�5Ǖ����A�4�6��*��TK�D8n~2�9���'�由�QFs�$]�;�m��(�5@+��un�ڛ�'�Jc�!����r�$�ڬ�ơ��������t�E��=�t�b���vC��L ��PD���1�̎U�PY����r� =��7L��ȓ�p�a@�&�3�uMW�K�>!<؟ޓ�3���z���j`�н՛؁	����[
&k��Ԯ���C��S���x�1��C!�?J��L�����@�X�O�ܺ���K�vV�'��N9ŉ��Hp�Q�'��_�$.Ye�Pjoo-sD��!O��3kP��0���Yag(j��U�ش��cO>�3����^��j�`͠��d�����&���	�\�a�+��K;XL�`͓�q󏓌�y������8𢻯�DT϶,�vv�]���>P�zꢵQw|��;O�F�ƶ]�}�amm:�`U�M��� _gP6B_�!A���*�{C�Y���ۏ��}.afHO�9zp1�1��CуULjb����	L��Xnj}�=t0Ud扇a�(�Xo�&�gK�L��y����=g��K��p�������|k��yWz��4��4G #��y'��J�5���?̈́�o��Gʊ�8e�����r���Y�JF�7X�0�u�G�X��|�p��=NNt�Dώ&h{�f/*��X�^x���p�&����3�C�޶Oz%ksƱ�����m��~�ŮN��n2ݕ�p�AUAB�̛o/VB�9m���$�̹�����Z�2~6�:�'p��Y�T+��{N�DT���ҙy���_�*W=��uj�VQՔ�H��LX%o���]�2/n#PI{�U'�HQ���Đ�~� ���= ̒Yt�w��9e[�l#�!C���3<a
���Z{Ah��igd�,_G+��\j"jN{$� +s��e���Qa�|���~��<+�t��17g��q^^X�v�8��fش��Ƽ���BV�����QY	ˡؕ���D��	�����{ʐ,�˨��H�4�~h�+}��(K�7ϕ&��e1NGL�P7m��繼k,�x���π�4W��D�_��'�A�P�r#��RV��.{����0�:~GG���wf=j�H��^眷���?��W����e�M���!s���Z��3P�%�s�XW����z�ӛ�АO�>�(����������/�� P�?�D�qK�g��,�����9X�z�$��k������bA�ɝwMp���K5�S����q�k�>Z.{1�:�x��1�D�b>�!qo�T��;L4=������>��˕ n܀NI�G�2�5?r�I���{]Ż콮�-�0Vj��Pw)^��U��,�:�9�04�ƽ8���Ѫ �<X�
8�;|��	�8�M��~�oˮ��G����ز�N��߇_"�j��%"�.�5��6�O�[N��V�F�HJ�]�"�`��g���j�U|�ƞ���zM����9�x��V��.R�k�2��xz������5L~�d���cT��a �V���e���D�#�݂������g2MhY�n��)��ރ�"e��lk���d���:t��K2��Y���|1S��#�@��Oټ����0���K�H�[���E��������:ږ&P ��E(gy�����#Q��kw��u8� >+�N�@D�������h���74F �S
��PG9�	Dh���i��T�S&_F�}D��&~��X�RIpp��f;���9����Ke�J�ϩ�?/� 6��~H�R�u�}��I��Qu�h�>[�?����D�wϾ���Q�p>�l}=@t�
�2��[���@� }I<v�Y�����| yz�d�@�S��uZ9��`;��O}W�K ��纪y��c����ݣ9�w�.����_]���΢�xȫ���C��·��)[K\��*N��i?�Ԙb}����k� ok��a�𼨚�K@7�Cu�f���+�C�.�)q2 �St 0M�.����Ah�"�	��X�$���Q�S� q$�C���3u��oh��`h�	�ׇ�\�U�P.�;,���SYy�B���Rx ����CLA<���ٕ�T�T&�!�H�q�$��r����
�����ޑ/�>x�G/� �m0���m]�1��y�wJ^�nػh�'�̬��vh6�7A�J6r��e��Ȥ�e)'ǥ&`=�mͭ�S:���)��\}s#��:�鳍%�	�(��r�"D���Ȫ9,�kK2�O#�T����VD��O9c��������X7��#���2{����#;�O���hӎ&CGD��V�����/�Ԩyg�W��J�ʕre�S���U��!�[�8V([1����zj�
�7E2)�g�Ȕ`>ِ?L������H�c[.�8N�������2T;��,�"�[��������4}wZŴW�6�6d�����xzǉ�lWl����$�8�i�h�-��wr|�.Vs�R���&�	�@�;h�S�jE>��/�%j��b�(�q���4\w�k��L����a¢¥خ�;&H$�D�5���0p�U�e��zP��Ҏ̟2/����@]n��F"��4�r�Z|��#�ez(1ǖ�x�>��h(49�͉<"�#e��`O]}�ݞ@�Ԃ���6��g.�FJB���&�i�h���}(7i3)Ì��ۜ��8�;�~�����mY_�� g�z����=�����u�.�v�zs ���M�Թ���1��9t^ ��,$�D��	wI�DJ){���b������9�olx���D�1�i�< '��ԁ��/��,E�'��0&А�ԂϷ�3������5��x�\)y&I�ُ'���5kAR�  ���k�!q�u��<����:7��T2�:�p|Y�44�c����у�1�ƈ*Zd�b�����z-J3�����i�ږV*�e楌'��2h�P�,��/v�o��֑#���3_b�Z�>~����`'�����oTmY<�Aܟ�s@"'�����u����7{+
�rh�J8aTfR�O��u���>��ܱ�i*lǅ`��b,t�&r5� ��D�<-R���Cb;������	o��.s|�r��U7!��Q���)���k*���v���S��&t�k/�o*3'XRf&�-4�>��|w����T��l��/L�G��Q?���JH;��٢�����G]�E�Z2�Y)�=W��;M[�2��|3p�;{17s&�M�e�Yߙ9ŪԁوU�ߑ�'<��/�5C&(^�����|�[w}�'�/!%H��w�
hn�߃�5`R�UK���*fN43ɂ_�~��D�)��V��q2S������^��zbBm�}]@O
����WN�O��(*e�vE�w�|�hC���_�c˅$齿�/��x{A�p��L�5y'u�|�u���==*��ֳ���Y%���+�*l�WcM(D�.o�㖟!^�g�D]�~��PH[��v9�C�N�+�~��]�Ƿ5ā!��#�������m�$rv���HӮ�&|�zy����o��S��b�C�RBlZ|.��[�/�Y�6p\��g�JE�p���"���+"�Z�Ω8�,&��WA홌'`����15<#�?��Sʳ*��E���P�I�_UH�q��AP�nU�,	l�v���͸�YB)4�w_�D_�՘D�?��Ev&�#;ctD FP/���k��`I�4!��̎�K��h���	'Iީ	�R����1��	��ռW�C����-h��B��m�GO���f��;W���7�&_&s7�C��WXY��؋Mٮ�0���E,����E�1GӀ[�b��S�GFHӏ32w�z7��WOF���ϒf�R�xG$�D�B��U�Ovi1�Y1R��O�(��U,�ΕU6�Uv ;�j'޸/�.��*t��|�VP<D��d�����{��k��H�7}��v���C�v��O��MU�-VtѠ�v���r+.�C�����DI���2���>��M��%d}��l�)fo��UR�ނ����GF��-��b���ͻ�D�l�*�w��A%(���&�&%�<ۃ�&��3F��Var3�}k/D��Al�$��"�i�\g˨0 V%b��m��kb�0�+S�X�Ks�2��y��1�v�{�آ?�����}� ���7�Ke	�Ip�ȥ,8��l�q�EW���[Q�e�kU<���h�1��z�3������`28(b�f�
&�N��WJ�.&`T�B�`�-u&G��b�8����B��,����G<J��Øړx��txM��'h���[��Fx���>��8������-�\È]y'��K�5��Α��y�O�7(�מ�ح����#�Y���2҆}"��K�^Msפ��u�8[���.�U���si�ܘ�O�����Z�(�/3V�%cT�~��ّ�ݺeJ�E�U~V�PK{��س�U���, �����M,��)���m<D���O�r�⭏��	~u0�)
��,��Onn�3�%��J�a"{�Yf��ѧ%��᪎7|�C&��	���*�英��]���!�8�:��,�ҋК��(Y��������X��mcM�j�$U�%Y.�������'E�q���q�k�1�,hg���lli>j��!��y�����+����=˲�����n6)��I��U+q�!��f������h
�ʶ��������[B#t�!/�
�T@|���+!6�)���&9�9L�lcZ/���������.f�i��]
�ho&:Q�9B}�=H�.㚥��IQ���pa�pa��FS���4xj���R�"@,�WF��Sc�L<m���.s��� w��fc��6�0��39��f6�J�:J@=S	�^�1�;�a<���sd�E�Y��k�b��ꦿ�i"����F?�����#���/^�+�U�#,p�R�P�/��,���ÿ� ��|�C�]+�J17f�����!��CAQ��ۧ����@
�ͱ��'P	�����sܢ^م+:K��<֊�������(��~�a;��,Z9���F:�\k�~�Es�[c:O��6(�_ ��\cTTr���_ް�^�P="m�F��+u��bV#J_�:$%�#f��G��(�� ҝ|e���Ғ��1�P�z&Z���ӻa1̿g�~N��Y����z鬘K��k���Q�a2�U��Q:L����L�S_?_�0~��2�;�x�*�K�la��УtD�����
F,���F[FGEz=Gq!�����H�@�eCU�9����4��>A�.��(�a6��B5��O�qh%X�|���_){A��u��KwF����3�!��J�S�d������X#`��#�zs��t�V��5O��
_Z=�o3G��d}�M?�2��iHpE�8,���"���V�֭+.�a
ܡ��ZU�U�����6����i���Ȱ�¿����!X�R9�P��VhM���(O�!͟��Bn*W"���(G�nc�5���c ��~���he��$��M8�v���9$m+�����B�z-1d-�b�l�2;@�g �+/���钰|Ooh[�e��,�e�S,������j�������QnJ�U8��K��j��!O��?�TzX���yy0��@펈�u_`y�� ����/	o� ѱ4_Nq�~��ݣ&LUר�ԋ��Y�J)1�$�dWG�u�܂���J�������J�`O������(f�.�$�� �O1��C��ƴ���[���j++��(��"(�߳��|��A}D+�(������}���g�X��$��0� �0������hHm���n��C��A�{�E��A�����@�T�\!� ���3�2ɶ�7H+ǽYQa�hۇ��`8KZ��w�����@���y�R�y/�d*��`_oJ>X���91QO���uE�׋�9h}��y���^��_{���J���I��d�()ɲ���]t����A�v�����y	0����T5
4SI��/c)��Kڃ�OMQ���R)���0�A��fmo�����iWuJ�g��g��8�`8�,{�k)ǁ��V��f��	[hDd^��rR�r=�G�|�Y�F'4��]3����S���F�ɢ��w`��Z���D��s����|k�u�O��k��@l�D���R�䑴�kگ ,�:[���y˯�]��QMN�Yj���w�lݞ�].:��>����!��/@�a1�I����m��Z��f����X_R�,C�;`��(pu+�P9"��מ��?��*��N^A� X�V�nO��c�{������Ч��7��^�9u8�p9�a���Ž
A�|�T@P+eܶ�o�b@�fHD,y��!,�l�
���+Ua;Vf�?3,��N�^���ByOWu^�vF:1-e��g��x���k;�/�,1s۾'������!�lB��< ��?{L�V>�s�Tω��tAڲ
���{Z���2�����ݬ�fV]n�����x7\�x���3mlΞ��;6�%�M�5�H%k4��Q�0:
�l���/s����@^�󩨶���I&\��:<��bJIp�9�[���>��`^>��@�B�e�-����ݾc·%��.;��BE�� �׋���d�a�!ށ��L.%K<Qm��ᾼAT�ƙ	an�A�B�������=B�8� �M�E�sl�i�������d�:N�Y��8ҩ2GI'��9�̹O�6(�%�X�O�����x6�
Ik����*`�crpy5ld��:�E����W�IT�t=�%��q�}r:��e��G���_�v%��[�/Ċ(�m���fb�q0��6捝�z>4�/k�i�x�BQ\#\&z	\P�C��55��O�0�xPe"`e�����^\�.�{�Ȫ,��9w�S(��:p�e��`h��&���O�(m��݌z� !Vp��@�� �����!Ht Y��4�S@0!\��MT$�Y$D_�(ZoU+�pu\zs�b�u��oܒ�ʹ{��#�NX�� �(���rl��B4�O6G2dx�<OQ��;�,�K�c�����3-.J�vŒ��Q��C��Fj�m�$-Y�ΐ��J��y]#���xvoA��&�nn]��B�`)���΍�6��b�]��4К�p�2-M@��Q` �,
@�o�|d%t�9�n}::���zu7��g
���j��HR���k>�A��X?�\�BE�.�-05a����&{�-�7$�� �e�1�*7�Y�hx�>qs����y���0+����]7?rq���#AKcKt ��2N���u�>���GK��bs:Y����^��%�Yn�@_aF-rb�rG�F�G�B�����ax|��r�Hq��R7���1�ޫ�jaa��٨̆-m*�	#�	�(l��F`+*�2	��;�JH�Ϊ�z఺;�SP��6��b?��y�Sȫ0��U ��o����b8A;l�I���]W�EPxvlE�qg T��s}8@�/�x�
{��lcG�Mf�=�d��E�ij���{�ӣlcϿ�ȩ�+&����t��~Ō�YP�o�;8n�u_���@8o~�ǹ�
�����*�\�Yq�ܙ�Pwƞ�'h��szK <������JS��`R;s!&z�m]�|yJپq3P����
����%�!D/��&�үZ+X>,i�Ci�+�b��kb�����su��Ȕh��h:�e]��`�"�̺��&]����~)����mBwaϹ߉�j���	 `�މwX$R�G�$��dJ^���V���*=�}�͆���j��z�WD"�z-�
d���k�4lX�uT��Vqhq��g�k�)���ͼ��er��[��"�I\�0�s*�y6|_�اTE�U`и�����Ԧ�J��Ь��f�B��~J��>���
�xc'̰������H�F���+k�_$�Z�U�R�$

����M��a@�|0˝�w�����M=�sB���o�7�2���[��`3�'��63��y`��|�<��R�ٴBTi���i�3x��
	����ƅ6�S\���Rga*�L�=g��!��[+�Va�f�:L�I����r+B��n�|�vzULnU�tWm������tR�����$���F�~uqc��r�C�6�gb��i�%
���Vd5r��kf������R��u_����k�*�,��Y�hڍ)�r��/h/)���7v��}p�8��x^�ےآߵ�f�0�KúG�3��l�q��`�!�C�UY��U�t�Y6�h��-�
���#��|��ߘ��`���!1L�?���B&,��vR�͞-�W _/m�Q���~T8�(5*��h͖P�b�P������u=(�-P���}����~�Y�r�G��,!��̊�(�5I�|�xi��EP;��!�8e2���ġ�6(떧�R~Pʩ�	�z,�kϯ ����Lrۻ�h	����x9��+,��Mx���TD��Z��BY�qn��μoA����@�_ѧҒ�v��J(";{�:��۫-}��x�]�T�-��؁�N+�f̡L��P���\��4��%<�Su��9��VA-��9����H�6iL��k�����Ǹ2l�i�gn�1�j2��l ���?�&�ơT�q`��,������B��E��)F�jB�\�t	��c�b�=1N��ی�C���H��|͢ �G1��<�B^��U])k`��L+��l��z�[=D� 5���A��+���W��+^����p��1�Mz��!��#�����d�ܽ�	�* #��?�_M�>�֗tZt��G�zC��c�"u�)��������� �}6 �v� Q�� \��r-
=�q���r�O����-7� BC�h��q�p?��s�?�	$Ш�}QR��9���&�B�Sw꫷[�H�������NB�ldDN��o/=G�������x�Zu2��/�O]Љ.	��®��X�\6�<�s�y�NIˮF�S��1�ED��v�������>*�J&7��XѮB����3�sm������7���?n���Q [EؙGn8�zP	�䳙�e��������𞕡��g�%ut�������^�!0S�.F���zpV�(�ׄ���&2�.�a��0�h��{��t���@c��c��	��)���t���×$��AfIy��5'�$�;=2���-�j�6�ﵼhj�O��)~uF���:�!ާV�u� !7�u��HR^szl1�@o�� �H�b�����/����щ��l�Q?�B��V�.��� 6�����"���&��eQ58�G���3&�k�.��Ϣe���K95�D��������ځ��?[c�j���x��h.j�Q�r�_���g�3$_T��w�혞�wj<OjΛ>KV:��n�id}��8^�8^ެ�mq�ܜ����p�>���e�2�ح^q���k^,v��S���RjB4�=�T��ێ����A)�yUnJ�����S(�� :��Ԟ��nxg��b�H ��,� �I�;�A1:�{' �P�}�b������5v�i��=����W�)��	�%�c\�y�i�3#�c�g�x	F�f�(���%H�,ht�Y��zm�!�~����3���9����ᾠ�G$t� ��	�#�=p/�=���a6P�L���]���Y�O '�[�'{��Ge�k��_Ad�o-�.鲝�@,�D�a嫾E�_�pb�1��x�F�9��v�.Cn�B�+�Z��؝0%���U�l98��+�)����7`J�*��X��/��a�PK��* ��cfz�_˹(���0��s3�t�k���${?� Հ!�����?=�{���ŧ���_��`��]Ħ�~>Jùt��6�0����p] .�P��6�S��(D@M��Q�;�*˹����(ut/���Ӎ�k@�F���@z��7L/Ʌ.�h���C�i�A0�Y�7񖀈`���*�vg��(r=4�,d���m�p��.�;��ɉ����9��z(;徳���ccdœ�(�T��ٮ0I����&To�k������Z���ktX��V@��P�W���vzuC�H�\����"���k�:j�:o����u]0�k�&}� p�+I�\��+mq��*(<����dS���b���V �,��~�Xͺ����8���8{#aӌ����Ր��!�(���I?�� �}2�[�_�0�r�������b{IUoy5MYD���HS���S����.<��:!��6Tݙ�;����63�w݅���Yh\rHY�
����6��\��n�'��S��LD6��(he���
CX`��B��M1������Y8(GLѥx�{i��2E<ѥ� �eP��+� ?�J����;	l!�p`"�ОO1D<.�Z����(�Z0���)�A��G1e��K�>Y�PQL�1�㩟q���029B��̛�ĽTǎs�r���L��b˛hW :�I>��[��[�N2ĕHU_�j��@�beQ5?
$��	���i�K�,3xPv���|�9d80]��h}���/q�b�Áyå��1O�C9e�I��]7�S�x|/�H�0��M)���b�$������XS���O�5�?4l�v0��*T��
���3���E�r�gִ����N���2-7]�LF����W��R����ac��(M�Z"�[Ka����w��~���	�^��]���Py���r�h�>�����m���Ŋ�������i@p�Z֎�e^&��D����
��+khk4]���0W3����3��=�h�R&��Cu)���_�Q��vt.���o�FR:�>���-��Y����]�GP�dys.�7���G��*]�ѕ�]) ;_f��tUW�!X�z�*0���k��ckK*��G9��뎢>������F#'{��*´���;N�b�C�3Ri)��J��
����	�����s��؃�E?�é�"�:��2���S%�;P7{m���U]�Y��.ܷ}^T���t�c����Q���#�ڲ�/"[�J���Y�>y�������_o����jV6���b�1�.\�!V�9��8�XF����(���^��Pر�.��wN�Z풑G�CU-������]x��K�}���(X�ˣJ����j�ݫ���x@~j�q��h'<�46@��!�ϡ���:`��3�b������x��w�!��7g�LYI� +�v��4���q�d�	��
n@�O������.�JiI��f3�N՗�M�G*��P*��n]�px"}�i�a�+��l�˷��}�;��Յ���S"�&s�K@Y���.&d@��'𕌖�K1IG�p��B�����2 �Y??K!9o����?-�LF�}�Uq�{�3�������X��")�񙧣H��ȫ�pn����?���kJ�|�It�h�u�]��rH��rcH�b���u�C�BC1�)cv�I�A�YJ�v��_�c��Z$��������A�&7.�?�Z��h>��~�����2\3��LC��9��B���~m��q�ẈD��࿁�/��]�����rzT�8'�c�}���iB�����gOէ��D�����థ��M|��y�g�]֮�'��i����@FR��ǣ���pns_\�jcH�ߞ��OcZ�l��yƫx�������h��� ����t�v�Y��E3�c�7w�!\OF i�^������CԉCº8h�el����e�nQܱ�quy����֬]\
����c���H��·��)>�5�U�((�������v#������*pͳ�ͯ�X�g�E`�D��8UH����\��˚���#|	g��5��o �$z`ϊsD8���!n�̑���%��!!l"�z]D�4اj�љ��FKfVe�p�;ؓY�ϳ?P�H,=�p=�bNJ{5��7R�]�'1LW��@��ͬ�Oȧ�O�z,!���`cu�.&���D��N7""�MG�v�Ǖ_���S�J�P�5�2}Ȍ������L|�Q��M@q�R8:�(��,fOח�v����|�잹&Fr��������(�St���&;=��Gj���2Sq9ˉWE柂�s�F�a���=u�6��s��+�{i���(��Q�zc޺z(:�R\X����{nU�ܝo�
;{${Y�=L����W՟��a0jO�x��I!�?/�SUBQ'�W�p�C�a��b��()���Chu�~Eh�nW�ؘ�`7�EJOQ�C�vY��TP��Q��H�G�ٰx��R2�j�穵�,�(g�؆����C߯8�k?;�
?K�&s��9�X\��D![f] ��������)�1������$�o��tB������޺��vد��5�}�aDb:vr�ɰ �M����8ܑB�ƖZ��4C��6��3k��.D� /�n�l��W�J�ҟO�R�r@Y�'��Ũ���B��ȏ����e����<Z���&�kz�/>֒6�>=uSӞ�����l0�hJ�SUI��x�_r��p��Hx��odb��yP��'� vg_��N���fD;��?S�<"?YU���9A�^��ܳ0o#]^j:�GL�Lj4S�<�h�?Gj�[��;�W�b�o<�8o��o���l�ʍ�X�7)�F*����KIb����͖�w.��έ�r~LT��5%w���A�d/�Ɵ2��� l�xh+�W�U����;ο\	E����r��3���n�$��$\7W��1�9�1�m��R[Oy"j�^��� i�S��H����m{��ُG&���IُZ��#�����Z��l,Qt
����������I�b:ia:�ߪf���������Z+���>�/�G�-~r% 7��|���Z�@�H]�D��e8�+O�F��2�筋���B��/����Φ���Y�XP��-{�W��}^���X[u<7��!������_)c��I�BZC=Y1���¦���3�[\q�f
�U��{���~�{�2��eE��Z�H���=^�A����9�H����o�����׻���	���w�;��}�E������L=�>b��rW�38���20R6)��x#^a:�\J��������LD_�<o��wy�,�s�_ui'h"��0:��#����ڢ�d2������]�Bb8�kA�[�~�ʀ��h�����
��vʪ��RȰ�mfo��-�)�����p!�Vi#�!��ٞ3�� �9��vI��خhJ�Gn��&�4��I��n1�!�o�pX6?-��uQ��s�6�&r����O�P����:�+c`�z+~J�)���\����Z��	�ڽ�i�VC2��&���q�l�JU^��l0ԃ���0DYvw{0�9_�L���@HL��*j���s�L1�}���ϰ��T���^�K�"~����4N4�[�����N��ҭ!�o�8�5B��f��ӥ3��O-�������nB:W�ب=&�GLhY������b�&^�`�q�-즱��L.��@4��!c��L��G����zL<w�|Hp��i�>�^�-�\�`>� �I�Iu���ՌE�M�a�r7�:��˨�/�2��|^LΔ�]ͮU,��<�*�%��ʍޱ����u�p��!��q�"F�%P��#֗�k�@<�聋tR�_��I��*�_a�K.���{��_���O�`|��W�d6�}<WJf�C�M*���&ۘص��t� �\��"����`p�k�54����q����Am�%B%�݋�P�0��"�(�z����Z���%IՒ86>��R	�ގ��WۆD7K��������2�V�u�a�w��EV��e<4��}xP5�e��U�(,�U���ݥ*��%�U����]�c q�u�Z̻��&�{ (&������}�i5�hs��ũ�h�) iL�,è
�nW�|�M��|��M�'��us�$�1�m���p|%�\�Q�y���;��c�hZv`��9F��	7ju_F����rD���E�0F��H/�돿HE-)�r��� >'X��B�q����˦�f�a+s�2K5�W'Q�sꐂ�F���,vQ�;��7���6��uNr�&�Z,����t��(�p.�.�gc&l��= ���.dz��� M(�W��$FU���
�ԪV�v5�E8֖�Zؓ�fQ9_tu�T]������tIP^�������g0�L#Z���tU���T=��%F�{��,-�v5�.w�fH���qN��h�ȣ�M�.��Y���JG����� 84�+#�M-�y�9�κ�������N0 �R܏z���A�|�A�4$�ʿ�Y�����ڶ����g<�z����_���`�H����b�0�� |�Eճ���kN�{�0v6����Ǳ/\7v���yĿ��s��R������g�|��`���&��S����9�[Ϊ:���J��dy���w����"S��_���fGư�NO��B��129����CI]�{.%`\�>�����f�&�뜍l�>�7?��G8mˆf�ҼzvV�
yn��#��R~t��M!�P������e�P��@l,�y�أ�G�5!)�����s��cz ��2]`5����,�1𥳐3�I���%~F�K�Vۼ�W�� @�^�������<��4�S�ǖh>�f�(QV �N�!*�D�2wX^YB7�~~2�zF+�=��鹿a|�4��*^q∳Ѕ1Eo�lHlU���Hh�d[�.��Ş޿�J�c��%��\o��<;���>���0lG�P� -KB�=���q��/n�FH`V�����4b�0	���^�ǳf���%A�~�ұD�&_�j���.&�n��W�oN��o�1.�;��V�dq��(�g,hF&��y����a��+�H������_}aj�����s:���_>�trƨ#�GvZz�=�	��-8%YX�x��^�	��I��l����{7t�I��+���}�Т����49�������M7����hAI$;���7CY��>8�vO0�7h]r��+]��;����v\�����]9�$w��D�b�^ep�Ԣ��+7B�+&�J4�V1��>�
�U�c�/�Zc�X9�֘6U{xb���;:0�
��f�D� it��Ϯ�%�)a�5~���bcL��r���h���Y��W+�ٰqh�}t5n�Gur����r����� ^0p�^��/�K+@�N���l�v�?w4wP�0��}�[9�%by*}�9��� ��˥�@gJ��~P?�I ���?�^1��(Umn�E���g�x���@	�ur��p�B�}�� ��b�j�0������K0�S��g�\��S���P�߲�,�*J��(��H�����
V4���0�
�������Y4a����8d�ϊ/p�a+��5��I/l)϶���S+:��v%��q{Ics��\NTC<(^ǭA�|B}��q�x�'�߳!aWE�acC�*q��{?�Q�|�yvD>tW?�,���FJ7��3����PK�>�3���O�W��~��6WDv����?�g}��K�F����$�B�aZ7-d0��3Z�}��h��*2��=GV����
�{�%����N���&�d�Ⱦ�s�$��Z��Tƍ6��)�)֜a����Ϣ���4���̑g�����2T��}~ݤ��+�] �ʜ���c�z�͹ʈ�2�\�'e���D~��1YuB,�ߚ�D�|��N�v�������]e4���d$?�o�qt��́��b�Ҡk�w#؏�u 7A�-�$lO�*P�/4Üd�Z����C�""�oR�V2�	Jˌq��x�r�e,�׾	����0]��������>����8l���Z��~�ْg�D4Z�3�&�)؃V=���Rp �|7'M��z4�T�����C�.Q6�{���U��S��Fpkdᙏ(�U~ř��F�sL������&���s�Z�X�����F!UIÕ�(+٠����� AF?�m�;�Zõ�#n,�P:��-���&F��,����G�����^�펬�nB�����m�!L4��JW&�U�&\�W���[�q-6�C�%΢�WY9����)�~��1e#+U7�R��D�t��J�/��Y�83�s(��'��^����N��I)��xejN$�X8|4nb��[���� !��^ �,a���KO�������	+`�q"����iSHޯ$o����ks�1���nw�xe`�/�r�4vzQ��AZ�,L��69B�u[ɚ�B�5sB�ߗ�ۄ�Y�¸��>�k���8I���Z-����g����9����9�R�Ȃ�w��������58g�㝻XN�lV�N0$n� 3��De7����9f�w��GF���d�*Ju����ViY�|KY�Lm���m��[;R��!ҹ
H��_Z�;[�j�>V�(���`1���K[0��Ќ�`���yc?&�H�JZ�Ҋ�W�;�Cq?wP
�� a~8��uF��o9ܦ��3�C�k`�b�ބajoq{�K{&�t�e���Cpq�P�pZS:�,^�Ag���NyCgg6 `�f�I8���w�_k-A=4]d��Dy���p��?Q��Џ>�VQ^K����'����T3�۠�;آ�C]$� ��l�ar�>�#�z^�Ix�-aơRB*�[�ݦ�1{׻鴢
%gF���}�Ӣaf�����jg�G޹|k����� x����f}7��gL��lѤb��nN�3��,�|X����)������\�5�;;�c��t�!�:���A���kB���mВ�=O������KD���Z����҆DB�y~$b1�����`D�֩�M�6�D�fDHW xd~e�0r��Nw�"2����	��u�Z�G�85ݺ���<P��nZ	���&�j^\7gր�,R1i�tv��v�9�潡6�k
��H����q��bR��jI�V%�f|_%�.~�%WRb�Fˣ����~�$���<p9dBj'�I4�:`�]�xQ=5����=gw�4�Ka���&�MpSz0��Yx�Ij�bsOF6J��:/��d��a��/�Pך�c�Z����3B�~��P7�-�?n�bX�b�¶r٘�� 9�=梊x�
��\_�ൢ�c��Y1pկ�Ӛ|r�ȔH���i�՞:�k.E���4C,r��Z�������� AP�[�P�� �(�A�� ]~4`f1��J;f#��`zw+�?x�O?f9H�ו�S��}��c��v�R�X��B��oi�8�dj#
��W�6:l�����Zi�({��jybB�b��D�5��$�d󄸆RR�J�w����J�[��,ˍ�Y�hxd�GNdgP�sl6H�9u�mPP�U��I�Yץ&���,���C��RW9��R�|GL�(�Eܖ�D��M<���t�B'CAf�<��Fc���(�����Լ.����A'� �Y�N�J+���U���3���T<�����D�<%�r�s~�H�p��2�������:h�/���(P15T[���T��I�UiDTkq���Ԡ}[�I5�Z���F�/�o�S��U���bzA��b,���؆������r����o��<�T#�t���#��{o��W���kwh`'ɵ���#Tӈ�;�ÄO~�zD��y�o������A�%�0%S�1�e}�m��@i��W�T�ೊ.P��2Ф�{z;��?0�
�4�BZ��Ch��'n�x�Sy��U8E��Fp�p=oc��.4t�\���3�}���5P+|)��価1iD�9̚��u�+x�F���>�8��3�#�������&��T����k9a]兪,��W�5�Ǒ�c7����[o6f�W}ߪ;t���3�42w���+k�2)X�?z�1���
�-�ƨL�i>N�(:UJ����Z��):�62��j��KGM���NO�������m�N<&��\�����s��`�gH�A�i7��ցf� 	��P��h�:"|��,f���P3>Zw��u��@u'��)���%�U5�).	n/���.$�-S���M�@|��Y�*�a[���)��,8����Qi'~d�*��%���n@ϴ?g}�,���y���tLv�ۓEҸ��+)�%PL�������N��j2Xu�98\�� ܡP/]�jC��='����:)���Cr,	����cG��J��}�@���D�>z������"Ҹ�-z��R��l"s9����
�l�˃Zz��O1��]~��Gs._|�m~���#IiY<��M�o��qw�^������Ϥ�a��w���1����iC()��]�f�O���� I��SM�Cjc�[�2���dSk-���6��/󫷷�?H!m���:q3m�N�2V_A�\�UQ@�4v:���Ps�+=��S�^ϭ��2�nw�k����/Vٿ(h ȱ�ɖn����G�=3:��$[ė(��X�6D��j�VS�ga=��U�6mAZ�fRѯ,�㭅���Z�d�ڱ�-�o�p�1�4h�Pҡ
�l`��u���"}�NB�?R��S/h��x���Ƹ��������B���s��
Ǻ�Vc��M3H�}�Sn�0+�^g'�=$��&Բ����� $���-t�`�l������Ƿ�,PR�������2�LM�ޜ�p��|���-L��M*ݏ`l���_��K@/9���k���	N;@�J�	�D(������i�Lb�>�3�����&�W���ɦb� Th�δ������||��o���]���Bt��̵>�3�8��D�ӿ/"6�,��)�s{�Ω4�,��Ԡ�[E�ܟ�	^�M�&�ez�7~4�ɠ�g&���P�V�,0�D�������ը)�H��b��z2�PS})�m3�ܲ�q��y�!5�Th	�<^j� �wg�=�H�������(0��-1"�-���D���p��h�}�.l7Qa��zrDAn�g�1~7i�,L>�5��=sa˜�Jks�����z��ŬӘ��x���=��6@�ݎ��J�u蟖��5��B���:�����>D�}�����7eSa���>��Jɺ/�1ײD@��ν%�)�Iz?NS�h�?�dJ)�S�,1�:{�������ƮТ�UD�8E�Ǉ��ۈ/��Ve$9V"�e�%�a9�t�pÅs23�ꇜFH�4��Y���yD�����l7[4<�@@���K
L͐��?D�k�MAzl=�1�sb����7���\����nԫG���x�sѻY�����=KA�u� ���!��[�,NG����G����zT$����.a=k�rL��-�F��`L�I@r��'�ߘl��v�u�+�)f�,��	�N���:���hKߑ����se@,/!=A��t}���Ӡ$ƧD���������������ǔx����W0����w��Ư��	�+��T�w��{��b�p�����_��@����\�����5�{Ҫ�O~�:
[�k�7F.�y�=�1�Q���������;,�6
��1;�E'����k;�3�Gj�Z���^2�N�� 'D��?�S�g���{��j��w�ZB� 
��ηZl(�@�o�D%�r�~�k7���R�+$�&Ҥ��f�N�kM@TX�����Sd$�[tG���1הp:�� �o�/<�<���P���>�'�<7�B%!��a_�i�<�Z��>B��B&՞�����1�ymMa��_ �?��V�U232fS<LS�Z��Z��ʂ�U��.�ɧ��e��.��M�G��m�Q��q|�b*�O���~����&�F'�A��L��Wd��ƨtJ+�a���g���3���S�t�?��asFǦ$ʪF���Y4fFN��6%ڥu�?�0;ri ����V=�@��E���c��V$f"
9tx�-���w ��\����.�n���gA�8}e��D��qJ�`�c�6�|���ϙ����?�a�?��9�$��f�X{Oo PU�:1��k7&UF��k���}�B1r�_�	"�g�����)),4��l�NG��՝����q~��g�/3��j�]?��`"�>ꍓ���g�����5�)����3h<�큛��ؽ��p_(�#\��)�,FK���m��Yu���}D
�AI*{���e13@zג/�,U$���1Kk�o���g<�ٺ
N��j/�4�����c��Jk��_�ц�u�ɐ��:��u> K�<�V=���h�-3�v�o��Fja�Q|<P�{ �����^נ����"]����
.qD=��j�ߍ�N�9]�mmt\�'ԟ�
�v�q��R8���ӄ<.껐(��IUT�������N����֌��d�11�Qh]���QO��>B����EXk�N��%!HJՙ�.�:LԮ����Ŗ4�ycx� `R�˻�����	B����Uk�b�qA�7���"�k悿4F�H�iӂNs���Z��}�o*(GGx��'a�LXc*1�9L~����%�э�:���Lap��������.���h@���؊5�]�J�+c2�0�}��%�"3E3G�k	V����6x5:_��U����?u�^�ժ/j����4��3uǺF���ey�Yx$}=��1qڹ8�O��� Ж4�	�'�?�I@�����.�������	������=��:<����.�#A�X�$�N�6�Vq�p�RB<�G� �@�I]%�Z�c��mV�M�M̮��Z"�����kz�-�\oo��x�6�ӯ�P6����@��j��H����x4'a.~�RO����g�s$�J���r�+G�J�WA��q��."r*7%���ynP?BӇ���m󚱿d��:�)h�_�P]H6|�0�K�}:��,)�����D�-o���u*8�1H����K�T�r
��߈�������3���Ŗ�٥�K����I����1.NRH���nNF	s*}�g	���ٷK>��V�����~QZZk%L.Έ�=\�xn��c	Z�+�b�`Qk$���5Ѕ*|��4<#��*߬��z2�'8|��Ż�R�	����"����~���Z,a�,��Mg�xn�WL0z��Q��c�{�ޟ��IC�_��poO����l�a�k8��d8�2g��a��a*1�2=lW�� K�$-�b٫.TF��쯋�<���vG�+��fS���j�8RW�є��mE���kG�f�mv[����"�Ⱥ����pZG���:)�1�[1�5�U4�e=<�����&��9�`~��B�E�'��q�p�aq�ȷ@�&�̵���%����P�u���09ɦ�#�{/E��K\� s�St5|Ӿ��\fB�2~8�����"�����T wz��'!÷��$aSiR
=x#����� �׾�ڠ��Q�ܥ鸎�}	��U��_5�,�w��F6�����}��<H�Y��G��!�_���`�6���X�,Ix�B�h4�W=[$њ(���0]sX����:���nih�:�<��\�W�50%$�`4��]����e%n�U�v>��QmT������<�|���?������x�'�0��HB+{Ӎ$\�Y\���SL�8��	�}y��m>�]�~�{o�=���q)���P�lű��|lV#qLZY��а(~E�UË����y잗_o�s�0;k;��R�U��'�^�2�U�l����H�a�]�z����%�(V/U��$�8j5g�u���ؘ���%�x%��	�|�,��!�]@B����lS(4im!�9Fi3=<�%���"������SٷIXp���I�Y0z�D��e�K"˴.��F0���D�y������ڦ��|<I�z�UDDe:4!Ivg��[i"sM���Gg�R�Z��̠�ĵ�!�/Z�2~������M0#��,��P�w��p������!�b˿-Aj{�����x����_Um� Jh��k?���OF�D8@#hm��}'�����g0�D��S[����Cun��;U�!�	g��3g(�H�����v�1=������|�p@6�4��
B�oW��.3�
Dw��`
��F;�@���'2S�#2f�H��՞}���5�I�-�H�ů�`��mi���"�R��p��%+kC�l/�.�U�j	SX��{�r���^/�����&k~o&]���Hj�u�7�JM:X D�&�NՇ5��-��m����=b����}�k��D�����Z�mN�uL��E���'��l��C��p���MK���HX�x���8%j�;�-��ۍ��qQ����e*���o0���˿�� Lqy��͒�>y�|S=��gC!�MdL(k���h����0=U�qY 8��
�U�C��[�ԟ�(1=!�u�sn��Hc�Z�LW/2�&��NI��!Kj���[\��0�g�6��	k�>�dlm&���������W����<P� ��\*<�%;�[(j!��
\�m�!}O��{�,������:R�Ga�>�+nV�7�FX���z����������ٜ�/���#C���u$k4^;�o�"�@���u {ࣨl��9�1B?ɢ$|Evv���x�̦�����0HbB�붔��J$�?�}!M��C8�X����D���5�+�IA�;�js.A�����	(܎�"����j�?i]���|3M��b"���dl�7ӛ��Х#�����Ou��t��	��+���z�5����a�#�X>��;E�_��g��&�>�ȏC�7%�3#����&D��C������-o���"(����"�GoBp$����b�?l��B��������؈i
,�YO���#%Jؓ�9�I�����h��hP��'��H��}�gq2XY���T5s��X�� ~B�n �T�_�%A '��<iew;�Q�!��.�����o��RDXk�����-~lG���P1{�!�Kݸ��:��l{���� Q�p���M��� �M;�8ޘ��Q5��9�:ad��%7u
�-�#����L�G�q[��ݯK�����b�6.���q7χ��eX�dz���qS����A|�%l2���6(���X���
P	�]�8A��~x5���*�c���%㲛J*ʪ�!x Drn/;��T��t���l���k*���ˑj_����g�b��������Q/7���I�̰C<����r��r&o�`���e�HVc�����cx;��V3�c���qQ7�6(t�M:�)��;�F��[�W�@h��l��X�eK�52���[�A�_�Gt��z�@�#�&���6��n�>��j�����j���]D��|��"��Y\�tЗ�(QGI��S`��L�5�N�y�	*x�O�-�s�Vx��Q��R��~��|�����W�`�a�*�qf
��Iյ�����ltt�α�0>����RBZ��ȓ���a5��^�h�Ŕ�$B�w�� ���Χ�h\��|�>o�3�k��ʭ�Sҹ�g��r�yd�} ���U��A��wi])0Bk��а\φ3ꭕɓ����\�gT�����.��/$�,t���*Uը/{��/�;���S!���M]�6�娢ɲl����D,/�ހL���&�HU�d��샂�I{j�2�;|-r\��j���'�0���Q?�Q]� �&Q��H	�F�D��%�Q]�ReM����α�%��L�l/���CcT�πkt�~��nv��.^*sH�]%,vs�+��E��6x*�5��/�}YV�H�P�S��_Tʬ�2�np�GU�M��#����JM�@wW0�v�Z�m=z�+ SR8�-��'�Az?��`�"�@l�`�y�lȻ	�[�)�[g���Z�As#b|�r�AӼ���<�ܠ��]��`jk��xB�t�c< �ϓ��<�SKC����q0Q��|q;�7�� X���J����v#7�Y�*��[d�r�B�jS|�K���wx�):�t�X=i�Y��Z����f��~�ϩ�^"~�E�0+-9\�`@U���5��
��=&S�������3Z�5����N|1}��9w�P}e���(��������V,5���O,���K���<~�gR���ov�S����D�I�]L,@N?�I���dW�� =Gt��\]ի�-�AQ4��^�I��E�$o]W3�ل�{�Ď!;e�<Λ���v�J�+KXǏ��Oe�N�"$�(�/&b��R>;������)�>�\��v�8|���I����㦡�xi�5�L��M�9<���l���\�GKt�a�vW�?�ML�\Ƞ���JeM���y�G���>��͂C�FH-I��p�"v�@uD��yo��!ty���'�G����>ù��u�$�\ފcG^.�S��b-^�M���D��� �l��bT�X�������Jl%в|�8�}�i���{�;�ڗ�ןm���@0��Ř�1�����Fz&�6��I'��ᘴo��Ķ鸘���IR��3��\w�Tg���0��$�ⰱ��&�����~�U�m��r��͔А��p���F�ǩX���y?��?� ��&E��3�qZ��~��z��I(��N�5U�I��5��� M���k����v{�u㔞3�J(ہ/^��n�.2|9��b�!t��>w+{�!������GK�?���č����*��,{����BَƠّ(�@���iH��nuA�l� ����%f<(s�����)�~6��/;��|�v�{@���`�����[*�ClRflR#mfF)�{��H������<�
j��ew?�`�xdɿ�Z �d��H�D@�b{�cRP��B�9�f�]2����Z7��k���gf@{8�7=xw�.Χ�y��-�c����$9�l����|ie.7���F�l6\�W��[zH��$�&����z�N���=� �G;A��p���Bx�e��J|��J�+��e�ջ,�
���ݦ����n�%�b����������A[����bt���r���5��[�e�*'�Ё�P8��Kq�1zu���ul�X��@j��J�E��a�&��I�l䧤��k�N`vVA�A���	�$���f%,;���Mf-�z�x�/�$6�YǤ�Cؾ�3������p��s���`oL�n���&�q|�k��(<WR���J  Ǿ��eͷB�^�Ҩ�=��E��Lf ������H&���MM�8�!<�b1m�q�¡%zɸ@��p�?ֈב+`26�;�+�Q��F���c3_���B��.a>-�󢐆�.�ʓ�{�"wզ��#�DC=q��4Ƕv�/$�+� �8 +��N-���l��^���8�\	%;�"׏�N�G@c�����D��teڄC��݂�I�U2%��o;{�c[/R���䚻v�uڧ�~o+ۘ��7���$��᪫��ԵQ��僽D�y�~��Q�~U=��e�I\�Z�*F�^M�?zQe�.N�OV�_��N�_���Z"�����G��@��J�M��#Z��S�6��32��w>���Э	��Rq_�X#* 1��}+��� "���3�S/lF�f��Y����&������L��Pm��YZ���743\�^o�,穀�*�x�����>w�?w-]��:*Į�O
(��>[M�CZd��C��6�!os���2��q�']銮�`C'υo����f+"�Sj>�$*��%�69%�i��jm��A�n�J1yo�����-��lQN?Q��!�(4.T�7~�(�%kl���jc| Ld
Lv����,Ji�(��D=}��"}؆���_���)�I��_1-G��0l�y�O��׷`Y��& W�z �?���C�]"Gy �>Y����GouC�S��i��?�֗v����6!�|X��V��3�\j������M��26Ż����&�X�V4ΞBEP7��S��"���E�8�f��ѻq�����B79qT`���hwUm]�A�~�Y�;�d��p�
ͫ�V�����������`C�d%Yt�\���|�|�����H;���v�y����+B��� �_
�,�`:W&�}C��{���[��a�h�_+���Fp�-Ѱ۟H�*^��C�h<*��"�#�i�_�{�e�r|��;����L"�����D��F�a�1�H2b�=�[/|�Oޣ�Eq6��K3|Z�9��4��@d�y�*`2�Z��G���غ� ����:z���k!G���vfQ:72��NEͱT �X�ۖ��ķu9¯����+���d���kw�)��a��*�з�����'�8�Q��;�B��{�<&��j)�z��~������*5v�:�9���N���BҴ
?�Ie���O=^'��[ �'��RA�:�̆j�L(��P���e�C���r-����8p=�)48�Բ�9���Z�Wl�����s��>H�( ���t�^���G�DX�<s<�*���Sb�ۏ�3�#��JV�!r�#�M��*؝�*�V��z>��0��ǰ�f゛8TT9�i=F"�* ��w�E�L�A�=��<��kI'�	o�"hp9hz�L{Li����A!�( "�8L0���5����$�y�[5�el4	��J]�|�>C� �$gV�9!�
c��r�<��&�Jf[C�Y*�t�oӚ��"��&ρ� �kE��,��z��ǝ�.7�bv4=skYpF� ^���*���o�q�ם�ϒ�Qf�<=!�Fhx�)/C7����>-��вvy�e����<@��1Q8�V��L�Q�]��}^>��-�}w���s����3���5�R����$����D�z��6_�LĈ�P}(M��纨`�>��Yk�V��WlIͼ=�ˬ�=O�d?^M֘V��B*/����@VУu����LCF)*�>�k�v
�H���a3�G�a|��L[SD�4��w��u+�s�.Kuz����2\�
�Y�S�Z��c�~M����'ȿSQv���bD�D�ϭ��A0_GB��e�&�2( W�ݠ�"$��Up���&�Y��F��1%[t|%��/m�ev�/Y��[9L��ݪ�-�n��܂:����xT�)��� l �,@��hS��u0�>ݡ?W�?a��Y��f'�M6}(ۂ��b���4�Xte�S�%�c xN���.���=V����7�Q��|��4��a���^�LZg2w�4��}�ḃ1����q�����i�g��ֵ�Gv<������t$T�2�2�:H�?c�h(C��~GE���}�}��b�r���&[7H���Q)��o��j4�Hj���n$��J�bl��rP�K*)d���.��2)���cDU�R���?���fna]�� 4��Dt�08�4�x����x�w����)x��0-��)w��}r��&��[r�`����k�Ir'�}�'��O���IC��c����¤�Sx��M;"t���f`+�i������)�/���,��d�i��RU��վ��k��?������T��u�BKT�$���~�A$�����Ō#eo�Gp��k_1Pc;{�ӕ\P�Dy`N�lQ���wH�=�N5����% �{W�\-�vk?��XN/4���m+ӭ� �U)�
��Xwl?�Qx	z�Ŭ�N֡b�t�%�Z�GZB�m�
d8����6��?�2���ێw9?$��܍�y����	�����	�ny��k�@^1�M��F�|�cr(����8(HC7���耭l�8g��L�=^�\�-jI�R�
7�����x���QI�_���%]�5����ƒ�.#�R �v~1��v�{���8�mug�g~��T�FUm>'���8�Ws�'{$�y��A�J#���K��=äf��@�q�r|�O��a����nGL9I����Uo������W�X�#���~T�E�t�ٌ{v\��f*8�uU	Ȇr�/b�����a� rv�a?��p��P�I`XJT����D�V�\�zȲ��8��ؼ�j�u�7�e�;��/R˥ձ��n����	<v!�m!/�	%�E:���`8�[�]����m�'�>��܈�|�l�MӍ;���~�Z�%�c)�-��_Ys�x(� ��s�-K�d���7�����3U�Y�ݣ*�,ݺ2�E7Y|�$i	sZ,&L�\^�ј˺إ⿗O�H�`Ԭ+��t��(���+0�l�q :E26>bּ�Q&)J����ۑ�{F�h�gi�6�����Gvl	���a'�U�zF��$���F�	�oq0���*�Iϫ����u �k�X�rIth	���J�-?��]�֛��͖�
c���{���4�h]Z*�Ͳ�9�/��Y�6��V�ƙO7$��b�V����B��ă	���E>�����ZN���t������¤"q����h��2�	8퓫���ۤ��s�7�����X���@��N7�Ix��>���*�AVaP��V��װr���A���?Ю�K"B�Ҙ�6,���r���ʝ&Mu�����uΐ�����)!�6��_^6�gM��c7������v)��H��N@��۫??�ak@�!	'V�e���3�ݯ�c0�O�n	Nu�$W"�t��l��.T�,jJ���\�T��~�}��̋bm?%�q���\��j���&.Y�-�TZ��#��8�7��h5�K(�ꢽ���x'�ޖ�E�uй�}-UUled�\�7�"��p��`{#N��
�߀:��>�F�[����K�����|�21�3����C�I?&_��B��3�������*�hF��Q�HA������:]8S���pZ�^I���En�3��w�KdԘ��M�4�k}���B�PL����%�Fƹ��8�!�u�	�n�B�����H�'YtT/� �e~]9'S[^��qSGPj���2�m��Z�)�R��w�{���JFz�9�׮��T��6�@s�7�C*n����7��4x��n?0Þ�9r⒗�ا}���S��A(��>n��pa���PEA�ή,hrg�����[�u�TfnP���Ԫ������]��?#_F�c?.��f슻�M������!�����M��1&>( �;x�j۬��-BRa�+ ���(AqIo3=�m��G�)$�j���qh)~˱ũ���?��+N�kn�#�G��v���a�uH�^Z���1���#W�����e]����+���1DN�wؑϭ�����΂
���}3v�,X�)�"]��tD<~�UC<;���<�ދ�ڙ��rf��l� ���_؏L�	$��ؼ�F�jv�@�����x�du{-��5�<�Fm�@�N�X���BCM�@��S� ~)������x��D��*#aI-�W��"�rdry�f���1`:��`u>O"���F}���`��ɴ#�$���\jL�
�<>
�䝒���`jDCzf_�)_��*�T�������/x@�n�?D�3��{ �P�(C��f�m|�,vq�~�q�S��;����z�jB���3fL�	�99��G��* $l	��
o`mA�K��[�/��f���tݾ��)ɜ�= `IB�O4��+��1�{�?0p��]$So��'��,I�� ��}��rأ!i/�Y]��.�'6�kŚK��6���n�U��DN�}��S� Q�;��RE�)���[�>G("����'��m�:�O	���5}��\z6�R�knՇF4#ݢ���)�O��+р�vc��ٯ��E�qf@�A���������8�ر��ֿ�L3I���i7
)E��M�8����
�	x�
d�vG�!��LV��� �M	��OBV櫌�h�a�VY�*9�#�Ø|۷}�LA���.����%c��sV��]x�R|0� �a�Oz���"L�=p�س�榞�����]09��7F+�Dϋ��$��$��:,��\������>��p�Cz�\Y��t�a�Y��<���{O� �{n�䟍��ҳF���ˍ$BVlD�Z^T��;'��F��,_��\��N�ݞ���Ө������D�ﳅ@�\տ jwM�ֻ !;Nb02Q�(8���P�����K�^��v�&��꓏��F�4�����⹒�D�;(R.�&������m���/�������vd�^��"Y6������Gۙ�C�%(D)���;�
����~y��������A�(6� U��ZN�xd�����w+;A�NQM�C�/���\��b/>��tQ-�d�����q�:=E	w,ihf���� r�%�N�Z27w�I����Wh���x�Y�;
J��e�%�r�3��&S�BF%�%d=5�