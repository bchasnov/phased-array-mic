��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\����q�?��e�I8�b�Ǽ$��"����ׯ1�V0���DO�B�N�^7��F82�u�	��[Y�l�`Q�Y�d�g��v�+���Jц���6�j�j�$�j��QJ� }��\I����-��H2���U����^�Y�	�N8uH��E�����w�^O"B<�(�4�D��eH���yg8f��;\�8��a�&>��t�܆�؊�U���k'P�O��$�ܬ����^{<
�3���;F=�[�4^���0gB�������lXL ��A����ҵ[V�xg�/�߷�����x��H��4�~x5k28�����3u2F�8�x�]���5��(��O�1����E��$GjB���<(z�C<4q��������j�XS���s�e�̊�ϟ�-�'��+ѽ,�.�NC���PB�"�0�bj���v]�h��Q��:��I��)��0� P�љ&�w���C�)?��q�G/9F���H�7R���ju���1ǥ?�����U�(�N�P�=�ۡ^�_�P&�i	�x�g��tj� =�b��C	�Ԙ䚇��CCj������ޫ��=/$)��GV��?Z~���n?1�Դk)|�� ���k���N'����0����ߓ?��/r���;�Q�-J;�k�f�s�*5i(m����z^�t�W�"uя���������&ZX�*z٬���絘/�e�;��b~�eZO�`6������ذ	YKr����T��[e���2B �E�%��.0�1M���W�*��iٜJ���b��s�qQ����f���G����w����+����tH�Âf��a��5�n,�#<޴�K�~sriSx�<l���G�������&&�B//�-{}�<0Ԑ��jr��ᘁ�]�6w�f�}�j��A�� ۪�K�n�����ܨ�	_m��$���o\4��g�G�t��}\\K �_R(�S�3=I�l��� �fA����Z��R�����_,��Ꮪ[.��@�P�"˭yc��Y��WyX��Y2������;��!���I���SZc�n��3Q�����0�ŉ�İ�aA_�Ö���U�s������E�ە��ps����
W�C 0�Ei�_���-A�2l5{N�7O��b>Z�R(��
rs��Kյ�g"R�"�!6.v�(?̻��UcO��{��Љ�.�����~�`v������4⏇�j�?�78�YD�t�|Պ��Ҵ�=���LR> w'G�#����-�p�-�(�i���=x�}���+�@�IÖy�)Z�+:|��S!�T��Z%K�e/<-�nVr��W�taS4.��n}X�����7�W
�d`q��Γ����3&�6bHƕ*���P#��di�9K��������8L*�hQ�ʣ�8���S=29��!��Pݪ>��+�Ʌ1���0څaǑ�[�&~k�y>�>��C����IO�a|b�m��y�'���sJ̿�,���ą��#�B��0��?��[�6.����m�Y��	.��ڭ�hܯB���������v3� �=&G�{���u��;c(uƨ��KA@ z)�b��Ͷ���~��N5<��O�}8�Kɤ|N]S����߃�3�EHQ+�Ϯ���Ԗ���d?���Z�UkZqt�����{Af1��=��B��w�������5�-�+y�g��E^Q��&Q�,B������'F�<Ū
J�	�	m7-�v��31X��Ds�C:���5���4^�)�S�eb/�+ϔ��C	.�~b��]�� ��h�&*%pҞ��}��iu{���ȷs���*'*�8� !ې�?K_@�O�jEg�����a��F�D��.�3��j�B�R���<ô�>,9:a{��}�n�Kz�[�A�����.o�������XB����s�ԥٕl���RA��$�L͞�P�6V�-҄dN��(C˶q9v��H�Xl�8&19�v�������L�Nt^f�����������y�B�&�ګ��F��2,��v��Q7O�%�d�&��b�ˬK���'�_�j�����pU���;�$�5� %��7ٱخ�SYDY�\��>~�1>���b�ז�n�K��m����qH���@(������:ka��~r0�t��v�$q���Zc�NNl��J����]�LkZ�X�$.�R����FM	^�������W1M�Cy�#�:{�wb[;�挥r�h-�s���z�=���hs���v7_�k�p=�
R���{�M�uT�_�ٌ�6g�2�����f���EfC�6Ԃ�Oׁ@��RK#�K����~�f�[�z�.��n`xi�O�޲D��(C��a$�zL�1��Rc_;Ɯ�g��#��(Q�?��J��u�G&��Taa�/��>�e7=�75��8�}%,�$�_n�:"�����[��/H1ާ�`P�U��`uц�d��X�T��|w���++Q�ܺ�޿�!�����u�~���\�H����&�^��GN���8jbʇY
��޹�ރ	8Н7ٖ�ME�;��si���nTzHij��62Ѝ!�^9��UIق����tl��)���7$���H<߉��]�;{��ݧ5�oސ'&��p+8����_K��u���@�k���z^
I� �$����W� ��p掠�:R��wW����B66	�!�{��%�:؛�g������`�m#�D h�]јt��dMCtBY��,�zy��v���_Ar���J)8..���<�`��:!/ߺ�/90�)䆩HpH�y��ܖ���r��[ߤ�k��3!`Ȑ��L��'�v�N��E7�*B�ȿ��Ŵ�j�9�+> �3�6��`�on��H��;[�2���{���y�+ז<�����OA)F��������5�,F����Iv	�&Y�C^�$�MqB���3ޝ2
��{��7�OmM������ǳ�"������QPD�s�������{L��T��1��W��oOŠCF�u۠�� ���S��(�'We����$�):tR�G��l��E���+ݍ8��I�a���p��h�5LX���v��/�z�����ى��������N0�>���I$�@�C�&0��fq�� '{r�S��D4OHx�����R0I��~�`]E�nP�@�еl�BY�aH�h~1{���is�b�����ښa�p��Y󲊧���Y�P�a���O�h|O,K�;"�����{v9�+� AgT��bb�}��MYx����e����I���TK�n�I��y!�)�z�u.5.JK{?���!:r�П1��IU���%��҅{��.�Í髨Bjl���X�5��dTY�8~^y 0҃��7yf< �U��u�8���*H��٨B�1}�/gU��'\[bzm׆�A��vƽ����8�q�.0��x��aAy��| ۆ�SPoP���J*���肀����F�h�U��܌�h%�mv�����~c�m3�?���U�%��+�?�c0��AzL����%���ewf��|�a\���V3�4�\{���:A�����O�P��Ԙ���%;����l�Ofo��-)>�sp��{��\���$.R@�<ڨ����mZ��GV�vP6鐁����(3�-�	x��]r���TC�	3���ո�SS~L���/EB���r���x��=�(�ۖ�p��u�W�X��,P(�\RHd
w=9E�:�C��Ԫ�BH��m���f�%v�m���ao�0]D��4����wR�\�tR��S?v9M_=9��*~Y�sќ��d�L߷�1������1����ˊ�ĵF�qg��ߤD!��s�γ�7�/����!��m��Nɚ��bY1}�.��[�#�k���J⽓ޑ����%���{�F�XM����9�4p�I[/�J2ɱu.���F�fo���}���P�@V�%���xq�
4<-7ux�-0��5�� ������u�'vTS� �4P�N���I�,��D͖�<>�0�ђ�n��ύ�����0o1VR-�و��n%&���A�g�N߹.�N�2��~�J6;�����
�k�+�E��N���u�"�ǸS�poIga�YK��?���/mW��P,1B`?>Q�2(���I4y�Xd�r+�-q�^�g���iXTl�������|�r��f݅�p���neT�ÞdB_�����jȊL��V�7���ϯ���a�i�Fs���x��j�âq��7�¿\ߏy}	o~�FyJN��9q�n���{�:����bHu��N���$E6�W�(l�ܚp�<Wk�L�[�f]k��KbxGߵ��y��D�!4��+�+Sk��k�!�*W�<�Ur�Z��Q[�n��@\��x�	��<ǫp)5.����2<7�������Hf�9ĭ�%l��J�y	ϵ~�O�����NC�u�Ӵ4WR��::��u�~��~z0�?�\Y_c�'+0؏�#�2�`Q�_��_�џ�*�ޘE��*�"�]T���!T�u���<byiYܷ��(�d�6����	m��r���YyC�	2l��XߣǓ��{CB�4�'�ȇ��3w�?Y�XǄz�"�;�bO~�D~G� z)��A�b�:��Gr!���X�x��[ӯ�7��H��j .�������c�GO��]<~�}�K�	p�����x�N���nE<��E�p��	�Į'��*��Ԝ\q�q.��zx3S�	�N(fe���1n���_8`qv���#�/I����$X1�g�I�dh�u&�]9W��!u𱀗Z{�B�]�+[k��s�	R� ��/���jq�����-��� � �0ł�ԨŁ<f��[{�O��a�R��>��a�J�4�:X�n��VC��I%��ê��et�+�ޔ{���C���\/�] �x�k��ʊ�<���}n1V�#f��:M���1˄�X�~�����G�PI^nڄI�Q��,��-h|�,�'!EI�Enң�T�=�x/��J���L�Yh�x�lm|�2	��;�c�d�Ow1vB��k'|вh'w�=��q͜�t�<Ú���[M�&��jB�/�G+��B�4�1V�v�W��!8_�{��&��FY{b݌���*��R 4�`-��aYV'-D����_I��ĥl �w�ag�d�T6��Խ�Yx�v��s�fT�i ����H���)�H��������/�_����gWOG��S�Q��M5�%#��>�~q��U�T"�g�,���8,�S�YF����F%����uLH;�N�a?o��F��a�V(��K��t������Rn͉���k˫��-o����w�3uY�2ֺ�?���}�m	�"�)%�ȷ0Ƽ���c��>pK4˱xP�녞U,�/z,s�#+�F���]r��^8��\SI�7_z:�#Kp��;ȺZ�5e�TG�:Iڮ��e>��
3��$��6:�9j�4���K�%K���PǦQ��0�Ҫ��U@�R��?⳦�����5�%��_�/M؀��f��5WM1�/{NکĖ�ھu�=Yl�Z?��*�č�#r�?7=�W�TUN�<­�W6���G��M���NB���7�tl��&��V.�kuP�kK}�00�YF����D�	��xb+A�yq�]rLZ�8LK�?��Ђ%��y��Ww��2+C�������x�p�(��Bg��M4@�����Af2�-�����
�Q��>�$Q���
`&'g�̙]���9�l�=�q�Q{)�y�B��=Z/Z���CG��YLˬ(�V��/���tq9���[�fz�b�Ne�`�ڥ��e���KR:��M���쉟�P�w��8/��d�Oy���f,�=���=e.�!	��c�B�$���/5	]�ڀ��/��ƈ��(Tf7a��!T��9&���	f����S��\�U�q��$5��Wwm!4�X2<��h���$Z�Og B�����n\�%�l�a�7t҈[f�6���b�����2���C� $}�M��%��J����; ��!t&�H1ɮ���k"�j���5(�t��U6�~|�v�ɏVx:���s_�Z#��0ׄD-׉e n����y��v����A�/91�6�Ѯ1)���&3��[��X��H�,6nd��mQeCع��T '$V�G4�H�Q��<���}�@�ܸ˰�����{8�(�P�܃�,<. �$ף���@S�ʟUi�#�J�S����cB% �Ԅ�5$�u����v9���u�̟�B��w���k=()O�M���I���[|��S;��њ�zoMHO���@���b�2���_�:'!I�@h�t�'�^�SQ�´��@�?Q���TJ��r!-��M3�ux������}R���O�&c&�=�:{|�[�:�W3N�x�..��.�Oz���p����n�U�[2��g�	8S��W{�+��r���l%6~W��K�]��IR��R�$�T���ldXש����g��f��TgP�JD���P�E��x	�E���Es�H)o3�ԯmE)[��W�o�U���Q"�]�uf%D�_�ݩ$���(�� ߑ��V��ю���W�K�q$������
�ԙ�w���|`)OukԴ�
ُ����ӂ![W��oc\x�LGE�5r~����r�j��9j��g���[�h��(^��D�V�!�p�T#cD�nr��Pp�c����F��k�h
T�n��K��~�p�'���S\�z|�:~T,�j�y�`�>�$ye��O7fp
�8�=�w��+��չ%A���9(����I�*.{��ϑ�|Uq2-�T&��FN��2/���C N��񲘛���]�"S�e3�B���y���IǛe�е�ѥ2Ïb��0Y��\0����7��_ڀ���B6ژ~�<*$N>���E�t�r@�GC���M��f��|n{$�kk�!�.U�l�t1����p��z,�	�J�8M�t܍�
���r���Hz��{\�+�uDê�؊3�2�f5�U���~�'_0��7�0 ���R���9�N.@)�V{���{E��W���9���6�Ýl���X��#��-$1Y^��ɵ��AW�mq�������
��>�Į�7�$4x5�s���>%Z 8�&p��f�§�P����-g���o_���Z�c�w꯹I��x������~Z��-�]N����#T����a���$��؎CO�ȵ�W��+�o��R��nq�oyy
��w�P-����*8�f��)V}-Ä́�At����{�7`=7U�F�K�Q��?P;�9����f��S�fi)�T��Yz��o�߮q踖	�G�u�,_�-��� G&���������������%bǭ���-��h>^��x�1��#���u���_k����g�l�@ڞ�f���4�,�f���'X�Z� �Q���Z��&��4�G�9/�+��mC��)�#l��>�\���J}��KA�#ר]Gb孇|Y���u�a�����j����QO?d���ΣfYM���ˡ��2�����8�H�8܆;�D{R���2`�3��6��g�R�L�O5o�b�Fq(�b�K֦rwf߳�uZ!f_[C�FP�%@�"G%P�hJ�1WgJlT��d�̙�X����	/e~m��9���1-�Y�E&a�k������H0$����w��+�v��l7~]����{�cv�j�l����Y� ��I����OD�8�RU)��Sm\����&���>�g���xԩ`�WO1�z�ѽ��������(�+~vyn��\��6�|Py��sn}!��������"_|�X�5��cݴ������>�W%�M/[�5�Ut2��� Z��s�]I�!{��iq*�� �*f����[�A�z�������?h�Y���+h>�_ΊU�$�]b�Mz���6�\|��Ov�%���O;=ajFBCss��X:�8U�	����=��k�æ���0���O���dL9����3�.�~Bt�����ڣq��ݢ�6�䭑[�V!X�x�5W���΁3��E��}s�}�N�0�t|�;#%2�� 'H"-S�,j�V�L>˨�\�ۚ|�Lpޜ�{�Ͼ��}��xvtB� ��OI8�?&�:2��7
�?Ŧ(v��2�����~�c�teű�7�u���d�$��ɤ[����M%:���
B%��s52JF^Ǣ��<��gP4��ץx���o���'��D�!����Q�ٮ���H]�]>�� 1Z�V\v��5���t�&�B�a�N�+��OmK�i��#I�&�Q�ۿ=�{Cz�ʢ��$z�eYF~`���{��(��P�yi����̄4��(y3^K����F�<z�6BB>�<��.vƟ��r������%��k��	/T��nl*�؏!�-f�"�I?#Te� G.�y�3���?����TLc ܵ7�zScP8�Ƶ=,���-G��qʎ��A����f��u�Z�����0�����i�hN�9��/�Z�v�%%/Uv��Rg�ŕ�[T���c��h�Zb4̟�������>��9�9H��HCX�<����ے���������\p@��R�<bmM��ߏ`ݐv����/(Y*TT���FHQ�_�g�:iy)}}S����.�:��@3�OS�@�{ႛ{wP��{���"�k�<Րr�9���M�(k�)/	r�7�|���,e�q
��O�Y�T���\jf����{�jG$'"�U�-�'���uڞ�);Q4aaH����їr�(0�툝>F���8�&"�?6��_�};H���>\:�ޏ��W�Faְ��ؗOZ zሼ�R��y��[�宔�.C�{�6�S_�Ot�=z����*-�l#�tﳡ�*��J��¶h3���L� ���'�d� ���(�m�ni���T! �w�{�Yx07����\����ڠ~�Zb_�Ն�al�T$��1��(N�u�5T�g���=|��}C*�M��O�Ȅ:pC�[�~z<d�	#WY�����'�L Q�����P�Lr�/n�f���p 'o76�%�a��x�������'[�����s�xEe�h�bm�(+6��I��`����ԧ�)�.Y��"��b4?0Tz �N�o~RS��g-4��WGPS�U�i]��N�E��9�4����mp)�� �LW�1��O[q��:��`���?RX��2p۔� �A�c�!��#'V4�f�=�7�	츨PUP?[���9�S9�j˴�mQڨшQڒ'�v�]U@�Tؒ,�k���_Q2����xJ~@ՙ���j ��~w�p�x+I/�ub��C�\�l�\d�������F�,b.;�TS%�/���[�-/����Zfuh�ܫLUPb�r��,���5�"H��1��-����Q��*�O��ǂ��w��f>�����1��n[�h.S+�	][W���:���Mr��4.��fg���\�{�G����Û�d^�w#<r���,�"+�\�O�����X�(k|�o��L)�C�=+����n��6�X�l��i�3Bq,ߜ�Ħ�
���2B� /=RՆ�s�z�g�4�:�ؖf$-��{;N���8����1��gI+��s1#5:��E�z���$�F�ct���>�Na�����"X|��m���F�7���l�]��e�~d�Z�y*��̛�)��~�!F�������.n��3�@V�]��4��b��B%�c�]S�h�����B�� �F���.*���]�ĮS��@�֔�T�+M�a`Jp4�Hi�*�)F���_Z����>5�Tg�&��T��oGt�
g�r��x��5̿�:��U��	���"5Wq��&��4��������U�����c�+�6��\{D!�<nk�N9L�{�����ķM�Ʒ���ţE`�,��We�q�-�iC�ʛ����(Ņ�B�R�A����lQ���Y%q�b��w��C�"����H}����H��q�!W���~xLzT �FxDC*��i���>�k�6�i}����:1z�$��"���b�Tu(�K '�få�bdȻ(�<�9!�=,���^�lu���dL�]�ŲG�/ dlP����/��i8����ŔE�+kA8jv�KoB���Y �r��{�ų�$�$R<0o��]lQ�V�T�U(	Oz�#H�K�Ʀ�js�+���]a�Fd�㍞�.�}��,�4C���'X q+螂ᦧl?S;p=�➁��e�-�d�|���!O2Mw���?C��S�b�T�=~�sv�O�b�`�C5�{��\3��_�)w���2�f�>ߩ׸ݢ){��,C���P<�R�e�x>��j�u_�ED4+�KQ|�Z������n��`IL�F��CS�I}B�5,X�񒪎�Ϡ�=�'>�4�
4C�	�6�1�}%hx�����q#�s�2tŋ�:V���_z�A{��B4{�on��WeH��]g0�0Q��[%�`��϶o�O}��d���K?nz.��)߄�*��0�/�l4ΈӣTd^��+��9@͆�´�ķ$G!�J�Ͻ�ԛ��J"���z��;�r�}摮�a
�T�� o�R�8���h&$��۰E��߸8���"��{�{袙�Ȩ�L���&�!����t��B�gqOO4�j����vX���af8X��� Ew�L��v�E����QZ�?��'
� ���ʲXygK�-�IM����R0;O7���9�+h,�1w���`�4O�]w=N�Q+a�^�ڰ����C���F=�#���C=2mH�̚"�z$g��f�3�&B�Wf"����A�������B��x9g��|_�̠ �a���)����h�����E�+�ߥ4td��)�cr���5B�@��O�MD�fL�m}j�`��l�~����z[�4nM�'�c������&~LO
��F��z¹y!ԣk�O�=������n��L��gV�D4B�TY[=����`�6b�bX懶׮�,mX����`.����<�L�D�H�9�G>�U��س{�;y�M:#�N8��1�;����W�#^x�����ȔD~*&��0ǋ���&kW�ƃ,7$��&��HU�M���H*y�??��* �pN4�W���u��10��w�H�����*H�Z�@��9$TsªFȔ���q#��ǳ��s(��Q���~�;:�)��k�r��`�]a��~7:��8�ߖ�B����V����]�:N��4!{g���z��cڈ�[3�G�Y�+�������S��3uN�:�~�-�V��7{���������r�y���u��cIͺ]yTT�L.y�k��C������`|���l�ii�t����SW竅-7�_��� �SI�+ע��0q�jo]�;$juJ��]�6<hX$��Aj� W�S�K��u{�E���Fɒ��~3���}��m<�]�ǩO�%9iS�%i;����阢o�S�;KJ*��.��Qi+� 8{�=���$
*Ӌ��nr�]�t�6���z�s+b�!���W�wv�y��i�����k�L�Iۢ/;Ŧ���62N8O��.n���Rg�J��L{6	�F6ٸ�։�m+�����p[����]P�|cc���R%?.�}���\��vkӕ��[G�9�C}a38[h����/ܲ��B������[ngG��Ay��#�zK�䭮�孂�n��������
\��1l�{t�ݝ.b�[<[�u�%�u~%
eplʹ.����C��a���95ӣC�-��
zK���E���31/���"�w'Sn���[g۰ؕB�zR~�/M�8݀�v�-���y�C@Ym��)����J6�]cO���� ��<������QAML��f��56�9Zǘ�|6Kz�Eɘq'��8�n�F"���:k���"�y�g���a�sj�#�RU�}&�ˣL�[GE㊖J{h�G���xn��@�ȳ#fm��b5����Z����L�az1�k����D�U�/�53��N�>����P����V@�E;݌I8-8���̊�R����j�\����ٻ��tK��s�g�L5JCj��L���)�\n��QCfE)*�$�m����1HEQq��By�܂������X�N��at&Un'�����L��Jg����I���#��	z��<���ILHJ$@A�Lu�c�Nk�̓�žA7�@��6-�:�D@��ù��^o�.��N�%��=��-1��0Q���	:c,
#M�:<�
O����`1���2�>>�`a���ʔ&�F����_�V! �z�+�"bn��abo�Mb� �LeP���>���,�o�\D�]b�A� UBS�w�~���f@M0�����Y��DRd�(w?�L��S5�����M�������Mf&��\��}��ng�"����j���+5�:  �8'����Z�%<+,����p1e��h��cq&�T)<����~�zj�"�ސM������vY��g���L��_��
�i��%jA�Q�5#+��x0u�L�$����%L����w�mA.-G���E3
��8����I��������:�u�(
�����h�_��=ݰ$����}�|/�qL\�����{'�p��3��?�$=��%��m�u��۰��R��}�����^�k��9!�ȨI��˿�y�v�W;�ll�����T\�jՊ(��z߆��f�N%��`�8� ^O�ԁ��q�S{�\�	4���%�2Y�	T�����S�L�D��I�M�V�ʺ��ؚ!E�G��R�+ vo�^��Z݋�>OKu��n]�/M��i}f'��|.?dӣT+R݆�}�g��;��B-v��������M�>a���VM�Y���H��^R��(��aT-~��ind�-�|SO����O�4PY����� �T�#��G��NR3! �(��ؐk�4{K��錖L`�՚E�j���<aQ��R��x4D6��X^ɨ���Ŧϭ���HA�d.��ڱ��+�h㓛'_�L�{�8��+&~��/8)���)fxd>��w�K�3�4�W����L��qaQ����L�4�_����3��t]5͑o�����\Yμb�Y��;��}�J^s��(�qN���1�G�^g�xqݩxQ���&�떩��BO�NP7�c���R@�):��Js�[1���(Lq������4NdBZ=��d;A^���Aq���x��x�g2��!��*n�̇H�K�3��tMEwh��tǔGҍ���V���ƺgV,~o
�_��W���f��|�|U��deS�no&���a���R$�x�9o�#l�4"���\���&]D�Xv�d
{�}�^��+�32$����.�Xm�9� ���W`���F묐��6��CV@�y5]�,8�l�c;�A��`;�m��/s#܅�.����_��R��2qg���~vP( �~�v�L-�m"l,��B�������it��؇Nr�n���V��~.#�:p�~x�ު4Q���_5��Y��.���,�9fޙo#
�O���������eÒq�|�q3�0_/�sl�A���Ka�K߭+�d&8��b���H?��B6Տ`L��[^��)ޖ�M	��U��Ro�5��z�=Č=�v��� �av]DQ?����al���9Ѩ�{YF��{�[�(��=���pZϤD�zv��fٲF<���z��i	dW̋��&�V��,j������\/�Co�������P/��;�l��B�.t�B�~�_Ѐ񶫾�����W��(���pv��]"w�O�'�?C"�(V��������]�G�ui�WFz��>�Ǔ�>޷Rz�)�6ʪ~>���8��\}�O���d�|}"�Oq>N�[���S�SL|��.4���y�f�:�U��8m�a.�ʲ^x{i7Fi"�V�ًk����5��n:����5߷�(}~ew7sdH�W�[�!�a|y������I5H�|��\�A��c���j:?�6�*��0�t�rJ4�.h/��CWٟˮ��)pgx�j��K��+WJ\���������Ru�ϞN�Ava���),i��y�@T�<��֖H�C�}��$� 7����.
E�! �{�ts�~�+}��|��$\���(��]�{�A����q.Gr� ��v��1\�U��k�yi��=���Y,q#wy��I�[�΅�gq�%B(�ܸJ�������:�sܩ���{��ި���ܠ��i�b�Bh��m9�.w��(m�<�sﲋ�������MEN���	S��?]���
j�y�,N��,�mtyK�?��_�x�c��.�h��h.6a�vHoe>ǸJ[z�q�t�X>���x)��p-���^������UYԦ)�9�H�#�U�!1�˟?�D��r�Y��*Y#S�o8���VL�29J�����Բr�lכ��;Q��w�u��l��F��Y=񼴨�s��'%Sbj������Ry��@�0��\��K֫iب�cb	z���I��|��_V���]E'Z^<z7c��t9?M��vRD���K�E�Bo9�Gkը�X�g�;��L�$ �Q�F�~ɶ��XE��o�8v.F�]���&W'��$T5�Y���N�f��&i�U��9��dz�c�ϑT�ko��ŭ������� ʭ6�Tږ�>�c詸HI
�R�uَ��B�,���4�ʚ�ږҁS�r�kU
,q�Y�8^Υ��,� �&��3qPZa{��l���vE�­�6Uc�2b�:B�(���%=���F�M"z�K�o�\Ų,�����n�}!
��t�b8϶)T��}�[ʞ����iy�CG�+]���;0��d��Ѱ��'���ܳ�8'N�k�1����)�EI���DG�S�V�	2�	^j,M ��fSʐ��������ٲB]`N����~��K#$��|�C�L�Ґ��x/I,=}�1|H�/Ũ��c�Cݟ�i�q�]�� ͉�IMd��Y�n���=f���о��|[���sA�ֱr��CX G��ID��@X"T$S-�S�FΨ1�t�3���̽*��Ck;
�
��c`�k��w��#s�	5�!��j���
#��c(e�
?_~iE�|��t�ظ���<�c�If0�;�A`4�<NG����~�&	p���]!�n�%�A��KXI� ���!�Q��~�T��(�>}"2Dx#ۤ�����i�c�]�.�o)�'h���/sʃ�r���p?r�Q��#�l�2��5n�+���g6z���P�`����.Яٜo�[��i��*ԧG�jZ|��[�Դ[����;��d����9#��(n�R�̵y��p>rƻ���V�8�P�/Z$�0�ȂLi����>�����/*k�
m���#0�'��*�-�WތcW)�Bom�����6���i�ơ��1�#�B�F���Z[l��\w�^̊��Bj[ N(ƫ,!vQ���ӡ��K���H���g�D��y��dFP���c�po���;5������~�F�Et�F@%g�Kj��s$��@A|ӳ�*�{krz^��oo;�t�������u��������I-��J�)˙�Z�w�k�O�e��rjQ�.����J�E�j�I��ϔ�c��[�h���j��c��� �r[��2}� ����s f�U:�_�X�J�OCE/�y�}���'�K'�ղq��_�QԜ�٣UV�\�Dy��Ѽ=X�.���$��j�e�� ��B�󶺤Hv����c�C`�,��@��.0���B�T�o�'��������v��#vB#�T������X;c���Ώ�82�ݜ�[��v�겄�U9��y9�{�jޡ��&��M06BpD��(��,�8���1��t-�̩L�L�(;S*�|0��G�}�cK!Y/�G����ǻ_9X�������������@̰ؒY�Y7vV@�'r� �m��(���N�R��o=̋��ؾH�45mC�vS���m���LDQH���M-�%݇��Fn��5F�	횏v*���V��7�d��b� �K%n^q#s��nY�=@��Q�F:0w�~�u.����Y�뾍��ްk1��L�C�]ҢǴ�uoN��?�]
Y��N����2�V]�O�y��*
��]�c�h&�s�!���L�#��Z�[����6�A]�7KxEQ�c�_5
-���	���.~��?������o�Hu�����'�	�C�*��Nm�X;�fe��h
�����3zR�'2��cpX�����=�J��[#[�S�Z�`KlI~���/�=U%�T�So7>T����l��_��~
@��!S��t�ݱ�s��9B��11¸��$�v��\�o43[	���m`�b�@s��L%�Wq0)��9���x�gm�k(kF�}��!�2o��3N��ڻ��Bl5��'����Vl�g7��=Q}V���gH��!�t,^���|<�i`N�i��.���0L8�yS���lzA@���J��kT�vtF�vb�ݮ)I�Ls��xhL��r'��`��kYL�`~�. �T�`ۯ�t~���s����˥�
Y��؅ Ƙ�"VJT�����<�b ���~-�U�M	��\���mwY[��G�iBH�D�U��-=G��R��8�0���R!��,ͬ
��靓����6������@�i	����HjL�l�df���r��k`�C� ����R	}:$�]��[��.V�z��;�\��ܷ���Qп�Q�%��ʎ�r�kY뎂2a�r�����x�oK��n��:�1���1,�Ov�WV(Z��ݜ�~�����t{���R�ў�p@����Cƕ:�&�&e���TP��ր@�� s���,!}��Ie�b��NV���l��_�[J����+6��̍� �H}K�¦3DO�\�>�����9�6?ͧsR��c�7@�����P�W?v�5�Q�����F�4����m9���/�f��@�hT���ΖM�ڔ&��$�����筫c)1���6�<dZs�s��*��x��'�à�&��l6vW���ި��������rǠw^D�Y7 ����r.���El�+/���\]o�3�~�|5ّ�ɋ���Y)�Ry�*\1�e���k;i�I��4�!̍�]���*�|V_�uDg�������Mof'��	���x~i.S��K��G�㓍T&A��7�U.!S�]��@������X�y�y��>#N}-�,���N[w��ה���.*[(�o{9
��&�1�ѤX��"x��j]�`J]�Z޼����WS*�C��|��Ԉ��Y�Vt���R��2�n�ь���P;�'��K�O�)�HW��0���z���F�A�P#�h��@�=�N���y���ĵy�N��E�#\f�[�\}�l���F��eJ�|*�_��^�{�40D��k�G|���@=&�#�����Ob�V�C�'�.!�)��yX�?8��oӥ���b&��2����	��qn�)�x�������Դ��xA(v�6� &����[?��hvdQM�&�&\3�Rj��F�GЎ�~�ڵ�}�_A�s�1���z'�߿Kܟ��//�Y��jƜ�$��UP����>��Z�
t��p5��k^b��H�k?�5(D�{c���������rl']���VEN��Ӷ�Fp��������z�/�۶�!֧n.e8���s�R@�^���m`�'�.8���|����H}�m-"b	:���悙M%��zol y���6" ��oe���fikN�%�:*n_��$�����Gj�l5t��n�/�,н��&��1��I��D���N<u����58�3�X\���q��!����Lݭ���٧����X]A�=��U��&=�V��8�J@�������þ@a�V# o�1��t���ki�g�q]�z�vC�(�:��Ni�Gu�'e��k�"ܩ�s�n�$��r=b�8ΒA"|J��#��Ha�*��J���y����*%EF�;!T�Nʶ�sa�KLʤ*�!�kf���/��`�r�-�3�{y��!�a�+.gQ%��J���ʐ3[gK�Ѭ4rcS���	J^?��F0u�p�0g�d%v���궧Iĝ��4Y:O��a��x2��P���hA�(t�b���(vJ��W�ڢR�O���n����6qS�b4e͞\_a��.Ƙ���ѭ��ɧ���7q���=d] `f�o� ��GB���*�<�eg
����z�Z�[~t�~gi�32�N2za
С��U	GBִ�n���w����̜���!h�iP#