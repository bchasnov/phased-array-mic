��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjfm~���*����Z�R�:Y���O�-��_��e~Ws���>�o~[��	>���IWA�+"����M�VZ�,΄�r�#���F�xk4�Պ�HLJ�Sg7���:��Sˤ ذ��̕�;P�Kع��g�5o�=lz����{ Жr(�x��|)V�E�v��:G*��#=&^��ܛ���������uX��rJ��w��!u:��A�Q¸�8�(,z���:�W�0n9��S/����}!���]�{�I(��S��a�q��/�}�J��s3ڧk����mBAEaO��Ű�Sjk��%�y���^�PO�t�����b����[����踛���[f]�5��d��g�3����6���X�%]�geL^ע��n(��T�CR_��}4�MFp���p�ݓ\�ֳ=U0���Gˤ�{�v�����G��܊z�}O�+�aC�[E։Ճ������,3��!�RҰ�A'	� �6dĎ��S}5�HD���}'q�j���A����Ww�H�d5?�8�;�De&ATG��H1����V�/)Cjõ=�]������k4]+s^���:4! c����OwI/�7m��8U^fB���R�qx
����=D8�"}7�������[r��VXU,oy�'QK����cq�K0�}��3�ʟ��hm��rp�OC�=S:Gi��ԫa�紗�r�w�迁�怶��>:��.3E U9�D��4��~�ۆf���m2肩!�ϒ�z"�������`|V_���N��
�{V�U��П4�b8�|D��y��E$�;�|G�Zԕv�m����2գ��2\c�#F�^m�T����(���v�P_��s.���^�?,�֫�U5A�y2���q1y,\�q��	E�J
�]���)���~�o�uy1AJc��H�(F$qy�"Ҋ���Û���r|U[:��)�o�MI�_� y��<�w\K����6w��¸W2��ϓ�P�E/��0�mAB0&L��	�S�.�`�$�����+�zꐟ��j�!��"k���:�N�0���;{�zA�}��q®�p5�/��ܗ�R�
��;�~�����ck��ȝ�=��~�7����勒jGgrR�Bܚ���
��23$��?<�m7�TR���v5oix��6T[����e��h�jx�>���R�j��5n����>�����$]�)W�4��˵ˠ�Cuvq�$|\%�|eF��A��i)��Q�X]ò���]새�K3�ښ2G���NO0zh��~b���Z�6�)�N]�L���Mo��� J]��o������ޓ~8)�/�Z3lҒ�<z��F�3*fmY���߲���J����
q��B�
�@��^�^z#w�.����Kr��#.�cW�P]K��]������ؗ�ū!��xX��Qx�@]jI���}�<bD�[�qzZ��W>N�s�˾S�~�X��"�{ّx	�a`j��m4Κ#���A`�� �<��4p�S�Yч�����S ��4��F��ƹD�q$]��`��sHl	ͣ��ҁ�G)��qhj��(�.4V ��NV�SSw���>_�hw��_���Л\.��[HnȁL�ct�2J�����'xɗ����d�����TM�O�M�~�Q0��H\9s�l_���^��ƛ�ɷ�f�􃀭7e�K�7�'M�폚���Z-+�f���s��V�=�}H��l:���.�1�\�f5�!u�٥^H{8����}@�@��o|Ϡ5��I�����Y�"(�#c���HZ2=���D�����d�`�ZUAT���NLA|i(�8P�(�!�;):�5�ߔ.��w�ahy��aF6��WbUli8�6�bkN�R�)�a���!�{?�9w0!06�e'�f�q�r��~̾�¢���J�
ZN��6�On�W���$�2�u����7^XVL�57ӄ�&S�!O�0w[9\�� I �5M����̀Kz���&U*G��$�|�@�(���'?VEڰw<�2��d�~�	NCGo/ve��G���k�ED��܋����!/�О��J�Ϣ.�S6�i��%)�3A1���3�	~8M�;f�?a�� ��a@��Y��<D�r�� En��ɡ>�Ǝ\}OJ�0.��6�	�y�TL�$1.�SÈ��S��
�2Ip5�d�x�6\��<.vL0$P����ҁED�p�X�U���ǧ�Pyco��4Fx�Ѩv$����)d�%�������M�kd���B�o�z`�b���:<0�ƿ�/�p?���w`8ŝ�\	_�Ax�+��3��i��Jĩ$�lBl1�n��qY8���/��"��nt�K.���\�zl�^ıqL{��8��vN�ƺ(r����El6����j@_^\L���ə5�`��;���Ej��	*2R*W���Es���*���?P�p�ܽ8�pp�d�<�Dyb�g9 ������Okt�g0!���w�
J�p��a!�˘ZJ�_�z�t�ih�K�W�4��T����P���j"��iQ��|���+��I/�9�o���nt��U�aT%�HE��d��}���$��&�&�	$�n�a�d��~"�q �3�0 Y����za+�6��=�`�dC����'�{��y�)U�'����+.���F��[���6�a��T���.��wm$�k�+i���6�E)|�2t��|�t���\-�q՟w�ٺ��w~?�Ɇ� �k2y��y�N
~dc]��[�;T57�m����K��>��iR��4G�g@���mf�_o砨``����k(�'>͛�ױl�̦�D�E�o�h�a���F!�Uo���Hd���-g��lÉ��T��{2,�v[椪���}B�Pc���+��^�B6	UH�C����!���b�L��2�ͩ�F;<a�*-�#�4o����I~G�,��=�d����Lv�u�Z@�gw�mxR98�cTF��Y1�sMʍ���TTʣ���3[���i�M_�׏���б�]U�;�8�W�`����gk��(Ƌ����B�
��|�6�Ia��v4L���r�R�ʘ����z$�3�^,�6a�<��y����l�G5 0��<��e���tj�qz��=��R#ᆐy|��3��Ę�v,�'�A3nrJ����?�U��1E�҈��N���ڄ�aN���~2�]����v�S{ی31�%D������ho{�WO�$���.,���NSd�Ĳ:�#�%�ƭ�yp�5<:�)��?�X�[�?���4+�A�Kֈ-]3���:u��WnK�`��\��JP�V^����N���m��~�6�l;^ԋY�.�d�<y���#��մ����<u3a���õ��J�t��>�P��&��+�?ﹼ��܌y=���t6A7��Uݝl�)��|��?˧ﻁޒ���ofL����b�Fn6���o��n��Yg�UV�=&�-�%��&��[�*�lX9f�X�#`Ž���{$����7 k�C�A���9�͟� n�{S���AƁ�F��K]�6Qm�~����T��\��'�99�?H����*�_�T�J&�sp���(����߁�Cl[}n	�^~k�������}lc�ꯛ^f�*�ė�-݁�8��W���!\d(ǝݶ�~k�G�4[�������܈22�����f��J5�T���e I�p ��i����E��Pl�ѓ������Y�_���s�X�s��U�_�ET��.B�+>���.`B���X|��7+H�|Q7��K!��I ���Ɓ�@Oa��$��L�nU����5�!�
�����Ǡ��u�k��ʢ����tO��w���`F�Ȃ��{7�^��w���D��)ꀞ��[�E�S'U��ʩ3�7L|��g���_9	�е�9�B�!ӱ޿/�q��%�!7���A�>�%�[�M�eJ~��-9�w�l��$�͝���$�Έ�TdGI};$є�Z��j����7��D���^��� ���~�A�`<��4¶�d$<63$�#�%��.�r�ѫ�{�4/\@IA�~Rv�{��{^����C�����vp�F��$e�]2�Η���>o'����3Н�P
9���!��ip���P�n�F��xn�@`���dB0A٣ڣ�`p�� ��Dp�,9gK��g�=P���]�|��"S�4�N0������t�R�/0�k�0��x��z�h/�x�B��(*QC�Ϧ!�'	��C�㪰&p*̽�G`ѱ<��y�	�H7�B� L�q����h��C�y{�Ϸ�~�CĖ�r�35n�������|i�)N��=d�$�w�4�/^3r%pbOEܿp#z ��_b� ؖЯ�F��\�ո��f�����4���t�	��0٪���j�� ���*�@?�'�,�e�aH���yr�b�|����r}����g��y�`��	�eQ���1����])Up�"gX�c�* �}ng��F��
!�����L����D����O#�	�%D��R�dn��׏���VW�^x"k�ga�a�Ś��uйɳ�	v��DƳ7^���Ղ���9�Ǿ%\�a����כ� Q�l\(�j����a�I���4��Kz�C�:xjy��\(G+~dB`Sٷ ��uz2�ʺ�K~���B)�BS���A�Z��Ȫ&��g�i���#�nKJ�SOB`-���!���4�Qԝ����e��ɓ�f 8m��D�ڔ�ڧ�y�i�_�6��癕jXE�i��=邹;t��2 cy��$KW���Η�)���j���Vf�)��#M� ��6���E�{�Mؚ�U�����(�B$�&��W��`|J� �ܭ�����G�O�\_x��ڒDC�]:���� X�D��J�̾��'���@���d��~�p�!��b}����/��[Y"$N��1YV���re�1����{6��FMT+�����-�b�a0���=���U#�SeoA;oB�Ҡ�U��`�l8�X�r�*yEs���@�y�<|d*;�a�<~��C��r��S�r�P�4l��*k�vO�P��ȧ��'�c�M�Z%�����h���H}з�/���Tb'l8�#q�?3���
g(�|�/���4ߨ�u7�o�J9F8A�� ���b�.�1vh��r�(PF��q������豸����������o"����N����0i%��O~�(P���I�.���h�&+X�kY;U��3���3BW�I�;ꖼP��~��fS�^� �j�F8���͞����M~�c��]:@=���,����)�C 7k+�xa(�N��[��fև}&�-�<XYŦ��5y�mxBy���,"�������|����Tl-w3尳4g�ė�}��`����"2���r��b9^ؙͿX�ܬ��c� �-#�:+��,����9Z�~�7I�Blu�/z4X���GH�2M>��Cْ� �:NP!�v[W]���P���EG�WﺪJԦ�+I�^[]�:(�mKO�LT�|RAM4� 4�Bm�䜰�2r#Z����e����Q�\�ꌡ�O� 5��"�ib9 @Hpz�������U1f>:L�@�{�����m�uʲ~�E��	�*d��u��F�G,[�3���f�L��|�g8�P��FH_��bLو(˥O���b�eE[����SxX~iZ)����)���b��g9�r��er4����&P��4�-N#/��0��!YM:ptTl�Wk��{����\�����z��>YM�d�s7���gI����ŹvH�t����F�LS279mgIE��	%MMU���WD0юl˶�#���t�^X0�L��`�h�*^g�!o�hl�,WI�={!��RB���l����N#<�t��ov?��E�z������%
���&Ӣ3_�c��ȶ�AL��h3�`}����\Wu��]���.vk)��Uq�� &cI��=�Q��խ��:�H� 7;6�\  ������}���v����e��W7���H�?�2��@��E{����|�M�Iȥ.��f��A�4+�hT��nd�t��T�Ѝ�EC�K�PN���
���e�p�xzCJXجHjOe�ׯ��G�F��a��a3:�ʹ��%Z�;��ǘ��	�d��N���eݝ�E����p��s7�:K5e�λ;bDT��4�!�j�YW�����لD�AS�o�W��1�o��	�,�/���4��p2ˌ�$(���*���2��RY��2����4W����4��~��d{(6�K
4@�H��e�BLv����C<+��S�;��D� ayh�
Gc�թN�$32޾[��R�N��b������޺N8ʞ�z��7I"���Q�y�Pp�Ck���\!�y,py֛\Jg�+mL����(^�+ɥ�'u�J��R��8��ͧ�!4K�>���]����ju%,l����ɍŊ��6g��ؒ��\c����$\8�<�*�q8jG���K$Z6��7��_����h�n.|������]"&�c�[�*!*��a�[]] B�7j�,q���_���3��¹[�D���� P�f�K�_�^�/��B�S��jG�t�j���(��	s��G����8c(�X�%.F?q�SXO�>T����g ��y�����B�:�+tO#f��s�Y�=~/�af4�Z��k�F�DrD�~�����X�_�m���2����^�G�(;���|���i�Q�p��!U2`l$Y�i"��n�qs_��_LNìUt��Z���?��OVl�v0P.-�n�>�l�{<ؖ!��z�sͬ�ǲ �$
�널�3kֻ�t����XJ-�H4�����Ryb�9V?�:�̳R�8���5/ ����l�����j`e�'������_v뗔�q��Tg�S(�<�������^������7	�������,���0�+����7I~���-F�����4���N�u.�*w�y�F}�:�3N���3�h��=��R�4حeP Y�G��>��:�~�jܡC��KA<P���S3bb<y<Ej�g�ߥ�������mC���&[j�w��C���*� ��p�?�r2_W�H��?�G�ޞT�? <fNs)B/��d��l��ű:�]�~"�s��N�sZI�WO��W��S��m�&�`�$?i!-{!X�X\�Bj�~��+3k��ȉ��AՐ�������U���̥8���+��mp�S��;�ݰ�����
�|�4o������u�}��P5;y� �͝�O\�1�G�m��l�@1�G��Y8�MA��8'��cS�g�\�M�W�츪��ʏng����] ���nl��1�Q��!�T�"5P�J�o��s�"�����=��Dt��4h 3���G5�ўu`��6�s�5��ʱ-fK���|(&�����Ը2o�+.�*���A���0l���Ox�C�B
� }h��d�Q�����>#TP˔H����7GHJ0*O��&Β@��h�HM��Za�M��RT��)���߳��t1zVݓ۳��Gl\N%�Y���v9G��T\��68��n>{a�J)�<d�'��mv� Lvbv̈!��A�.aX �ӏ��qʚ���e��8��f��2����IS�hmf8iyƝ�M࿛R�÷	�\AñP�z�h���a�ĝ="fIȶ{��{���;2�N�<���� ^����fڈ��D���޺u�YiF�;��
y.�Z������R�n�BQz����Zs-�:C~�}��p�J��BU����Q ^����f|�F����ȯ������JÌ	����S�����q6�K؛�jf��dd`�T��z�V+"}��
��̠�A ��ZZ�:s'�S�r�m�g��mJ�Pш�&|�9���c���lg�z_!a��S�A=������VV
q�>_ө�g'~s����R�-�g��(�k�tڿ�<,����H�V��ڵٸ�|k�����F��$f�^����y�CBI����e�ش�!��ݙq�>�Ƿw�$��|��^J-�م����i#�s�qSD����V\��BR�m?�R��e�Q��t `�`_r���=w3��	�Fay�D5FƧL�9�Ȍ���#�z'RG�Ԅ�O��J%��X����3צּ�p��[�~0_�:,D����a�熧�R��F�x�9�������I�%%f�WC3�@R�;�z�Mض��:"��D�8�ZYKa�[���w��qgr4j�%�_U�mLP:%q�Ц�QOY+}I�-r]��0�'2����<������{1�np���f��FƖ0d��;C`Cq���g��`���lռ�O��R^�H%�c�D�����KV��5�����W�qu�'�.�%�杵�ߢع�)Tn��e.�گ������/�T�2B0�����<��.=�i��a��@��&��l���Ƈ��+�,���IOnR�'>, �f��D�z�Aт/�/���-b	 �̴*��Ͷ �F��*Ead�T&z�Ň7�J2����,`A�S�~@)��L�l�l��U8�4ahp�0g�TTM,�d�%����21j� ���F�Ø�����^��M{&;Qrc"RL�2U���{��<�/ǘio=����J*G�����x����@"���b,�_Ac��H�2� �X��b߸Np]�#J������#:���V_����܉]dL5�^yt�����iO)51z�p���#�J֧�8Qjlo�~�-�T	9����U�5�WBK�֍�m;P�P�)��_r��K�f�s��W/�tV:�?->���k�oe���=���!�/�Ǒlg��� �?%ח�%����Lu���,S|��f�y��z�h�q���E��jΧ��Q�zz�~o1���{�����'�ҋ�H��E���}m�X�fB�va����#�g�G�Kۀ[k��� Ɔ$�+��M�(_i�pN�,B�b��k�~��������bW�X��6��yb����·��0��Q�A�-BP��z��	Z.1�\�K���U��K;��q�0$����:�+��2�^�J�I��VFU���[	���*B1����W׸��g��y:��Q ��Pܓ��[�0B�S6��*���O4d��Z;陷�n�оؑc��Cv�}f�nO�GTx��]@����"���x�P��(X��I�܇���Р����""���	X��K��� %v��h�5��	�<�8Xd�j�O���Q�a�ݢ&DB�k;����Ç"j��a��_IA}�!Aμ�-]���}$�6.�=��GB�jݝ�H� �/U��c�����.�1�.6�����fÊwT6����2��䭐 $̫��H0�����6&赬��n�P�|�x�M�6��{G*TD�8��n&5�Yɮy��ʟS�9]Wu]�Om&_�FV�7��P���O
�M��J MF��tT��.���z.�y�q���(��5�"�`"�7=*F��[% �o.1�ȉ�z�W��J�G��7�m���� .�[ދ�����'0ϭ���Lbw%B�����+�+��$:����&!LBC3胕�_	���i�+�ֈ{�����Q?�����|����lYi*ޱƾJH(ܻU��ލ!�"Ce�����b2�C��~at���V����;��t9�{�}N���}�S�&����a�_��7��%|�[cPr��Pl�|}%����8�^��D���P/�.6����_m�x�,��S�	���1mWv\.��&cW��r���X3�H���������wU�.q�ǡ\߄���v?"��#�kl�Ԗ��2l�f������Y{��9�P��(�DYAߩ`i�,e�c����	,7���P$�>�^��� D�^O��Ac���^(�C�ܯ*~@�˂�b1��N!lsk�3��[�K��2�%!�d�5VH������P��d��_=P���i��4�:&V}�f�{���?�o���d��������w�^�D4e�/o��)�D�8h@�{y�H�کw�x���A�[�:������<��k����@���Ţ�C��)o��W�0H��c�z�g1�C����Ͼ���|��Tf�E~��ǜ��]��l,s��J��(���>�g�8m��$˞� �O�{����b�Ia�Y�]T9���,YO�Xq?��yE�Z�r�-��{�;���;��4���X��E7R�:pWMhV�`��'"{B��н���oH	�"f��J��>66+�E|�m��!~���܁�BK�-b�pT�ߜr�)��6Z�B��մCo�v���/��c.!�p}G�`a�)�4ݽ. � Ҽ��R�T[uq���j����)��`��m��y,lp�������F~)�S3;SHt��g��"��m����m4ꀪ�"��o���H�\�_�2Fa�^ɋ��~�{O�3�LN&��Kф�[X�A�+�:���i���S��!5�+�=kU�D��-������p	�)��*�����u�����ϖG�ţЕ�h�F	�g_=>O��@#����rǙ.��.tٜ�ôS>���k��%�a�� �!�oO�
���Fſ<Uk����G�H�����!+�XJ!��@���k�r-�j��q�y!�_�r�a�筊��MG��"�휞�5�֮�Y����kk��v��3��g�g@m&b� �WM����積$y�J��zZ/��I2	��1�P�c�*L�����I�0�2F��>�� �x�����\Y0^������/��2fb7�w%U�Ӟ�l7��>����h�Y�7���]�7D����8@� 7�"���i�����ӑ�]n��b�AÓ
�RO����RL��BkFǅ�z�t�U� �t��@rAZs�%mNIL���mІo�vP6ZN����7��8��$I��p`���K�bƹ9�Y$��ܒ�^��"�1u*�xd�6�<U.":K��e# {k�á����>.U�ܥ8��Cl�7�%g0�B��a�JA7� d|�.E�@�	"*����_#i��fH���J�����R?��T��P�Q�n�"κ�.���[�Ee2��ל{v�+���g
����@FG\Aۍ�P+���^I�`Ƨ:�mY�s����E
"�o[��^�O[H��3��V��E�[�n��@I�����/_���[�:޹�^�-ڧ���8���Wjh�NI{盢�ue��*��5)�nm"�ц��󚀺I�UW��CÜ����@>�BZo#FV�.n� Kֺ��_;E��I$P*���cܴL���m
��G)���G���CS�Z��:�:��Ac�o�U����i��#����W�����P܎�d�4���M��uy���3fP�/�I0���9S���ՠW{�º)O��X@�<t�2É�+|s
փ��\�n
.�v1
9�9�V�&��W'f���?9�M�_
������9��%Y&y�`��	�۲��[������X�T�I�I�#3,�|�J[��}�1�6�0��ڻ�b����*�i��!|%����}�*3�������z��\���+	�B �V|�6��)�WE���Ϫ�\@�%���"����5����1k��i���C�ɑ޾J�@��7�P춌6����+l8o^1J^ۖ�鄸�j����$��-o.�:�[�0�%v��tK�y�������Ì?�e*�u��2�ɸ׼9�i��k��u�#��E:�_������%� ��&ehZh�Ԯ�������������~$uP�a�.���業��5!�'ej��Ǡ�l�fXÐ@hP��P' ����gB�_��Gb����G'���a�M~�����W����nخ���p����r�vv�bX١�j]_�1[���&E��ӣ���6��wGn�*K*:�}��	�d����!��E�t�i �P��ʁô�`�l�����/k����c��e��M�{�]O�Q���u�f�Ra݅�v�=��F�XЕ�ƒ��c��z:�3!�^�6�`F9Oԏ�����͗ʇ�b@��[��JU!/O}z	�;�QTV/e�yz6MCgC�]��~�ꉝ���n��꓏jɞ?v�]��=YL�]]:#�w���|wD��@�?pv^�t��~�
�0|/���(n��Eкc3�p�#�� ��b�!����,���`�9�A��GU3ɔ��E���0K˕$�>Vq�M��
q����(&�d-(�N���?���8�~Vj�=g��˼��\֦G��7us#�����L�����Z\�SB�&-V>DjVc`���Pe�^�K$�}H)ʢ����!�ӌ}2��Ir�x#R_ F���M�����5E>10����uw@P�}�~ꜞ��d�~�rS
$�o���1NA:��U���&ട���k,z��wŷx�%
z[��V���=��h%aQ�re0t{�[��0k��0�3f����;�cXdh�`�X��3A�9]y��p���D��"�*l9��[��j���9)���3_�BH_)<�z�'�wD���׾�h��-1y�סz�4�.��`��G��R�����=C��P����y,!�kVA<���L����1���^����K2�m�6ͺ���z�<�M/�M��u�s�4�Ɓ#L�Opz��n�,��A�%�=�\�������7�3I
�LX������~oo}�����=����Q�}e��۱�e�e��y��}f}ך��kId>Ԭg�b�4�x����qm�0��k�\�R��$�j}�ϡ�w)��_�5�r�mƮ=��c��5:������ ����b�x���gF� ��]o{<��t�^Z�ړ	�Do�E��ҩ�O˞HVH��8sTH��ǋ��N��9� ���>|_�%s�5^��is�^�~����0|����e��q{4o`�3�6Hv��_�\o������Q����Y���"���{Hۉ���V ����{��Q¸����:���\���ծ���i���SO���Q*��Z��y����0�ipMG->x \��{�3X�zm���a�~���9��-���H�(D�2�Η�7�$N��RNp9�իPJ�BU��-�+B�0>��� ����mxJ��k �yI�[��I��@a�k�w�����x! �YH��4��-3�v���� o�����߭���6�>�KK�TP�9�w��cۺ;��%��"�3;{|�3�s�{DH�m��Fh-�򸴀M������Qڨ�횘�?�(���7qS%�r��F�r(J�6��)��N�0*b҇������?�術(��CWj��V��Y��l�q��'��$�yqQ^��~�Iu�N"Z���A�D9ucܙ��2/J;�@���)����ᗦ,�f������W΄��{iXA|�Z7j����\C��˩۶����p&�JM�U�������!4��I"��t�_����$��6�܂7�3P��D�D>���t�0���ѕwQ��$���A@�L^�$1��0d�<~5�4������QeK�'G��r�ټ?��J?{��l`Y�n��c2آ`17+��)��X�ai:l'��^�c��=i����n�gxs������y�B��ޒ;�����bt�+���<er��|�p<1'�6�PU�G]�On��0���E�A-��F�m��һw���l'%]*��5ܾ��Tm�@�Y��]�I~U��<��oq|.j��	!`?<�"�Lq�k�`�ף;;�����œ��8h��>g*�wŌs������hU#���mP� ��m�?�d��X���P��s׫;�(�̌k\ˡ�0��|Q+^r`][����/&�YZ7[�.~..2���3t0z�c��ir���ډ]k*u�3�pe��Y�V�yag*/5��Y���)���f��Jv�����Z��~�!Ĉ��!øR{�<2��3E�u�򳞥C�\��;ڤ�I��w���Z$}�:�E�kY=�5iA�n��&B\��hΠ=/�t�<M�,����	�G���)L��*�|U�-�]�7�F��e.Ym�O�P�2�#_=Bo��Ŋ=,��j(C�g�O�l��f3��Ļ@���y���e��0ً�ѩ���V�t(G����T[˿Qb��>�a�� 	�`���>V����*EMA��,��>Ay=��z˿��|0nC'��)�Ù1(b����:�H�O��ߢMZ�&���h���Ľ�0�+���2秃}Rp��3d�A6�d�[(��n��=�������3�3e~�<H	8�
bǚod������C�g�z,�&���4�=�;�pL�sn���@��/�����ޘ��5�eǷ ['���($&~I����a��Ix����4�N^NPzKa���G����=5]��W�L�ܕ�����n;� ���ڽ�[�ۦ�l.�a8~B
Y��PB��e���D���^N�V/�$�J)��{ɐ͡bpj�2u'܀���,�k�g�ֶ!w}�A��[}�0PbA5]�������37�1�����x`~���-O ?�D\M�)����^�v���2�H�és��w7�Adc����^+��	Z�U���A����|��>R�*!�1 �����]S!���Y5~n�� �Ɩ��b��5����/:�;�_�S� Gs2?��'|{�N=�B&<��K�@=M�-��<�d�F���M�_|2�Û\���:����<e�{#�u�Uĭ��\�6Y��������
t������V�Ս�z��`}��R%�9�쟡d�j8��7IW��$2���Γ�K�{�Ƀ�K����f��vPe����oݢ�������?�[5����ʊ����KAx.q�hy�;@��a�՘�j%��.O�K�����ks�:d�o{����5��Z%(��M5��VEJ�_w�����t��"3ʣ�������=e&,nw����l�CΚ:����Z�/qʙ⹄���U��@�������|f,ftclke�xx?�w^��4I����c��ۥ��Q-C0��-�K���_LhHud2�+Y�,[&T��&C�+/*��OZ�a���M�ˎ���"$6g#���MwB]e�㭊�p`���(K�nh���L�����W�v�S�7>>��\��\��~�]�5�o�(�R�MW��)��x���\U���ҼQ��a	�"�}�'�kH�p�_�P�Fq��7�U`}�������..w����&-��;�+j�=XZ���� ��b�^�0�.���J�׺++��}.o�v�<3ٛL�%3��L�q�	4BH�<����BqHa4�~�V����� �� ��չ��xԇ,�m�m7"��cQ/)����)f���E7����$C�_�5�m����{�ֲ�N�b.V��d��B9�n�83���E2��l�)-T��V&�N��!�(����U�9��kG�EL#�?<?�5M4X�����������J4>�y
#���`&��eb�,*�z5t����!�򺂣5�W�����o�-�C��c}4��n�o�1��y� ˡ#�q��Veb���9K&e<�"�_K�;��F�A6#�G��Ʉ��Α��3v�6Sv�*¦�\�K]$�_. �g;�q�T7�Eo��O�=؃C�!p���5�	��i�6���
��%R��΂0�c_�����·�nEZ������tjE�����| @f;g�%��H������aB����m��
��c����,x{$��},�M��D�}e��KMW�[�#ֿ���N�cG�kֶk)NxҖ�&��5�!	�7T}�|A�֋C��n���ϸ֡�z��ËۂG:Wŷ�t�ϓ�ڎ.%��hQ�h���8��YP���y��1��:g`g��� �����d򌮿ϚrqW�g��y���<�[�M�Y��>baΗ"8��b�+��/V�v���`*�1s%] 4v�7�D�4Ys
6�0 	�j�n>2E��]�=�7�7�L��>���F�n;�2��L��&����)���aܕ��v��[���[>H�k�+�T�n�2(pk��i�t# ����i���� �O�ñ����:eh�]g�X����h��'ێ�>�Z��7�u������0��| Z�+�D�� (��z#9w��on�!��D�i,N�YW��.wO(�ȕKW@#[�7��[:8���4�Y�{l�����"�b몞_.¬bI��L5_������'E�����&�)�jZv����S��m'�Dg��Ϡ��i5�i�@�8�٘��H^Q?+�#7iC�^/�(w=ܠj�o��8VWn��>Vm�X������q -慃-���'�9o�@aiJc��z&����X���`�oc�0��[�f������-�~����b�r�����e�df��u����������������E��3�S�#qh+Ͳʱa��1�w�F��r5´f+f�_�4l�)���2߻�ع���I�~f�g1 T�I�c�ط�h�ڽ�w(����$h�<�품~�c� (�1�%E3V:��"�*bj�2M��&�1�M�E��Q�+�#͒Q��S��c@�G9�> ��ʉl�@ؾ3z*���+r�s"MAM7�r'f![nI��P��'.�4dQ]��0E?�y���$���>j�������3�~����x�+����,i��G<X�Q�	�iѭ�5���  ��
lhp��l%� ��@R���m��]OL�hjP��j�s�!����b�;v�`)�%+���v��+d1�����]lF����λ�<NM�&�0@.``���ڿ�`Do�)�/���0��6�'���V�(�z�f:��"u�#���2sʎ��q�j��zE���Y��-�W_[m�v�y	�@�04]!;�=ĿZ<�;)aU�Bw�V�)�p�s�;�����(��կ�:f��0��� ]�d]�S #�q��|��:��%��YUZ�T��ُE�.Tf��B�1����e�O�sS5�#}��Z$�tu���W�qC�e�1��;��F����f�����j�*�[}��i����A���t��Yw.����$ �&R�+���><����4�Qռo��f0�j�*B�oɒ�i����ilm�9��>�����9�a�X*�+��H7��I�	���*;)?~D�D��CP3)�����`~�As�ߦmpLE\w�c�ʊ�!�����'�OJ����nU��Є1u�bcrN�_��G���=�D)ì:��b�d���XJ�?Dt09l0�
��a@�=��m$G-�4D�լ�
6��%;l������P��s�S(��S�-�#��Dҳ.�����������lx��/�哄xs�KI�L� ;nѧ]��ъuS����l>r���d$7�?����V0p��ĩ�T�4���:r�v�3�w�dV{`瘣���f�u��P+}^�ޙZ�@�� ��yݸNƛA�Yp��9ϒfM����Mȧ��2�}VQ�~�<3,o�[վi5��xLYO ���>4o���t����G�w�7��uU9�"�!셬���ߡ�W���'�������ʒC튼�x���l%-�ˌ�2��p9e��WY�AC�.�������4�u?18a�b�����*9��+*���~�Vgef�fS�Ľ�a%��2��w�Iy��@g���Q�SW7ֹ/�Xo|�d��J.�����b�]nj�M������=�
�h�`1;M���7����H��#��$�P��)q�n/�����=������G�a#�n��/�#(�n�Qt�l��w���剀 Ͱ���â��g�_�Y�^W��DI��J�"z�Y��<dI�kg�$P0��^@�~�s��!�*���M�2#p]fާ�X�[{u���I�$^��U���c`zv�V¦Xx(#�ў������$	��l��Q'�J��?����h;�\�+�U[����Z�C����;cw�j�M�}���N��*��a��'6���r�%ews���閨Ȩ�u�i�d)��|����jBN��� b��P1���p���2⦨�p�9�
~��U/Q�r1r��,6O�x���E�M���K�%J}��cN������bK9��,��K���,o��x�g�D�Z]ap u��8�sZ����87k�Vr�*�]b{�δCz�-u��M}�T�X%��i�`����-�.D���j%��+�eiK����^�\�K��"i��`Ȭ���&&��Y�<]_r�V��O�����wX!�
We#�Sa��>2�e����E�Pp�}�A�]]�pE� ;O׮�@/��C|���d��"\�b�{�(�K�LH��? �����g������5ր���l�����z����10�?���'�%)�RX�qx����O�2�U,uֱ�u�ɩ�!%��|��Z��ITt��c�RǕ)�0mO�'�є�ηpu���H���2b�~�;�ӕ�}��7�
c{�<��a`���#���~�FġY|C奅�1���pZ��]~����#$�HZ�gcc&
�Jw���7��yn;ECY2<5�~�"o�$z��`�eB��l�s���(y�l>xY��	Dl�M������RV�|�s��1��1͊B�[S-�:CW��4�n�ʵ�ʇ�w x'"}��Z>���)�P�֪~��O�d�Js�h�Lt��WnQ�1�W@��?���B�].D)1�#+���p�o{rb*�i��lfwA1@B����D�	�`ڷ�$�eb���̃131~����:;��n+�lQlz�?ΡL��9op p��R]�����ۜK9��L4�w��Q��l�� t���>�@����Bi�M_U�����|�ţ @�fǳ<�βJȼ[���yF�ٴ��@!��hw	��WI�y/&,S�~>FA������8�vUxjڄ�E6��7P��}ޚ�8�7~�[�w��(u 0���y"^�»�*�?�UY��AT���
Fo��u�0a�5?o淚�����d���>q�V}��2�`7N]��0̊��0�;��T���.�F��B��8�����Xh*��i�=L��ɴ:��XƧ���Oڦ�y���ʘ��J/��_/���X��<X!�n��e�:<�01kp4���z>���s՗��+��b-��ܧ��V��Z[�h�j&�Ϻ��F���"�܉sG��֒w3F�6_�J{W�=��$n�W?/.HC�	���U��ŀV������_w��ī���<B>-���J��c��5 ���I��I��B^Gnq�jزci�A�:Ji�j9^^��a<w#�=�=c����AO�T��%ˉ���H�;�u�"j��
O�>��3�|��7�i��un6�A�jر�-fs���*i�!���gLu��Ը��� hY���X���)S�Z����`3`��0U�SS�d;_o%��w�nMx
��AB�;�#���?��;�F�3m�,�6������ɀ��D0�b��g3�pn�ej�t�L��*��3�9O��#��r�zp��I�B\ �o|P[}�2��3�?Q<P�ǈ��6��H�,�Ŀ�ū��vj�y郂�K	����V" �S&0�GC���[�כK�JLLn_C|/A!�VR��W�"S��1��Vd/�����i���3Q$k��~J��2��q�7Z�w��+�%t_��L-LI�0����;�i�$�5��:�-u����:�9��y-��B@ʿ^L�[����J/�H���k@�x� ����1_�c�����҇���M&\c���#,ۄ�;���@$zs2h8N��I�2�����g_mw�=���Cc��7��X�F���+�k�����z.b�-##h1����a�T\%Ň�ؠ�� �Ob��D�V��b	��� �t"Լi�2*_�Kހ¥p�z�֡�y��C�v��H���=H��k�%�p�D�{t�:�fAٗ��O)�0wq�3�V���P��ٝ6�PSPS"�C�2�8�%ضA��s7��.������Zq��
��Z*H*ٽ�'?�*cўPi�߼���w�}���N4z�`Fa��r��GMc�R�Hw���nG��]6���n��`�!]c��X���s�{kl�#�}X`��M�0f�Q���}��2�t��:S�r&��t�u�謅f�4$��N](h�Ks�b��+�K�k;@_8(���j>
��d�sm�5�[�dC��;v��*�/᭵δ:e��/�#	U�(�.�N)7��"|֎�2��z,�@KM�2�.�$Q���-|Ρ;͛�A���D;T7�"�4��o�akr\�v˧h�&c�e�ɶ�K6����L��|�|uAtpj�μ���) /��*2�u�V�z��5S*���)�������Mo*��(w���:�ǀK���Z_�R��e���Wf$�r��~�zK$U�	���u%ly�d�.jl��������+V�H�=���ďX�HB��}G��v�������h��.<� u�#o��D�4����#������ w;v>�A��7u�|�,8U�^'�̔�Sm�(9Vs��d��I��S+���R��iĴzADx��$��I��]��}[��>t�J�oR���;��	�������'']X�9��a.4�IU}����� �iA�~��N�92��C�i��JyV��;��a��U�Q_d87��*�z(�Nj��<Ķ	{Lj0����6�vL��y8�V���c�#�'�=|��t
�r\t��������Z��a�a�T߇C	ǋ��j���UC��S���~jV�R��`����~�@�ܱ �&B�g���A���۸�R�x��3���Ľ�&n�x�%�H��/ ���`P�E3�JtmI�nO�pE��d�'r�^�r0)`�#�0�U�_A^��}��ݞM��Tez�Jj9Q��6w?��Д��>�l���n�$@�����ˆ���>��D�m%�	iT.e���@�N}����S<��q��蕩:�C�?�$���
���!�H�>���s�)oǉ⦁�W�/]��0��ئH�n+h����Ct��g�A�����&��Z�^v�OM�����9��Yҭ�W�I3˱mxtE#��W�S���n����8_`�R/�̗o��`u�Itu�l��p��I+����Aw9+ɛSXA�}�]��)U�ˇ�2[h�|�^Fu	��S��3q�=��%�'ir��}�!��'
d�	�����<��V��,�w��>Q+RA;�눒f:Er�.w+W�e�ж���+�6��P�Pl�BS�l�Yy��!b%��<툣O����6=[��d_�b������
�8���K*�,D��C���u�<4�f��Co�����.�:�j�MͰX�6=�hQg)�65�Ʃ�O:�󷡊��_;����⭋
V	�o���2�BK��ʡ`ܻ��蹅w?Z���#�h�m(��w?`&WD|�LᏒ�4�w�$�� �b�N�p:+ر����^FN(�*�\����B�-Q���$X�>]��U��qyGq?��xR�bms��AA]�Ù�D?{|�~�ya��~�@%���h >kmTS_�WrzKz,�����={^�{�y�[^!����zn�>T|�e
6� �}L��f�������~+���Z;B�ڝ����`�9���w3o���W�v4�Q`9�dU:G�7��ȬM\O3�_UhLɊ�j���M	 �U��- '6��K:���vq2�^��՝nvR��%��C�;}6M�!)*b,ۡo��*H��1�	\\퍔�m?����F�+��?h�����X�.�X�=j�����2�2�X�3=à��UZ*�r��<j7��L!)���Y���ˬl�Dp��}�\?ibi�e��V�	���"h����wP(��g/��р�׿?����7C�y[Bor����rb;�����9����(NA����tN:����	��s�>r���]E�Ҫg����n��GI�퓆��돔L�尻�U���,8�&!_���#zo$�a"D�r.��䂼�(��J5D�UB���O�PR�p�
��G�G��0�ɕ���`��m��!I����[����#{gk���^�+訲��ͷ�=9 CT����j(�z�F�y�E�e�s%mv�b�*_ng�L��I�5n��"�)ݓ��4��7�XSd}Z�"`�^L�\�<��<;ʛ�DU��qF��^1�@[����?�\N�狟�\-�B������D��[�UY�ܹ��!�<��t���9184��u��fM�� yb��2C�ZK��+ ���j��j�|xi,5A�ٓU��+�nf;�d,(J]]`rZ{�-��X5O	���͡�O��z��aV����/��D��2��v[�Q`���Զ�-�!
^:��w(# �M1V��H�v�ۨ��6&�Ǖ�([���Ռ��y��@CE)�ѕ��+�f[��I�Ԩ��|���V�bKZ��m���_��d��������������.�0��� %���|��X����΄H|L)��TR��C2ӲS}�d�=�2�B+^$���kG���p��w�f�t	���%���}���c?J�Ħֵ�P�,��g["՘�ʖ��k������bڼ��1:.C~I 4�#lƑ�`�|��x�e[�S� Da����2�����Ta�$��I�kF� QŃeǳ�M���%K}*,�ްv�iUV���j�Ix[c�~ޫ�`5��2˹N�L"�)�l;i*�d��ɚ���:/))� j��Q4�
��{H	%J�zӻP�$��H������p�s��,���;��B�I|���������������$�h�[���ӵou;��t�<�/���8J[�ĕ�2��˚S�t�98�O6gX�#�D�%3��qa�����|������ϝ˿OI�7��S��m���	�j��4Y���3� �h��"Q���a������,[L�S���Z��4	B��S��uSz��c�x���]��U�B�}��|��4&�-0m���diREu6��%9v ��Qd �3�F!D?@�����XF���h����=+kXq��� �r �0��@�.����yb�p��������x�Lܸ'�N|O�XRC�>0-��ӈ�+W�6�tU�	�3b�5jp�W�e
<�C7�1_���d������� ��Q�P�ܢ��ڟ���D���=_�>L����.�Rc`1�°)��0�zf"'Ru��Ԛqfl�N����(Z���@��t��ɦ���KI��R����$	�Y[��J��3��Jeo$#ZC;��g��?&~������4��g�x�V��وH�rs�\��	��P�I�(n����݄����,��Xި���τ��?-�C$CyeI�3-�y��0'ê��A1�Xzҋ'��\�aop<TC�>_�"��V{��@ˠ�;x�M+�,��}X����Z��)F��S���vL�E�|��qb�e�����'�����X0XƇ)^�s�����cv�U?U2��%h�Q	�O�OWo;�?�5��Y�?BmD	v�~�E��1���G�Po��ު��St��B�9]?�?�۴okf1���Bi���g�A�S���<��0�72�4Ӥ��"E��=6I�9���S\��x�e/	��g���Rk�_����<�	�XX_��V��[\o!d�,hCs�"�6zM�B�@�1Цw��"J�,]�I�§c��]�n�il)AڢԆ��v����߬[��1���˖���>������L%&\�o���*�#��┮�@�N1����;<�pI�C� )��6h����$�0�LЏ�9˦`�(������B�����:Ս��J�����}�W�iV-�uܒ8W#��)��N���A9cBUZr2�7�5�=�5A�=]�\�/3�I䈱��Fl���z9R���Z7�%~��=�N��Rb�F���O|X�E�E,��t:p��a��\2�R���Ù�AL���ֻ>1{��㘾ˤ�"�\s�Hm�4�gZ�`�Af!�2&�n,�>��T	�.��.p�6��,�.�OjO��f��t�ab���S6!�I��O�f�h��J6�2��vK������-֕`^
��(���1�3	����,��Q7{�m��^W��<6��O~�����݋{
_��t��Af�r6?�K�{~��HwC c$�gq��l�\�Z�/5.Ͷ���[�.#��������l�i��	��ǂ�����c�ճ4�������W�ªHSKXk��O%�F�&CH��+��{�CÐ�:J��؅$ �*���j�p��ѦӁ�g�֓M�ą��V{�ن\�Y�e;����;�Q�p/t��p�F��vf�`H̄Ĭ�RC���Ώϡ��c�J��J=��630�K3ҽ�X'k�gE��yiɌ��:D��� Ӑ=����G��?R����[1`'{����%�9�f�R��=��
)�?�WCm��Bo�3T*��C��K��T'���MhK|K�=�}p���m�X.���_ ��B�MstJ�������HP�EyCx�VP䞐�1,?s����@�,�[��q�54:�X�d��!�m@ɯ��Aa7��2�@>��2�RG����4�p�Hv�鲵�V�w���*�� Mk�f��T.�.cs�O�Ƭ��	y��8��.��jk(���Bv}��ɓ,��x��"-����l�_KL��Y�����ؚ����m�Vm�m_H@Htb ��k��#&6Ɂ��Ø5�^��w!�����w�'<ϐ���1u��1�IҶ��b�[� 6�q�Ӱ��w=_��s��w�=|\��]���=^H�Z ���ǩ 3����"����Z0Ρ����"���/��`��\Q�) 6T��'V���I'"��0+m{��/�+g{M�9�W=�_2��/�j�=:G��-z�v�����$�&}�տ#-��plt s��XY�;#�n�Ҥ�.O��|\6Dj�6��l �����2����,6g�Z��ZFR� m(�y�<�B9*7��)|&���i����9V�ԒTF��]�H��z%��gUc�r⍒T�z�ɼ��oh�
�~n�� ^�s������Ҝe#��wo�(�
��&m����0Zi�b���|D��[��A���M��d��0�������X)�U��V�'�~�<�^�wޡ)��+~�?weA���p1���;d㴫ޢ���v�����@p.�
(�n筇��
����ـf�+G]R2&R�/��-	U�s ���nÂ�s-�=T[�qM#�i�2���Z����f�z4kp%φ9,ɡc*���~����#�ex����Xa�̯�D.t�v�CL�����L��ǑXScz��$Sv �KyT@�������gV�2,z_����i��i�R}��
[���>���U_�^@}�LB}2ͥ8kHCäc޵�^�eMQɋ
����6�M��aj�/vye@�٠�^/�9��ݼB�#�H���B.	�ګ k@`z���-39�H�d���)s�����NQ�t����v���\��Ҙ�ߴ�X��ԁ�1��Ŵ
��r��"��m��y�Rq�k�|�?�}7U�D�a�"ɛf�\�RR���^b[7\�z��iX~�B[ߴx˗�B��yD&,�כ�8#��Ta�<"�6�<�m�cg4����4u�>ZU;����<B���/��H�Hw_��$2�s���.ǢK����p�YpT��"[/�&���C�[�8��S���,g������pU�.�E��G���!�S����N|��b3�lp��譿��־dT8{2=#Y�<a��A��)�."~���VhVë��I8�7�̉�d���Yv���0oj�Id���sD��dO>Ԧ3�x.SQ��E1�����\\oͿ��fH���� [MW���ї4v���*+aq�0�!��tw��ߦ��ߘv�������H�*�1.P������gb�0M��Tj� �?۵�jkU�U��-����;}��o�# �'��pw�<'���_KD�d�y+�11�3��`�ߺޠ������iOKJ5�����.VT>�u.ظ�rÿ�6���p�O
T�!�6��ޥM���&�)%�F��e -��0*7U#0��/)s�P;5?{|-�ɮi��?�� ���)���/����� ֆ7���f����-`"T?<)l�l��HVR��kit��p�v�6Z}n[r�'�ڕ6�A�O���[�*!t4��m
ͮ��?���;'�ֆ�B^N�����+�BJ�T{��<��ܢrz�1q�\�<��5�껌��9.�dY.�&���"��Z�7Ş��)��A��*��<Q휜V:�׸ u@9X1��/��/�p�hfA��ij�O#��Q��3Ҍvc����ƛ�s�A���i�׵������ 5P�4J��{��ㅜ"���$�Z��i`O��St��܌�Ps�$i=�:������N�;���bW=-��8k�c����ת��_��]ݛ溉
�J|E~�H���:QCgD�%�	��@og�(�����}Z�a׈��M,�"3�_��67e�J���D3�)O!hUQ�
dr��,jz�A�ت���:А�A��}P5u|�Z��=�c�X�(�˲�����F�_���#X��ߎ�>��9�Ҩ�/�'�����h�����j]a�[X{X�и:$���R?�UЃ�|��	dؿ����%J*
GBъ�n����#�����Śr�ţ���,]�r��L�Nf�#�r�o�rߚ5<��FcG�1Q��h)���ƨ6t�3���k��R�m&�Fj�-��L5�(�Ji��O6�b�)���~֜vH�}}��(��� �`�����O8���� ��%�u��c+�pւ,�V�[��6Z��=\�����e�N�4��O@
�=H�QW������S��˪�m�N�v����*B�w�0�Am`>A��GܶP2�)��]`$T8p�e����u�\d��{/kj�s�[T�)GD�[�Xa{!x#���/o��G��]A��1��N�Fbp�e�@S+*Ώ�rl[CR~4���4�y!�i~|��Yw�O��L��j@\�`�3��ټ!3ͻ�f�?�
�9.YA�@'IH�"��n���1!�<��J��)�vt�}�R�,�|����$nfR5�D����2.�C����Q�:���c�;~�q@��GZ���ф