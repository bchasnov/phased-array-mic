��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�]��Xȭ��p�oȡ�;u0ީ�^�)�>vys���2{�L�~|c_Iy�K����-��9!��\�Bi�D��{�Ԣ��r'T��NjH��ဣ]��9��|p���4dտf+����ؐ��7&Qa�z���m�ࠧ��3`����8s�=L��4�S���J�7�h��J�3�_�������p�t_3�ѹY��S�!����_-)�_�3s&_.��������
��������r� ��+$E��J<�Ӳ;�Q)Fu��7��yʋ�C�eTc��l�jh��o6������C�#"��W������~Z�^��3��p�(� 0+���o_��?�����L"Q9or�����;������� �IYlPn�ˡ0���Z�9O��.e�IY�8��ˉhQ��?���hb��u*�`xM��
�F� x���t"I�%n�� ��}������,0MA5y��3Q�XI�����~ɻ�-9�VBz�	������D��B�1Bwr���um�4�4n������q����#�ϖ��P�`��s���O��6��X�0��F��4������.�[�9H�� ֌���K�/Ti��A��G'��0��@��*���Ϳ��B'���p��s\����;MT�>�uA���'�Hj����TAc�׈*[D�!!��|�6I��|�y(Z^��$��y���h���פ�ֶ�"h�\o�_�S�ހ�K�-, 6ݴd��X���;������2��)��슛���h�e�ff�'�D�|���v����(`u[��e�ϻ�T`��cx^+��_I�S/�*�q�P�Z����ܗ����S��(��gd׽�&��P�we��@�{�>sVJc���A���.�(-p2�ܵoN��=%�=��ę"�D������������wg��������b�T����!?�k�%��G
;c�=F��o�� ҰT�n��b���3���� S��_��x���<��Q&+n��y-Xc`;�җI�a %����M;�T�/��+O$�T�|���԰"]��[K,�����$v	9�\d�|�s�0O]���0c|�9�b|��"�xU��]R)�@b\�a�e�����}f�^�눝G�]��@5o��ɔ'r���C98-
�þ��V��������0i���`	=)V^�t�'hL��ԑ� e��^ʕ��|{�UY���ěm�x�X<�=��
�Rj��V����Pl�}p����>Z(t#G�I�g��o#H>:����,�|zN=�^��aHw�b?Q�0�Y�0|e�%��u�坜�j���U*f�g��O��7K�t�ݸĐ����cI)㵗��o[�H�C�_+����b˳��.�d�8U��k`�j�U�Yg���¸$�~e�9޵��iҎ�-u�.b����O_�_�؝%�_-S7/���M�3i��yz��*���إ�Ȗ@�G�*z_p=6ٰ���H���	�wf6��mH��h[Ȓ�o��1�U��� I�T��|�1.�סt�}��{�RcǽFH!�d� �x�I��:ޙ8q.J�
��~��g8� ���Z�h���
\�ٰ&H8S��C1��� z;A��;P���:�����U���FB�.F2መ�N!�|͜�x�	!��JV֜�cw��.͍�YHxJ��e7W�j�eW�ǔ��ʻ/��+���7�.��{�~{�B!ഗpĭw(�)Z��bX���5���D��&d�y�ؒOcfF��I�fn�;]���5�7�2�0��'Bӵ�{���+^]�M�O�݃���+H�ó=0�߆��X��0���rg��;��{��^��k�;�4(�U�d�T��1&�OAjY���(o�V����?F-�\wkGeY?x(��a�.g�*����'ޢw����XZY�a-���쯿s1��}�5�\NLO_0g�ٔ��gu��0<O[��}�hB����p� P�K�D E'4 ����z��=huvB"�p��<Z����b��J�H^8KT����ɔ�J��Y�W�XBWS�HK��r�	���	8��v�+�ao98lk�8�u|Q��U
9���eg�����80
���W'��= ��!0��rEH%�:���i�(^c��xU��	Rx-"V:t�P5!��I^9��^��Łv���33O�I� \c+��`$�&��2��A���K,�)n�$�����oV�Sm)t��W���X�e��*b�й��J0Y\R�TL�03޷Q�/ �h|M"Y�&���O�º��M~2I�;N�����u��Q.FN�P(�����އ��cQ��ϲ��~g�o���l��W��ArϜ����T�J�8f6P.�}K�sg(��p�!�t����־�I��%G�R\��r�����L��=Uq�I�u�i���G�l�$̷���ԉ�u��i=2o�����@��>�˳�}C�0��KN���pt�>�x4�G��#V��[K�/p�"��+W;�)+�3�#0�'85h=	�zE�ohon�-��� ���W�82N�p�e�[/6������cA\�F5��S��V�-�e)N^I	�8�F�rTu<�ڿ����c��c���ۂ 0�N�4����h� �2�i��k�;���]���j����c�=��C����qם�m$�?��Gy�|���g3Eq6�RwAui{�Ft���!���c�ԜeN� *>�[��Җ\������r�N�)8������.\�&��m�uJ%�S�N��4�]�(;�!�5Q�hZ�iJ�G�����Bۑ���Θ��|w��9�\D ��>K�EE:@���6�Ag���<���X�G)��@�V��V7�2J�"q��w�R�FAM�(_�`)�g��{�JY@HJ���'����C��fe�U��r�A�qwD���� 9�9`��_T����b�ԹM�����q�_c�'GE��Ȏ�`J�a��e�->n�./)X���F.7�h��II#ޑ>�o�%��Mv�������W7���p�Q�@�6�TBs�x��$�'r#~�(��b�'.�z�ϐ���^��L��ZƱ��	K��|���9����_�����-|�k��l%��-k�����N�m�J�ￜ<��_�X�/	��S��W�q^7�2ALw�������x��>�E!>��(Q�_fK�S��Ox��55�%�����D?���� �9P.KM/'[ёJs]�i����-3$9� �rnw@�c�N`��X�8��_�=���o��#g.Ui81�hMt38d�������;�[u��;,��Tߋ$�Ns��΁W�(1IS���� 謞~��:���1>������r�z��*?�0�<�ʽ�ɑ���?  $%�¡����9掄B�ǟf���/q��vA���L�: :=�O�_�� �Ҙ9��8 (m��?���7WbZ"z�����F�xqVý���	C�moM��gN)���-�����u
Nv��'	.�ȎD�**��?��Ux��ph���ppH��NUn�,��hHj�SQ�t
y`�'�M�Yb��<s9��$�s������Ϳ���(M� >�Γ(a`�w���]ԇbt�.1��'@�Zs�%[�2�0_� �|��c�۞N�&q ���'S�Ǚ�Wݫ�cz��5YuenϻN��o�ІA澱���o�J?Q�HF�/F���\%��ٮ%�%���Z4D6"L�a��n�?{��-U�|�Q���,�^�f��I�����(2i��R��L��z�S�P$�(U���K���~�r�p*�԰���%}�"D6�!��9��U�\5�GwU��`23Z_HȄ�!J�
��� �J�@7>ɂ鈽ϴ��M"���  gu�?��B�Ʈ-Jq�Nڔ[L�S�t�%jʟ~v� ���K׾��y����ΤR��ͺ9��v2uG�Sz�a�UG/O�[7��^R;�:a�yfџǥ�`�L��ڀ�Hhn�o��;��E$�k#o�L��Q7�RWᅟy�v0�\�`�hv0��"�I�(ԢȲN��'Y'�t�Þ��Zα��7UI�i6r+ގ��ݓb뉜�{���=�L��v�M���z��mZ\��.�,��i;�-��P=���A�}C)gL�x�@�O�bk6�G	p��xRFm���*1�yw��ң�ٓe�%5uIJ��7)G��K��}�O*	p��P#�s]��+�������9�bޔ�'Q 卩��`���L}�����.���<���m�
���Z"ragO��q�!�]ÕB���GE;�8p���D���h��GE�> �����ܽ�(9�h�M�!VA����UMH����N�I��)5�3(���D&������)��'G��2����}��������W�"﵌v�P{9��O o �ʞ�WikN�~/w����X �Y9p�,"�K��<�SI��qj<xH���K�o�}����� 磥���*wGNS<%����/�e��6����XNKd_u��cD�C<5j7��� ½a}�fse᝜b��g�2|/$t"��u��ݲ]5h�8DH-�E[w�'DG!�=0�$q�����;E,���?*�qj�oêy���v��(�%,��HHT_���z3?9%��t�a���G�u�hY�E�s��q�g/(_�>�ҭ�:fQ<q�kDK���ڲ{K�E�SN�Oa�
�B�LH�鶲�`�����)ӣQ���2��*X���,/�f��0	 ����5�v
��6�K�lݛ��9�#�� ��  3�a0QRo�C~�Uϖw$���\*E�5G@� ?�n��<7�7È��R[�\�rj�����: