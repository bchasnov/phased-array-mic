��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>b��z�P{��|5-`����'\��}Ho��ns>e�:!7�ѹ�A���9	�g5#�=�K�8:���!���"l�!���r0W!�l�%��J�Gk��[H�+��kOa��dI�x�\��Yq]GDX׻<��ڸ~��;�G�	����v���,v���V7�m11��Z���X_�w���9�hVE�Qn�#��f~Ѱ���^��D�$e�F^zfkhQ6�TƀU���Sfv��&_X́��\h����<a�6H����<-�Aq���$�UO��Q�}S�v�[�	��j޲��!|_�5+	����~���ؗ�P�m��R�^���ᰪ�a�-��D'R��3�F��E�RK�>�܆F�p��l� �4�w; �d��1Bv�sn�\s�JU��xJ��o���!b��_<����� }^p��/��f2���b�~���e}����W��3��QeT��Ykǵ�����T����v�!Zt�9����ax.��I��P���F� ���MU�5%N�����+�O�f�].��ɣ]o]�$�ɺ?��$��%OI)�+�#P���w�i��%@@���3?���oh����V^��U�����R��v����$h@H������*�A'?	�@��%Φ�&�N��C�,�^��*h$u��14�k����oМ��m�n�Dk ���d�i��̖@	~ρs�[�U�"ĥ�|2����5cxX
��wZf$�s%���YY�
x����CKi~;D�t&���JC5�!GU�+��ɂ3�#�i��t�
�5���C�@�ҳN+7�o�} ���d?�[#/��JhQ�����D�������M�����Lۄ�v
k�� ��!8vM�Aڐ�x,e|���Z�d�$�{%�W������k�q��L�Uz*'M;�
��x�|��4����C��դ�KE�������)�%��<�1I�-*]��s��h�a�$�5������I�1��"��&��4p�G�J۟��a���ܛ�T��'��g���ݦ=�^��3Y����9\5��f�#	���y��r*��c�.�CB7>88�'�+�^���5����+Vq�47^-Fc��A4�a[G#��<����ՊL�����!�|�\�0�F'���tγ�N���L��2����ޛfcw��c��98I�0���m0ɩ�T���i���!�vxn8u@���Lݰ�[�K�
$��9�e� pl�v0�W�\���&�~�oe�B�}[?���s��S��C�I���q��5�5������%<Ҋ�>M�����D�S���4�
�Le9&6�Y5��m,˯èm�(�Y�4ؗqʳż�g,`�ːD�w�c�<JD^�Q��'��ñ骳��&T�#Cb�R`�|�Uʲ�q�\D�!A����D����"�v�%_����C�l$�Jc����
,eD&Q�b��|�U!P�N'N��YST%_�� T����9��dl�+/�-<��9���A9��|�.ZB�����^�E�f�o�b�9���휍V���T@
M�5�8�Y[�N�[{�����[w����qW�^j%�4K�i>�G|n�yb�����XɁ��� z�^a1�D܉�ȲJ��SiM�6�͌�P:Iyo��>��(W�w�)ӌB.UqW/J#;�V|����S�>TRa=�����C�,䃆S2��_�y���0��w%�3�B��S*���cY�˾R��]��5E��|�f����y�8h���[1�%��5R"�p�y1�]���*D[��kuK��ֲ��w��r�C�|�h��G�c$������_b�[��N`v�(V_��H}���/��Z�V�~+`�_���ODЋ;0��9G��{Y��g��w�s"�-�
w�d����Ѯ��%f)�_ ��I�S�դ��	ڰaв�P�U&��a��ԅ�^�z��RȒ5���]�J����k�I���4$���)�)S��K�+
��"?���Ǝ���dWcĐ��*�!�De��G�̾��2.�Ȧ7�N�f]᛻rYc�o�Ɩ���15mu�i%�Ԏ��� ��g��l��_��T����+8t������i��'�I4��Oq�H$-�'d�;?�lh�C�Y854�h�a�,��}���m�
H���3���\��ߟ�����D��t��N�ܑ�S��.��:�!�̋g1�;7|���R&j��m��@o{�М��[��Lw�w�~B���aX��n�u�"���@���RdVvm?�4��٩.(���0�QCu�Ys���ډ���W�k+�UǏ�T��Zid�gQ�;I~2ih�6V<S��[� ���|`�ct��v�g��]�Zz���������=M�$"��Λ�<}��,r��M��FnM RKۄM�++���'�,�q@�>�k�OU���:nm����a,��:]}+i���K���J��Bc�*-[Q<6Y���O�VX�G�;���Z���LVJ?���|���7;f�Ym\��8Xzi�v�ƫe���'�s쁤�`�A�wf����	�ݱ~$G8ZW�b��V"mW�p�t��6��G1SO�̭ס|�ʨ����TO-�g�RBR���g/���S�Tf�j�Ɛ��8���Z�0�����@��Kd��m�CF'�QI�q��C���>Y�%�u�۪���dQ12)l�	}/�\$�`Rz�+\�~�t����Y�)�͹2�foԬoP9ڷ��j�}���V|���&��̽z�o���k�Cj$2}��+���rn����_�&�� �~�
A�eJF��7��#��?`'C�Jo�J&%�U�v��lv�~0�Zۃ�3���o��נb�Y�[��&*���#��I)Z��>zG5y��ƎS3��O�Ǐ#:�p?�r�ck�W�]�ȼ%�H��M��2��:+��  �A����A�s�m�G��u��~���y�0�\-�1S�[�$?"6mܱ����ysA�D࿾w�$P-���i�`���-Ӡ$�23fH�	��A����3����sz��4�I��/Z���^*a�ϊ�L�P����@7�éjN��r�I���y�I�!����!A���C�_���*�b�����Z	Z�->�M���Y.�+o'�Ḩ�e�}�N�d�-���i�\W�qp�wUs��y��~@���������mx/\^X�e�t�z)���?���H��� _�@��myV����j$��"&�1X��J8�B��o�/�tB�a^~P�{Җ�.w�lQ�\u�v	�!�0q��_��D�ċ��&ֿ]%�	���ԨhR�L�ŉzsm��*�\���7�A~3�po�u �OG�6ە@�a���GO��gڠ`O��;l�u��?�M,Ρ� �)\��ݣ�O�B���"�I#z	]2�I0ݺw���y}��l"1��|1܎�Ča�|��D'����^��ͷ�篒Hv�&{	�P�/�B��\�T��vq΢~�����'.��=<�H�ؑ�h��{��x{�Ts����eNUN���;e�t�.�!�ul�+R�8��Vhvm1�h�-��1B�C�]g��mx8���W���`,s`B��۠v��HskY�7V�.����F��l�nO	����6$��; �5�����)�/7W=e�b#ɬ�zl��W�2�ƻ�W��o��r���E*���o���/Z��z���0�y��� ��UMv��l?g���ZʌrX=�yQk�������7�M�.�e�/�VKK��㘢d��X��k@��y�"��*�%��A��.������Ύ�G�Z�Xǻl�~`Kr���cfI�ڗX�l:#0<�Ph�U䟱�X��4�B���`+�u�Q�'4C�:N	������{8H�zl+1�2E~���Ĉ���>;#EU����v�5C�!������?7��=���i��$K2�?�i��ȣ6�8����Q1C=���k� ʌ�"�Օ�6QA��I���쪀�(S���ʯYâ�����1���۸�� �ԧ���Y�(Ѧ�����հ�i��š�=�T����8hl�� xۓ���k����8�f�]��E���Ȯ*�Z VBz�c��p�A�Xe0�g��n�X��$�mn�"��G�"��J�u���m FE�7D5m�n�����E~L���U�!Z�F���t����p����|�_����{U�-��cZz m�W?�4~i*O�����C�>\_u���߰��u}e�Uk�i�vW�%�X�H\=#���GYء���ctH��rMSΡ�^z��ȳ�D�tƏ��%XG<J��l�~a������B	[�]=�/*b����(R�V��f?�ן����S�nN�D����k\Ѭ���V�'��ҝ� �m�4BJe��4�Ց��MG�]�B~t����H�x��p�blF�Uk�h�T�����G�ӏ,` ���\������6r�`��/�� ��)���E珊��%fwߔFG�2�?ۚ�>�T�'�Ez;�T����Ft�#�0�&i�K�ﲞ����DS:���X_o����y�
��IA	�֥��VD:5GW.C�Œ�l��4��N��u��3Bw�����W)�͢��/p�������D��k����i���.|�D&N[;WiJ������u0���� �s8X��A�C�v���ARM*����H�O�X��0��+F#3{Z誖�>A���#_
"[�S��˗���x }��Va�U8q��|�I~�W���F�q���7h񙿽�#}��+�d�|}Ti�8L���xh�f=c+��F'�!p���<�լ���\���k�&�&�Yo�fg2*wh�AI��k�G�@����y��B�������Miޔo����/{ȅw	���D��TQ���5��w'7����b:ւ�
g�[�d]���Be�l��ܙ�f��z��1VR1c ���x(�7�v��r�&����\1�=K����M���87Ĩ!���zK-�FM��&���'~���r:�揖ðN	�EPNjb��֠��Si�)2Py*�}%��]g�M���򙙹#ؔ���[�nm@�C�)!��z��629���|���N`���!�$0QpwO:��O�6���nƝ��/�z�#�Kk*�O)�w�B-�~Ѽ[K�=H��.B�B��V2i����h+\���d*FO�L:s��T��m��d���
���G���@j�҉�y�����=.����؈��(5R���d�-��\��>{��8vVJ��(�!O�v������g?}8L�����;�D�ft�	�K&�E�p`.p$mX7�,ɯ���ݑ�3�Ő8�ȬON	l�I6o��M�����
S9D� ���Ґ�@��Ș��Yt"�q"�Wy��dl!hH[a+ S3�6$Z��IJ��R@��՞��.�ko�zN���5��}�v�dX)�7k(�f�Ġ���:oX/4h�B�J9�携g1��<ޣ������B��;�n����F{������ge���Ilܭ>��|�_	鑨�dE��`-�*~����m0�t��!pGf�O�Z��ӂ��K��j&G3³ޅPR�>:��v�E��t?�|8db���uS>-!1{�(��?~�a޳��>��It��������i�g
d%JI�Dt�X�ߓquRf����F��̬Zt���@� O�ĸ�����y9&e�z���/����y��L�Dl��{I��1E�Ij�E���ڛ�̮�s�cP�	h����Jm���c�n�s���b�Ӥ�4�'�ea��B�//����P�l���-+�I���L�)C<���/��^+Vsc�m����`����[�r�/���q΄�I�Xݵ�:�N�P�$���r�q��a���U���-� t�ε���v�ʥŰCtk��~f�p����Y���\�����M!twe���W��H�)2�Pׯ�T�����u��>-Av�9脨g�6�!1bA\^�L���&R���c�f
<�;	�S:�4>�S�W�qB�b�߇cӐ;N�F�<�qP��gIB��H��6Sx��@'L�T�{�����gE�H�-b+�.�ٳ���
�A���v�u��K/}W,�מ�g�[r�m[�l�e�����zu��bgfD�.Mm<&Nr%�}�Cl�gNo- W��s�M�8���L�!?ɢ�&��pl���)X*-r��.c��q�6^�Um8�f�o0�]�&�qq�v玲-�:h���od��r|��z�U�'缂w@�w�)}aSU�p�!����a(�ga#P�Y���b(��Zy�JP�ET��DϷ�+��>M�!8��nbiWu�#�(/��~��#�'����K��ϼe)VA�h�Gލ?G�����