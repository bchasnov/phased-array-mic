��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1���e}ʲ��cg�t�ϙ�a�:�KR�%���ݧw���ȼb��{��2Hr�Wr�����B�����?��Z�8� ���x�
���M�����(��x0�E�v,�t ����e�O�~S�y_��t(@�:�_A�o�AR�'W�My󤣠ˈ�Z�#�}�X��*$���TA����2�M�!��_��6�z�V'�72_�F�|�L��ְ�+�N��CG�;B�-�nSߔ��	kW�4���7��e=s =�}�l�ĥyN-\>��쩂�&�䛙f�JW1��R#A���fg��In[*�����WxMU=� !c����P�"���VE[��*�b��7+�8@I��F�	��K���`%L��bv�?Z�>��$�,�.��'_�|���d����lz�����mD1�L�ެ�1`M���3�)��i_Q4ѵş41Fs�Y/@���"(�i=����|��yyv�r>Ţ`���.��7�'�Y������x�sLR�3,҂y��6[�Z�*pǡ�%m&A=��dן3�Rè���(�̻�W����bȻ���E�p�*|=�(vF�R:~�V-��A3^�6���t����������ܦ�#���~�������G1YH��{?��X�A����t��dJ<*}"Ř�$�E3ߋo]	#��D������Uh�f�\wb�ݶ� ;��'�e�RQ��'�{	�0*v\a�q-v��l�k�Pp�4�ޓ8�� �!k� P'�1k�'�7+Q�DFV-��2�2�.�Lt�=�4{i��� u�n���x��+_;��%Z�ЃU7A�Gї=�����)�F$+L�8i���y��u��N��Y^%�k��n�>��p5r�������C�cN�D�+'Ym�vO�	��e������kr!tΥk�'8���KȔ܂���Y�zV���9�Fl�9/<��ܟ+�
�S���.V�ӆ�zX�E�e�96w�X�o�A��e�/y�į��Nu@��1ʿ��7(z�n�ﭡs3�U��R��c^Y� XԘL��iI?�v���4����@$��B�ϥ�A���
��LX�P?��:��/���u�|Z�g���H,�#>�)���۟HY�6]����Sgv��kݷ�ВZ��D:M'ɜ��\RSӁ&-�T���<o�jj�"���ĉ�M��x�p����_����@�{��M��2r�W�V��~�����O��zG�D��z�ZK��S�=o\�������P�0�q/tI�1�J�lv�ƙ���p�o�"3�5��(N����}����z������OJ���d���Zd��Y8v����J�\'�uqH��6^g�g��l�-��2���(<�O ���h�J��Yv[��䒦���������7CE�#�!M��!)>�18�z<M*�A��7z��5@��V��5]��n�܆�����us�B���M��nא!�A!��1��W��q��k�̂>x���F�ƚN�]�-����-�c����:h\�p��ǩ��0�,�{�ڪaW\� B*���i�WQ�FM�s ��Ð�]���u�����_����вꆇk`�l�@T�j1��A�����YL�{I��*��E��YGL4�X<��0��{��p�X��ϫ�vD-���KOZ��噀z!.��F(ڢN�B��tp�O,�iR�E�C���S<�e�Л�=��LSV>1hNK�]�h��փL�%�eǜ���tʂ)��*4����j7��R�Fus9���A�!�&��AKO���9����/���>=�f�[2��w�y��9�o��-=�Īh�tܮ~M`��o�#�Zk(sPG�$g@�;�=&�ދ�2&%��&ND^��;�MDX�[j���=��D����?0������~r|�J�w��N� �}�������A�rTG5IX/T�B��T�q��ϫ �{�e:�5&6WA�{�vѧ=�Z��v�s�j�|�s�*��D=�)�(v�㤈�ƋҜx�A�.D#��**��?��p��O��1H�PIڭ?���#=a�����(E������*,w���35�.Y�J<�6f�P+L	�8���(MG6d�QT��Y<�Cዾ
�O]�~�*q!��-ܛKFw$�i�Jѭ ,w<ˋ_���#��ѼJ0p@xx��V�1�e{�xFw޺�MH����2�2�P���n�SF<�uD ����������m7�Y+*�����3vv: ֒?i��'ĕG����v���J��s��;|�(.3�^��%="��_9A:�x�
�|�2��݅�Q^�E�ʿ�[���l:]�����i�K�ȝ�_<��3ĳNWv��\�7=j���ʬ!�	O3��2�Z}�����f��=�Qw����<��� թv�-���;r�?�p,�$�G����l� ƒ�M(nJȺ��h,.��$����*dӤ�l�ܭԱ ˰��y�P���g�	�O�W�玜�R�?ٓ�LU��c
Y�)�d�D��P�U�kRE8ln���߆=�|���q�.K��.!�DP��P�g񁀧���H���&�dC�yS8�	3�#�̒V�$��˙��sHhQ���B��<�j��Q9���U�S0������+*�6���"��!�n�~�&I�ٍԟ5c9�BMpΟ�+[x��k_��3�|7��ۮlj��E����;k�(�h%�z|�Ǜ@�QK�����,]'Q�I7;frJ�ɭV8����?��\tK���M�h�.s����X��2�
�"���>0�
��W��3<�� �$ ��n?�D�>�m��]��()�)2k���y\���_]K�� `�3����k�=~�6fD1�u��|�=����R+Ԥ���Q"ބ2�dG�oiXo�����J��ʢ=��rkQ!ڳ��������P��G�V��z��e �0h&�AW�$jj>�{����"=��V�@��F�H�LX/�7�>&jü���ה2��B?�pPy_�E�7l���7B�!��Q��q_����bV�*��$�DI�dJ,��V����x���6,r1n������~���lI���*�C�Ĕ>E_�����b<-ϙ`nX���ܷ=uv������3"r������N���gZ�=�0!������M����}��Y �2(  �����'�ؤ�]e����]f�c��C52dW;��yLK*�M����
���l��8pu`7o[8�l���۷܎������l�V��@?'Dv�H~ڤ����ח�b���$|� C����@���ň �˄��uo"�X�b�e�_��8�K�q��p������ ��P�(�����Qe��#�A��:���W��V{����իF�� =��4� �Ƿ=]ُM�OD����p�-�LC�ݍ���Fc��3.Ӻ����#�'��{�� �;(��v���2}����U�#�a@
\�Q,�ŭ^���c�~��C��Ao�$oy ��y�vp��fҋC �m7�l�a�s���1KHkHw9Μ.�WNcƥ�T7�es��FA+F��Wɗ�w��R#��|ɥ����O�N���>�/qjP[o����r3�6���X��#H��kbhnz��f����W�4j�J16�	�����tern��^PdWm��
�	��YF%�I*��D�!�i!-.Y#J��n�������(MҌ4��Lze�b�v?WO�&���V��dˆ�dlfyX	�R)�/q@�xY��mM)�.�1�L;�f�:��	�������ɣ)� �l䝖�� ������E�|V9Y���\��Y�|���h/��v����N1\�¯q|Oy�Wڬg��������@D�X��B;��Lr�$����|ҁ3!�%Ԯ���6/3Rc֠���%��>�a)�@5�I�x�MԺ+�+d�A�s�n^��or��#3>u|���f@�4�c٣���=��߀�؄��s��܎ه7E����V�nj0���h�\�d��H�&�T���A�Q��o�J_�][U{c�m��}�!�n��2�b���R�`ML��K���l��� �vu�%Oڳ�X�Qe�%����v��Rj�8�qWR�u����3។�i�.*�L�o��/�;���{����o�Y�V�Fd������#7R/��q���\
ZSJ�-�RG�{��+t��xߒ�Ŝg��@Nkڋ~��U�U�,������k(�nBE��Bǩˤ�IA@�cuAx�	"�����G`���
�ʸl�j#f��&I��}��Bd=�_̓��A�Ɉ�u1�h�7t�j�"y]���;3�����[���G��X�3��#L�:��~з�o��a+��	i�o��[!���p�m l��n���t��i������EarH��F3Y��srV<� 3x��5�{65ߌM�,Bc_5(1:rT_j==6MGN��P"���<6O{�	�ȶ$f`8gW2���D���Y��i�w^|��C1�8��C�׍Vf��^`�5ئ'�V���&XYq���;���k�ל����[��w�/�lo�ν��ASÿٺ��&�2���c�b�O$�P�I�l�-J��:��{ud��n�0�(�����x�-r�Ό�Z�i���N��^���Ǳ�g'և�{O�[yv��/���,�{�B۰��D�l��S��K�N`ȳ0~��p�y�P��f2�aX�Sf2��K��Rm�W�?q&�y�痤h�-Q_7���F�p��������bU���ƹ�Fo��,3�Gl�+ď�f����!4�~�U�s&�T?���3�?��=/��{��H�s׉{6Q|e��F"�1SN�Q\*ح�7��[�7�nQ��j�����n��M����^*� ������]��<�?J�#-#K��Z>1�i�����	F�'����6Z��9
LJ��Qv�^���Y������5��u|x�}:�0�?<�C#�4��J�����0;�N���
\E�A��*r{qX;M�%��9,'��-���HR��U�80�:��Z��1%��=��� #�X��9z�'|ތұ����@J�������]G�6,�G��*5MY��s��d�;�Ks�����.�뒶_�9�U
��}`*l{o&�!��A�H��'��[#�~�+<��>9�W�BG������m��Ѫ��[I�;�"[$�G��FG �ȥ���_J��*(��#��k�^x�ȸX������n�!!`���]�U��}a�.�k�iS\�8
{� S�e�*6qe�#V��H��R��
X���U�my���&a���c�������2�˳�@4���I�z���]HI�`ܗ�-�8�T\�������*©R�0+��ԍ`�\�Y�U)9	��Z�0	�6`��u���3!�t� �R��25k><���FGpӖ#}űN�5�+���/��C�*�7٧�
� ��1Lh]��o�q��:&Θׄ��zݷJ�"�](�2Jq�/G��[��A|Dϭ��"V7�F����>�$=Є�@�RFҵo�M�ߔ��������E�A_*:x��p&�֜}Ҕ�'�ߝ�7��[P��>�ӓ?5�=Y!���g�1|ߩ���Zd<N�B�7�ݏ�j�d��:AYa��#�`�oW�S��J;l�%�P���?d8̊p� H}�郰��;�*�V�Y������� l?r/�[Sl��(�����~�0���.*�e�A����(	?����Ҡ��}�Ff���r;��h‴>�����s�����>=�ɞu��rmz{ ��������)���$x]�G}�]���Z+Z��==O	��-�˩�g�(�\w<%v���f_c>��Uİ��R~��>_�� �݄t�i#^��f�����򙑦~د��%����'b �<��tpփ����(�.�nTf�|�J2k��p�8�p�%	XIB��
�I���+��ѱ���{�L6E)Q�l�w���M�Z"�z'\Q#�28K�����H2��oQ�5W�5������J�X%�U��T�SHE��SNGy*,ؕ�"X<~Dc3Ք�7�-[ox����ƫ��-?�(��ht�#�42��+j	GA� �0;�����6������~����lU� Ww ������LK�9!4<�TUҕwt�:����J����۸nMW,zaH��E	�	`�o���O�x7�{$���ݲ���v�A�0���o�<��>B��%���
�y$v����)8����2Bh���U�Kt1\���[��`���X���6&V�dW�tL�I���r�F��d�A���ߪ�(��mk�?oT;氆z �GP �x�R�_�;�r�1�S:a�	��y��%2g�J;�]��6���RJn$y���t���KJȗE�P�3�`�,�L��vS!�x8�n�Ds`1��%�XH�F~W��j4�_p}[oZI��mBIBf?�d�[߄�"t�Y $�6`�B�]C~�o�����ɲmi�hY���!4ȴ6Sa��H{Z�gi�	7<l�y�I�ۀ����7���C��-	��`c��b�Jp�K�ro�[R�d�Sb�`���C2̏�=��Vb�����7���2�� ���F�d�I���~��D��ӻ��tk��B�	o|B�1��*�Y���g�����ѧ ����'�R"�(���>	i�sE��$ؾ7�Ȯx��Bz��Cdf,]�z���07����CQ
�ĭ�	b$z1����ˆ��]�ǽ�U���/�^_�A���@���Ɩ,|b�|��tȉ��6������r�&jF{�y�?q�abp�/0�ag&|�A�"Jf�E����{�a�R'!\��m�V���!�4����F�f�O܃&���_+s�����(�A��8rn_�|nJb}����f<��h�������pK���i8�i�fT:n��^�CFckc����GS�qe�/ͻnF���! P)�;�>Ź�o��m]��y��ȫ���i)�~�h����.�O=Ww���t�|+aS�d�VG�Hw-�JQ�����0��e�Kǎ+���PC'Z���O�5�8bl�:�`�����q�xզ��|�PhY>�qBQu������-����tw���k�;Ol��]�o��}�*xX!�ɛ�$]X'�ɒɭ�@,y,��L��4���	N/�Wv���{f��_c߲�y4v�_��

��+��=J�G��YZɫ/vG�k̫b=����i��Ӡ^�*!��;0H������lzTv��J����T�����N�e���[�Xε&�n���ҡ!Bg��Q����o`?�4����p�\���ͫ�.�s�o	Tg:UgD�lfy/���*�k�|����
��G�%����=�.2X��U��qY�r� �R<�qK��%�z6�4�,T�'��P��,�tv�1g	��y�X�a����#-�`�E��Rp��q;��q��j	i��5@t&;| ��Q��Zz~�?�n�: d-�>�/�o&%���SU�Jc�F��9
h]r^.W�ײ��,J�N�]iJP���˸l��*��1N��A��>�,�K#*�)��Ǐ��#�BB9r2c��2dK�������u8�A�Ƚ�B���x�sꦍWo+�|p�QӞb�p�zp���B�zI ퟗ���j'�}�5d�9�'��Yl�$�B"�` �m	���Nn�=��Vr/�/w|,M��`}���ka��F��=���R�p���N��u�"n����@�w�@���G�yg;���ɒ�e���ɴ,ZM�2r5;�d�q��aj{4�6'0.¿�E1EC�=��M<{����֑�L���X���5�P�ʽ����bh���}�������di��.S��ujQ�	��o�%T�8�9y�[׵̽��h����+�������:�xHD���*�[!�$������b��|t7ڼR]r =�%v�!����O�����ݳ"%c������N���ן@��)�>c8�ޭz�f�T�� �.c��"����Gל�͏�J�s�Y��R��ͪomYOy�8��Q�)]��M��@�5�	!�C��%���с^!<$��}�/�>�i_�mR;�2쫰M���e��NS��^�;~��q��C	�9n �-1΍��>��Χ��5o���,����P2]����q&
BT�ՑP��8=J9�U^*A'��d{*ޕա����nd���m���ق�GsGU�u\�,#T�q�	�g@ޓ�ޒHO��\�vZ3`�bQ�F��c��,\{����7Z�C"�~��;�iQ$�V�hk�,���1SQ�G��pX���8�KO�w��"i����(k�n�&��A�f%#�,��ف���s�}���c�Q��*�/k���#��ڰr��NR���AW?��,��@�/G��3D|�'(:}����+�֮���V֫���vXL�(�7���1m�7�����{�$���h}�͚��j��Zl[q�{a���xl�D�@���� /vMq*5�G�-�O�e5�M����� =V��B�G��!wuK:��R����J�W�V�
������|ľ�hj�U[��M�W���S@�����v��'�`��p*�Ǻ��0JL
�pg����fR�wq,�_��ca��[�]3��B�����<�s	~VL��,JQҐq�S,��ņ޶u5a�\|�3��ޞꬄ^P��R����4��jC�	��  {O̀�c�ߘ����nC���/���%V��ؾo%����>��&��t�������ǪL�XE��Zu��6���j�W��y����n͂��2�b�#��_���C9R����J������r����SmXt� ���Qy������� D�J�i��_��痜	�C2�"�?њ��ys��9w���NI59��ݣ��U����Kca;x�:"�j6r��4Ը��GL=������}����Y,�?�<�:�z�wu��ll�.���^5U�-����]&�h�Tt�͢�Qo�@��m�`���z�9'��>����&�r-��H�5heŃ+����b�<g-i��_\��(F��Qi���kuY�=�V3ي2'{>�2�:�|��0m;�>J��{]hr�p�k�B�XA����B���K$�V�P�&P�j%	] ����߫%���6�La�<ƕ(6�X�?S��`ʖ ��4��`eo��6f�#�ݨ��Wζ��ڒ�63�o�v@����|@[���׉)s�h�mǞ��?�f��`u$�Os�]�b	]|�8��2_e�:0?ƐFu;q�$	�0#�۟���������j>a�J� �ڊV(��jZ���[`�p�zl}���M�>��3�p|)^N`3(j�l��&\ͯ^�8=P��+��^�+?�,DS'`��m�al��s'�����T.��<tϞ�TK�P^�#֧H�j�^;#�����Kکe��^!�i�'t[Ȧ0���L���%0��QĖN��׀^����è�"����ߛ=��[j�g��<f�:$U͖�{��b���kj�S���%I�~x��a�0.MV������~�f�Le@�C濥�(���Z8��^{Ӑ!P��7ލ�W��.�X�Ez�E�(��*�0q��n�՜2C�;��#�py9ٯ����zU��q�p��?�g���l�{�'��D��b}��T=4z���-�*!�zh=k��ğ�'��7J�OJ����w�����[��6�����s�{p��p4PP<l���=�I�u���G
�L�����:M�5U���ؑW;/��?Rg��b�����[��/\�%yIe��G��E�0����~������#f Tu��g6�2{vD�e��4�� ���N:!�&�bT��~O�"]e�$���bbv�^�Np�?�>6P�/I<�W1�i�!-�fӿ*�,�X
;�ϐ0��-}�c� .���ʅp�e��p,�7�����6������Rqm�*�nĪ��0ڳ�?/�`�'6���*�s21�v��l$��]�?Nz� �+�x�X��=�&�ݴ	���1\}����3(�1���Y�� ��Q���I8L|�I8_�3�?.L�ت6S������W;a��A�f�T����7�MXDd�`����X�e��~܏�&�� ���?nY��r��&{�P�'�:Ϙx�@lDə���}e���>Z���e!����.�-.LG:Ϸw�^�b�%<ḯ���������y����v7�����
6����x۶:E/#)��e��}��n~E�:�OA
f2ڱ�h���`W78:�)���]	�u���5��Vչ'tǦtZ'�xg�W?;�*81AM-5u��כf�P�/O��5p�V�Ăk� g
�k�;6���R����Liz?�L��)+���ZC��
�"b	N(v^����0�2w�H����J��@ �@��&��|͒�ܿgS��j���(7%��f���R,T�{'4�������ܧ������j5�І^�����h�����I�����h�A}�����������	�p�찀�+�g�i���bh�f�6�f���i��k�J�9�(ֳ��U
^��0Cҕ��{hzL�jwH�t΅��O}j��JK�S:�d�v��DC�Ņ�@z4$m*w��Qh�V�Zo�y^�{(ih/�/VuI-F�j��l�ڜy~���x�B��6*��� 3U�?a�K߻v��}�Y:/FQ%>!ۑ��q��w-���%R.��^��`��$��&z%��W�t�'s�T�Z]���4�l*�;�����*�v�gΘ�K�C�H�3��렲� 0R��2t���c4��\d�l��S��;k��<���|B}熣���e56᥹�(��@��⁓�B�9�H�9�b\�xG����ۺ��Z�
d|݁��$��r;�PBq�#Y���GCF����@~��@���I�;��iG�	�[�P	�������Ô��n%��6��4�N���J� D���t5�>w4p@����1��Pc��ک���JA�#�ϳ}���AP���Ox�cI�x�ge~����/r��{�m�ʚ����'g~ns��"��C�e�y�5�U��(f�Hc&�3��KL=�$V�ej�)�0�.	x���g�yu�2'��;���&����:�b��VӋ������!�A"�?�����n0��/bA�� �f�Θ���2�1�j�C9�%Z^�9'.
��6�&O��9��2l�p�w��*3v��DHR=\���}�C�gR��q ���K�����>t�2>�4&�kk���|Q���c5�o��&�ߴЩ�T�:b��-���G`��K�X�-����f�0�x��s��#� �N
�n �p� L�sZ���Q���#�T9A�5����
1�+&G�GB�G���q���I`��-��2~QhV7G@ߖ9�3��}���/G^x+�._V-��j�ީL��'�Q����`�5�sa(��ÙS��!�H��4Z򕲗���������n�4��&����b��ѵ��"An�m�x�r|�IoD�!Ǘ[މ�Rr��W��H6Zҩ�b��ϩK�x����%����W�+V���?ϵ7�G,=B�_�M7w�_��UVW�d*�m< SX�#x��}�7'�9:�5V�D�E��jz��֏_�%3�)�%�6V���0Ugs�%����9t���|L_&K�-9#�#ֱYa ��}�vZ���q��a�!���v�}BTA��hm�uj��7Z��d���Fi��`���mi��R$��y>)��E�E�!�sIT��=�KTP��<���뷤K7��o�̑}���h�vQ���kGJ�ׄ��� ��\�}pǺ�p����i�JR������&C7+�?�>�&5	��'ܤH(����@4R�j���sC �A�q>ω��A�
o� w>::�L7M��BL�W��+�o�����0CҘƒ�rԟ�'ae�^>Θ�*����< ���.2���D�=�>���<A���px.�N�:1�X�O�m��7�\��Hɭkz���xA]B�}��r���b��E��]�?%��ZP��n���T]��7f�����q�3"[���P��zaz0r�+=��oo�߹�}F�O��Ҍ�=7[��|o�)I+�Nu,�h��ݴ�1�U+V��V��2�5���/�H�v��"��
Mt�!V�I<�M�9XDֽ���?:Egj�.[�}c���a`�����Y��{
����"�7���N8T��aY��q>T���Q=Y4���x�� ��N/L�Z�;�Q�	�nL��=�Ot6����B���,�v�jm!qK}�|�%v��`�&�����C��|3�s�/nHڵ_�nDf;���Qv����s�L�q��g�*���s5�B�|��q�?�
@;�1�����'
�yhPY��\�雏o[�Rs]?������T"�pA�o
��0�M��}{��`���ٱ���.����u7'�کI5����ԊF��=��6�%�{q����>�G?�[oB]�W�4�o���U�a�Iv��X�ɑ[��m��UIp��4��B������4F�n��:�H	8湠)uo�f�Ev��Q:#ٖ@�%tA��j�-c�W~����(D +���v�T�G�/� �J~Oh�DaM7�/7�ܓ��3b��X�a�>l/��.�f�3�V4���q��~}XӁ�t4	`��؄ʱۑkޝ���_��Sx���9�LRv|E�מ%�-'7%�Ύ���:�UMGR�3�x���l
�g��dpL)3���p@��J��i-R���j
eo�g ��,U��d�s��ёeR//�G���;�n�[�a��1I�C���$���N4I�B������(�T�$>�(e'�\+-Hl�T�#�nё�N���҉]yeg@�b �:��j�[`��w4�������0�T	�J�#��I�ʵ��Y��Z�~�
�S���'�?g�$�N.�K�9S����,�;���ё(�q�%��)bB��q�
5��
��R��i�5���%�m�h	� qL��6A�����o��Ծ��d�*�e���7� [(���?lb�������l#1��:���'�F����K��?�ٴt�7��F٢����(�e4��b0r���͖3T%�*.��e���7���`�*��-��?ED1�Q!H$���ӝҧ��UPRݟ�U\���:<#�j;��ٛ�����|o���	���i?	�^ ��?��J�i'�69nT�o<���^nc'�p˙��U���\�,�����ƣ9�Q4/�G!����P���|�xO�#f��oؿ�7 =�� ����F����S�TF�j�:d���Qh,:�V�|��K���[&�}S��˴O��rezv�dSb��OW(����i6 ��$�>>sx��ɨH��O�>#_"I��D"O�|�*O0N���C$��7�Oo�jХ�6�:\)������c��e�~� ;�e���7�2�2y�,(���e��ē=�f�&���_�0&]��Zh�Dh�<�Cli����"n��5(p�$4�/ż���2;�K�|E�s4�x�b�����{/��v%V,�:��T-���� 0���
��h�����n-L^��wkë%?��}c�z���,�˃=�o�Ծ*�[ǋV���Z�f�rL�r-�C��D�{���=ͻ'g�q*�垀�u/`*x�jZF0������˼#����&��{x�.��y���N�����E��fr_nͳ@(���`��Nbr���w]��v��6G *��Tu����1o�۶}�+���c���xH��R03�h�G�P�G�"��l����c���7�5��&���=2铃bT8��uT^��5�����F��/j�ԕ�(No~�d-�(���5}�b`ԑu48&_&e����;��OAgH��`:���UQL�2���=��%��<��1aF_f����C��� � �ҕ;W�uF��C�c�;Y�p���e�ѷ�}�,2i6�䯿b��%���$�
����<�|��szh�4}1�x�*�)������m6��2d�Y��b�L��Z�� jl������c�xQѳP����f��i=�I`��R��;�t������f��l����aʌ����"e��Y� �>	�ɦ�zL��d�.U�ڸP	iR���"���N�H�������ǔ< ML:��˟c�K&�cq�t��((�G	t�DW*��i)(�@T�54��n/OI	\Q�3��?nA9|1t�y�C��͐�K���Ў'��D�������4��l���Wf�)	�a�-�4�+�Ω-��F[�֘"@�-3�`z�ph8N8?n��^�b���S�@���ޭZ Jm��N)�&mW���ݼ���U(|>q81�Ɉg&�<_CQe�X1 O32me)R����o0o��V�-"�3��,�@��:�W��8K��%g�Q'�5{���_� 8_}��H�X��q�mM"�,u�E�D�䍾*ߍ�V�@U?d�!=�d�����FũL��!临R��>�{)���wp��F��`����M�b��X���� �=��7� о��I3z�q�^|��;E��M�5�O���B�~�F���Y	��$��Կ����H��P�Yo :�v��]j�-$�����O��ҥ�wb &Q��T5:���A{O�H�Ը�cD�Z$
s�/(p��'vǗ�M(7�]Z�o�=&�.��T�U�R'�B�9������e.�+kn��b6d����RX�H��a������L�i�@���m"��L�a����	�C�Υ*<�`Bl���f�'n��k[���{�@L��Mq>�K(�^�2tq�In��h����`շ؃E���H��Cz�u������/�07Ս@����t�.̍����ӕE�d}���<���d7m��i:�&��lUfÝ9��oV�W�+S#�u}���|*+D�������tVD�4�z>���!ߝ���Im�͎Ͷ�Qlwe+]O_H�e��@�Ck��p��eDļ�8�j�9O�3�_�(�^� ?���"?���X���g>R�˙~x�u�1�U���]����ڵ�`
��ECJPeZ�1�<�w�c��SIqϩ����@y���������(q��בF��-����\a'��+/+ne�r]~5�7_m����׆�\���n՛H���QSd��i����{#��Z�_�zzD�9c��ψ�B�fɋM=Oo6}�y�b�&�|�nf��^�����$K(���m˪-��Zտ�J����>p�J����4tn�,��(�b���ڃ�3��Y\U��eӫ�L�C�0GSɠ�v�,����3�����s������/:ዑ+ %Dq Y�Ď�̪>o?gB1���ʆ���C�ջ!DD�@#Z0�+l���H�����M}�۽K�,��g�N9i)��+��dEC���V�*�B�gtn'�z߶��讴(��ɑ�����H�[$+�s��ҳ�)�ev�§�L��9Jpt�s,��P�s���R�&B��^�K��4QM1������P��,�D�'��Q�d�DM���qu�xƎ�<��҂#�2v�5�����I�vY�L�5Nx9#,?�a ��i�E�H�Wx%�5g	+�Ԃ�C<oޒ�޴�F�>����1�7�����e9����r�-EP�4������ }`�av=�5�3���9���G��4�폘C1���B����p�X���'�k��hџ.#��2��D��xW)L,�
��,^0�_Z�� ��,>2W�R+YXN��꺼�l/U�%y��%�����ȼ������Z`��ܙ%�rY�^#Y؈�th��mK�+�f�Қ�ov���X���D!W"�>��L�����W<[��ª�;Y�5׮��h_��X��ӃOV���l$����9�h�g�5��ek z!�F�EM��෠u�GE��e\k�^x�,eU��IA��!kV"�W#.shz^��AC�*��Qʂ@t��Nه=U�˩��,�琘06یgt��f-	N���*��h���kE�VaY��:ɡ*F7�Ӕ�r�^�4�wI��~�@Fd' �c�{����M�/t�;�TeY��3y�L��^��q��`����`�>
wmV[��G�������I�MDA�\������T�u���m�	��P���sVH��d��n/7q�ފM���\j4�S<�O(�Ĥ]���D�F��N}{pi��	4Z�(ދn�k5�܎r94�)2�M���塯��r�[RZ�����H��1�PgIrr �ZM�����uRN�0J�x���U*pCWX0��_hʴ��-��1F�uG��7Þ��ʽE���5Y��yX���'��L�:W�%w0��s,X]�rz�C9�Ρ�t�҃����4rb-�ʾ�u���H�[ o�-�� �g����w���{j��"������՜$U.b���T�.&���7�䗦��dJ�������6�k���r�����љ33QCp�E�޴a�-��[Oǽ��Y�';�ޯ:��d�p�a�6�������=4E�YP�bi�\��)�q��>��X�S���5�k"C��:H5@��iL86��"�޲�����  s��@��g�[�x!�H��_�� ��'lʟ4�D����� �z*���q>�#b�^��3?��_�rV8����<@���`��u�����T�����j?oo�=D10@�3�!e��"nC%w��J��&�oX>�v��<U����.�O���	��S��3u��}�kv͔���85^�q�Bx��Ƽ���I�E��Ǟgo�C�끧��C,�RD��=�����\S|��P�D�c�L�)@���)K�W]I��4.U~�&��h!`�E�"�
G@&F!�R2�r�V�Ǧl��\�~��@�٭���}3?]�Jt��"u�~#_�Y<%Cv]�/���Z��D�GR����Z��V43�up��,��l�P89�����`.��h����c�C�2�P���n3��T
��R1e��z�!%�h���g�yY��qF6­Y��9/�2�� �q�t�U�a����� ��d��_�12���,@§����
�)�l��!��x#���v��܋�>z����Cw��%�7i�����}l�N_J��U��pJc��8a�i)����J�Ep���������l�i�o���+jT���D�v���� H�̭��۠���@�N��.4����nO�������b��""�ɭ�Cc�\Z*����T���	t�ОK��c��3�N���ß�=LD)_9�`�ސ7��S0ԯ�NF��Y�?���^��P����/�ɮ��^���	�$C~r�0+5�|�C��[�o>�V�̠����7W�������>���/69Y/�7�������]�B�"��Z�$��UD�����2�&3.�^�x �:&�oR�i��ā{���>���No\ߺ�!�(�<!�
af�����-�)!�@�\WX��k���DO����*������ѡ5IV��t��[^��#N��.��q+Ѕ����t-9k{��a<� i$;�"��'k�
M�;���{��sH���XW>y�yE^�uQJ��S���� ���3�#EZ���=�٧��ܩGo$'���R"GG���������bhP"� ���Xߣ��ſ�f�b�AD�1�-��6�7�����)��k��)��8QD������2��z�����LD�]�ک�,��g�b�\&��^)�F
;��,������� �c�ƀ�[b�w�'��%�@-Ł-���T���!,�P��z�������-�����%�m��'X��8������(�����M(g4�j{1xry��j��v�j��*L*��j���:ky�.�O�L
��yokPV��B�7��i�]+2�)i�f8�-H���������G�MC��'�\��=C)�o��b�b3��Œ,g���劭B<��|�*d�c������o�����y�s��c.Z��{���k�d1�*ux�C���+!;/Mk«��΁�i�ڋ!.�tYo�MQA��L> �+"�Q�1��g�Ĝ�A
�y�17b��
|f~<�`��"&8� �Ǳ���=\jl���pT\e3�9i���R
E�eUS���1�;V�f���t��V5-4��U��s�yv�"aCɌ��C�.�յ���@�s��Iz ���5����z�G��`���-.CW�4�|`�]�P��r�]M�}C��\wjӱ�:3�%�����!���j7Cȗ��[����/'/��Z�z�J�6�AC�{��G���Q��$�C���;�QH��{q�Ud;�J�5�8����M��+�%y-��&�O����A^� ���YX����(
Ͱh�b}���r�2F�7aiu^�X�51	LC�Mj�w��U�aT�c�J�R��߲&D��Ȓ����w,t�Xc�T�%��a>�$n������_K}�אJ����s
1�?},����.KV_e�|f���#C��
ȳ<
5�^��I�I=G�"��S���օ��u���U�ݢl��(-� `��n��A�l]T�G����7|�K���J�U	�X����/�wӪX����ˮ�6�n��!0!�Hx2�w��J*���l��g*#ڭ	N�<ܒ(w�ˑ2̠�K�Z9��`{�J~��8�6(�]ڽ�1]@/z��sT��i!Gg� �2���z�P���gqpë���=�iH����5�ILV�ż>W����V0+w���~�L�ԛ�{��釶s�Hp���VmF�\�g�36(����U�����bu��8bF�����m�j�tm& T�aFK�"���3�Α��w��A�rn~����y��#�?������q�$\*�v�`z yc���P;��d�[ԯ-0��|�Co�x��@���M���fr����!i|Y1��jꗫj����)���4���G����fƙ�;	Y�����u�}:���#��D:�}i'v1.)#��_�j���c���MȬ
ٍ�.&X8��	�Uv����c��\G��9�$0İ���ܫ���Z�[���̯K�9L��y��.� �궮��Ii4�����iU��ˋ��Ⱬ5�O�h�u��t-��c%�O�����0"���z��_�X�uB�Ք�g��Vc�u��������r�3���%��=�����Ǒ�V�I:��j���_h�g�$X-C��������'�ҋ!�j�̹�xo��v����v:�Ŋ����n�An����n�#;�Rk���D_�&9��2D�уt~�R�>�$�5�Zc+���9�h	2/��U��E�}��O�~uy��HHgy�x�,"S�T����8d�Q�7.�3�!p���;�,�P
���+%��;CKw�`+�C�*�a߽>�E�Z�C�Q~�5 �W�6��3�j��(:� GO<�)�E ���휠q��/ ��d�7Tӡ�X�	�"��6Â�ۭjgF�C�ph����̇�#%4!��J) ���Ge��}��.��ywY*�(�I�BV�&����3��A	�ҩnW���G��j$<��%@�4�7����� �M�;ӆ��J�vE{za+W�9~�i�퇗c��:�J���q�m�D_�e��oP��8&�d�[�!*����,��[�-pl>����ץ���+A�:&őXaCM�H�_�&,��ȸ�Tv&7��,L�k#P0����H�e�/\{�y��WR�I�@�[�y�Vh�ċ��im+$�Qf�Л��k�27�ƥ�|���.}����ԭ�)%#�t`;�&g�Щ<fP��m���T���t��X�V���tX�C;k��1��s\��۞F^`hp够�=�4���Q�;Q�5�G<��R"�b��ش���%���y���ѥz�"�sENv�	��Ъ-�>�?�!���Γcܓ������ƳS��6x�ւ�fG4(|9��)���2�5����FH��Y$�~���*�E$>�f>���N��é_���*��79E��[�����2���XA��i�5a��M�Z8�V��kS�Nk�G�>}8Xw�=ș�/A�UK�CF��>PJW�9c�S�9]I7r��s���@k|ZՐs)�.~�S%�ª��Zs;/{�Y�-����j-��Ȯ)~ס�r/n�>Y�%CLlx�ʐph��{@��"�O���,�Ic�-�@q�k���'~�X�C�&{��B+��o�s�A���]^�/5���D�p�Om�C�uh%�Δ�ֱU�j!��9�X�3l$���f���Z�;l7ߘ@��%���d@��d��F!3�.,c�wr�)yh����ﳖ��'��15���r�HC�L/o��ZQD6�EYŋ�B��BPKT�Fz!�N�s�-va��;��c�ҷ+��0|T��G(ʳ=a�ZA��V'�� �����@Sg�{[�wG�H�_�G��]�Kߠ��"A�G=������2K`�r!��z��H��P8CP�[]R1*ɯя�9���Rd7���ܒ	$�<����X=O�ՄM��?��V���@X֠�������i�[%����Əi7�B��?�B�T<�a�n�]Ί)�;����v���g�$&�4e���
�_�3�/��v��	ǅ;��`�+J���ćj���Y��t���K�,�D[�
G�C<:<�>J��_��5.��g�G�K��=��eN��x�Ź�4�k ��'z��d_G������4� �tٜ�>�Y�k`����b&H�P�Y��s�	�$v��52vd_��pF+� {r��H`�B�{��.�R���e0K�=�B_O�T:�-�7���n*�{M��>�[)L��Ϋh<��k>veL_b���)v"�����gb��|ĳ�]�Y����O�(,�FAu���I�E|tʄ_��!-+����9��I�q�����iz�|�{��߇�Wy�ydA5�x�8�q	��8�a��&yV6̻�}�|7�a���!s����#��=��2����g��'fu]T�N@a�t��l���L���������"DiQ�C��E^F ;l�m ICK��j���oO;�/F6���Ϲ��K�cG����)�l�N��c�=�*�_Nj����#�0A&e� ��x�L����K��#Ex
D
�l�J�ǅ9�W/�����1+�ufm�a�_���qL[�n�o쐖,�~=��C�Ï��G4�97�7������V��g���|u`w|��3䭦G4}D!5x������vO��|��u���"*ϟh��	?o5>x2f���Ko�B����w��R����g&��Q�k�� �>��ܱ�����y��5_G�f�i !"����F�FŨc&�Ych*�Xf'����M]�ݞ~���`z\�VR�Q��oɯWwt���A���d��g���<"P�E��L倚�$(�m�y@�؈sz#���pD������r%F��s�i�=�ᾙ�f�}�1���D`�q�'U!&�wV��^2C��e���G`�vq$��r�of�g��r�g�b��4�\[�����tcI������R�kBE��}�%T=tg �4��F��>�@7c���v���`E@8�:1�LtA���r8(̵np�̀���T��N�?!�d,��B<.��/�ؔ�Ӌ՗�#�p��Xc���ifЗL���ٶ��R�ų�8+V�DN�ўq����w�]�y\�e��Ů�7�'�G����
�����؞�?s�O�@N�¦
���AoH��i�=1��ʥ���+$�3�9YΔY�eo9�iƩ}�CF+fj��ô�<�(��]M�޴S��������;����%��E�X��.H�����O��(+�Ek�@������Z���u�᫨�re몢���ϊM8Y��o�6=�@
&�*���r�I�D7�
X��7~����W��hFp�&;Rh:x���0�r�D6ɔSVS�iU�����H/B�@x�!�Y �ֈ䒦�#ێ)���� G"!l�!�o�2��o'�?a�*�%��X���jREM���jUP|0�RE�^cg��,hxG$1$���4�#���,Wg�����%�����J�4^�v�@W�$�i�OvaW�ʋ$�nw��>�#��D���Il"�O�+����o`�y{_��˙+~�N3U�u��Z�D% �;�tC,�U�f�m��T�iB��6��A�z���0���=�-Z�QvK�=%E�^��w�6�N��t�2�u�%2�Y�/�e�p��F��{D��F��t����~�����ؖl���J�a�K@�P�]3��P=R��vF-�����I��07��~Y��e�����T1�c3�o�~@Խۄ�3��������28��#x��
�+S�r�ΏX�&���	�kH����I[���?d�7"� �(���#�|�G��'�>˜�����܁CoÒ`T݆`�5�ʃ�x�����"�]��Ȍ��9B�yТuЯ31�K\k�=������1��$oe㥏�'<Q�m�u�����b��Z+��+��E~tgGG��*��e�Hd"eo��_��z͋e��Qᦑf�L�`�r��$)��W�����u�t�4�~1  �)4tT���`��ĖO��`(��1�O���I