��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\����q�?��e�I8�b�Ǽ$��"����׭�m��ܱ�;iR�%~~�T{u�q<ѥ�mu���q�d���w��N�Dt�+���۶_5Oݜ�Bb{짧�u �N.V�����2D�U��Z���5�t�d mp�� &�G��Q�؃�"W�Ĩ�F����WV�J/ɢ0�ps�N8Ţ�E�9�ݵP Y�q�OL��ö��A~�X����W���bn�/!
��&�A���M�x�q/��&+rC7ЏA�Y>@)̣��"�u�-$sZ]��S�`�ɳ[߿G.	�a��e��b"����.��w�o�,Б�<��GDk�G]��Gi4BSS�A�����������e}�)�'�:�s�n\�F�Q_�45I� �"�r���Y��dϦH����_�$M�V`��5~�45��	1E���ϏV��])�SY@$�`I3?s;�X��ꛒ��s���\	c0����%����j��8��B��\ڑՌz�����u�����ɂ�|$��ull�@;p����̓�ou����wnKx�d�_�[��?vQm6����w�H6V݃r��W�E��&����k�U2;|��>]�T.`zw����7RA�0�f�|�I-����V:=sg�o������A�+�~�+g���0��\AB	o5����M:B�99�:�Fj�v��B�A#�g����#�r�����l~�V%��M��3{ϗ�>ɱ�f�4R�E�Q
@�u�A����aY)��' �ۤP��yeवP��:tTK)���`�tIo�uy�:씻.»���'i�7�  \3�؊\��il�+޷N2`�ɗ�κ=�����ApQ��ɼ�U<�ω�P��S-���}�Y/�?U�>�9p�G>��Z|*0.�%��f$������D���/�_����-��5��Z������"hh'��rYќA�Ί_�|q%��R�m�*�3Y)UH�4��%e�{l�3�^Y_�7D�dR��s����3cf�c��{'�L��^ rL�Q���FnxG��A0޿��蔤�OhO�=��X�w����	&����/ҷn��,����o����*�|jk
u����s77�c�?d�Dx�=�U�T<�_���>�/�a������0���+s��dg`s�/���v��s(�y�͸gI�bE��j�����<~��ITA�B�ٽ�]�"E�������0��>�u��(Sֹ"��4*�W�Bn6"�:���iV���&��?@�n�P��!.��}�����]�b���_
)��������Cb�N��xJ����)�T�z������Y.���N���6&�fM�y���E��lzē��U����p���,�N�`�h��̊] �c�*""�z#E �+)v@8��WƧ��7�HJ"W���aV^�C��G�ASOL~�>��~�U˕�Nە��:��/(���Ca�ͣ�������{kȊc��
	�'�����E�s COH]�s�?l�6�~>==�����360��0� �����h$���p+��Wϥ¸�dE5z��ߓ�3PJJb�~���<�⭦�S��T?�o}��m�*ZXZ�K4�=
�0��<w�iV�!D����^Hn�#����kF#�R7�LT��Z�|��J��[v`$�V��&ma:L��������� 7�zl���4���a"\fC<��+�XN1��tC�V�w%>�����n��j�#�83�+����Άx=����ۋ:9�-֛bAǲ�G�&}��(R;TT��{e��*Jm�7�S�V�P�/��{�/��˔V�M�K/��;�����s=�y2eMFd?�V�q�p˞!��b.� o;�6�w!�E��M��wQ��C_��z��&�_se��W�P��K��J'�
"�����x�ԺMz�'UAa���S���/����O9������3��oa�����g�V%L��]����������v���M��\S1՜����7��3K�9�T�i�$�j~�lWa��\4��k��C%��]Η9
a�g���](�G��M��x5TB΃�IR�e�u���iFH���i��QN��� ��Fd|�#39�����r�o�j���<_���Vh�!�e��� 8^]`ރ�{%�4�x��ylp{t� {�{$��)
KE^Dۯ�2>��5��t�k<b@����@|uB"p���'%��ٚ�W`��6�Q�v1Se�轳��ٚ^g��W+�hh`�c�w�����CL�2�vY{�����'�&�^� �{�ߴ��S�6z����߯�]Q�p:����F���`#d'��,�?��_aQ���5�A�Q�p��gE�� �4u�5�z�<K9%�Z�����h���4�� ��t����|ғ�Z��&b��ʤ�u&\ځE��P����cs JA�����F�*yI��A�����!

���:��Zt.{K;ҵ����L���5Yb$3�Y��=2�f�!z~��D��EpWEP>s�XJ�6X�W�2E�̐I����La���%�~���ka{;J��1��y�&�(�E*xOq�BJ��=٭����E&Fy��d����S����4ۜ��|A�Q��?�A�b�:�5%��+V�0]�ad�!j�?�"y8 �����#8��^Q��*�z��EN���Rt2N��˙G ���n��K��M��˺U/ap�ʃ�Qp��dS�`��V�MRA�Я��&��F���q���!R�
�`e`�`�w���_��0(Q�-W��վ��9�+�=���b���]l�����<9d����PQ�IӢa؂��:L���|���Q��ړf�>�,*b�H�@ʻ2Q\������4��5y�{���ke���sz�i��^t��o�\{�ۀ�|m!�H�z؇������F��V�Ũ4��M%�ʠ_��:��5�x��
�f�� �� ��n���x}�;LN_?8u�ޚ���D�U�0y��!4Ss��!�y����w��얓�	�)q� ��7yW�Cѝ?�qɐy,=����Y"� ՄċL�}�Pc��|���Gb��z�j	Й�=.%���.�:�h�'��)��:Ě�f�p�5]u��m4	2�
Y�n��K6.4&:A>��_�@�z�{�$>�~0�eo�]��A���ߤ̓�\ Q�pwe�(�r6�Q8�2�=�v��;|5�%SH��'�v�(�����(�]��a�Qɞsu�XP�����c�n��7�`�3@���7�Sq��P&`Q�X?��Ժ��}��3��R�'6e�@L�^7H�I3��\r=#"���y���#�'M䩾�������Bu?;H�����;�=��WŌ��`mR3a|��WXP6���������D^��ï�Y���b����p{Yǰʲ��\��ԛb���� �R7"��1��2X�Y�s2�BH-�7�/��M%�[#���RL�������sh��% ��(��#�j�&wؼo�๕S�ƞ��]˘��g}O�n(GE�M�W�Ȕ
��[���|*Nh�Ub�_��F�"�aA�&#���`v�{��|���i�W�>���6���M;2/�n�������t�C��>m�'�bO�6�������h�_�h~�dv�/�r���٥G�|ƜOb�nRL��Â����C��.���;d�{}%i�-V�4�_����±������>Vc1m�!�RM)rV��}4�����,P���X_@ɖ�����Cl6�U[C���'�'���UO�>�[�eR/����ˑ���V�Pe�x䇫�YC7-NY-6N _�!�x �΄�}v�Kv�����c1����U��}#W�"��.���qm%Y(��v���łO@5��f�
�`�ͤjZ<8��T���=Ǡ�K�G��I��j
�-����7|�{rHiUH�m�.r����Q��N��8�\��(fx:�'�	�����������M��U�}�x,�:3��:�һs�����M���#Y,�c��1R[��1�W.���ư�b��e�!l��M��ՍL߫�B+Q���:��Bn�����g	$��MR�0�2YE0$ё�\�^U�kQ9�H}<��� ;j��D�����,�|�#��s�M˧<RgBa{��rQ$A�$-���]��B<oYt{�3Z��"�uy0�{��CO�X|��
�.�$�Q���~{���W��M;ީi�f����}�5��:�`�Q�^��,"�?���پ�xZ�|���9roKhĝW�w�S
�F<:o�ݒ	�	qH���/��L�ޥٶ&���1��ߒ�K�����`�x��+>�D�g�R{'}J_��r ��]
aÍ��2Wk"�pL����^�����b+��D{�@|<o�v�Є��a��y2����-wwo��JN�a�8�Kͯx/_H���M/J4��|��<�`�s#Z	ES�?h����h� �,BkK�E������Ǝ1̠C�!c �B��!�ǿ�Vb��܏6ϔ*�JD1�1A�?�" (��n���vM��_��eJ��ҏ�W״Z�����8``&�IH����O���jL�jm���S~��8�����Bc��J��x8�����H�]F�^(Y��լ#A�+S�r�C�Ǎ0��<���+�!7�W��h�(Խ���GxR8�(pS�-_(���k���1���W�/ل�,��5�o���E+ Z�P��Lp:�'�/���-�����4�^Ӌ�ħ��_�V�_$����f7�Z -;�?k(439��_�i�#	���l.@91�l�pGxRk�wn���B��a:a�\���u�=x]`�BB��֏#&�Y��l�fbN�}���$E~+���VEnͬ$@����5�b�φ_	FZJ+CS�uMZ�����2�� �1��2�^a�ѯ|�Ae `*�?��?��γh^��{ɶx���襎��B����1�W�/�KI%G\�775���݄�d�H�Q�� �Gx��\���>h���6Kԇ.���h*,�u�{*.��r�T���cV�F� e���� ��p�6�37�N�{�gn�,�9��� $�����C�Aӳ就 
�����9����]a���fve��ԣ��e�	��B���F_X�yF�t�J�RR�P�V��ߩ�V�����ݐ"��_<�L� �;��+|=᜚N�N�)���1|cO��P�㻔	�I�������� Eĝ�M�����
"���!Iŭĳa�����gV�ԳB)AB/N!�˘:]H,x�d4��g�7�����e���o�F��}�N��9��3 ��e�;������G~������������Ġ^Ob/S��*��G�*=��2����_y�"3��|| l`���c�;pk��.�D��zl��(u�9����Taz��Be�#���*�z������y����'E��?k*�	�Mn>��&x��~� P���5�9�n	�:YM��5>����6�_��e�DkH=/n7�M���VZ=�\�y�ߚh;)U�$\�/Z�}��]6dG|ѹ�W�˚�e�O�%��oA>o=��N��?>�d.qS���ׅ�C ��y�:_�_��$ꅾa5�I�ʢY�8Q�t&��z	��n� g����Q'��M+K2�� _k�����ҷ֗���%yV� ��$f{�c"�#�~��c2������S��}��	f���r]�2���`��@�eݶ��:t:���ѭ˒'�}��<�,~i�P��m�ev0ث�p��E`��N��>�9�o�&��9ߐ�鲼:�R����/v�(0C���sq�V�:{d�B�E��Cy��d�WH�=������Z�c���=��uvKP%_e�n�$<�̶[.����,��9���L�g`��Y#�m�u�ϾP��D�J�(R�.OxΚ�
����% U�U�.4�k�p�4��J�hG�#��>�:uL���wR�J�5��H��t��f�bI|���C"�5�m��ף?K��WO��te����Z涼�pa�$��s���]���#�� G�����ne��ᖠ��lc*�nYI�4�_��1�6M�=���v�(�=���5�����o�wBe�~�*x��(;�;�K�.M0
�©�I]9��j��m陀&dɰ!,�~ܢ� �G���:@��I�=���d�B~0
�0�-Ij.�F�X_5_�����Ռ�	�l��y�cx�z&&�WQ��ڀ��
}�sI���A�5 |8Pl��(u*�q�JR�x�wf�ܒ�\�����jJ���`�'���x�ba�0Q㟯��3Q��Nd�l'S�dh���2��GC�]'�^��ǒv���7�k�w ��੡��F��6/1�Y�$�����_�)@�e����Kq����A���$s�gk����E�B�e���#�f_69���Xe�������ص����fF��VB0�J��F�n`#
`���_��lIO�Fa��D�W^��ʙrZv���A�� ��Z����n��Yiu�㉸;�BM���UV{�3Q��3ǲܭ��]x���V��Ѭ�i����m�U�g$h�T�j���V+	ܲؐM��.�?��<}U+��5H+iV��e��Ym��5���d|ܧz�����^�| ��2Jd ����Z��HΚQ�c)l��S'B*f��-���g+d)u�8(�먙�R��\��ςQ��;L�������	��JC�Ʋ��*o���L�8a��.%w��Mv�"8�FB� PH)�_]�,6)ĭ�CC��yq�cd��h�Tڋ��o3���߷�Fu"�Jڟf;n�y����������[�Cqxn�v�2�]1��[�:�9׋�.7~���G"Pc#~ۼO=�>�o9d�Cư^I����(!�j$���a�C�w��wß�N��_�`��i�ȇ3�0�+�G�ݛ,�x��@����!�n�׺]�_XjZ�n��Q���9��{�����;�Y��r�����/�8w> jrp��]��IU�ۚ­	��x��T<ӅO(�|�+q�X�
C}�b�\��Z�}�?O7AЊs��"i� ��Ͽ�C�-�������v����]&����Y+��dZPDb�o�̇��'���x8Z5зo����+>�<��^�`�J�Ֆc�0�y��?R�����c��y��汞�}ւ�d���4lZ�=_��d�u샕,���Hr�&�~�e�or�L�������Dwͤ�cN����[�'����ܢ�×����@E����p�W:���̑Cx����W*�Λ���ï���9i.�XR��o��9 ��%hVG'�?{���c!���W����/3�.�k�DF)��VT��أN@Uu4z����7S�UD��k��`����y���|Ԥ�c��ʺ[6�,�$�`�Px�'UЀ����e���8L`$$Q^>o�A	�c>t�hǘ��ׂ���П����(Z�8�ǌ^l�mow� �$��*��fY���n9���!(�:�Pt����5k3�>&J����>=�#l鎔��������s4������@�&dGE������D��Ѫ,��~� ��k�+E�H�lތ���پ ���(�K����@�@�½y���n����"��aT0�B	���e�,�=���k�āth���CZ�7�O�>�A,CW�!�L�kn���z���M�JE��$�>e��gR��g}��I�-'�R�1��/�?\��kh��ih,��6H�,'��=AS��㣪T�!\n��Q���+�4������\H�P����<�2�r�ڪa�0�0�p���}�J 3��+�L=?)5t���/�z�P8���Xe����u��sח��;���<;f�j>�/L �"�$�� �+�&O���x����2�?�� p)�񎼅\�[��5/t�XQ��Y5e� 7IO�����B��d���El�}�$w�s�J�2N=oSu˶��3���U�s�U$��:V�>YG&��NS��4&i��v���R�T�����}��\pIU|s�+)�H�'���m����A��P�Y�f"���& �z��X[���tJ5e��de:[�ލwŪg�hغ�|����Pl�U�g��e[����ʷġ'�w��op��+��/�<�>���Č�5I�B�0x���j{;&q��M�!L8�I���7��O��<=c~����S�����ݢ.�������cI<���rݍ\�]<݊�(��Rv�SH�(Dƭ�e%"I�c��`�j��G��L��]�l���^��3��T�4� �q�70Ј*AN��B�[1%�#��nߵ���戅�e���U�_õ<��a��K������;�U�F`�����?;װma@fG������C�_����rI�I�����)!p�ʘ*u�$�1-pB�_��Z�'u�s�;��3Z��2�|�r
�����V�z>�gЌ$X������ �������m����5^	�V�T�굻���)�g��u�5��G�^]3^9�ĳ�2}{^�y�V(2����u>�>�vroQ�\�?���0�T�k�y�3�f����f1 �EI���~�T��`�3�ޖ��Ln�ܡF�a�O-g��o����T��:�����p�oAY�V�<ϛ"��s��Gu������)=qw�L-��J���wf \��$�����Th��$�h���������*/�*"Ҁ=�014�2�n�"��[`���9��5��������'�A7���ehO���l�J��kA즈��PXm��h��Za� �(�	�m�����S��Ry�y��?�$S�p��L"iwf�OZ�8���_+�A��V���%+镹�?mk��s=#�W �D�]"+2����������������<��9-��jv(2&�%a�0�L��X_Oi���@8=���I��u�m1��+w{8�k>~-������g9\b��C�D�s9���g#)�!~�l�^��*z&L�E�؆��dt4��P�(��P�v�����Fp�L�enX�I�^�1�f���R���i���8�IWtIGt�3�����Y��1.#d5A����������8)s9S��5�$GatE.XRb���;}O�1
w�꟏�J[��Nc;j�	J��
�jﵴ��A�H�tb\�]H�FT�?���0
��C���Y6,�*ϑ����`*�S��(ݖ�qKm�����A�LQ@OgR�*��!�1D�Ie`a𻛂����{h�l��o�@/c��3�������`��!��cWh��������|\�M��;�()߾>[�fH9C�D�m ���C���:�,j_�������p��"����2����l��*��S�#&��@�����#?�Y�.��h����N�{�����e\��~Y�}��YY�4����N�j	n����>�����CH�!��Ls����WP��/�^���h
��4S;�!N6Bi4|�ԑ<���d���q���^V֞�y���A2X���y�크3�G�xL�q��2�H0;s��A�+���UJz����j�l�K��K�2�c�A���$"=a.��6��#ݘ��@�D�jo`�e�;�6��2���U�C��Q."d}�Ny}!_��A+<�@|�������Ư�	k�b��R�Ow�[ ���x۪�ƛ|�rF��1]~�i�������t���ص/9�_[��K�{����N��UMҬÇ�+��_juo.&_)�|Qڢ�!:�q^|�ݠ��:���8P����V��+=�`'�V�;�Y)�/NV���`��k�V�|<d?�4U���hb3�� �����l���E�b̿O�x�� �h9�)�P!��������u*O�t���f�-�k����������G������y���p��������|<�7Z�BF�R�_��P�����/]V`�zo��@p'�Mڠ��i�f3GS�R	��D����ZV
����u�<��1,�0����D�N��H縨�y�z�K2�W�����ey@r�g�q5+��;��z�pZ�8��}�1�q��?I�γg�J$��H��8_����#V�p�t��5�{.g���!����Z���b[{ׂR���t��ox~a���u_T����%�?�������^�N�8�
c�Wޯ�� Y7������8�a�/X�/T�rK�C2�,�o�Ͽ�	}�G/��ݶ�|��1�����
��S��ѝD�Oa�<L)���/H��_��Ŝ =֗R28	w��~�#�v3�����i�ܙl��ڏ�D�1C�;��G�ͫh��_�(�'���L-�n�aJg[;�(���6�#�7���R"��@�8�9�WX,����OUe���Jȭv�8��� ��N�둯����u�rA $�HEU�0�������lbU�lEX��X�뿾�$<�Q�Y��Fj�����ʻ�{D#T�2��(���q�;�?�G,^1����y�J���CWJ�xe����ڟ8ze�y���ef�Q�u��N7LX1L�@�q��j ��Z�b[�T)b�V�	2R��0_��E$*��l�v��X`�Eٖ��U�m����"yad&�@m-D�E"��s�J��_�`~����2~	��%�H�<��QN�z�5-��l.� "،�z���c|!.�I~ �zN6>�_ɥ:�W�;��ƽ\�v��6�9�D�t�����=o��{�Y��x�K���}��	�Ϋ`4�2�6n͵��e1'6-�)t$�����]�G���R��ž��t�M���ņ��&rEG:�O�7��vb��Ċv���������M�Ot�޵m�Ј͡��j�X"ٯ�I�"z�rM;!���/iݭ��FމV�!J��&�w�S��$�&p������
�sc�A���ޮ��-Y�1u����`�_J$*$d�\<Bo�*j]i͕r�.��p@X��U��J�P�l��C���� �H��m�*���A���-K{�ǹJa�=��f)�%�^��"��K+��_/,+���	�:�S)YhTgr�����9��YwgtWy��髳�g]_jr�������0�+L���x�.���y��	<��\R�Vvtc�C��^O��3s�x�����|%`�Z�\2pd:a������M�-��cQ.�΍[��.���ڎ�q��l" ;�+}�6Hϯ�
s��2�d�ȕ=̈��uhW�BW�^SV3+}�P�)��7f���J+@����Է��he�o�Tv�?1\���J�2��b:�	;�)gӿ7���D�{���&���!�#N	�<iS9��â0~�X���MQ�	΄'�J�a3�,R���So\U5O�5������&8����1(�	b�Qq"���&]XD6�C���Lcfm{P/V40�S̞��	,�za$�s�7� ��t��6�B�C߸����̦*�V�1�٨x�"����7q�وK�����>�J�=�9,ʅ������������tǎ��9p��sF���x���0 �o���s�UGp���.�W�$����{��`���j(�R�P>�F�	��ݚ⹕B,���u�ݏ�c�\w "�.�$��M�;�VN���J�	���썀W����E�~�=�&�#���UZ3�q#Y�;��|�;��t��Hʬ��X�ޛ?�I3�NYnR,R�b!�k/L�����?���ַ����X$�P�����5Kw��zB���])9����ӳ���1L�"�2�a��g�U	���9+�F�-�5.H�B8[=EI.��Gi@Pp�x�I��W��z��os�ǀ`OU���W�ԕ��Ϟ �����qNW�1�����)� �3*�T�#�����tn�ߓb�{#��-k��z4oI61�v�h��RC���́B'z��B����H�)l\����H��e�:�#d�m�K�^T��=~��b�s���oE!�!x����I�8 �CxN��h���`#��v4�d���X��k�_�o�|9yА��=�$�9��uBݖ�x0�_�:'��}��]� y�oV�����G��G �0J�Ltts_R�R4�F���>lQ0O^bX7��T�D����Qpd`g���K��=̖^�Ϝh7($���/��-*TFl���	�����8�
!v�������>ESy����,86��F�2�����Vmt~߬������v�����	�,�� ������)๦���
�$�'Y�V?Z⺣�%� ��g'�A�am��9���f���/�r;��IGIseۍ��+$V[��S��A6*ބ�ˊdL�����Z⌊Ʃpgo?fܴ�t�!1��*�t���v"L�,nx�������r�T�m/ �$�-�� ���ubi/W���g�u.ϟ�xk_$�\S}j\���a �I${�������������iw��� D�&�v��#�#�[�{�Ǥ�^����*��$y�7R��q���8u��"A�%z![V�6���-�t�4�JY䉗�
���	3v����?�-�H�i�:R(����D���hp���%)ҍ�i�߉�*�l�}���?�O��UL0G$�S?�G����T����g#'�FĞ�#vǛ4��ߜy��s�FN�X^�C=׼����-�'Rĥ�s,�oR���o�>?d"Y!�1`��\�m�ճr����]���� ��(�C�OtAMș�ͷ� ZD��!��%��S�������W�m��1��*�@��S���],�M�g7��n���7H72|m�-����/O5j�_�ҿXK}����pѣK���~�诩1�m���\�{�c���#Б_fE(��ayHY4?~��7j(V,��`��i�A�o���i�`ɒ�(���G|4X�0D����#�{�{����R'T�JW�p�'ۅ3�n�8N`p�.���Ġ��}wO$��v�Z�I_(��J�Zl���U���1�\V�|N-���Hpt�
���_
T�Z���P���n*�|zC�?�����a�@@W�$|�H�N���]�(����R���9�~xBj�GYF�����r1�E	��GVU*�=�{�cꜩ�
כ����!.` �x��GQ����F�����/���vTe�ͺp6��v�㟙)���5�����M=��.��};Pt]�ͷnO���4ɋG�}���O�Bs<V�+1�xe�%:�#����)!�UY��A����s	^tA��wP|[�f���V��]��N��eD8|𣨿kB��?Z���:`������	_�ywR�,�L���V)nD�k���4����x_��j-�8 12�w�i�]`��0x���M�햟T<x�'8�VJ�)"�^��J�P�^�r(Xzl�WO��뉬����������_*HJ��}]`'7K����i��-E'N(WV`��dt��M}�]�\�	c��D�3veT��r#�H�	�<.�i:�����L�D�����J�5|�F`�,�h4�
���i�p���t�I��K+|��8&��~�A�_yV��+�5��g�f�*�'MJ��vrd<��?�Uc�f>�Ec�<ꐲ�Iv��Nj����<[������d�^}SY����f��׿��M�XMp�J�0�umX�p{�ܪ�)R[s�;������viZ#ߟ�A:�a�1II����`�)$���V�|����R��#Q� ���@��#%ڐ�x˵��5dy��;d�w��f�-��t���4�H?��U}�J�ZY�J8�+�A�&��~�¢��i��
=��a'23��v���P%�(����]]o��#��U��S�H��b�ϑl�3/{�﮵ӲA��* v�
�^�t�
�iW�zT�QI�Ў�@}hKD�)�O�n%�_�ԡ�T2���TH,G��9a+2t�=��<�F�%l�+�7 �+��'�9
�,w��P�8�-.��Z!'����:��@�:J�g=�4��t߀���pQ����Ѵ/���Y>�����r���[�x�qE��k@0)d:�س�(��<�X���Ј]~��P��ф,�_!���F�0���wI��ָ��N$P�f����/�
�L�RP4�;��y�D��\�]�Z����)IW:�����d���/�8�k���E߲2��p�ܤv�-P�LǢ�c�LX`��r�Y�81�����P�ؿ�Ń,МgTcb����yo��cu"��<����,�LOy��NT ˰|'�҃���-��t��%.mF�[�=v��@�E֒��{f�3�[���t-�Q���}�����C���;����<
?%"��g��}YhV����p'��he��;No����)eA 8-i/�4�`r.�Ix�&�L҃*�XH��q^�c��!�"4�"2K,8z����Ip��J�2є%�}E�Du���}5���-��h�Qm�"�Q`w�'
�~5.0�C�p��_�,�Ʒ6��5��:d��v}�y/�Ia�cx�l��E J��b����{�I%Gص�*W�1��M�J`(�ʃC�O��MP�=�#��z8�G������̂��GX2�S}wӤ �~ �i����v��T�K9�mQmA�ꮻ��~1Ϡ�^�����_�'�����3�o0���u�X��Y�6������_F�d�$s�-�4q4�(��.BB�oP�(���yA<���O`�lp�:�Tp[�D*Q�q��4��B!ZU�k�fF�E�J�1��m#��q��r+"4vǆ�\G���&�H��SQ��N�_�����.��H��|N����<S2	1��9��[���� P�#�����Y��닽����J����7r��G����\��	"�k-}�T(\�n�����H�7�!q��e�*�)ݰ�)�rL�,�*D,�a�ѡ���=)� }��Pc7A�5 $�%"KD��5A^q��
�)����;`s�;g����_��ze�!���zXlw�7��w��+�z^�8��h�͋�a��`#i��-�/+��C�R�^&	m�wrXS?�s�?PB>�Vhrï
0�@��IX�E���?FNv*ß��{���(0�wseJOh�h�"�������T�g��x�wa�N��c��J1ʃw��L�8��r��zpέ4m���y�(Ȅs)6{?ʉ���*�!c�K���'�h�5K� _�b�UE�oV��+7��)������茌g��Qo��#�R���
����"�z�7��}��J�ȊK���/\5��X�c1�V g~gP�\�x���Sᙬ�<���u��c��,Q���7�p�ў��Jgb;����>e��91�La˼J$�0{�x>��e����w����]Y`����+5��h��a?��B`�y��.��Ō���x\м��}�5�	}��8G27�?�"5FZ;�����?���t�\�KUW���)��?'��/�SA>����eV!��$�8��\�Σ��]�WyD>ؿ&Z��� �ğ�W$5��?�����2
TiT��O4)}���rG����N�HN׬�g��֓��Uq/��z�����H�{�꜌;�ըzQ	��;r��|vnP��U��(��[�k�bSDPe.q�l��W����m��t@����k�Ouj�|��|�-(��jBU�R6-���+�BZ������ ̦�_�e��l2�8{�Y��^����܊ґ����U��{�7jo���)�w�h�]��8So�gJ@�X3X�eW:]����vY-��o�%3�jn�c�|��S��s����PG�$S�ݑ�� 0ԅv�,��՘<Ȯ�����I\
�y����n"�Ʋ�5,�]n];A����J�5~p�S�������	'����d���bp7ZW�z-�l�QB�Tnj9V�$(�j���ㄯ}�Cg�*t ?�O֕_�g)-f��uѪ^�k���rA�]�D��_?���r��#+ ����,/#�J�����]�>�|�Pyf"�(�3�8�������\��}b-H��E�[ou��濣����0�pC1�L���$�],�!<5���s��?���		nP�,R|�j������N�H��v�O���M����\�7`��D
�Q/���I2Ά�a�ޫ��N��l��V
��a�@*vMs�КZzJ޲$�?I�Z^^�'��b(���mp�
KGɅL�R��#'I��?Aʣ��@�\�Z�C ��Yx�4�W�[�:�ʈ��j������g�7h@fi��aEɄ�{������4xr����m���K�}J���o���mh���<A�Mv��>bg�~�`�ќ��#�6�<�ΥDd�O��1�� �I�g1b�����	�2A��ǡl�"A$�w�!��ip4�៰\a���|��u��N�m@o���$ey�c�9����g��<8:�x�����#S�Oh˵��Ȣ��>�v�8ZKr���שi��=P�8�n�:�,!#w8V��{�v�r&��<�I͋t��E�J긁�w��Z$����Fp���B㲪]�e����t]���}&e��40�1\+<�-��Z�nbF��DR��`��{)���/�x3-������A��(��i}@�"�/��F[ȋx&q-� R��W���������~��I�_9�|!&���n%%�S�[M�#PAd_���VR�	���I��c���R�w�R�4-O]~l]���X䆟��O\Q��<��P}A)��	3��4Þ=6_�G�D]�
���5_�n����1�R�B|W(2]���y�$#�B6��w�� Mt���[���0��V8���?��˶�2+q.wW
M���h��Կ�;;K�2$ւ������:��{Q�+���USx�T���"!~+#y\H< ��D�xCH�[A"0[����2�����F�E��r�Ψ��Z �
�ĒϨ�c�ȂG=@�d�WY��4�!r�t�e�e^��	� r�ߔ�yN��^��:���P�TY�o�gB�g�ϙEz�O3���8T~��(���*���v/8T�B�����")���!��%���h`jՀh!nXZ;}�R��.I�m꩕�A�S�����N|��$��r�p�#(ܐb
Y��$��"Ib��	R��8���U�9����S�\�{��Y�e�٤���9�@�@#��@�M\b .#yu�$�G��%�&���?��4�:�VR��O��Ɠrc��m��t�����t�+�5����yOm�(^K�cݠ9Hb]��N��g\W��/�2է���@\T� [�4�[0���Gl�V��앝@3��|�P8d�䢗<��v�:^��<�T�$*�"n����GEuHhW��C���~�~�d��{�9^����f�����	������4���(�q�w���A{�4�Knme�Hj��n�a Gy���A��Rs��C�O����������'A��~��3�	�vgҏ.�#����pa�����r��"q26�pf%;��������ePb�z$��μ��ֆ�u�h[�`�Qk����.U�R���'
���}�>��/�:�げ}�ք� JC*5�,��p��/h~���bdT<L�*[aڳ{ṷ��T��@m�e�=B&�cu[�D�Kdί��eXgOcLhx�����$L�sUVb/;�)�ᦈ����w*Ɔ_�5m|Ш��<#m0���R
�Ѵh��B�9q����#�k2A���&N��*.��}��K.��������e�V��}u)MY�w�� #��	%��ϋ��n�׈��>?;�ə�s�/�vӉϯ��t��U�7#E�D��	�~��)��q9t�D͜u�k5���I����R�F�X៵6'w��i��v�W�7 �]5L!�?��ɫ	6f�b���i*8˲�������B
�\=I>'���\�Ĩ��g��v)O����
F�9�#��H	�I�'�I�_�(��X�<���A�7Q��d�����F��� �����!�1HM�ފ�+���y�r�w59��(��6��k���7C�D�5�;�&��%�W?Z��>��[�-�+� �4G��|I��Dl�+�Z�F���p�>���ot���	7���/v[`�ѻ瑷UL�A��t��[�l��پ'�y�)V�M���%���C�����-2qIR�'�V��<vLX�ߪK~��]`V�}�0tqO���u�����#ܩ�eZ`q��3�_3ű��d+���O�3�	C���������duP��2�ɇ�8(Z���$���6�y҃����'6A#2i�6��n�;�ƫ�œ#r�������{�
j�ozv��~����_���ם9���%{���IOx�@5s��f�yF;B�k�]Np�^�/�-�X��f��T�=����Si��mc�8���������5$R?��˘��o'//��]le�g�w�<L!���4w�ǭ��\�K��B�HT�y7�0�a����07B��ܲJ/�0�H�� WϏ�IoU��qe��ާ�������ʇ� �K��i�ʹ����wj	G;u��C���!�A������.(�U{�1�5�ؠ�:S(�?���ѿ^Y�Ac�
���$�J��Є�%{��K�5�9$��A�L*NZ8_�T)�&������K4Fƙ�>�F�g�$���ϸw(ė�:ى��da9�7-�h'GO6L������p�x�J�#�؝��#�#�������0������K�<J3��6�D�𼉭aj�:�����GY��|�_*�(�ȍ>�'���Ѕ�� W�3X������3�g�-���#�A~��p�|�D�-�ޞe��{5Y����������/],�\���"�-�XȞ�k#f��3��=Ԃ����C�Unk�p<T��/�P�1�#��i�9Mw���.t0R��Z*����r�<����<��"�{�Jނ��۽�v��a���hE*#�͍
q:�oA�ŧ?s��3�?�ʽT�TX�Vw�o ��Se� ��C����{�Λ|��ۢ�&�� #��vK���&+b���"+nN_d]Y]i�-@3�����*���sd���U�k)��瀢4��!�
��:�o�*���íѤ�������B��7��r��u��yi�!�j�
����u#��e�Y�} 2RM��SD�Gw,���#��fh5�쥋Q��BD�9Ø�(�w">�f�&$	Γ\J��g��Tɳ�]���6��_y2� �7�f�9y.��9�l��w��x��c؎����{��W�B�`���`D�N/��K��	D�4�`c.�������a�i;�ؼ'e�B�J�N�i�ɭ��x�e
���`�5 _)0$�l�*��!R�#���*��? ���%�x���T�}�;Չ��Z��{��D턍qxj!#@gK�3�\(�����i	�mv��GRYp/�|��u� h\U��%�-TJb�>���q�	��q�PghY��̩���J6	���H,Ζ)D����F���ä (=�}����~�&�֝c��dU
�0�n��\KJ{���E��W��_����{A�)'{���	��IÎ�_�ܷLOkB��K=ْ��q{1�֢�XU%j�'����䝓	�	�AW�^[����_�GpP�v�Pi��T��Jq�W���5V��l���t4��!��d�nA犺,+R�*��M�X+���d�D(�w�?�������G�����?|L�6�$7ob3�z�6o��d�G�e'�G��d�a�5@�i�8�`��5.����gU!�4�H�Uv5�^|�Ukm[�7�ٞ�������_�[6����`�k��D�:7��T6�D�색����oH����i0t% �U摢r3�/g�BQDAR��9��k�d��ү��cZǯ�� �D=�[��擁(p�7u�����-)}`�(4�.&f���ɟF�w���'�GѨS��gs��*�5�o�Sؠ:Q��Ό���b�'[<k �c��<��^�f3C������)]'4�/�8]�`�K{��i/�\�%a�x|vu"���{�Nn�Y�Y��h��K.ڋQDJˠ2�[�ˊn5Ne7kQ���YCM�8��;���O�aI����$Q�6]���q)i�c�̏)�/2�U
�
��#ł,��ý)���%���N��Μ�1l���0�:=��8�����[�u�����2Yl�LI휺�E:��V��Қ�������lL<��Ղ���ͱ�~�9lX�5�PGU�2����Hܻ��#(���C%Z����֐�g���+�:�H�*	�x/\~{0��(j���	��#��Sp'���2L�x]d��t��Q�����-%A��G5�hT��rhV�:���c�3�1!m�'�@-�(y�&6��C��Ưߊ�Z��q��/��7���T
���蔼|��M��œ�x;f��ڳ�h�t_;OрG۲:�v?0����01,�҈�=�%J�"��.��wJ���#�:1T�&;:)'*G��xJ���s��p?��Č|�h���1�Yx�+
ڬ��{��B��a�Rt��a���H����;y�ڙ�4�.��i%J��(�l��a�8mC�A��4��t��i-@p&��M�{"O������)6"I�D?c��W^������!|�T(�.��:�P+�`m�XE"_��zi(�ֻk���<kk7��xRM�-u��n�?B�|��1匷��]���q>Ď�]�Ԏ��my$��>�*�=��]�䏱03B�%�����=n������U�(����g9���&؇�s�
O�Ƨ��@�y��|ݟG}"	+_h��]�A����H˙KG�A�/�'~B�+Y0�`���٭��B���Up�f��뗪��;� 坂0�h}��@����~"�R�cð�������w�S�C�'���!���sU���)���%7W!���.&Uc��)�S��Ul�2nuKvƄ�4ܷ�`l ��(�/#<F���l�&A$Д77>'n�Ee[�ݖ�*B�p��^(�����J���4�k
_�G��m��%�d]!(��Z$�>�fɂ���$ｌBH7�����������!�*�~Է)H����%R��jd,�|K�c�(�Μ[�����_��}�9���T���tO�Bf��b]����L�`:sR������gp� 6��^4����5J$���I��K;�2���e1=��l��v�<t�}���ky�-~J�,O� Lo�X9k ��Z�T3�)L,"%\��2*��r�� !�?%�ǭ6=xjoL)I�����}��L�'kv���w��Տ趪M{����jL��7��oy3����=����8�r��ZO��Yi֩��<#�Y�MV�^\n6�������0�! ��i0;^\X�6�R
��?g缋d���I{vF�_�r��i{�؉skʅ�Bj��}s��,�4ć��Ы�-ӱԇ������9F��.�ir�S@{��U���f?��]/^��㝊�����걙��D�����FfQ�T����j��G�4+خ�C��0M]8�5>PV��N��F��<˥XsI���Vi�BjeAI�13�
� a{w&����I�4*��a>yU����>��̝� �s��/��!d��c�[c&/�����VB v�-+,�#��[k)p�����d�s�Z�b]	H'C]�VLS|=��#%�C�"1�<Pf.:�A�j��ދmsEڽ- ��~�Ɂ�q�^�ᓔ�]��h�|=lUO ħ�Q4�5Ǚ��YL���¦R�mŎ�i����K���:�\tj�G�Ȗ�q�R-��������D9�p$��$� ���:�3?SgaP��"1�D��f�z�;:/�an'�x񱌠�LϜ>�Yʍٞ��U���d+::�^�3ڮ��k%���A-�Z@w���}���q�cg�_y!�)m�-K��1A��	�E��9J�-�[Ⱥy5���ȣ�F&�DT������mV��KN��۟ڽ�������aY��2A�.F�,o�B���q�Jww�|k����Y�?+�́�����0���D��nv�P��S&�T��e�A���H��,�.�<��Q�
i5��
�0���@���MU�uE�k��.��cͧ���C���m;��%�E�Z@��������s�d�p�Sہ@���[����*��]y6���n+�f��	\5�v�b��q��[��o���/� ��P"��˛�Ģ�׋��
�wp�Wx�Qn�M���(���"8�e=Z�5�!�Qn}�0�I�:�`�w�������@i4�?w����^���+�3����n�!���0b�o۬q�
E8B�푤�Axa�jj��U7(��D'�Π�X��S�3d�C��ߣpQ֫��Y���*AB��Q�%F����*K`_�K�V�h�b �x�wxU��� ą,��C�﹏b����D�`�(�d,��=�z�I�"i�{���A,���I'�p��n�,ߍ�t�떁�N�SZ,Ywd:�r�\�`�^-���DW��ƁGf�C�BnP���p"�\��l�Yn����F��C�X	�	���P�r��d�N�Zp����< x���Cro���Y�Z�54���������eX����hIpM��	5�,F��K�ħ˵>g63��}�BA�k{ o�-�Q�U	@�?.����Rs`L��A�oo�a_��a�jT����bw%:�@�x�P����S�FQ������w�V��HC���d2�n�=����@b�z��`��˷��8T_Y�~�t�
�x��Aň9���ê, ��\#�Z��g���޺�0��G�R-3�s���Z$T��E![�	̲��s��.���UYoD�-��Ȟ�\�����<gaX+yh�h��a{�(%O�rbc����c�'�u��~�����8Y /y0�^��AQ���ڞ�ćy��y*A#��������F9m�H{M�x⻺�P��8{��Z� �n��ˏ��}A�����5d��ԅά��ak݀�w}:a,�%��/\�5&Z;9�k������g� �n`�dU�����NaM��n�S	��+�߶���
x�������5��w�vk&�y�N!(��l)&�ά�1x2�gU.G�0![/��,eI�
��QkV���S��'���m�
���s���l"�o1 ��#��J�SJZ� ��+?]��G��܇W�\�*�<]*ppġ���{���t|�>�g� )u��R�N�ZIRU�?E���q�tP���,
8�xJ#[" >� ��/��.�ܕ���aփ��o�q=%^ׅ��w#�;�0w�-��ceAs�L=�2��ck��ٷZ\�3�ur��M��+� ����)���t�aے��5�=�Ww��+��4C�9�¸�Q�@(V���J ��I�X �\�������a�2<}rb��~&�\2����l���(W��Z��+����tNѐ�?3�ZLq�(�X\�z{-�U�ҸC6p'�ٴ����&��X�5�<�����EwF{%f��������X�/��@�Aq�Y &�y��M�!ݬ��5	hn�����x|�7�����BI&NH�_0��>j;�mYг&pȎ5�	�xăw�&��۽k��e�bTq�Z�߂������)�.�8���S}�del� H�G�d�~���(�K��?ht{��鋮������p������<��/@]k �rd�C�4���yF��s�|(��˵� �w�HG���m�k���m:;k�ƒR�sv2I>wu��f�%JY9_!�3�%-�� g���f�Nۂ�G�&�[nMW6���=Y�'M/ yV=��hа��&܂q����E|�_���i=@��K�ܤ,o͌��:���J����H.n�7��V���V�p����7;�C�&_~�	B3�Fc;�'�yg~�� �R�{u��z`h~
����l}=ꆑ�`ko�콝��|)�k+ݰ������"�� 
#<��Џb�mN���}i���Zø�����(N?�Ȗ�;Z�
7̘pf�EɜЗ�ΐa����mz�(̇V�5��L�[�ә�\�s�f���a��%U '�T>@Fr��6-{ٌ�X��L��v��l�Q��Z\G��*�`���4:Z�	��+qU7}�֕8���i�˗��+J���Ł� |��̀��V��ׂ2G�&C?�O�Ⱥ1'���}E6&V����<[����Xd����ӕ��ܢ>,p�n6e +[[V�,s��y�p�}J��(d��5�Z��>��{O�o{�DX^0Gt�5�F�R=TR��c�d�!QUMB�n��T-��֢\��B�t��-�pk�(>� ���ѣ/���w��^j��>��]����-�6�}����T'���yF\E�9�	̾�ݐ�-I���-��M��iN`�$	�[E��D�ۄCpZ��]ί}Gn����I���>��]��#�gm���ܟ�u�˹�0!�p���8O��_;�6;�Ҁ�|��>�HK@lxuiV�)��	�&b�Y�CdB�5��+�nQ��$�yz��\��|�D�|��*��5|\�[D>�*�p��QCx��F�#�:�=5%S�wZ�ׂ<����|��J�e|�'�J���%�X�b!�
!�2fY�V�]��9���JzC)Z���ۣ�kF�R}����n�#�B��Sbx,x�_���j��Ik�r�שcIP1#��"2��aB�w������U��њ�敮�z��nmHY�����o��+ߜ��VH�P�y��P)��;f�f_G�a��� �F[3���<�W����~z{��&�B/�HǠ�S��ʻ�ٝ���Z�i3�=1Ғ$
�0�
^J5=m0���5�L���3�j0!=�Z|]�l	!�����3�o��fK"��@2>�Z,�.~�G�=u]M��U�%ھSH�B2AMZnO��4���Bq�2�c�����7s�!���Uӕ��N���y|-�u"���sB�o����|E.�c{�|�~�]s9r��ǌ��f х&@�Z�����9$��g���>�n�5��#���Bn���m�8��Vkc��M%�)d|�*��y�ȁG���%H���
d���YH�n��0��8� �y�3���[��\�߳<��c�[�J�P�G��I�s0߉�ҁ�7j�Lx�c������Bk�=NI��>b_SB~�X���Hk��4��	�Q����&q׫��P���#�� ���.�i��S�4��R`n���<���,n!Λ|�W�XK㳲z�ң�Wh\���ݼ�����>g�mԓ�uf�Y���E��3h*�T�r>�|�Í��}�@ec���E�ϧ�}�b�����1p��i�6�J�_`9�|~߱ѹ����іu�*�j��]<�;)b�����H�V���*��q��xScQ�TSΔ���J��\��v۾G���ZSEo���RbX|@N�8d����V_.q�nx��5�g��-lևy
Ez#��Z�=O8,u�\�7z���hF�6Z�_m��ʪ���Z�%�� ��6�s��L�eNvC��d%�W}L�����Lގ%�_V"ߒn�I� NIG��c}AeJ�t�_z���p������5��:q�$��EeT�=d��)q�w*����A�4F��n��b�<U�"�n�K;3� �j�;O�]�ޱa�_�a���eC|L�slsl�!Pl?����}kM<����ϯ@<�!_�ޚ����aX�s����$��L�Q����JJHW){Uflc��O��mcy���Ƈ��I��f�
��n~Q]�S��޷���=T�S�Fw�)�Qb$�y$�jVlI���0��}��6�O}�x�Ѧ�œ𜬺p�����2�8�2��y�N#L�H�����}�W�[.,�z��ytHc#86^�7�T�/�
�D���d(Q��IXը�T�cjQ���ײv�ډzkX��9$��m�oZ�3����U�q$�TΎ�2����:<���_|���ᥬk�'sl�"�S�)۴�>m�B�ئ���Hj�t&q&������ZjҌ��OZ}�IlF��Ϛm[��γ��R嬼b�s_��{|6�N�V�++Oa,i��4�3/�0'��_0����G�Sz��P(3��Ēbu�eȇjw��c�F�{/��m�Ckܜ�,�7`��T�.�����3�����7��v{��R<��x��4 '�t5�C�'J��Q��@CU�'�<�8��5��c����� H}�s�2�W�>I��}\��D�^���e�e�(�8�	�6$c�	g~�HҾ��	��7��ݽ��K��~���(Ƿ�ԑ	������� �2�6d
	�<�����V�ot���+W����غC���H�������>�"Q7�"d�4�qƴ�5+��,i�I|h��G�Y����= �f��mI�[��,7A�?3e׭��B�-���)����6�"2�-T㶢���������Y����Y��[]�O�z1�?U��Nn�ّ����	�P?�YI�@��8�gW2��Iuj�Ғ���y�f��"R�LL�㝘�q��d6�MKi�
t�h�YЁ�%!����Umʋ��Y�Y£�PF������bd/��[d�m���T���z><�
�������}�UI��J�u7Ak����X�q������{I��nɣ9�d�o/N�wvSosz��ڟ,/߃'�%�L���W��$c�>SL���)h%�>��=��_��rc�^�ۄ�:���\	O
s)��쉹��Y�VWb�GW�ߥ^�����7����
WL�3֙�a��]�"�����=LK��{p)YJ�2|L���ʮ���=c��Gy�P&=z�1�^�j@�������C����v���Ab�r�F;Kޗ�_[@�y���,�x�i�$aSe�'n�_@-=TZ�7���-��S��i_����
	~�2�iV"I�����Ls��'�Tn�]y,c�w3�ƾ^^jѴSF��K���	GlB�&h�(i������I�2x3?0Of ���V�e��i�߃$���;(zLߙ��z��8X���~�~i.�8�~��y�삏���1�[�A�+�"�V�L��M�c�3�O��I����鯏4>"��r��"k}��ۙ5�6�p�UiL�2=h �hA�����uw�*#���t���j��=S9�ю4e�"���2g1s|��׆#�_]��7m��-��5���$�9�����$gN�>������x��!��K��P(��J��}2�K=>Q��������e��Xgb�e��θϻ�=�'<4�H�Bh�J�ϳ�;5p�2AB�ҩ�*�x�}J&^�߸) ��Pz���@i��^Q�-�os�Rs8_h�E���j[�Yfx���)T7M���\�'Ԣ��	��q̤p�U��$�� �;V���
�[��f`OTc�y����|�l�h
k ��oq���&��n�&s�; Y����EPe㥰>��?�а����sd9L^쎇�3��8��|U�Fp�zU�-����AHB��':&��+w���2*����qu�1 �7�K@���6!����(��#R��|u��}Ǵ�j�r)~�g�ၢ�*��G�l6RΊ��2��pɡ�7����ɱ��OF	*�4k���Q��" ��/��P~�t�a�����������*��
�]*Fb�����mc���d�d4|رW`:J�W��zB��q��\�N f����?R����S׻��j5%�r�]$.��eȴ�T���x}�Rc"�)�u��F,%&��� mv��΋�)�@�s�QIf~;�]�ǧn�!P�K�_gz�G�Is־W���u
��$2Ӂ0�W�펠��b��	�u�4CW]%롁g�tQ'����I�N��˕	)� ��}Oc����L|P�Շ{�=)�n3^���sy"�Ĝ�PLhX���9����nx��C>��V_K�]��E��N��/¯)N�q�{=i_x�^�%P�H�	%�3c�QA�[�K���\�+��B�Ti�8g��8K�S����:0d�⿄[��=X����rm���(n��o5��^y�~2il�L��omg����gw��`���!�)���.�&-�A�s���9߁�]�A����a���ړha4��!$���g����M%n�5X���q���a\�V��Inv_膚Pm��Ԧj���)�D��P�֢�m�?�,{l:�q�V] �>r������.}�FD�V����_�%���w�w�̰��}�W{:�W'ױ�so�Q���)uum��P���%&��2�����G����B�E�`��W���0��b�+��mo��55<�)p�6�=e�\Qw�La�塀���1���=�֬�lR�/aR�_�S%��Y�D��\��H4�����3B.F�Rh��ЏS��##�����4�Sg�-�n�-��,RQLT�t{�Gby�Y���LF�h�<&�^|�lMÜy/��A���j��'\�,j!��M'��1x:��y�Y=M�����U�C-05�]����o�B�J剳���"9�	�i��Xl5't��I)SW��0�MP�p�p ��L��M�p�2wF�.�_�O�B꫼�~�������˼�E�V;ų������|M!�R�qأ2Xv��M-k�&-\ľ�>��Eų<5bn�Bpa����L����Mqc��r��k�i�Oa����ǳ�v�?���)���O�wwQ"���4N	B��!$tk�B+�X蔺?7�}��Ѹ�0hs�*| �	�t� !f�p�.A��ƛ�O\\���T\�G̢	G��?s �d���uE�Ny:T�1�ϔ`�o[�߳���]t�D�$>��֑�'�Y�S���/ܝ X�Ul��Q$S��M6���x#o_S������V�^�(�����sU�"g,:u�������1^	+\�;b�N���I��A<�.�m�b��*���&���s�|5��FH\^B.��V�J��H1�8���3�a�uٍ�<�"�aH�1ڰ-L�TP�Ȗ�,xwWM����ڔ6m��J0�,#��eR�VN����p�X�<�)�R9b+W�G�o�)z!K+I��$8l��8�p_
-L��d��H{����tq�[�o����榮";|-{3B��Α|���9gU���ph������R6|`6H����:��˻� d ͏pEё��&�]h�&]4[!�?>c�t�"t1���z�HE׎�Z4�8��H.��8�1o��y�G?��DQ 簌�rU����F��Ш�A7��%Z��̣�k������4�*ӈ��2	'�+��s��[���O&��$�,��q<1s�ҧ��{�Oh{�x:̙2�ɹ��<e� (C��u�^�5c�(q`75�
�V�U�v-}3�8���@ew{n	8�v�m�kv2�^�i	Z7(ø��R]�%/$�đ+�O�G�#R�=F�w�tfQ�i*�ή���8z�Z�iA�>T\L��2�A��@B��0��tWb:[9�'L�y��L讪�R�,�yD��*u�����?�FƱ�u�����Ub��Uv�WM-1��17�o-�ҊTy$�F��p����I��I��'�2Y¡��=հ�Z��n��Z�ՀԦ6$��u�C���F�`\]!(�uX�a�tva��T�0Kلbl.�[�B	Ţ��v���s@�6:��	�G� ���|g���[�80��E�,9� <&����v^ӁL�!���pd�U���o6O3��,���p�F��].$r�Rx��YJ�&� $@6�vo�8�l�m|M�a�/x��H�s;a�Ֆ,2���Q�#�|��>19sz�ԗ)>q��Z��_W�:ȇ^�>���{{�误���
��
RT[Z���U�2�.͠��U�Ú�/�@���ron*����!��`���O�戲�v8K���Y�~�R;~�;#�}��?��$9l랪7��Z�5h"+Ȕ�y��&��	�^V/�}��X�~P�$�O�EEOcw#ʏ�o���ɼ��q��{S�{���)�[p�j�,�/�H%������y�(؍�I���J����cڏ��L�D@.�&Q�!\�ⵃ\V��[�܌φtDU���!���D�I��k2�h������r�R��y���P�3�f��=z��L��*�����14&�J��+�]���o�m�-��Nqy�+� +~7Z�^�<*\ek(X�T�bmg�_P�{��4��I��)Yվ/�{i�"T� UXea��	�8p*9|�@�"�M�	�SN@L�"n<@��+�h8@Y���:gT�a�	��Z|���Nq�鏞������>��b�L��f=�`�F��ŠkC��vDэ|g�EhW��U߼*�/ח��r��Q���xS7����0_Y�_��ųx���*T�'ܔ��J�B�e���kd��� W
h������kK��O/_�5�$�~Z��t�/�v8�l�?�(��eNu��_�3�{�Z��99��B'�{���(�8�x����f�N۱U�W��1/�"X7�Қ0���w�����>���b�x�ݽ��kE�\��p *5��=�v������7hR֩��ź�O����L^����Ě�sk�&%ٟ����r,K~�����P�=`�R����X7WA�-k�ˌt�W�Ht��\pa�Z�1�����گ'���`��%V�V�#�ص%��f����G^�rk4���_���˦0%EZ�(D��Mc*#{̵��I8
V��
�j[��]�։$�VwE���5���c�b�	��n�D�c�pHnA���Ms��W�J����Ϳ~��Xf�u~^�v��D|�Ky�?,�D��͹}i�X�tii���Ԇ���H���(��|��E�8_���Eɞ{h�e`R�W��?��T'�80�"2�����C3?n�K@����Q�eD���1ú��* Ew�=�	���bTD�
鰱O��7�wt�bXx�`�5|ߟh�"J|�f@���_�"[��|t�y)�lrP��\�Y�S�X8~��I���X�?I�ӱ	��J̗��""��� �="���9�O��������B�Ћ7C�ƧŎ���x���K������O���9V�ޟ���ۧF������ ������#Z�'K0kU�s1�]!��4���/�n�a��T���ɂ�
q�k��NQ�,��ûֈ円��]���ȝd�%���Ts\*�%�':���w,I��Br�w��@Z`I�Mί>����0+��
���Rӓxb�������J�bP�b�Ͱtn�˴�����ٰm��=q-��t`z�����J�(ݢ�ʕa��w���a���I�$��W�h�R�ÞP�t^ƩkSr�U_3�x>�On]͉ߍA�+ -����V�7���̋zQ�6��E@��rD����������ƶ�s��8�%�l��'�8��dOەU�w:`_�i��W�+%jD9����늁u^� �W%{�j=�>�%O'�#�����������%�Y#,j&e�wH�а`�M�%�����~�_Z��Bǜ�
t�jZ{[˺��2�FK9%"��_��9��%:m�	��a��w�q��o8%9i���\3z0���a��j:f�e�ah�0�Έ�X��X�\g����ȱ�.��*�p�і�k3G?8���?d�0����xAC�a���y�߹���=��w�	�/ G(hm�Gol�B��xh��r����}Z�T�(�B  �&�{��K�a��}W׶�\4�0�����7��ݗw.'��SCBnP\Ε��ɣ�L�~���Yuz5�"y����S���K�K�;	;̎��a�mҡ9.��ʽ:���UD� \�h
�*�	��u��S�榼��]&x��LCIdX{�[ޝ�*M��2=�/epX�4���v��ϝ�������� ݨT��u!uwj���[���~���R��k�y�q~���W'M�R�����9eel����lB�,�Q���|���MW�PW1UhA�fU+,)��8r�|���
����N�����Y�/���p<:�@{)������O���m�O�Z�x�/�ppyÖ*^"2�mA��@����37F� /.�B��4׍�t��Ɖ)�MP( ��D���AƳ�!�wk^�zS���?h��5DWSF+���77�y��:)�> �\���WBB bj�"�����f�:�.��o#��]�����	��/��/_h��R�*߆�1�k9����إC�%���)��z%&���E~ԯ�9�e,�n�7��^�X���R��N�;:ɣ�}�38�V�f�R3����:��S�:i�N�m��g�7�خ�Ě��Ob�+ҿ��D�'�h35��$t����7$<S�I^Uz�YF��49�J�7�t����c2�d��A����O��a�:U�.c�4��q]oV%�Twl8�r�,�/�aُ7K�����P
 G��QQ|-_����M�L �:�0[c�f��x��9]������o�]Q�]�5��"a��V��}W%c���6�2��e۹�~�'���+zGi�>��{=e��'+���Ep���#.�6k�� e��Du��*j��	ɚ�盛@��H���Iy�i��������r�xb��r�	3C�#�3��wS�+�or�1r��f�T�"�'~n,V=��#�]����ǋ�#����\�-���;����R#+d;�$�&�"<�-��z$�n��u;E8�_C�_Em:�*�5��
y?� � EYh?Ё"u���!T�����戮��Da�a�+�9cVz(Wg��	�Q�1.������e=�=�v��j�W�������9�Z�1��ʇJX��^���u�N�?���9���������*��r�6�aP4��߸ѭ��}(���]�*��Ha��t�V4���d)���Ҧ��F�f�����9������9��
p�$�&�R�,��ZA \� �
�g~������ZCcD��@��ßb�=��}K�L�(z������̀;���	�v�mdQ�W�͗�A{��t��"V_�xZ���O������� ��K�l��������_a��:�i��5����ҡ�W�|��<Jl�غ����X��������6�nz��UC7��2f��>��s�c����F�w?�Ej(�9��]5�Bi�dA�Ҁy�&��Lam��E*�<�����d��[�h�-��B���ݺ &�%�t���-��ɐ8�J#ë���E�����
4q�E�#/;c��qp��_{�L�(�.�r�H1}ರj�(J��H�Ș�yL�g�N7<)�s������+�u���񁮢(ΰvpEL�i�L��o��ۍP��3z�!|��<fn���a�����gS:�/�x��ň&�(�����I��2�xڐ3��q�&k��Hl�Ɓ�#Ny�Y�]÷cTB���F�(?bfD�F�O�r�'\�(���5V�
x�MOs��Ȥ����y�9)sI"V��I�������ـށ�)�����H0u�*��ȕ���j	�����Ԓ�;���K�J��en��z���/�r9%�z�����v9!���=��lY�پq�hO�1ś����!�b�X=I��J�n�N��&����.Q���)9?��69�8��/����`��؂�?�,�c���{����0_��n�Bm�L����z�%i�����Py���P������ӎ�+��M�e[��ć!iz���m�=��{�ђ�Wo�f8�Yu���.i�{�s�7eTx{���U�?�(�RY�L���P�I!�����~1���$�(Hi��S��x�b�n`�	���J=����r��a��~E�_�{��_W�7!}q2�\�tYO�������p�� ,��ٰB	0z�D���:w���;Ip 5�mV�����s��o� C�j��ڛƵ��u��;v���x�PMR	n[�KnϹ�k�'�H;??���
���8_I�H�ןߣ�\�d�2l��J3����,����E�b[��1 ��1��<i���JRo��-᪹(b��۠�i!��ݩ�|Qc 1�VUM�خ�v��=O�g�Y�Q�0�F\�@ (l*��˾d��r!!�	����Ib~�0~�'U��:��3>r�_��뫄Q��!^d�s���9_���{����ə@l�''��H�#L:�*`k�������xo?����P[����OoA�I��/Hl�1�I�ڒ��C��X��·�2��z<�(��hR1�C����댾��_Rާ�x�0��=k��Z���K߼��w9����Y�����~*-a<�P:��e,\P�61�@$��E՟���9�{�B�c\n��\o�3�7�- ����~��GB�F��4@A����m����;�U2�@�ݹ(Y��qU�5�-�uGʼ�v�G��C*�;9��ʯ_x)�; �OE\� *�8�v��Z*��%y�Dj;�(�/�ܛ�C����0%�|���[e����Jlґ'�#�]�Ӏ��Rr��e��(>�)kVk����Ӏ7�i�^-�y�7�8Ӕ��v�p.�NkȽ�~�wb��?�M8u!+�,���!g��/��gg6�h���>o�n�!���0:����WG��zL���
h?���U�֡Z񻍑x�P�O��T�-�~g������f��՞��5����F7\��*d��j�$���Q�������LX�t`K�~�3�M$B�0?�k��:�u9�c����z�4n�`��T�-������u5��]��L2�$%tnY2ן%S)`2��d��{*�C]p���M�a��#���ݣ�x�ҵ��;!>Y9�@����lU_���FӞ����k0�6��ya�ĕ��CgC"���������$��N/'S�C{@��˖��@7D�`�ͱ,��� A��.:՝xq��r����1J�oYjX�Ŏ*�u�jV��Y!�ᶆeB`�?�����*����ПW�<�J�����c�g���u,"���gE���+�SB�����,c�{LU��!z�%_��T
Ҹ�G�ށ	жU.'�[3󥯅.cxJƌhS�/tQM�Ě��BZ��n���͎7dJ�ιY��`#����rM�vVɷ�&6r��1(�~.y�!TX��?xLF��|@v
��>��O�n���CQ}v�P�a�>4�+�1�(H��J���|�N��
���@kQ������������V�;?��i��\ͽ B �kv�5� �k��Z�����N�\�S�I�;�YίY��
u|��:�������i)u=�?��Э�^��=R��LVd=�xk��ҙ$6�
�F�S��سv�Q�E�\���{!s���)q�L�ȶ}���⇫̱l�I�U D�O��Lz?s��y�]��&�����?�A&n�7M���oMF ���阍��C�tq�,B`�=�6R+`�؝)�N͂4jH��q0av�8���G���(�.2YLoB��dj��6�{h�;������wL�@	��E���D� �
�� �8DL �-'	\�Nl�ob/���exdu�F(q�uL;�1N�q\qhT������~X�j�|=��	} ���#<�t}XA��P�A���>��9S�G]r��m|�_�w_��COw{ʂt:W�jb\s'��B����;���~������M����<�%j�4˜��LSI�Ps-T6k���Ӣ9�bv�����&�`����^���q$�..���*П�����i7���P��N&;�&4��f��M�չ�yj�[��'��z&�YJ2NZ�G������4�Ak\!����˵a��E�蚈6Wlz^8uJ{�ƌ�[�b���B`�:R�h�R��rր�U�R7��~�܍�Э�0��ļs���xAo�͊�$�L��r���-���'Θ�׎fkcϔ(�� �z����,x�/dOGT����z�~��!Xn��v��b���C�B�?��h6�K�$����?$>'^���d\#���7T�3�ú�s����	y�P=F��QG�ͦU�62�M,�G��	ѵ�.��]�`�s䃩G���g(G���ד����j1	
��f[vp} O�����"��G�|*�}����R?C�{2�r#�t��=�]Z?iG0�3��j���(���6뱰�c��h��ִ���y��bKU���o����������f�#_oHxʫf����9M_h�楷zI8��~G�M�|\�����0��J}��}��N3��v�2-���p6F�{���.g?�tL��m�
�j��Ï�F�87��޺#q�6z���xM_j� ����Af{�\����_!��*�h��G-�a��W�������&�}Q0��8S ���Eu[���ќ�/�ϧg�*q
�}8v֯#$S���]��˷��r�E������E��x�?2� ���ͯ��F�ju��&գٿ�Znm9Z����"0A�!KO,�ޟ�k��1JR!��\�[�l	*&�ƛ~��rp9�<r�H������(n���� ����h]�w�:��ߣE��Qd�Dd�Xǭ&L��{�%��MGE���]���{��5�r�}d��}W%f������zs���@_�$��5�n'�(%�����u�D��� �>nuĔ1�n��#��+�As]n����Cf�v��z��S|O�g�bYl��͐�1����Q����x��$�3��+s��D��+�(�R��A�36��40� 
�t&��˜dТB�b��f�=\5umeB]�k�=���n�ƻD�15ҕ��!�SY��-���G��#��@���`���'�e�8�LF����=;eTu�1��4���RT�i~�����=����I��		ϩ@��2qm�/�!�,^��}��,��2��[nE.M�V㭤�}���`n�[�.>9#@/����m{ц���:ѫ=u@f�����vl\A�Ѓ�Yz̟v.��J~3!��V��*��P�������ZX���ǂA
������_wi���YYo�������̭`����)�ts�{,�Mu��&<q�F��gG��E袍QH��z��Ҋ  d�u��7�/��QO�~�FQ��.e�[��a�pc��hZX�GM����铔ؙ<̑=��J���J�^�>���C6���<�T��xe�S��^��%����Bq���_Z[�X���C�W������İ���QA\mZ������G�~n�U�8ՙs���;K�-�9%G�ԋ�z��<�o:��"�V��2�(A��� �sq;�|�vG�o������p�����5�|��wo�$T2<<��д_������5�sS3>k�Ta���y���B�%�#R%�o��C�����^����ɠ��^Ў�ӊ��?5�6�d�8��X� ��g��N8zȞ<Eu�Fm�#�AI���������
�r8��U�D������6�'o�7[)��צ��/�`Z !�(���t�+���V�<�c���$�?|�3�p`��ŝB��K�ޔ���h�u]@��J����P�;�T�;dW�GA��T2q(����[�{���*̀����`��Ͽ���wK)����Ƿ�l�I�9ɺ��r	��������`ȅ���Zv�8.X=��Oz��RL��IM�)�]w��A �gw��Rbj���
�X��mo�,�C�$���"W��k�B�Z�$��1�R��_������D7�Mu�B�0	�ww��>��Sւ Au�5������)���i�1G�
L�ܾ��j��ȣ=%��o0@��wH��<�q���1����2{��Ml��"����Z���%=�/X�S}	շ�{�4(yIaM��H�b�U�Y��⢘8�����szM���6<��w��
��~E�q����e(1�+�<Z��3D�[���g�J4N�}m�,g�\�X�S��1����;]m���+�`<|i=�������c�� �N�B�9�����k�0�u�+����rK&��TS�rUF>��[����u�Iw���7r����;�&Y	\�G�E���ႁ�����Ck������H�(�̪� c�0�OkǠ����NM�B!��9���N����f�>m����,��L�R���B��j�xD�p�/��{�1G���ڐ�d�7��1�L^r�3H[�.�B|X��b$�.�Z�)���.k2A���`>�&�V�y���IdM���2�Z�4��dϻg�~+���ˢp҄��է�0�7�S>W*�O��;m�֨�T�g>1��O���j�������Ve��$�]x��-��X ]E�H��"giT�p3�i�hD�b�OŅ�����7p+d�4����lm�<�P��rI�Q��^�E�&����0�۠G�	�*$��|�6�{0)�����f���+��2;Ν�9-:�0rV���[���/�U5����'��l"������.]��o3��5���Q�R�/�z���HJ�d�:����kD(�W���J����6l��0@j]Ջ��>Z��bf�:�$����P�t�Q�>�� �Cm�J�6x~Y��!.�[[V�U��c��
��� ��#ۚZ�48]V������Fq7���)�^Z�qB,!�Wi|Zy#�*^�������X-}g���	�%��X�EҴ_C o;����D_ú��q+9K����[X5�)��XB�+X��@P:��� M�h?h�;QL~�K�Q�S�`��2I�e�]-���I�8Q5�"c)iQ�6К
X��E|J6��9�s��AY ����Zdz`�B��dh��\��(Ó(�boDfH�/.���� *��!k@�g��xX����ݷ\�+:�y5R��6:��?P��<L<�&A�%ڨpjh�G���f���e���H�A��i~u
��7;�\?�
�%tB��tg+>���B���Ea�Q9>(9���a\�[mqIM��NF�"Y0��d�3�W��;j'�,�+%��f�?��
�E"r��q��34��R:�|F��;�/��C�i{/_�d�w��{�p�������wU;���f1�Ϛ��~��ؔZk��Q�޸�V�'�]����t�k����B��$r�W�Bu��/�!�35"L{|����/K��D��|�0�JuK�����:ӹk{�7CG��O�7f�rW�M5�K�-��6?]t�aN��#�M}hh\~p��2аP�==��@d����4�nC�ӱ�zi� ��U
SA;i�`�I�ރ�
DC��C�����GSԫi##��w`Z���qM�L��lʝ����1��V�r�Hr� ^#����9ˤt'<��tߘ���I�[�ֿZ��R��������ni��޺d��z&j���q��Vg�j��m��.��zӬ�?�L���>��q�7���J�k)ܿ�!Ͷ��VyV����)��L�6t� ��
񝏈Xe�j=�V��uJ�_�6�{ w��� �O�2�~B��2JW?��ѱ>Ӹ����M)����_�eZ��(;�cy/��v=�tL��V��f�:�K�U��h���~�(�{�}��u���*�S5GU�Oi��5�o���s�IH?2������j{q����0S�B[\�ES=d���Ű�ΓT��K�/ș����2yjsD@�`xL�[X*:M}'C��<�f4Q����A���L1���mq�^�Vq�U9j���v{>�L�m�!�������ى�;��+Co�B����֓�)P�P�����:Y�AG��/x���wӂ�9�S9��w�Ŝ�K;�&�9�wH�2��Vʲ��
��~�����w�+?�F@�w ��o���,]= �I�ƀ�H�K��ȸ�������H3�2VͶA���ƾ��߷���E�9I'���M�����	�F��a�{0�-��ծ8U$��C��ǻ�"c���1*�3P�3|��%�?
���Y�KJ�i -������/�ߣ���o&��8�7�����n��L��t�/#J��<pk}G$�J`��뤏%�����u=� 8��\��6��(+Aۻo?
a��I��&�>u�@m����o�- ��`����'�%ma�oI��^X��帾���A| �z��ZՏ�`w%���Q�̖.2*���E{��J�H�	��8L�=�x��*r�B���V�dj�����fL�T�,�TS��,�/ft�}sq�e�ZC��
���(�n]� ����ڽ1M����cB�5VaY���O����z����AJ��H;G�K�!�*(}gvp�BU}*��^�wMy`���ЈwIx^�ɵ�ikK1rLjcOX;�����0?}�*��~a�Ѷ���1����\�"�.��.	]K 7u�����f���[2�NiV���,��!{�-�m�
8s���SH��_m��[dj5�Y~U�1[x�FQn�V����3��"W�����H��Vv�W�����8A~�Zm��*$�-�dR�8�ӊ�a�8���2�tR��ZPϛ��x������ uǄN=;�5��c�䜁�ۿ-ͨ⣢;2�խƥ;����;t%7�|�~e�Jq>�B�7�i�-h�X�Ds�<w�ߧ��Ps:�9c�!
���G�e&�̸�rW
���!s1�t��c�w;!�51?<#i�*2��Vx"��`��oj���B0 ��k�2j�p���}�ʹ֦������"f�kY�OQ"��Υ�~7{Z���1�� ��]gI�o�F"���n:�v�ǖU�����g;F`�}�d�S�D&W�c�0�W�e�7YNb461��L�	����Z���V]W�{]�#f.��%�|���a��?�u΃�|����w�+n���{_��q�S��WqS�ƛ��( �M�(�:�'��j�ĉ��/&�F�yҚ�	#�ꪻ�´Z�Y�գ��f���6R�-�j�&έo�OR.��㽶�vƄ~5"j\���L-h�=��n���fg�!(��8���)d�E�ץ�P�<r�%��UYR)�~���ǁ���Nؒ�� b-�߻���C����-��E�I���`�>����W|�)y�YH�jI��~���o���	rڙ4���wu<x�Q�\����������?lH�&�nNtt"a���'uik2����Q�Rh\ ���K�H�����X��K���V3e�A��ׁ��|H�&�Q_.����1�>c�b|8�s嬕؉I��Z!��*x��,).��%y��@N?�9�0A��L�١�5�����/~���v�5{�J����v��a(�M^�x�t�m�vH��P�4��/d�E��j���7t�4�n�/ե�U&G���:��(���T���YRR0۲^�<w���w,�C]�[�!I� ׈%�����	o��Be!��)�#���A0�ˀ�pK�ѽ�G]�f:~A{	�t�3�a�H{=&n������J�#F��Ĉא�+�$T�r�.ryc���"Rv�{y�Y^��q�Iő�� ���a����"|&����U��ڍ��t�S'A����s��Ʃ�b}��=~6�0���AŻ"k��Aq7��o͕	 ������1gg_�<ů��M�!i��՛�h�uT���U������dm&��.���?N�[�]�>���B��YD��p�5�5IV��2��Q�Ƴ�����c����e��+0��x(��f�al�d(�}d|���dR~�>��N��A~��z @��D��~��Y���SƚG���XE�Cp�:�P&x'Λm�N�,l�6L*��	z�T	�׀�{v�%N�O�hb�?�j������TL��(82�^
���E��@����Ǖc=2��62����oۖ��"˗?'�T�1��U �Kg�T���|�_����5�1��i)����J❘1މ�	�<f4�"���]�R	�[���'ܻހ2���[8����-)��P���Qʋ������k�Q�7��A��>�~�W��o��C ٛF��Jz�����n�J�?��,*�z���J*
*�Բ�=��X��\
�����= _�0apqV��O���,E�@���i�:�yh���Y��P������П~\���K�_D\v��*ShG��j6���p�=�Z~݋6c�[Ρ0�I�z��(^ul���^���SKE�#h�:H�|-Q�5LOx9�g�Y6?뗸SX�o�.�z�A��mnj�=a���@a�(O��#�("H~J�r�3�^��{�&-��:;H��W� Gٮ7)l����N$u��3���>Y�G M�j�'�k�<Z^,�N�ı�0, �X��S�`=���DV`��iJ�y
�a�QR���!.P�R��-�?� �cxO�W���#�W`�:��Y�l�<R�@{$I�CQ��	��	=�)h!��iޱop_ƞ;O�|+�p�	 �?c�&�A)|4��O�uf���S��4G3q��Ã?O��̵u"QP(�+��(zC���\��4�d��^#�8m]�ao2D ��.@c�(��H<+�+ۘ�����e�M����tπl�t^����rRa�OЅ�t{�Q��)Ȑ�%��}��G��ͪ�L��@�r�"�r�w���- !�V��2h��ER&FG���aFr����<)��崙�vΨR_��
��6���_������2�+���OD�k�Jil�|$3�����B�E�N����҅�G��a��!S���{�?i�#/�+�j��1��KR�.8�;�e&u��m�ʼh�u�IS��^�?JF��*����v��vk�ľE�+f���.D�YoW�ܦ%�pB��0H��n�I#|��e& >8�%8�z�hh�j�V����Q�� �)���Ā%O�����$����b�N��d�[+�j��"5H��t+�9��Ъ����@���nu��N��7"��j^<�9��f�/�x�C}�I�T*��?j�kX�q�U�,��g���1`�U�'=��G�ޞ�m9��3>k ��7 �3gW�]�P,�{&CѶ�O�-�{�����ՏBqi�f'��P/����P�)�Xcy��k:; 7Y��W*)g�%�ޜF/_z>�#&̽
 	��=���:����;K��1�tw�"�-5��ى�6G�K������X�ܗ��������a�����P��:�|6�su�S�"|�2,�o�<�}\�ĭ>W�x����x�i/P-��7"^f2s�.��U��w,?�3�? ~�&X�k��$��h$�oؖ�6��
�w���3�f#��%���&��)�g�͒�e�v���a8���XoW���X���ur��e4��^�E�-��>�s��h"������e�0�~v^�mI)�N��S#_�C@5�-�H2l�.�*eƨ�����ǫ�hȝ��+��ZG��I�!;֣3�He&Eh[J�V1a���ߖXkg��Ьlx�g��u$s�(Bo����M�YO9���ɉ�Y��
��8�=�g�����B]�J�~�l��F��sh�(�[��'�G�r��}�kK���e�s���)��,�o6��� Mu�\���s�E-�������U�W��f�����2����WC'	�e{��@kd�fYoe��1��m�u���W�i]W�r��6��~xUV_G���~z0�Q��.�Q6��r�͘h�!��K'�gS����K���Q��=�^^@�2���o8���#�+�M�+ۀ��f�eF�[���уD7d	d��~:��X�u�J�E)����M+ t��k֧�=]z�7����t�RT��7���7�V#�{���Q���S�9׋Cf�V�g�?��%�PP���� d��(gm�б�;ԅ'!IǤ.5,-�>�$G�"ݝZ���1�qagS����,8�l�Nn�ٕ�M�E|�=�2cNMk3e���P��>2���2
8+��RDɐ~��[�w�ܞ��e�4��(�Ã�,}�D��*"���������7_x��\1�IJ��V�b9����'Ǣa�ǁC�Mm�����n���UM�#9LĢ:gD4�3�x���2���Y\^���9���w��D.EQ�_Gj\�'̞�x}���ų-3Y��~�38�c�%��'r����h[�^����-}v�75����o7�.Vu���̋l�?�Ñ�[a��t�o�_�q�oH�f�Zg f���o�-�Ӆ�!����\D[��`������
F ˖Y�t�
ڴ��y,�����`����� N�t��R��c�k��K��}!n�_ͽ�I�p��f����
^�Q��&h4hN�a0l�L86�_␿��z������J��x�
x����X6%^k��ŹN�2���V5f#�I֘5����ޕ��O�U�Q���F��X_�k��G�ꗭ󭑏C��ء/�Lu�J�Ō}���H�� �%4��|�y���J����A8� 騚#Mn� 
��2�~3�}،.<��۶�׼���Zl�s��rvʫ7����߃ ����f	��̫!I�]�~M�-��Q�ޢK�e��[5N�\)o��w�4%R�rH:��&D��
&Հ<�:5e�T��;K�筂���E�N*��X����^�����-=^֟�l(�y|��I��VVJ�j⥚��#��s��'i�D����ԎN9b�U��;�Z�7��̧��pz���E��C�o�� J$ m�w"�M�0�x�k��	�	!�|���[D&Ϙl��f������	��x�k#���N�L��z��}Vgf�4�I�oԋ%��xPJ�ae�jw���1��UGl��+��9�;k�T��)�h�yN��&��-.xv���h mx� �f��l��Z�1Seq�̢�[
5�i���7�e�..����t?<��'�/gÑwO0���ZZx��,B�c��8�2�ڰ}	��S�S#<p�l<�@�k�k�b�����UXʒ��Y^w��w��S4����E[�wU�����{�ך��񯀍@(�~�N[�����oW]  M#�C�?C�O76e�e��H��B�2�m:n�gK���p���pw��ȧ&ٺ�nX�`��P��{�8s�Ov��+)<x v�vY2��37�~�6���&�����#����ʃ�rˀ8S��ڵ)	����bEiŞ�cW���W�8������[%�o��1�l��KX�T=qx|�b駆y�lQD���S���/���{���I�Ov<���-}�ݘ05O��]虏{)w��Y˳���!x���!No����[���*����ŭH)���:�ԁ|pdZ�2��7���{�85���Iu\�h�i�.�@c4/�!�41�&㐁��z(���[��G���gʦc��B�;Fh�rwU9~���&$����	@�;���@��Kވ�I�v
v(�+�}���]^����iZ��<���'��� m�@]:��b��Fц|"�I9%�W�Ｎ�1�"V��;��n[&��U�4�79��Y�ߺۊЀ��4ja�|Z�S�;���b�rK�������c)��f���d3�r'�N��M]zmɔ��%��(�H2��kj�S����4����P�3�ٶ*�|������x+coNE��l�ȓkW2��?���5��"��N����8y������Z�3�֠O͇ckˤ� �ןj<��u,1�B�a���osI�*}1@h���Ӂ��+�D�c�ed/���E�4�-ށJ�ƃ�tfГ۾�5��TM�[�u��ML*^�W Б���j���*�A��(�J��.\�{����e��P����vc�d�mn!XɭZ�{b)��Eݜ�	MӌOO�������-T$��j�[�[5޺�S�1��F;>������>�ɑ���c�E��f��	��Ķ��G�0�J�8^���*����R���4�(Z�M�]]
-I�\3�����*��H*�wn(z'8����A��Ke��U(2�S4=��L����3l�Ӭ�S���;l]��|`����NJ�}eϸr4}1LWq^|�qg?�!>}�RQElp ��<3�S��d
B0��'�f}S���K:����{���p�-�ȽK�o3�f�F�_V�B`������"�����@��P��џ�;�@U�3�י���;`��!�_l�u��'(6���I�VC�����k��/����p�r"2�TUb��eП���=K�R�os��M���ggM��g6e��ez*��W�z�C�0ͺ��pQ �ʅ�$ϻ�z�S)��g��%b�}+�5E���AO�N|M�rӂ)�
\��:9R�+@d�P���C �y-�W|��%�l�x�LI�����G��GxeG�l]4�5^y׊��5/�/9t2RZ�#�2��x횯č����b�2��}7�]̀�ݽcf�l[6n���D�F4�b���n\��id��!���b�?�4t��ٖ�s����b�G�[�����������L	@%v���*��H��U�3�A|)Xy7\�q�K����w+ ��a�^����2����{���*�^I8�
F	���ׂ�i��&S�2��ʂ]��T��1�"��DS��8��* ��f�V7�+�B�e�]"�O��p��G�jK�;���/�2�]��+g!.>�1�s�7c~����p&_N)	�D�"a�P����.��o�(n����s�ñ
�f�y�b����guj��|�JD�d|�2Kʗq��8;�f�5���L=�ヌ
��$Ne!��B����,�*�%�tK�LL�uk��)�������S���'�ܧ���&��;��-0�����B(vc�$��cu�\?���7���cZ��R�,��0�`�����7����+�.��4u�~�P@|ѠҴ=���C�JNyi�E�wGr�gS��'���v��O^�Y
����s����<H�� ,]^m�sk��Hw�R�ߖ�������]���`�����u��f�<A�Qla��i��+V�?���9��M'KA&�$�r-��)iAE��t���!��o��90_��y���N�^t`R'@��Bf����v`qeO@�k'wBG*Tf����y�	��\>}�
��=�����N0;�e�޴~�ʡ�p��$���sa%�)�:|&֯7I\F\aX��f�N��`�Uun�=bC.v(����a�WX�������}�5RD�����RL�kq6�+��2�&Lv�\��&g�Wn�(�� ]q6P;�U����s�M�C�7w��2_�F��{���`�̞֕A�b�$���'�Y@c��O�6rm]X���ߊðr;����SK�ed)|*#�5Z�떛Xâ�m��/t̲�aM~l�4h�8d|�v�J�H	�v���V�[�� �����2(�AA8�m���~��wW�p�9��Μ/_{Юi��A7��ν$ R���aFL�.@�x��C)o2���POz�ÄI��JX�i(F�`V�n��,Ny��6�-R.�E��n���}���������
�Lއ6��H�u�W�s�pɏ��+���M�@�h �H��8�0s��̍�Dv|Jr���{C�d?t ��a��@sܢw�܂�O�n��J��xYM���@�P�r��V��6R��0
��Zw)\[�̟t��z�#�Q͹V���;��-�EF�!�{���a��#g���ܔ��D8�¯UI
�Kj({�8L�|��4) ���z'{���ׂZ:*��ǧ���4t,	������[�eK"�1yYnm�xY�T�M��p3�u���	Lu��N᤬�f�mJ߸�)M�E`ߠ�g/
��d����dD�d�92|ⴠʕr�a�男TM%e��q����99�6�%�����젱�У~�w��ݜ4a�p���u��?u5��*��2O�`$���͏����Y"R:�L��*�����0rb��ڭ���'�x}d�ZC�. �����[4���A?ə��*�[���O4#�r�	�Щ�������Y�W՞Ԏ<�:9�5���6�t��Hi꺧��ۏ�V���rr�J"�� e��S{�<�Yى�#�����0J�]�K��hhl�1�𱑥��z3u�ۺ�v���P�x|���@#���S�,1;����I�>H�G��^t�s̧39O�k�f��@��Iߋ�再�xZ��!���u����o�ꥰ��Ќ�5�H��A<1��p]$���*}�"�J�n;��n��͙���sa���r �z�,6 �t��Ƿ':x��}Uꁗ)�� ���?۴:2]�&଎LF�����Ϯ{���_���l��߫������������=����i�t�K�P���cRgt�u���/^a��L�CJ-�ɘ�S@�����)����YH�̛ -��c�^����߈��=i��y��0����@��T�k(��;�چ��&��9����$����"���"a�zҺc}�z!q��_��Ent���Ӳ�a!!��W�c�|@N��?��o��:3j�5��9|~�30Xj�R�T&פ���\m*�ӡ؊A 6�7B��=3�d^��g��=�wK��o���v ÕLϭ�Ǽj�\Z1�g[����B�1�������>1�n���v���O�vg)��ih
�h���u9辮�Q%h݀3�V�M?t>�3������6a��L1~?Y�{��������E[���~ ��>��F�S���e�)-w`S�Bu2�
�_�?��M�������Zf�b���\���/��ˤ�Yڥ͂�	���dҟC�͟G�o���=�E��/D7�RM�.����~>��c�^��L�"�0b�k,CƙJb�n�"��c}�e���ё��R�ګk4+�/we`y;P'��k �V�* ~5�c�bFyNӅ|qW���&[���u6�(sGM���v�{�`�l�w�)
$��]�j�<�[�m�7��<�t~=\O���������^��,�d��_�sd�߭IۣA�w��v��a�k3y��������2�O<K��Bdr�2����)�/�yC���֕���}��h_!��X �i�IoP���8d`�l���~�az�q�:�P8�,9PO��ˀ�p����u������?�y�PD��3� qC�S�r�A��jad���~/}of��F��ms�{%+��}d�Qw�<�L �]�؟
������@�R�:�������p����$��E��G@_�啉�//%Y���v�� m�t���t�t0pU��CS�[��I#����UÖ���b� �J���3��Xx�B�K�Ż��v�1�R�2J!X��,N�~���Y�W�񣗕�vt�u�^�<L���IiΗ;���O��J1�� (v�����&M�9��q������,���[�:ŏ��	D�E��3@*��?��h��+�шK	áL2,k���!~b�g	 7��=�	�	q�oM��}H�F��^@�{�U�l�ҏ� �Jfc���|��j���	 �5c�2c�1@���%!���$P�R!ld|=	Ձ��b���h��HbC��Թ���-[Dvlf�n:ư��r�4^z�+dK�p�[.�b�)]/s�P�M�mǅ�y*I�p����k�5����Wi=�X�-����`K:����I�@~f@�꼉��z&-���3O0>|a�R��;���<�\��K���Ĩ6<u��)
�L�q�f�@��M��(��{N��D.�^@[>؏ܚ�`�x��_��?Cl�޸;���շ�'�f�2�-Ǎ24�q�ɇ� >��ʁh���?/۸����Co1�,�/K�{�����U��ןDRH���fe ���e9+:s}�0E��E����%�2~�ϩ�K��mG�c��6���5��aME�H����Jo$���.���.|��́5�_���Po�ꀤc��Ǻ'R���]塯���!�y�3x3�1�$H2GL}2��Z9h�[�g�b%�������K�=��V��h��.37-��@�ЮZ��<����Wf��F��~]�CЌJ1�|�標 �,TH�J㠊�)� ��y��%���E�2��*�����%�#V��-���8�j\ss�Afz7Rg�t�����"�cV�ݲ�IM��ܤB��!��O���1��f��	Yv�J9;�\{8p@tP+���Y�5�B����ϴ�?�/�ZT_��}V���"�J�W g8��t/�a�ؑJ9�d��8��B=e��;L��C���ql��S�/�IՇ�z����@!�>�g��X��<t=<����&��^$�����L>������*E8�w6&4�(;Bv*Tk��i�6�H���I��8BUU�Ő7�=]�sgs1��+Ǵ�q���&ϒ����[uE�M�n:�Y.��(��?�V#Z��W��� �r�h�/�R������Q���w���>k]��%Y�'��I�I��S]�� ���oc[�����K��%����/8sI�]z�B�M�q�&��/��^���e�{�Ln �}E�p)|�*������W�@>3�H���<L[��|� ����aL3?�ވ[}cZ�m�q�h����,�����U� �&0�Z��[FV�X*���o��N��v�I���Uw�� �D�:{8�Í��N�^s;V�m~�o@�E�[��5�b7�4r�4{��n�3�#�Ӵ���Gy���(u�ON��(Ff�cd��ߡ"[9+#1�$ �C�[���X|������_i"��K��fݧ��� �w�����I;�t\��5|��3�g�u����.�L�(t���� �β�`|+d<�^��}.��	0�دm�7O�@>wCښB�t;JL�5�-0r��9�L��a��/�$ Զ3;~�Y�bD�9R�Ȱ�u�7���%'�i�θ'� ��P���t��E�u���/���-Cv-�
�4DY��L����T�*�P��~�QE�6 \&*c�$��-��Hp�󦎍��Y���]E���-1WlWe����$O/�ңʩ�!�8>�*��G��B�|���&'����?� �J�7������X��,���HVq<w�o�����lڥ3�c'N�qa�mO���"�$��x�W����N[��I�P���A����(}�z�ѯ\n=�A9$J�GAF[�pL�1h۾�ݾ7�\jHpͱ���!��C��֓����k6'�TJ�M�ʪL����s6:j�<�[?�=P�Q@<��{�C���s,`g9Y�s�"x�����/Я�I{#]յ ?�B������i%��O�f;̊��u�@Ttu��B>"��M�!� 4-v�B�B�u�����_.� ��o��E@���yl+�Ca��gJ,������_�b�\�B��H�Ϡi�qE	[e���P��_�7Ӎ�4��N�ǐY���[�1;�|���n���`���*��Y�TI*��Gd�p]@,{zhpF��&����!'�����������1��_�*Y�{Z�����{@��>��o��)�VLmC:�� ��-��aq���g����K�� �oH����'�9!��r~ ���k�8��\PM>����ߺ��@�M��K��}������9���QިX�\�Ci}�/�L����h��ʭSѭM�ڥ2����mշ�#��bL�x�f�QBR>�c�%��:��sn��1A7��RJ�E��<��� c�wy���j��1���[͉j�_��9��xN�`�����@7v{_�1sD�ƭ���:��&��X��M�Mp_���C0���@������	���@��r�$z���4"2��L��y �8N%�G�Y¼h7\�8�Y�� ��s[)�Ȱ���諳{����FM�`n@u$��Dռ�6׵�jxڠ�;o�tn�3z?��â��|�,�-�bC��B��v�3rF��P��j]��i��}m�!F,U��8S��o� ��o)�x\5�|����2I�x����]7��q��Z�ɗ$�vgw)GQ�ؓ�nB����t(,�x�9� F;�����[����3��
m�y�v���J��ҟ�+$��n���:�pu��Ҝ���%�Ɋ�����CCDtd�N��"v�������x�c+)��yf��i�N�������������@tfM{oڵ��Ҫ�v`r�_�֍S�<�I�\N�w��6�%s��秏!/ա�6��Y��mt�<��bh��׉l|<�u���2�wM>�oзU�2�ӵ�F[6�t}�$X��t�2�'�叼��6�8���>`�K�2?Ǻ.����%a���ݓ�%�8V\L����R
z����PŪL�T�����}=F�v ��}\g"��v��3�oѧ��X�*:���kb�V�=���G�zm�z��z{kQ-��p�'��]��X#��<�a����r��/i+� ! �E,�,���0}f���q�jN��~��)^Ņܖ�\�+P����		yT?	��Kl�%TEi������Om��#���\��.~�P�R�Bb�gyy]���'���%q�=����O��,2���!�]d��"'K�L����P����?y*��}M�r_���R�+'�47RǐSl:�<3$@���,�<g����Z�ˍ}ʰ ��$	NzƜ1t�/��\�����,�r�#Fa]�6�z���|��rL>��v�ܲa��*�{��		��-.��"hpB޷�׏�\�&?��C:��!�m�EI�̓K��1	gT�T��ܜ:'�-��і�^��jw\�H#����S�=�u���.�l�[d�[P��`���J�/a֍����wʟ�&,?�,��l.��G�Gj��_�=�4Xb����6�gHwc�����Y�ya��2���[���<�b��,��� n�5N�Ag�] _e`�\�3S2
���Y��h�!ܲ�Z�Sc.�NL���|�����<�����Rt|�0�&N���4x5H��p�5� 
�H��v)n4	s�EP
�n��a%<�?��������nv��V)<����±�+����jj�]��ʋ�d:idN�u��� �c	����+85;TU����06�֍v�"h$J@K���BaGg��CKk"r��:���ySV��es`m�lP�2ҙ���[��L!V?�{x��[�'�N�c�m�/��dW��q�j`����L�[�vM/r��e�����<
��T���{���A��;�������/�`��[� ��%�;�~�pb��kn�`�S�jP�.����X�8�C��i���N���]\�aw�DOC����p�6\���/� �0��-zc:%H
����]mQ�y@8��nj��D�O	$�k���=��`��7��:��}��'��6zC �`��?�W }�t	>��-*a�+b}74L�P�:󦞖,+��.݊}NZ�A>���A���x��f����u�៪��������^~��^n��+�o����܊�1�>6f�`�� �Q�4߾Y
�%�$�໸�WG}�e��#�	"K��^�=�Tn�a�jĸU=W���R�p=Km��@"j�_8 �E!���p�QY�M��a��=q�:�y�-jy;�-_{����H�^z/�{l~?fi�����#o�V��+A�>M�,3u�K�-����[b�׃n?���t�#���d,䪥����uqUI�4��;��av&+��:�V\�x;��=�!7�DwuĻӐ����X����ⲬњƮ-Ήu<I�|?���]���LhJ�-��������h��Q�h@�@f����=`�M�r����E��ĉF�<O��k$<�]��$ܞ�Y�4\����)�w�Rˍ�J�wn�Y��U�e�Գ$R�}�_�~]#j|#V���WH׉E��#:f�i�΅��n���� ��I�ڤ�DvaΙon:��š��< �"����<f����YMd��72Y[l��)_��P�H�eu:�]��WݥX�RMp��Fً�mx��Lr�{�i��!��;x��|���ݖhi�\3�� G&�T��jPw2"�V���K��w��b����C,����_�^����Ӓ4-�,%�g3�#jO)�W'�.��� H�����x�tbN9�躅;��
H�Q�P������#�;If^:h)�FU��ac���L�vغ{�k/�7���[���AE�;N=�`�G�BOF�9�E~1�{��P�+���\er��nփ��D�;̑t�Ne�K�+#(�CI��KO���<	���u���E8~�ז���v��s�[�rQ��J�B�J*�l�,ۄ�[o��ER��sL�%=Ўx3ȌC��2�u����*�=�L�O3!_�6r	��n浊`�����Ta��W%+���@`)ܟZ�S(i�&�9g1�a�.�iX���B��D׽r��aԒ���oM��61�+X���+�<���MJ� Z�p���I�A.<)�]E��.ș3)N#�j?��ir��N<�p�ޏ]�t�t'���Yow�k.��-փX1Abh���$yJ���
8���)��\hztU����ܿ��RCgz�}
��`��܃!�MQ��-�U�m�{�eT����k��h
��ʪ��!f�Eu ZG�q�X�5��m~+"�>x@���n���({$��|S�(c�q�Ƅ�٘70H���e�fE�:��i�c������v<>����;j}���Y�i� H�I�����b�gs�`���Qv�z.������@R����C����w������ԁ�+k��3��N�`�Z��D��+��ϧ3�K���Uf�����i�M}[�L�������;��sUR޻y4C� �>��î���6��~E��X��{�{ޞ7��B�g�_P�Y*8��sw�H�b٤�afQ<	��8Dg4��r���!!�m����5�/� *0D/oX���,0b+/W�QF�MD���~�h��o�}��$�OF�u�"~�D�wҦ��b,WB5�b����3��f��C���U\"4nf�Bj�4܃_��;+����R�8yc���:�I��^{��4��t@�����aE	��sF>R�\�b�U�G(\Rǰ�e!�*�h�0Toe{�.�L=��w�m8
�Ty����A(UF=����zN�t�k�1�`n0T��b��T_94#��ۛၻ6�����+G�dAzc���d�'�7��;wW=jѭM l����X�k�+�Zї����n�w��*�㧪���R�!wW[#*PZ|��=�UF��n�;�0Z�~ 'Y�CLȭ��v#F|�Ժ��$f��2�4���W�1���+~�L�>�w��-�Wy���uK;�h�(��,j���ja��r��`����)lzo�*�1��A"��C�V�=����)�s��p�V;ПZ9����Ɠ��γF����c*��spE����N{�U�g�G�#d{��m�[*s�~�z��-�>Q�.���x�)��υS0y�FJ�}˭� '�?J�����d����&زV�z��C	����Q��� ,�����j��4�/���p]��k��%m�P�K\�i��������Cm�[	��mB�O�7���픶N�n�KA��#��g�UYJ��>��!�}�c07ʥ�l�G5�Z���F~2V �qV#��ά�9�`�U~����
5�U|�|k��Q2.ǆ�m�1o�"��W c�����Nl�[8! �ݖv�:0Q��
��n�
��"��Չl
,?���!���-H�r�.��\�6���Z�o�s�?\��$�3���i��U�@r0ލ1i���ڴ��$�o�)��#L���by~r3��,**l�u��9�NE�|6�c����v<B��-�P�/7سoF3z��Yx� �.*aQ>t�&����.g�K�.����k�"�vx~\�nP1���\�ƨ�`)�7�G��Y�S�$f_{�Lb)�4��z����O�og5��Q�%KT�@7cJC�T�����z3�q�$��b�J>��i2� )��MA�?��b�t�^I �'1D�m��۳�8�1|mS %��$環�y��,�O,��."v̮��tX}^�\��-}�c�:��G��o^�[�֘���o��zM?E�BM�Y�$�zf��oFf9A䄁�/��昧�kh�����h��%��t��[��e
�]:���IBo�s��ҿ����q_��,�G���wR1��J�䳩�����I�^ڰPr\�^V���b��D�K_�EMq&l%�8��{u3/f��� D�/*�);�4�E/JO?X��8����JZH<�P� ��1�(l~�[mIF(���U�{k���+��R}������C�<�߬4󒶌���TYE�VQ��7T���nݪ��"M��&���gt����H���
I��fuZygG��S�|�����.�+hE���������1c�e�9�d:+�A;��݂*��ͣ�3�^ɏ��~,B2��?�����ሹK7w�O�i���BZ��#�/l�<|�A��J��Ev����/�Y��'����Wń/�QV�l;մ�ƅ���
mtR�YL�)t�Y5��i�v���H�w��l0�W����L,"w��q\kd�t ��g:`ܣO�JY*��zz�~n��I�Ӧ��Bo!��g$M>�n���^�� ��I���3�_T
L)�'5�����-�}�ڽ+��Sݽ�I�ȁ��E�9�����)|����~ ���u�'��yUc����jn���<J��?�ݨ�x��c��X�hf�OQH��x���${�cv0tZ���������iև��EwF�+,҄Qr��r��H^}o��4 �U�:�cw�FŚ��	Pa[-F���,d�8��>w���Ѿ5���q�nE/�G�!L#0�s��n(�Gn��%�*L�VHی�'���Y��Rەr_)G5��[N�;C�+[4�#��76�h��y|�(U��)VOFٶ`�*730�pޏ�]	��1�.t�LQ]�P�8t�S��,ȉ�/��6�˩���~'�ө�9G�6q�),@�̬���B�䒣.W��R�%��@�'D==z��G��8u�2{DC^�)�)�<R�-vm�f��(��9��MU����H�.�������2g�7��G�[eWT����|�*��ݽ��=R&*�eٿ�ucc�YՅz�2j�Ek�lm��Q9O����@��Bi%��u���ӟ��^ߢ�X���&�b���9��������0�7�ϓ�/~�_�6[�)�.
�X��w�[Kj��'�~Kb����Tn���l&w�9/�Y3��iQ����2���òٸr�$~��U:�n�_�о�Xw(�l}���!:��ȧ�*�����V6��)��'*��gr_&#gĶn���E��2i�/��q��'ԯ�����Py�cp�?�`�~k��9�P��Ť�>[��#����T��ы�d�ӡ9T��»"����%������D�W�
/�3���y*������0���n[�E�_�v�b����&����UL�J�^G������E�V�Db���}�)��~����hK�^זO�)݄w��EcNA�2tiԣ������,��
��J!��z���g~^f���)�k��65�����7�xnٔ ><����M*�;��H�l�6A����їF����[�<t�K���O�E�*o��	cR��ySy�w�
>�,�Q!Ln@8v뤧3C$
�}V���~Ri'�
`P}����B/�y�>z6^Ua��ۄ��s��I�K~vM\ zU�'���f�CH�B����-N�J���9ϋ�C�� ��2ڥ��%D�]ȼS��.�Ɯ����.>� ���
	�,��歜<(�E�(|/��O�x��d�5Q��@g�ݎ�`�[,`<R���#"ioۖ֔�(�%c����iݦZpUl��_�*E4 �ߟ۔�.���+m���x5��|���|���Y�kU7���.d�3h3����"ɨ�)�Xe���3�z�?ZF4f�\�%E\1����_��I���La[��<z���m���M�]D/�<����p$1��H&��g���P���L���J]��> k)VL~�б��#��$@˵�;�V�B^V��oHy����B`��_n�K�0���5���tx2+Uc�\H3�����%�=�R2�6����mR��U3p�ݚ:yy�2~%�L��� �$w�`�Z	y��$�BD�(��?~xU���| ���ws��R(w�4�F��ub�8���uvQ��KϚ_˻�gV�4�Ӌ��1�,�D9��a�a���S�U�i�Q~2�`����E�oqټ��U����]l1I,/7���}e_k��/�PX8�۩���V�#,V,���=++�6�|)�S�v}�u*��G�Et3q�����]�� ��O?'}uDr�e$ڧ�N�>�?w �c(J�V?g ,c���Ƨ;&G�x�e2q�
E�%���l%�����,�N�A��uT�"|��Q5{xQ�������­���M��`\GǑrH��z�^zI��u/����3J�q���a�W#�0�pY0l��� n�	*�&������Ө�W06�������(s<�|)���̀���&gnlSF{6E��.�6'�Ɖ�<�;�Őc�4�է6<0jL��*a�MzN��֠L�4�0�S/Pĺ���E�k�7|1:O�@t�3y5�f�a�VL^	`Ň o���٨�gp��4 ���^LRݚowL�<����\�$C�$��Ô����A�Y�VGŌb������3���{��fj竤_	��Uء�1O�W��b\+v�%��I���̒�����]<����{�)���y�d6.��F�q��1��$�T{�(�U���JQ�Z��v�l0aYJ_E�qG +��uL�@{.��cUk�kL��Y�S&\ a%i�ՊU	T�T��n���n��_�3z���
$NB��n4ن^�� ��~Rf��}����'_��+��r�~6��5��t�ٔ���'�����j���:�A O7`X��\7A��҈�+,����Z�����ǐ��'���`�qL��m��+Bㄛ'��[l���s{�B6�����XJ����6u&__tS\��0�U�g]C2\.T�3���٣�V:Ԥ׵��xX��zA�-�͠���Y�i�v�k$V�(|�)�N�B���x
��,���ބ��`��	}�.��7�D�\�mR�F嘺��7�̚�TGk�X��d⯹L9�.0égt�0������Np�I\�Cp馎[I�R阖3�p�g�"�b�g`�����Of�i�_�͇D&V��&��DuaS͍�U�8�4����"�����x�w­�����?�"Bÿ)n�n����ڝ����z�	�7�'~;���7�g�.��y0�jI���Y">�u�������KPu�'��\LaO@�g���� ��6b^TEψ����A�Zٗ�Hr�dG틬o>��<_�k�Sl�f�~�`>���ŹST�36��׆ ��R��'3BP=x���yM�ߟy[b���X����-FK@������Ǽ)AbR��gJ׍v���`>~9�	�)�<�A ��h��{�aޘ��*�Щe�� �^�I
�(E�A��uٽ�o?�H]�7V��*ܯ����c�r�XٟГ�dZ����i��p-�3Ez2<�`��Q��Q�� R�a�p_��$G���m����2g�6���n IM����X܂����f�����o^�"��z�/[E1���_��G�y�*�0�M��W��ޏ�*_M��J翫p!`7�T.u��|!Rwx�c�:Y;N��a\Xb
�Ƨ��i������9�R^�)n�ZW��A���M��ؖ��bU�+lT�hv�2�ǌ$��/��Og�fnZê��+l��g��ĉ"G-�faz��yƽ��7v0���"k,�JY�����o��>3d2>�#�����]Ϙe���mO�9��qS���.,(�K��
)�;|�:��~��^v腠vճ��ڱLĤ�L�ɢxqJW%��d14�4��]p���8�F��j�d�h}�5���OxY�rۙڏ��� a��"��I���]�1g�o\R<9�X�X�aySK�(��0g4t�Jܨ�9����5�����T(y�Bg�E��*���������v�D;��#5�5{SH�� Ҟ�
���M>)���)���6�٪����.�KW�Lj%A���2H+*�E
2�����\N��z�'�'�4M�}*�;��B*z}m���b���ucM��J@��w���	�!�G�#�`�P�W�1��8�l:ĩe�=���w��I�I�ɑ&��L���w�F�W��2����sl2~��N>O�q���L���Ƕ�,�ҵ��󑶷��J|H�_59�g��,���+���7�S��C�aS1r�r���������5�I�N�L��
Q�7����p���6�Xm�3���X.�S���aEZ8����#lWY�����ICX�p�{����=���Wy_���՗b��(Z$���	��h���p�b��0ʤ�(��-����V�?[Q/M�WZ����^����	.���\�s�)	n!̄LF7�v�<�*u��ML�d����<Θ����<�^��&I���@�I(���|�fS~����ʓ�VI�*<���*�rH\T��=#�9ݲ26댔��6�N/<���M�Z���xpE1��6��)�����j)j��$��B�N�.�Ul��E�I1�B�c����]�߂n�|��,*�z0_İX��0�ӷzM3�}x5�n�!�FV�2��
���y#[���BQ��{�HԺB�eg�ʷ�HˆJ�����}�,l,�R'���Y"��0FXի`PYh�D��O���o���
�B����Uo�0V.�4�0<���Q
Ȩ.�B�IU�<>4��-�7VQW+�C�Ca&�S�Q�fxc|�אC�"��1D%
{�O2�ђ�(A"�<�|��ئ5.�#�+ �"�ژk]?'
�C��x��:Zji�4�<�E��ޥ�˂&l}�}F���"r����Q���ݠ2̙}��ȃ�JTxo��Y�6&Wx�:1w(=�	�S��4y(��@�H�j��.W���б-%��*��a����z}ܸ���ʴb:v�րuvD��M��P�[e��Ls~��h���C@&�enq#>�Zd���A���>�~䊍Hޤ��+�#90�o�2d�>��>WAk�4Yӝ��?�cr ���S�7�6�|
�)�h�(ѿ�+�(���p���5q+�x�b��6bnA�wϰ 0]3�7a/�q]j�g�S����Xn��+���"�o,��&�z��aK4��{�s�{ ��`�Vj�Yˊ�?<Qp`��1��Rb N���@As7�'U�ʢw�1��?�K&�[L#���y5��4L)ݳ�5!(��Lb�Ѯ;��%����K^�)�Ĕ�I��d}=�t���D6<,;t�i�,fL5}��k��&4�aկ�5�f^�w?ͯ,0�}q<U�)�_kJGwT����_�(����K�@���%X;���V#xC11�:L�\]�<��W��y�="k/�1ּ�X�$E�#%�`�M"���5_N�N��p$��5�ɟ��. � �x$�}�X&B:�°���RQ��H�~Ց���E�W�NR鲡y)�j��ЧF�F� ��D��=3fmm��<��ܥ[X7�m�-¢����˞�a�F�"x�>�1�4��jI���_&cO���j����il��M'}�4�� Y�8u�+�����z�|���16��%�,B\�����hY�]���.��l8��W��!1I�N Z�R���΃�ֱ����d��3�@[d��TGa�1i@�mWma7.�i;�8:s�&ݍ虋S��#�X/:�����uq�,o��ޭ�9�@�ģ�	V �ҡr��%k��}&ۺ1^���d�3efL@�م"���h���)��\���Үjo���,$�,�� �ǒA'4E�	����:H��c��x5�?7�YB�S=��ڦ+�	����1�6�O����O��$�T�!����#�����8P��'����nD.dM�Wގ|��<=|�M�G���khu��.�.��!;K�rM�~�X�W0cpI�T6}�¶�ya��q�G�|:8�rS7������8T٧f���AM4z��,�7_�a3����\��Ʒ�(sxl��^�f��VW�z���xW�oN�Q����c��\%�e�EVڨ9N��p7˱�{��Ș0���������hT�>�	u&Ĭ�_�y��1C�m�6��οr�U�ă��S���էU�B��n8H�E;o�����x
�O���ǧط.!��$H�"�?�^Oε���M'<���24/��*�,bi{�,in%t���2;�۞�0H�.Qd�d}���
� �ҚXU�L�;>nҎ����8 �?x\�q��A�֬Z�!���x��͑�H<��8�#�A�C�[E��� ���3���Vn ��3���0T�@]��b���qK�y����%�n� *[�Ή��$���<\ �����(Dt�s��݃�!@�DsqE��~k���fG��V{j��H]�l_FO�8���#��Ͼ�0o�}6��}�u5#B��Ƭ�寋��.�=�N�ԬȾ���t��i����ř�?�^��<1�����/T�mB{~��;��U	�Ϙ.�C�	�)E�g���^��@W2��0#�ڝ��h� ��I~���� ���EGBU=��Wk�.��W��~%�x�o~\f�*Eh9��K!(�6g�V	I�!cb,�O�ʴ�M��'�~��Y��T�m 2
�9Y��RX��{����3��-]����w�im`�9�*�V;�2����L&�s3�L��&)��*T*�w����Ps�/ӧ4i����fO�`�fm�ùh�SD��Y�Ǧ/�nm����N�4*^Z��݋|����Bۃ������V�j�!_u|��A
ӐR�w�'?WygJ�]����n��ធ��+9jpV9�M)���4���L�)Q�A � ($�o#;s��P+s�z>H�� �-�Bz�;@�0 ~�����h14�N�DK�ds=��<�������M�#��m�Z�l�T96r��<~1;z�S�����p��]�٠d�J���^�44�0(���b�bU��?i�n_=���^)����̓z��Y��M�财S���}�U�U\�-�ՅO�%�A`�meEmtDM~J\�S,^��vջ��I1��ì����I(�Z}�K�Lԍ�]*�\I�V����Lܙ��"5�4��O�� �� �=�*��ȹ\�����(x]}�������Ӗ�Mn�:��wȪ,�h�3oIw���`9C[	LB�/�D'I������˚oGF�֍i�/���g��U��⃈�[��u/g�l��`W6�AH� �K���c�w�K��+X���O��]�0�e��j�0������9&��#w�@&���Nk�QF��9�J����*���,����Մ������*�[Ig��ܖ�MRLR����<mă�����;_��-r��%�B �o���|�3�W`@��h���y�d����J|L�.�-��,�����)3A����R	�W����.)�at���;���O���vC���������9%��F��MK�0{�z!�P���t��P��oIqi��.����L����t˕��!�t鬚���6��RP�rI�`�+�(�·é��p�fɁ+~��gTNx�{dst���]���Ýq�=�w�����[�.h�9��k$�v��|�������`�����T+��_W?-���B�8�?	�w��!N
6 ˔Q�U<S�R\�~��=���(�b��������Z��u�!<�8��bEr�n��:Jb:{+C�n7�ꀷ�D�&9`M���<���nln0Kϱv'��:�
�;�4Bzd:�)	.�σ��u@�����~��i�9-������G��@Ï�I5T�N,X�5�hS�� �B�9�c5�}�"%ͬ��W֙\�$�� ��KA�{[���-�'�+0��\P/�����':z?)�?�-��G�sݸ(��$�����ssmwĥMϗOy^=�m}�4�o��O.ު֍?��J.�K�̸R ^����=	6��[�8�,a�.�XT��:� ����rd0��&��e�KY�s	rE$�M�Eμ�V1)����n�t{
�<�!N�D �i1&����<�tWvyK�Y����Q�_��Q`9ب�p۲6�7
��+0t�>D�߅s ¶z˾��n�%�r��X2{!*;H�$�>i���q�H0*��F'�T۲{�t��;p"�Q*�(�~%æ�J�?�Wy��}4ֿ��ʓ���j^'⚋��<�֎�'�ܰzI=�o�n44u=$Y�����f�Y�-�7��9�؜p�!}�K�Sd�h�f������t������U�W�٬܂Q�)8��z0Y���nK�|���U��)���W�S����;��TR�B�q�G="1oY��oea.
8n8�A�|�c~C�t��T���on�]��*]���f�e���E*[�T7���Uߚ���nMƋƓI�Q���9��z���Iu��6�8�p�[f[��>t��J�����>�`ܣl��ޯ���I����_���P,��fhu1��Ԛ�m��>�ETC_�i)�HfZ�\ŎPxJ9�� d�.k�:�(�'���
us��hA����d�s�^d���8A�b�<����n��يI|U�"�sŠ�k��l'ٞD+���5_-e�/�.7�&FT�Ü��P��q%���SP�lFM�"2
�1J!m�Y��.0�����)�]`�����~D\��B��,���(k�Q�����i/����mԒ�~"�q�ܿ\�2t͙��M�؛��G��UMb&���En�7,<cծ�8V��j'���� )g��׍*A2Ib �������L�-/��탙]Sl��Ph]���<�1C�@!���N���}zmCͧ��dXQ�w�5^�l?��@�/s��GB�QZ��5��SЍP2�����E4����4�Dz˅��ϵ*�y'���{X��$��`��4m�v�+�GSr,	tL)�Dv�f�c������WR�w�Ɵ�i�������on��֏�9� �� `�p�)���q&�=�y�l�����j�4��÷PZY��:B����M��_�e���������@� "�JG��ⵚ�cL�����nL�H$/��6	�g=	�ۓ�RF��Sr�V�����H��Xޟ5<���]�FI�~������R�E������0�{+��yu�+�s��p��]X�j����Z}�Z�	���U̓��t/w�F{7˰�6(�z&|����M�)�t^,��A�e���q_�R��^-��lU4P��\A��U�Z2��g��FY�99k��Ϸ�+$��A�Q��׮hF�m�.�q�g��U��ҭP݄��ڵ��xity�v)I�xҬ�Ddx��~�9y���en~}�ٰSIzzח�B�C�*fϥ�(����k�nC.9�]e����^��=)]Zx��_^�G�z�����vL[.�ipSa��J��HU6��� �cv�s�0n����������Uc)��1Ǹ.TC�R�MP��O��3R�QR�J�5��;+=��Lv��;19�.�+���2� �>c�b\ ��~�!���eG�6X��!m����a=j�ǉL��rJ2�4N%�k\�sTU���gnS��>Sw==�M�q�_�?��P�C.�Z#�ܚ�pKGA����q/&F�f����G/��1	�Kj�se����0�'���p�ǄP�7f�[X��D��6�'t='�Ȥ�7��f�"u׷ ,~T_FwCi�6��	 H��S��m�}���ʂ?���t0�͛�#���|�w
��#�t������z�FrY1�m=o�89�qƽ��׼�g�R��=�/?,�2�zrw�B�}��Q"��	ck$��xoF�(�k��_�ڗg�oe��=����ܧQ!	��F�o'Y���f�I��z��ʆ���eP�YZ���Dr�?,�Kc�j�=fۏ���<�&�������
 �R��̡���1����}��Zl�9&n�䏠uO+�|=0A�$[�3^[Ϭ}��Q�����Ԏ����f�+Z0"� W I�yE�TR����B�h��*��ҳ�V��dD�6e	�ns)IPE�����U}H��I�L�}���D�'a�:��ǨY�<=�����	��_�A������Y�'<�r6���l�$��Ǌ�1;�����54�t�h���x��9�d(g�Uak�&���k(-\����蔗��~�+���x�e��ǣ9��������d�|�W���=���.k2��	�V,�H�$f oZ~�ml�����/�.qj�U����G6�����1sR
uRx���|���Zpꤡ���ӦZ9�e�z΀�E%�/l��r@�P!��TFΤF���P�&Ж>ڔ��%�]����97��6�+���w4�I�$���STV�Pc�)`7n�3��ث��v"��]�}�@�_��0O�9(�IF��6]}�pwr�_p��1���~#_�clFeɾ��ك?�k(r�sڄ"o`}�d7H��Np�F��Ÿ�����imYʣ�`}�$]n�%@3�_����D��q��\��m�*"�^���jL*nӿ��ϊ�:�Z�3g����]��v׾�;[�!���w��Ӻ����\m�:o�l�6����B_��h�' ��[�;ކDz��x�����>��sb䞺��������<]"4�ٛf��=�H�lƬ	�m�-���������j�'��d&/__��ՙw��r��>�Ȧ�#_!�O*�n�+�)�o��l�8�1�M��8҄x��΢�.����-�T�֎��Q���,#H8z��c�4�#�_�6~r+��ٹQ��;�ܢd�3e����v�?A��2m-������� V��,%����̧��5��'��5:����%����vU$�uCW��}�	��j�7�A��03��~Yh}��8?Ϡ@զ�Хަ��&���(Ҙ�e�I��v�ƫ�H�p��q�H��O��2�W�@<��i�����ո��\k��?݇�m<\��^g�ґ� �lB��c���!Lv��h���wh����K��9��4�z!�D�#)�'����È�@����P~4�l�ȷ�[@��о'����׭w���t}�ޏ���=����l��$8�+,"D�b��m�N��ݨR�|+�Y[j���h_�Sc�f/ ���=U���̃�R��x���h��#z��q��4�*_��H��˪W�2g����BX���LC����)���Ր��d,G�n���X6��j�B~�:����㍱	�n��[����f�!=J	����ϗ�of8�2��j���I��ٲ[���*K����������\���!9+��U�b���м�#�-�1�k�	�C�lB��j6�oTN{>���l�F9e�۬l�3���	#�É��s7#��KHp��:�AE�s�]j��~�<M��{��e�� �� J-ln1D#F����g/F�Ic��Ɵ��L�&Z�o<-WjH��M֭Z��^��B�$�̧R���,�D~jȜ(٤��*�~�C1|hR���5�����pZ���z�T[>�TP�`^��MO���梞�������+���)F����J��5�O�9@ͩ.��ڟF�P~���VP5U�p��&�R�o�b��Z�M��#��1��D!J4��A���5��;<�������<�eJRu�q'����:I�[D ��}��B����UȲ�]8�akz(��B �]�[)��w��CsE�3�D���>��E��"��Y�G���2�T=�L�ጊ0i�D�I
m�̎������ғ#d���M[��.T3�z�Y��!CPL8Z�Bݭ����.�h�Vz'f�^6��x��t�nq��T����� �&�B�J��5L�V�ln�W�Z*G�4i�~zݡ?j)�]��^/�����{!��FT�x��A�"_Pᰟ���ƆDi<��^����D�>��V�z�5���=q����i��ѶX���������CҮ�G/��TV�>�k=�&�?�8�<��.�A��7"G��|��e�W�H��Ca��8���m��!����SD}���۵�~�.R�z;p���Qָ6<��Z$̙GyR�2�g�6����I��5P��m�6����f �h�n^���~�(7�K��Nm�Eߖ�
�_��^����N�����z�w�b�6X;�]�)�^�>Ԏ�(���;�/��P�8*/�
ڊ͏�<��@��v�ͫ���D��Lqc�숄�j�����+Gϛ�۽������� 6�l�$$rrt]"H�R�������qʳy��Cj��_f�1Bty�<ȵ��na��� �$��V������Fa�뀏ᓙ��%�7q��ә�ޥ��@�ۜ�U�0�̆�\�/U�]��
s	�K����'�Hs��9Z������b��4�9$���X< ���rG��Tq��)`�w�.7��m0NA���[\�}kW��2�c�%
G��ŋ�*��t*���y	��
ڵ=�۲O{���-�؀��NG����v���8�O� �i8Iko��*u�G���E:�T��B�9�]�:<d�w;y`(�T�Ԟ\�3��!w3�ƺ�&�|	Rը�E�( ��t�����V����}	�hԂ=�P���8�\������06����	o�L�� [�0>S+\o��!O瓬�.׬��?�=�@�:�	[�"�˦v͹�krru�o�:g�aYrC�}�V��2��!�n��{MD𡎑�8��n�F?-+��ɿ��ɪ���,%�����v="R'fbV��t��i�����O�s�"���o;�n�w7����������P��.>-�]�x�Ŧs��R���ֹ�w��k����yyvI��m�1��慿ܑ7g��t�q]�`C�o�z�}OX�o��ȥrS1Y/f��>��>�!NVFeN��%��Ql6Y��I5@�!
��K��������i�l6��(DCE
\k���p��Cݫ)�NZ4�����$jq��Zx��6S���7�d���~}D��jO�ѣUP�2|9]Tj��w�Ԁ�A�Q�.[��[��`��=P��k��:����j� �9)��O�D�ʏ�
���7�ڷ�[�Ξ,{Ւ�s�3����������@��w�qpd���I˚����H�r)��_�h�z��8hK��C�7XY��"�+�zw�f^It�ʇN��@i�Q�R�����s�x�ecu�|�Yp\�ͬ	�"���$��^��ѿ��s���g��4|�ܝ������B�T��|KC�y
����58y���j�̠�8b�b����n�<Duш���d��`�R�Df�6R��d��V�o�X�5v¿ֽ��&�3�90�H�@z�;6��2�kW�)��Kr&�7��
��y�e�R3MY���WG�zj@�Y�˓���u�'��_8|�"�ڟ�[�.B���i��E�#yZ)(^F$�4H�<�5@�@V��=�~�2�+5a{�(��~#�x)m�yk�!m@Gg1��X2L���{^�����`7�P��bŸ�k�������[�;H�����@��.�x�
�ڈ��VOr=mk,�ݎ��(o@obN~��)B:���ó�W?ә���`�n��O���?��_�LAdQ˄�h>�w]$��C/��&�J0��H���ux�Q�
ň*�h��V��\n��V� F<vf!��3.[\/�o�bg@�3�Y%�.��I�r ���[ޯ��C���ZKw�Ҟ��k�]���T�Ո=��31CVܨ����x�Z�P��<�0��6b���V� h"?�v��,E�в�ٓzJ�3}�A������L�'�#dP��:6Y�	�F{Jep�V����4�9c�H���E�>�x�*��3����w�޻A	�9��:�j��,�Q����K�QM۱����'�	�����(na�1�B(�n�`�i�q)���Gk��7@{�n2V�k���J-���p�]]� �.�i�$Qϕ��\KIF����!�i�pRt=}��Ǳe8A���.W
�۠�}4Ӎ˴��;9kd�e��n�!�<���V���@��D��)�p,�d�t�������t�̘�X����f�e�!��h(jB��E�W%��0欕�G���:vm<5;\H�@f+eHp�����p����xQ�G�i�jo�B�ݢ��S͏!�Fۨa�[�:�WD��~j�i[�Q�m�OߨH��%��WY��S��6I'��>�b� ��O��� �H�[��Gm7���z�)&���
�C�;�/on+Yr�I�2�-�^ 9����	2*�k���_� ����!np� ��?��j~N*#��ܡ	����6E��W�^�f�r?�tO�	��e�kc�'�X�|GtC2�Izz�q�8��Y	���N��7T�����&	�=X��QO�k��>���fzl�Ea�E�ÁC��:YKp�{�=����w��?I�_��s�1��
Tw�l'��$��՟+�̀�+3r17.eQ��p{�߄_�k�4��Mh�ҫ �k+}yoϞN�,jD<!�h��f�S��ۆ��iBL,o���������⟲�������K�4�I�<�2�A+a�O'L!h��D�hm7El�v�����4kO.�� �e�Y5�'��4nw��^xl��$���|�xҵL2s|aQ쭨@�kO�2�L����P2kf����B��r�D�y���������j����U��R6�G}6D�;^���fx��Kj
���@pDXQ%U��ڎr��[���'�=fn[(���Ob�W�MQ�3��s�5��ؠ��0���l�P�BvWR`$m%CSm;��;Ѝ���bو	ǩ%F��8�}�W�]�Z�S�������x�O���6����6�����vY̈�25��Nx�j��ϻ�"N��O�������K`�������qx� m��E ��@˃�{3�)6�d�G��y����0(L?�%}d���V���Gv@f�᫆�r���=''��	G�����$B��'1��	Ñ��o�+���D\��M1��2���\�h�p;z*�?����c��>���`�L�tDS=7*�Q!�S&�F|j��舭����9�)�!����?�*�]��ob)s��8�͵_���yvD�8|L%�q��@W��߷�y�C��{-񝑺U�v�6H��n���?���%���@'�W�D�g���8`��k�.�B�B�u���O"�P��Ѫ��K���F��{�Jj�NpL-e�v�3V�@$*��qA�_7�! �2ӡ!��{e�j'��Z� x5ӘӞ�0����}r�~�<B&A�6Խ.H�C8޲���  � �)�n撮�v����0��]����!ug&'�(���"P5���[AS�,��{V�g|�`�x�����R���@����	p �n!�Pb�m'�ʎ/ٓ؍�Ө�Z�����t�����Z@2�b�GpZ�B^��|3�}G����I�"���7��Mf��Ap�֔��0�ҍZ��G�cA�:����M�Dd�im$�Zt}F3�S���&beD	��b�D82 NL?��ˊ�(}�쐙���x�k�N������*>=/ؖ��n�;�>�F�1�-C�$2�r�\��qpwRiEկMl����
�]+x��7�	7'��˨�IWY��}�}���f2t�w���Ƿ��Z��T��|,:$StZ�q�|���.>w����uF�
�>s���-?�˪�(�$X�]xD+�}G;8X85?r�~݃�|]C����?�_;�	�1��F�ۙi��p �Zl]�E�=����V��Z��]rО��� X�����%�+��u;���MO��A�~J2մ|�b扬�!'����#�"-�H� 	.�A�v�4�V�!�'1q`L!e,	 9�����iWj��uاv�}�@���/�O��9E69���=ܲ_��$]�R��x�h���XϚ���l�nO�^QZFr���IY�K���2��P�:�!����	x|_KǆH��}�ɐ�)���O (�����pq�*�PgR��f�^Q�{�%
�x���G�~�5��O89���ʆ�,���s��^�&e����
�Y��V�Jg­�,��,�̊p�R�Zp�Vp������H�E��ͯi� rL��c�#��3w���|�'~|�Em�X�«}1��(kE�����^~'(/�bX/L[�� ��#E���ǘ+��s��x�/�|�b}>1�������z�?�Ɓ��4��lwT�Ɏ� ��=�{jr��"oq
]���87�&a$�2]��'��d���e�yyM��H��E�Q�cVj*/���b�i���R�J^jҝ�a�zQV��r9E�=��;�4�3��}�T�loхd��˝������I���[ҡC}SjI�'K��u
=S4N�W����8#�Oj9�+w=O�5�؎��Բ\0��ZIS�i��#䮵�gVy�C]F ����v	����K�5n��ܠ������V�y���qt�ܞ-��������˧&w��~@]�M�S�K�+�����.<����:�|F',N�߁[���^:�-}�J�:�B�=�^�S��P�E�� ��\oO�j���������Y��'�܌?��d���r�,Kx����Y��j5w��r�؋$���O�#@�L���W�zx���g�*��,'T8�ÿ��8v{P���/�/Nη�L$���4qgc�
a둜���j�Y&W�6q��Mі�����%C�w��������e�Q\(�?J�<K��C��r�`Ԙ�-��^W��T#���E�su�|'��<��`Qw/����Ù~w��9��־S	Z����Hl&��0�[�������\��s�@B�\A!R�a�j!�׋M\��ѫ's6_�i�.�&FhAQ������
T]X�&��@#�ym�!��I��j��*1{m�O�%b�̝w;vp!@���4�"�|��C�%uH�����1�p�T'[Adf0��=��3`rO��q�%����}S6��Ύ��)Ӗ�V�~��{)��F8�bi�0<�Lw�9�`g3ӣ�4�p�xZ�gr�"e��?�{Z���%���;��XX^h!#8�w��e�X`s��3�o���x �<���Ɗ����x���z=U3D6�1��<`�q�1�w�J�i������ob��Sx�z�f>$貨���Η�Ͳ��Md�l�vm��:m������(p����E�d�u �����X�(�J�2� ���� �V"�r���t3�C����E7���$�v�i�ݵ������a�a(��Ό��3�A�/��
[��U�E�:�ͺ=ѵ���+MՀ�芲\�C+���T��I��8��������6}��q{:)�n�ʞ<[�t�!���ŠIVAKm��e�,�9j"��7PK:1�\���{a�y��.g����) �o�`.d����}��G;�~�}-n��<5|�ԃ�s���̿����Q{�~@�ř�%���� d��,�C$" Qi��L���-��x1;���\Q�q�_{���L	������%��tC����vI�%F�b2 G���`�`ل�	~�=�������Rtx�|�4˪�`G���Ǔ�ƞ�U�rMYM!�8"�o�����X��<y�3� ZuP�\���%����Q	R]�������Ʋ�N'��^D�\�!���,y����� l;��\���/6l��xH�y�3\�5���6�M*�kiޮ�b_�_�b!�_@��Qo&���	�${[B,��E�E�!^W]e㢮���!����(�H��EA���=x�`���lu nF��D�����Il��
]q��G-6�㒤d����`��>��Lu �~�L�l�p�=<������@���V����7�|�y�Y4���GF�S^ɝ^�����j;7���ć�sk�B��	�@j�j��Fo_��Zj1g�����ӀX����{㊎u�R�U�,���6��%����}�ٔ#�B��J��2�e�"��5���j�-b�<��)8�+�{��J:�/�����jڇ�f9T��ǎŜ�J�>�o����z=�=�b���I�p�s�`�Oo�I��tPޢ��VV#W�]���G�+�` �7�I�b:]d:��wY�����x�^��g��רYK��w�< { ��{�β�\ɉt���G�ЈL���[���� ����r��f$�7谝d�|�]�j͗Ks�"Ħ�ʛ-���U\�����[A�A��pչgz��|���)��Z.�*G	��2»v,�-}?�v-͍��^\�!��'x�����_2��Ƙ�.�m��^Ӄ	b��b�T<n�g�VN���< �l��g��g$��Y��>����1�K�ׅ��Lˊm�}�,���	�`��?�m`>".U��e0�ՒL_�U�R��~o��� 59k+���k�
��Wε2��^dD�v�-���*.�돰����JY�����͛^�T}�=-{��ƙ��X7G�t5x���Q�Wc���R
;�z�#��h~b ?�=�a���7� ~�2��35�7 ��5��J���.��'�D\�#{��b`��;��{k���I~C���l���GгOQ��Ч�&ɠ	ۼ<9�`�(����jC�Dc�}eW��s[� f٬�e'�0^d����*�wi�<^t�>|&���pY7��/��u��^���������t@nv���N�L��q����98cx ���=R+=q�'�:�ban݆8O�k��8n�$��d���F���-q���n�Td*t��yZz��)�C�ڰ#�h	~��&���G3�[�Б�L��v���)Ϊ�S��y��{ߋ�ZlJ^�3�<(�ӹ�q�f�`ȣ��T%Ɔ��K�U�S,)1�P�����%ER�8�6$<)���;u:���i���]�:�C"�� ��m7�O^�����'K��>��#���~���;}�#���v+��}�[f��|G��q	Kǀx�X((�o����G�EeF�\�x���l�k���1��m+W%�2}�q��l��wI{�1����m�0׸��.��^��b.��,���r�Hb�b�ͼH��?��ao��xFKp��(��=n�6rӞ����#)i�/!r���<���0$��z��0{��&L��ϔw]f��rO�$^S�d)!�
Y��f�S�Cg�|����%�]�A����m�>C�� q�3;�W�gJ�x��C3�G�x���Y���-d�Y�/C��+RX���7zc�*�v�Q����)8z�s}"��H;�//�/��/���5H�	 �����c*�6���P��*��Oa�21��nm/q\B)9�`��7P~�0F� Ћ{�vi�c��w�����\c����� F6d� ��E�3L����r�_���"�G�)�ԝ�v��l��L��]�چ�`0��,�T��'��W+��3>�^1U[��&]h-���@p^�خ�9�tշ�]��B�Z��?�_���C8U6R��E�̽@*�Q) Ѳ*����ʠ����GU���ڠ)chU�c���0^P����~����A_Xدq�ܣ���_	������&^��������Y�p=3Erg�붋.p���u�¾ ]��JbIt����(*��,| ��`y��j�ܶ�z	���v��_�z�ޙ��5Mg;���J~�^�c����<�n��y� ������zaä)�e0�^Yݽ�m�ka��8@H��D��i'	�7�Ƅ٨�SW�[,ퟍ-&o`4��1ڂ�Y֙FѺ�ƕ(�c��3���� ���SX�T{�W����fI���|����x/}KH�DZ����5���.���a�8�a�2K$�(��F�;�"4���:{�.u���&�AO:��Ӹ�g+�]Is�
��Y��E|	�i�Sn���JI��xK|?��i��MX�7�uH��V�gLAߠf{Ւ���\y{6W{]�*#�Α�NG/Q���׸囥($����� �<���Fg.:
�R�������VY��ھ������?h@4.	�VI������Ǐ����׀3����m�\06E��3�q�-��K,d�[gs?�����+������LՇ9n����<��|���O��{�	�S��YbT�K����jmE���Α���6�T���o��s�X�k�����n�\=���s{����Ju�.iZ{S�ss��A܎�I�=;ĵ�c�-��%�dyV�鋸�BZ��_�w��$�߮6���4�S�*��)H^�.SDx��d�����2J��O�m���u�D/si(�ɳ�3�t6uqX
�&^m�NSe�{���*8�!P#��DF��X�`��d�OS*R$V�x	Y٠å�ތ)��ءO�����|;?�:@Hd���M�[�	�F��<�����(��M��FM<$v�$�,�F�24"|';��6���m2@�]o8rZ�Ku����#�'K�W��.���|�����Z�����#��]�LO���Y��-���l�ٱ��Д�?��nD���y��"�3��BI�%�
!Hm,(��i�2���XG7(Y{���O���q��1�:k?�v��1����<�9ʽ�tr=8���l��֐��������肗�t�:`�\��b��
�LF�R�8�Cu�CC��¤4�7��j�
�;�V)S�z�0�weR��C�����]��sAІ�ōCN)��j���*h^�,��	ۦx�!B���O�@2�؅5�����/��g8
׊�1��w�5C����i8t6��U�Ìq��x��v�z���T�/el�>=���L_5��;�T��)+���c�*���
���Dv���#M�P���Jq�W�Zàܒ̯d褹�#��\�'�j�sy�F�98�P]Z&	��F�����u����A�zV��gID6���ߢ�"���걆g�dAE^	1r�УL�=V/�����ܗT4�sa�2dOM���M.v������F*�b����P�岧�c$kd�"�o@=rcD-�q�0�L��~�(
�T
PaS��K���h���f�Hi�P�9���6D�%S��Iӳ�~�C�h�%����Uq�B��/��!yA'R�d6�!�s�lEL��mzǍ �_+���8�`����p����Ǒ���׾_�����5V�8 �R�$�P�Uy0����wC�	kC���( 1nkrr���9��4��qf���U+J�;Z�a�]XҤ��E����+\|%W��a�&^ވU�=� ����W��D2^�z��>��s�h�E[��x�҇@��
��4y���%S�K#�����ϐǰ�P���M�Jgֈ��ſ]]pێ����Ψp���E��C%�1�
,X�^<���L��fXU/�%�5J� ��ߺ(�6X�=�/��y�G�
="?E���,<�4>���=� ��->|�e�w�#��:����#��
�u�8w#п:����VL����ޡ����S�fS��=[Za�u������: k�v��Đ���0�VT��ԧ�V@E��V��
�F�rf��� ݧ
*q���(�2����j���c75j��
`���RV��d$�$������j#)�@��}�=i6�������'0>W���f\��f��}�y8ZY(�>��J	����I��a�Ľ?i�5XW�ߠ �b�� �G�<��J��j	$�۞�m������

��0�$�}:.9O~z�x�U� �2<ʪ �����C���*��D݁�3����D�V����x��K9�o~��� �so������/xk]�>pǁ���z�cp��&�T�$}ڂ��8�*iFu,~�7q ^`��W�J}_�NN�S�Z���������&�}��7�� ,)�ƒ�$2݅$q���H��C��'���"���g�i�9E����b��-3�4#��F�K���:u����t�$��>�ز�#�∽����x=����2����>Ԋ��`��BE1ʀ�RzK� �_ߞ����j�<�`����|8����or����X�{�'��j����ξ[�3�ؤ�j�6�W_��z����?0sPQ XjZ1{�Y�1���o�C`�.�_V��'��f�sP"q���[�+=�1�a����l\K�:���[�3�Y_�ڌ*��6	6������ߨp��Fd�"���� jQ��
6�rUq�[�n��� '����is�lO�	���O�%dY�@d�,��)���+u#�O�n�j��s����(H��&=s����(-�/m'Ì$�����y��*�>u��e�pW �5f�`�<��ѥ���Ŋиb^E{�c��p���ݖ_E���q��Z�'HZk���J�0���	8�1��q�I����\^��]�W�?\����ޖ���?�^!6��G$�*�)Yw�,p�J�8o���>��(B�y��2�v��0�	^Ы���j�[��n�D��"�d�[N��W�&�]/�h�R��B.	ٕ*��,_�\y����%�\���+�Gt��' o��~0#�cRg��=��im���scA��W��zY�1��j��q'�=E��eW�j~/I�$|�\fk��H�Č�����Fiw���a�$C�OӦ��#k�����P�;/���J�5�ų���(6:'�r�w6��;��W��ׯf1��9-3� �7b��ڊM����Q�2@���ލi`��M�(j�Դ����M�r�ΐ�uM�J�;�L����Fp n��_=&��V������GM^�݊J���7;�|Ɨ��S\��W�_�LN��������KN>3��U��0K�Ƨ���<.�f��!��49���K�J��$���@m�D 2��K@��)�f$�	ZE�Q���E����:�M[�k��SW���C�wV�~��S[�=�����d����߮D� �cv�#bO �C�����h�c,� ��!J�^0l'�`���,�@�l]�W"t/�RT���؍�����4֋{�����ye|_kT�cujX��;��K����l�d�'g�2��7����+��D"F��$ؙ�_��ܡ�j�W��Q�"S�s�l���hqc%�� T���0�t�~%l٬���85"���b| ah�5�rd3��	����@9�Z:�߁ &t1�Kb�����L�S��b�o�{�S�9p�&'֏ж*�yO_�� ���Ϫ����gxP*A~����[q~�K�B.oز<$�,,KU��'�OĿ0�*���%���1#�i�s��̮m���u=B��i�d
5M⁫44l!ȅf���E��3m�q����B{�z�=!��`��*%C!�ql-���<�5X�J4�M�ui`/r�(��E��g>�.1�t��>@�OD������@�����K[�l�R�йD;9�XG�g*sS���y�$ML6f�pJY�i~��Is�}H
�a���������9)����^�f�F-D@��/GZ$�2��B��*����i<�<}$�e\]��)��S�l�i��$����%�W��i��d[%��n��to�%Y���[���#�ɓ�҇.ޕ��ߗ.
S�@��c9�#���b��g�ź�G�m|O�hN��D(ʠ�����k��ҽ!�@�O�W�n_�Ð�k<.�(�3�B����l,7_?���I�t]1Hٰ$ً�sNc�Μ,���z����&=%3`c>��<� ���q���nC8=�/Q�
��W������p�9�L��Eᨺjf�F��GZ*ۦ9���Q�
�TH���Er\�g��uWs�!)��%N�n����$a�'�|�ȱ3��A�dw
����j=�̾�谮��
w��R�/8�ܫg��ՠ���B�u�}�:}�J�f�,��#�hN�̐	ɪ�1�M�a��\b�c�ų�~��wa�֧Q#��(����c�%LP��ԈMJ.y���[F�,��x!#Q�;%��+��m���5�'���Z��_�4�9��T�s�Cn��pE%�`�Ҷ3J14Eӆ�	��"T�_�~(M�%�T�ǵ��ڣ]`����7��OU��.����M*�<�E���NsS����4��8h4"�����,ƅ'p�p'obo���@=4z�.nQ�U�*|���P!z�b�E���{[��������Ww��ʵ��Z�p�o�6�+��ø��/���@�ڰ����e��a�K�Y!�>R� �Pj�@`{o�^SA�3#~Y����ܲWKY��Z�À��������R'�W[��G�V����ō��Z7���5��jҶ��؈5���N�|.��By��E�3Ga����������	��o�u΍�W�$�=�����Q�
(Ơ F���c �����Id�
\�f�)��8" ������w��7�MUm�%��brB���������A�їX�ѣmb<i�$`.kF����Y�a����x�<څ=�'�G9`��)[�*�_[">.���=�j&�Sj<y×^������6�^�}���D�p_����܀�?�>�(54�����d�����?,`Tٺ�����D#���b��ӕ��Ni��L�Gk���V�����uPV���\�F�N�1ySݷiu&�=��v	AW� m�*�[Q�>.�C%E�l�A�݄�d��c.�����1qG���e~U�F�R�������1Xr���=e�o��ԏqy��U����������)4���)N�%{�¸�b�vP�I[a��3�aWQz¼�	G�Be��͈��N;���KA;�k�i�g�W(��U>�C��J#���|zҫ�pš)��w�k�o��<��=��Mn�_�2p��J :�Ī����M|p��y�������|o*N�#��ǭ�̸O���M6e5~�<���{����4����$�gCJ��L��~)_�;�9!�����Mm�h��Tk��OU}@��r�;��Rb������Tw1�?R���C���F��c�.!$�3��Z\:�KM�y۳T����m��:]����a��3�D+7F�TH��1��1pԕ����-$v"�4����é��a!�J+�]V����q�d���}ֽ��ɭ�U�Kbf����/4��P�Yǻ�v����}aQ��A��`9]~z?��Rfp8�����	�hI��L;�Jh�l�ʖ�2 �W8�����V�*8������Q{kZ$� 5o��+�6�[ ����x*�#);Ġ�ʶ�J;/g�L��Z��>��t�G�rBWrF��OO
X�A�'��ʃ�����0���!?$u�S6ol��j�l1
(,ۂ@J�c0����V���`�d� ���[
�Oi�>�@\�r]n�e*�{�����kT�<?L���5���\��-�0�^H��/u�*P��riZ'^os:o$7Y81WB�"��^��H+�:�� ���15�V]�bW�?�9��p,Ti�Ks5RiYR
~���:��gX��Y���VB�I�Ⱥ�к���Hu��������E-mk8�jg���j���v��U0�v��	)`�x��z^�� F��sL9~�;���h��dp�*fR�,���j�\|�ɒ��"����ߘ�f<�����ЬZ9������E�Ɓ�����P����߀;�2�kED�wA)�0��[	����Ի����\w 2�"���vƒK�f���ƍ� ���L޶8����X�g^RR&�����j�RH�C��m��t��|yߗc0RC��[�!y�v�Z�Cj
�'sޚ�C/%�`�Ab��ؐ���t�UOaU���\�Lc�������ks��P�InZ�}U��ޯ0�d��|�~ZD]��-n-&�bv���.��l0
d|Ѵ�O$�(��P��o�)�ν��uscW:K�������F�Xv\�0;�g��Ԃ	ؤG�m���&ѺI����$35����i�>z��u��>��6˕��U�/[��"X
ʾ@�s�
��Ժ'z`*+��"�|O��I�p���R5=�Y��G2�*�����8��FKS)SK/���O⫇�)�$Ba[`7	�ؚm��UԮN7�|��T��8�Z>��Y��^�DņF�Ǹ�+"�R]�馜JG��f��+��1D>�+��k�e�;�	@^�H�l���
G�F���x����"�����>��"��t~ݘ40��ȝ�T�2�R��F�o
�m�o b�WT���6�8Iϩ@����#N;J�	RA��t��%��v;y��#>��ёт��ݭ����?�&�M�k�%5����5��{�Ø��x[/�������}=s,�";oW��{�~��kHiI�9%�i�jP���U��3��|�������S���bԂ�}�y|������4�Koz�$���v	nF�ib��V:i^�ˈ��G5"*;=�ӝ�2!��9�C�\��h�x�n�Rzc�]��~�O]epsD�.Sk#�i}���"�����)K�U�5�UU�uU��]�aM��YR�5q�%WSU��h��6����(r�v���HZ��Z�*Ng���:�L���!��x���\�ʵ��[?�i�e�O�'��y��#�rsA����V�l����F������$d�P;R`lEX���H
�ʭ�od`-i�i���5����u<��
��+R����:Pn	�%u�%��Y�Ђ��L���gˌ�Šǖ��f׺�#a��`H�
O?ĵ�O�A|͓A�]��Gnj��Iz�O�R����8�������:BI%���\f_�j`��*�c�(�m��u�� �[�m�|��"G���?x�>�R��q�h8�_O=3�ȳB�����Ӣdɚ/v���L�re�V�?B������昼 �)�΍6?���6+� ��~��[Q8���o����{���P�!C�|���zo^ƺq`z.���ׂ}�N��4�{�
T��ٔ8c������`s�>U��Gn��h�YEt{��.����=�b?H7���ԯ�K	�N��AD� &UU4�!��;G�@!�jP|	��i�M
����k�0f�!��?R�3��V9X��mx�T��g��R3+d.�Ǭ���yT8AV���0�=�7��[�%�f�d�fqEo���N�XD��q��b5h"���>d�,+R�X�|�Hco";5��v��v-_I���C�60�P������rN�K�ctlP�7�ýa�;/�L3���b��V���T�9�,��� 2.�%\�����_x�����xm����5E�s�W�p�p��0��z���4i�n)�R�`IF/��9;'7-w�kf�<<V�i��T�xx�����}0���	�%6�� 8����m͒��eE�������(��</d����
���7բ�ې�syNF�nDK`�������M�z���F�mz�zB0۷~��X~k�=�/��vW��!�?�Hg�M5l�پ���o��t�U�;��U3����<ݐ���L��3�c`򎲌L<w�B��ry�"J�2Т	�Y$�H��C����u��Z�J9t��J��tA�1����-�I�j��(�Y1 ��فz� �8��0ow?�\M�w�)K��=⼥[�w���f�T&�Cds��ivo�#C����3����xG�<�ǳC�ƒ W���ʍ��-%��!@Tg��i�C��2}T@
-��A�\��5�Ͷ�$m��%P�>б��W��/����O7#A��=�t.����5�Ix��|m���XV�s}ҷ�W r��@V���re�Vwֹ߯h�( ]������ns#o�j�H������L���,s{��ǁ�@tF�[z��'�rOR>@����(&��y���������+H�^��V���x��gU�l�xs��*��r=�0s�}u�F˻ҝ�	&���|����,���F���!�/�k�둫j>uar����ܘ����#I#Qa�ժ>7���xt7t��&�ci��/�7�vgh�DNXzV�5�]�:�4}�;!�)/&�LP��L��� �[})F<h�'��?��|p��I�_W��\VrfWq1���|̥�ǟ�������E%&�z�t7s����� |�L$�4<�nt�G�]�����_�٠�6U�h &&M�wd��r��FҌ!c�rDT��؃�%��;PsLg	,�	9���z��!�Dhn]���xF��u�J��^pM���V�QZ���O��NZd8�^������ilXl�@ߠH:���ֱ�Vg�}�,�"����n�Mh��Y��;}L�GIFr�GD�kѨ������Ԑ�Y�d5��1&����4�V��H���
;��<�L��]����&W�~�z��v�U��m�.������������H��k
�4܌V�}��Տ�&� a%��(/:�A�}Knn^^`�lj���|����q�S������_�Z�l�%��q�U_q��,�%x�M2�X)@#��CQ�C/���3���qfN�tTyw���]D�{�Po>�x����~��;8�����aD� ޥ�C��h���F�E't�C�%Ed���Im?}�o�"���'n#���ފh�z��䢽�iK�Hn㞘<�u�Q���U���;����i�s�|�X��]:;���[?��潵��Dd�wۧ��k|S	%��v)����F�����i�WQIDh���[�ә�	s|���=�t!��u(��]~P`����_�ā^���Xd�Ƞ�	��y����5Y $V<Q�[ ���Y��Y7s��'X� ����������G����we�ީc�:��V:��Y�v���	�x�q@2 ���`�6]����S|�+�$�G�T)���>+ob��V����ܸ;d���उ�Kd�逌nj=��M��� Oע�QLm+�8�w�(;�Ͽ���ah>�{Xl���Pa���X��GS%�G*�;�LJ7l�#&g�V�Ў�����F� Pmx�J���!�]�خx�V��p�n�Fw�n�l�%�ۯ2#�V�Puq����
)�.��2F�`09� jȷ� ��O=��·�*��"F�g��2� ����T�4A�pNB5?��-�b@Fb
��gͫi�L �s�w]$��� ��EZɚ�/���2�~�tO��L��u��SQ�'�^��KD��bg5�:��i;���C�����ž��Fܴ�HV(�����:˞��O��=ڔ�h��wΔ��R4R�gg�}ç�4�7-֖� ��B`�'��M5��s�to��g끰+�Ez\��k��i�=��7��BN��-�,%��6�����M�g��X�w}fc(���%A��Q"2?�z٬ݨ9������-����Δ�*O������]P�~ਹ�9L�giO�5�Z2\�Dl���G�W��k�/�#�խ��BP�z��s�� �	�Y�>ׂs|�2�퓃,�2JĊ���t_�{�Ƹ�Iy�P��cң^6l��R�{�_4�\;1'A<�����Z�π��iIk���EC�U�����m�)��Q����e�7�(7v��zMY���ݫ�E�?-��-�����i�؄���泲�M%fI�x�FhͲ����s�|B?b݂iiN��hG�&��Ens���R
��?+$AO���W\�8�H66t�&�Rh��+-��AaΩ@����p�!�%�3!�G����+t��&�	T���@XC�Eբ�����K�*B���F�����%d_ֵ�cզ�����W���q��[�����<.źN3W������,�rаY0 �gr1��"3��$H�(=8�{����A5�P�]E�\̹!y[��"�'�XL�].��U��?L�DZ��ЈOB�⪛�Wp��z�5b�s�����{L�&�0��	��e�������H�^e���6��+gS��#�w�~J�tp��F�\.����=Qz/��\
�����W+E�>�*��i3�Ҙ���,�����h-��k��"_�6ny۩=���v���U��9�����+"]��HmO����N��w,7xQ�]M�A]C�)1�<C�1����+y�M�^��rl(��e� ��&lF1�TS@���LD3A˳��zp)�X''{3�%b��4y�V���j0TSF�bL�@��8֏��mLE�X��mw?.��ؒ���i�ט����(��݁���jmd���a�B>J�qt���؂�&ZNY�%���
�K^?�v6�FlC�v�E@
����:^�th,C~緝�,q25 �