��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\����q�?��e�I8�b�Ǽ$��"����ׯ1�V0���ϱ ���u�ӿ����9����-�~�a ��?7e���:�n�1����P������2�k���j+b�_G��+~Sz`fy�|�`'ݴi�*J����#p�"�0����aL{�:��{�ʈ��.���P�gt�B�S`^�RF�$����X%�ft��8�N�����Aٰ�M������'M���V���de;�ܮ\]��G���8(ș���K�-���m��~�J�Qi�A��m���-��X��x��qc� �t�ϕCૐ�\�s޳I�te�0��>0Cj�t�	�-�hc!*
��I��ڸ�(7��E�_ ����D� z,��������o@���[=ov�e]V��YB���u�j(B�v��$7D]��HA;�\��x�痓�0C���z��s2 ��T�vf���Q�:ׁ~P9>J�]��j;5����9�-�A`�r�r覺��	A}����������Z������N�ef����،hY��1�R%�  ���t�*��h�~�_r�N�eB�Z�XҠ���Ia���NҪy��{@��*��~��MH}ݲ�x�I�>a '	�x苃ؖ�K�r�����<>:�S��׋����-���Duu�:�U{����l�`ɍ��놾��Ш�'(3,Će<%�}l�1y�!�������	u�q�2hhǢ�o�V�����u^@!�m�/�H�.�4i�]�gW�r�Sk�J��&Y�Z�b<x�=b��'�<���rRM�"g�Z%�ޭ+��ED�V2eT ����S$�?�����o��i��������7�|��
���E�o��*��*7g��&U�#a����&�|`��������"���}h�Ф���-�?9R���a�O�j��kc� `C8$���{c������F!;{e1�y��_����5�Պ��^�(�gď9|�Y��I��"��ǋ>^2�k?��_o�P����d)��7�E*Ϲ�WM�i����R 15��:p�5L���eI����t�{2.�5�Ч.6V���P����;�spi�\��'�{�(�j-�঑"��j��ú��6��{��J!�qg����UC���3��U�e�8Q�����a�,3\�G�/2c��{��OA2��T���CR}~g���/���[�h'�ZR�ֶ(�h�<������u�ۖ�^B�,+��<gam/�L0� ��mV%��3,�[��s["SF|Ri`���]�'����~���av>�]�݇���I�@��A0d����ނ]n���L�n���L?�& �dg4��<��}�-���
z��B����t��@n=h�kܙY��ֱ�¯&"Yϳ0kbyoX�v�5�s/4���Tlw�%�%8�>;����G&]��n,)����֧vf�3�=dS���������z���Y���EX����O���]%;ʹ��Ʉ�'��L�r������f�$ɿ�
d��q�`���8=iZ���!�{������Q���͞��1���}�b�ԣ���ݬmm�ĭ���ad��f�XF>Gi�F�H���X������{a,��UF�����݈�b�Ae�I�Ae�s��u�S3�5���Yy[�s0�9�-�H���'h����K�����9�d~��
��%r��V��;�o�&|9hr<��!@5�лi�����\a��E^qA� �i�G����z˲��SmZ�&I�C�)�X���k�W���с��gF��'xg�Ψ���`��1S�͗�eFwֱ,��=��cq�:��A_E5�I���ƚ�TT�4��R$�� �^ޡM^7���w�D҉.���>����$>�v��u��e�|�q�P���ܵ6z��+6�C�s��k�z��ͭ�G�ң��|v^Of���)H]�;(�ڊ�A��4�������q[���l������YƦ�c�l,�g�y����27:�I�1R�}E}�1$x�.>톶0�̅�2�T��lQ�>���o������$�$*r��ģ]ߋ��?_n=O(x͍�e����(U���5��˲ sW��s�S�EF�8��8툉���Lp8�`X���#g���ό�A�-�e|*�� �n˼�>�sk��<o�o�LF�u�@���UZ�A�L�bAY�;_�|xyp�0"K�?��$w���'�a�a�}L�74��>�����>���@�n��p2ە-���dL��s�&�x�3�ݳN�k�ֶ��m�d��ҫH���]�0�D�r�>��u/�[�u����2���G����P7�N�l݌��CY���1�h;�R+��r´FZ%q(!�c�����9q���-�%+ ��(/w�5:�1��漌�,��̢L�rg�B��@�"�ٞ�5���f�4��-�zh��X�Eq~t������	��m�dIz�}x:�支��.g�|��ͥw]�A�\�{�
D����N���6������MJ�=�Po�aG#f���"�S���X���|V�������>x[�U��Y�DkNv�|~=�����b�il�{��e>+2�R�ܛm�85'4��٩�y@�7�}���F�=n�u~�#�1k���$���
}E�<�R"�&�П���S�0-�`:k�R޵��l��<3dZ$��Y,j_k*"��<�IK,9sM�|6�����P�ˍl�dQ.l��0�Qє�qv��o��$yD��Ǩ�b��<ͱ���Z4��=�X���]�q0�������Ƙ4�?(�g&�����˨�7���X�gq;RO¤)��َ5��ϙB�����@&UB���[�u8�0ܕ����?;�{�:�?��z���8�޼L93�F���q�܂D8S�ӕ�T� M쭯u��VW@`ɢ'0v�L5�g�?�r-	��9��ƲS�♯h���=iMy#��x�y��;����?\���#[��`?�eΛ[�]�ݹ��=>����)��FKF}y�}:�E��:j�2���d%�VG~4�Iy�8�qE��	C���X @Cx͙�=�誣Q)P3ViD��G�]Kϰ:�.��3����~�m:��n���(�������j~tL��� ��c��>��G�#b�z�ze#0F��U{���ht�5�ɳ�x�̐���~a͘�?��$١�PM�C5�VӁN�b��jc�UM�z�B�ˉ�Ib�mz���d=Q!-�O�����ܗ¥�j�6���q&��'��)�q��6�m�6�s��$�e'pT��N���tjI_�<ot��b�\�x�L�,	y������NTV%���nJ_h��ԗ�4���+���-������l���.���p���V�n��8{�2����k��k�CҶ]V!!n�J�Y=uc��6�E�hhN�
{),4��S,�6��2AG�33�c�B��v��Mw���K�["h��G���d��Q�?"��SFֶ1k5�Z�YO8o@E�| �L�lN�1��4�$�%)�"�ԕȒ�U���a{e~��L	8�fl�ջ(bW�F��r�"��F�1v�ds&1��J�+Q�%g�����ŧu5+�(�r�����>Y�}S#7b0�HgX\��X��W^���o"2��m�J{.���"�=qdV���Yý��Vo�xEu��c�nR�G�9(��¼�}��]��AfJt+�@�,�ZگL���]�v�9���|e1���!&��8zY*
����Q���ķd�r���ZnE�f�ЗE�w�\Ք�����3�Ko������T���o�ߟ6D�\)�bN���J����8�~��1�fdb-�8m�Ab�����>�J9<vc奾2��iŝ�Ӓj_b�%-�
��c�Cނa�
�oQ���v���(�8� 6()X��<�2��'�R~�H�͏�HR��)ӢE��4��S渓1�B�x0k�񳡷�FO�G���'+݀F'�H��|Eb�d����tŚW7 �M�~{|<=��Y�x�g��B�����%����Y/+�w`���)*>y�C�Ȧm�N	m�ԩfԾ-gtHx�r,^SWx�l"m�j���}C������9��REQ�_>�i�2�!X9��4An��}Aڠ�I]ۀT%�������x���%j���2|X8�#��u^�����)�K�����FG�����;]�s�f7{V�)�S��g�`n�s!����8�޸
C�þ�,����}����T<ճ̀� ���	d�V�l*�'E	��x���P�U��L?�����Jwٲ��)�;�����k�_���M�G�<spV�:��,�b*{K�83��
�����֥D���072�����U{��F�D�euX#/�9[;�딃��I��h��0��1lw<�T~�)���Ѿ���g���K�D�Va��[KXX�D�WE3�4�%.��B�矴�&1�T0�?0�m�y~��i3�ߤ�U�]X%��=*�PR�cXc<����xgì��^���2{M5�^��pOxdlq�ކ~SRy�,�!�Y��B��ع�vt���a ]y��d~�p�K��imܒ�k�!�fP��Gg�M�oF�~�TF��%3AB~�n��EJ��ƽI2]�}]}L�m��v�Vy.����lM\F�����F��Ϡ.���x(�d�&��j�,��9������<�/