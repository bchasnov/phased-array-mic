��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\����q�?��e�I8�b�Ǽ$��"����ׯ1�V0���n\��ՑV����C?���A:Xr�D���)����08g����X�#�����O����Ͻ��F�敠X�e%jE��@c�Y���ir^��<�	�!_AL��~q����	]W}6�2�_�C��������FЍ�m�7
��9bd�2�>��|�G3��޻v�nI�~���YqT���Gb*Z�=�Dd�h��UI�J���M�=��G~IB�W��e�>�W�^ذzmg���D�/ü���,�Z�!}_�e@G�d	["���-(�� a��<�0_:�p�&�$vl����=�ǳ��m>z
'�yc�����C���kI\|�t����L�|�5T��vXl^�N'x�y7	���;��\��H�m[R�b�&X)0���1��+���j��1C���j~k����kw%&�;T��Gl��I���]H��9��G����5V�R���,m�����'��ڛ�$m|���1m�x�C�A�I�#�멘̲L�����Z)r�����`	��׋�}�Roc���{-f'�?D��
t��U�KmD�	��ux�(Ó�.ȥ�n�����ۀ�Xa9�mV�F��B|b \����G��Kh��r�։mY#�)AS�z^���Çr�����*���|)�<Y��L}tdv�v@��CFq���"�N̴�����I�?����U�&��LM:�"���f9��?�>b26� ����&����W�E�~m��ϽZ\^.��[�/Hش��
i��(���Y,5�Id~kC�.qf"��yI �o'��s.�CƖ�]�Z�iu�����8_X��C�X�r'w)o/a���S� ��b
�v-�I�C/�@�I�|�_g!��Y@͏��g��Z���Lʈ�o�Bg2�����˨t�I���3���Si$l��d���N��_�lF*coM�8z�t:[��
��=���gY��:�QTߗ*��\�T�D�*΢3ĺ�~�C	]q,g�hQ��m�T��}{7��M���Lۍ��Oʇ�Oa)&�$�B��oT�58��5�YUX��@�
 a� �����.v�a��#Z�_��Qt_�	�Ƽ}������T)E,+0g��pN߷W6J��Wg��	��c{8v�ʔ}��J������XT�a/�t�ȃ/�^��f����I���sȂ~�:A����mV38P;d��Ǟ��;c�3�#��Q� ��$*����URFA��vpu!B�g=^axFp��о��﫳�.�|�2��JB����Kʪ_��s3�6�<�A���ƌ'`�.�ء���ƍ�@Q��a�fX����pB���ܵ��HA�T�n�*���wƼ ˈX��;&�Yˎ��~%��=��5g�a�}л�2�ɹ�0� Н��x���U�A���iz������Sqƻ���fD�P�ȫ�����^�������8��S�w������)p�;m?ѭF��K['�5�oN�ݞ ���&�͊,Up)WQ6!]�� r������ߏ֠�9��t8uQ��H��F"��.z�����^���%���h�+��%���Y~���"�!��j=���8?���b"La�Y'�\-w`S�1�y���؋��Ė��k����{��&����ʡ4��U�Hv�jg��������jZ;��s�ȿ2Ҟ�z���T�`��Ԏ�oõW�}@[�N��̐���}����S�Ω����}�nBƚs��/��er�b�NL��.��bj���TI1 �Ͻ3Q�iu�9�#
kp�ɮ�
a���}�Bq��}XԢ��x�t���Ѷ�F�����)�O��{(�C8�E�[��k�/�2��E�����8o�i�i[ w�B�N	+U�����v%�3RVǲ.I�>�z5^�.���ݍG���ޝD� ��,���˳t}8Ƞ��P��.b�}ĝ��{
��"����;ӯFt��]�s� ��Jp'2Ҽ�ukZMñ7��g\�\|����I�D�<��uʼ=;l�p{1��n���*v�m�YP �1���N�'%�sE��@n4П�x�1� ��3������*?tO�R��"˃��L�jwC4�H�������m0mݖ&�iC���G )���W����&����[o��#�	��=�3C�?���m�a^P�\i�+�`�J}���k�����"�+�X�c�!͛�;�y%�.��6�|��}D�x��C�ғF_���UA.��Jl��0b�Q\>��A������Ub�E�g=�P�QV�}w�i����2��8����u9]E�H){�nI1�Z�2�FDOռ���c,�F�4Y}��#A��l��_�0\��lO�KU9{�f��qx2>J�S�'�G�L�9.�c}�7pc���`Lb��r�B��İ�$z�sV�j��r�7���Ѿ�:d5��y����'�Yg�q�V
�[ k�DC���(P��bYt�������E��-������d3�|����U5��r����K3RkU��
g�A�)�I3��;W�?���P�7�"��ۑ}Wx��-��{�L��oh&��QҰt{��]���s|������L�<���&�j���Z$�KH�M��|�=8����'��f4<T�3B.�-ҎIQ�d�ڡ�ɪ��U�/ێ�ɕ�:F���"�*w�s���7x��_�<$����@�uF ~�s��&��t�Z���Z$�10��Ⱥ��g.ʦ��8��� �u ����x����P����W�'m-���#m��j��ø�J�4�+g��\բ֌��J��R4�au�H�7zY��_�m}�bnD���Y����ʴ[}P��͸&A5!-w:�U�˔�����MR��j�"�����@X��:pf[�e����R�b������J�ܠJa���f��͔��E�+�D��g�qf�I_�m�U�r���K�9�V��#j���E�`�3���}Q��d�8�@F�R����DB��"~�B�K����D9�2�����;����%-2p��螸k��ޣ,�������-E\L���UX�.`�n��S�/����u��p��btgX8u?�+kK<
��<q�!�ʒ��
NkK�P�1F>h����H<�륦"���[I�2S>Q�M�
���aucbB|>��˻�y�Pu��3c��r�s/ Z݀�����,\&���5ge�@(1�3��R��/tb0Qߴ��C��I� {�����|��6�;]&��'�C�^H����w<��h�>L�����EEm���h_z|ȾY�n��3�uL�U����!�f��sA�ư�]D�u�I�K6�5�>����)"���*�E�2�����@Dh���
�Cb�o��FxS��T�t����N\0��JsH\�p���XF+��`q�Y:�f�E4�ked��&�_�f�+KB6��x����o�qPC�`P�.oƏJ�d�0�q�o��	����������[Ǝ�XZG��nQL�:�;S'�N�&Z;Ϳ���P�SJ�kW2�چ��z��-ӭ�٠�%���d���|����ii[�H�x��ʇ�@G��_�*%���{hZ�bCv\p.�M��~ ��*a�l�ӕq�W{=�yb��2W[�%�#� ��uA�]-~��Y��7#��[�|0�����Ft?V����@aNq2x)�a�=�����@׻�t��oln��7��Gx�8��+(�7��� 
������i�&�p���x|�\�8�
�V��8 �2	�3��S�����P��M;�z�B1G�`7^/�e���8\*�}5XR������,N��j�H�5��M�w�^xw6=_�
9E�2�P0��aS���6� ��Dd�2궽8�s]���M�����Q�e�KL���ì;{���E6G�󍶅z��(Zwi�����癫	��9�[�^s	��� 6�6�V.]���E\:�đ���Qju�,��ؙH��K��6�-a�s1X��M�8"��o���m�F�2b�3�S�:�
���^r���c;I��US�|�0pt	
d������fj��u:o3EŶ��+ܹ�͝)�,z���kͯI>a��IL ��Z�}K��[bq�&t�߄�yL�2�.f������g����Yͥi���0m�2GjB]Z�t!{0��S4���3.sK��@�[K�����,8M���)��|���]qS�̭E�8;8���.���Gڷ��/��ɗh�-'ϝ�i�Bp�2��&�%�.R�kإ�Zo:������6�����ZZ��n�F�n��l�ω�7�9m;�@�(�3;������`ͩ�W$����L���U�f��o����� :��`�0f&&�:W��d<7w��2=	�ŒP9O����'/� �\{R'e�޵���$w�����b��)R���Ӎ�?�/P@�(����Ť(�L��lŢe��������q�g��EW�ޱз���ӆ���2=�a��p�i�G\�G���=GNEě�O�I�΂��L^�`|χ�<� c��OZ����3>?r�[6�2��?EԚv(�� h��έP<bxN�j�X#L�.�����e2M�钆��~@9�aCAP� �br+k��סژa*6�r�P>Y'�F��pڥ�.����&��#�O�R-нw�)D�6�%nx\1o��Z���D��W����"��RS��=�݆j�hj�3/� ��rv��pς懅��o�ie�mb*^cUse
�����F��o��5��H�5����iJS��)�Pň�(T&� s��Tt�cN�q���z�ï���q�WY�X��|5���*���@b���ؖNV�A�̦
3f�a�G��<D@���2AC ��j���r�������Ka>N[,Ǒ3�h)��$�B�kQ�
j7��:O�h��A�r�b�Թ�b�3��u�3@�	0T��Rъ!웲�ݿ..�
q�,���&��}B�H+��P�ؓU��Uw5��B����A8��ٲ����A֖�:ǮH"���Gi����95�a��b=�*�`�]�<�W��x,���zbe��{��n,�h\��o�2.r�v�f���t�t_��Yw�������W��v�h�L�����C����&".x�+��:�9�d��kz��6h̚��>T��a�:���c�B9�Ƿ[�]�Xb%&�d��.�\U�=����D����vJdPfd)�����*vv)�8��~R�H��������x�� E-t�E��dˬ����{Z���X�0�z�����a�B�0���� �����T��a�4���A,<el�{f�q�̅~�$�7��4.v�Őt��Eb�	G��6���%��nX�C5m!��д�9��^Jx]>[,ư�f�x�Ա��w�R���7��敂ڲӈ�)ш�ڮ��DFXY����#D���z޶@��&g܎�{$��'���Y��3qE����{a0��){�3�Ю>��S:�J+��&N/����'A�~4�	~��1� N\^Yӷ��9�Q5g�|�x����|����8lO��E;q���V跕�e��z�Vʚr�?�~�n0u鈜�X-�i^0zVlv�iu6�rFΌvb@�~�|��>hr�YZ,�/~P �l��QX��h}�TO��b`"�󴥀�&�����@��d�҂��/�ɮ��+�c��kW��`�E;Q�o�~?�e�p����r�hzcb�B$n�V�A�Ǜ��1�b9�}Z�V��������B�	�	׹�G�H�m����n�j8S��OG��;N>:u�HN�uQ�Yj���[?�m?��?xv\����1��(��u
P���}L)��U�]Z��Q@�l�c�*�Y�Nq�VxD_L���H�	�f�����(�����XHE�^F��0L�=·�j
t�L((-��^�#?���E�U/��:��K�9lg ֒��$T��b�����qZ&���pq�U	5l�9+4�
ՉQp�U~[�8	��;���x.̚Wl����h�S�m���[�����n�Np�_��ӻrp:�4Q��d�6$�2�'3�� Y�=xS���]��i��3�u8l@<K�����i
:�!���ຓ��Y�C��y�@�P�$�"y/ �B�q��O�X��b/S.5�\���[.J��j|bFīތ�=՗�h��9@Jh�@���M�8mw�t�g��@�"�#� C������=�L����Cܼ��Z�Lb��BE�TG9��_�3e�_� 7����<�&����"��D���zj�
e46M�Z�w�<��Mt��"l��+K<i�|u{�X�ylc�}��Y� ǞW�N!����=	����&(�-���	;!X.�`���Ƣ��ٍ���;L��%|��>�b�G�"d��\TCj�,P�0v��M��\y�=zw2�ID"�.@|�t���+hY ���v8�4z���MH �/��%<�V}��ܨ�uA��@ ������M����mW8�Ni��;���}0G="�ޭ
�#v[�6�+<�|��Z�^��B EA��,)�DFF�Z�B��P �\�бɌ�u�'I��H��3�|Չ$�+Mm1���*�+�A��ە�p�+����$�2I���̍������3@�/�`�F)�}�k'P�(�U��LȒ�Ņ�5�,v����X�<�S�P���\M�~8�._��TB:Wj�!�-�%f-���8�t��-vG��	 ��`��y�r�X����{�����.!1��P,�P�Zw[�kše:�?��3i!Ր��Ch2u\ǽ�L��\�I��W'�SH]V����ho�V��f�N���^��J��1��:���N>sS[��^$pc��d��|�Z4��3~/�G��M��s���9 J�&B��ퟩ����Qbv�J��I���1'G�{r$˯�X0q}B#H�4!��ht�A�y�h�{b{�+�3��k����4ŵbdYM����k��nZ'5���d��+��B� v����ɧ<�szFl�A�
���tP��U$�!yQ����(�5/����0�8|B����K��#��(\��Fz6a�1V�r��i��jP�ߌ��ʰF�}��Js��BӠ�0�z�V���2�n����|P�j꛵xiS_[>Kkyyܩ�[䦸�����˯�q�Ƕ��QI�6o�&�֔HW\���N�e�~(V�CSKQ�gJJ@.��$�]>D�X�E��!�je]�����%R"XmXd
wO�hD,<�{S4����9��Lk`hS﮵=�_	��[�Ӡ�X��}q��!� ���<��(��"S�����f�֘̄)�܅T���#���ܦ���Qdpس�����Z�xX'�ƛN�=՜��������<V�	� ���ʵ�4}�L)5Y�(k2O}pӱ�M����l+2� ZM�85������"7/�C�$�SX{+�X��\A?�J��ZΡr�* �@9sF<�J��
���
�T:�l9f^59���f1�t0��UmNYh���ªɽ�ߧD��?|�o`�si�k":Ky� ë�Y�I>�kQ5��?�h��
�z���OeeU�JMIM�M*��Ǎ�y�(���D��!�>���]��K�c�x�Oj|r\D���9��s���k��bv@
�;���zwM&|����w����e�ϱ�9:]U�m�G�:���L����E��u�DG�Q62W�Dg[�Y��<*�`�X'����4 ���M����I�鱝~����OPp��0@�r�l��DF5��-�����C�Bڊ��xH�(pP|4���pL��g�N��:��W�O�p�1Lӻ[�tW�(r~�Э(e�	#N�Rq�(e��e6vC�Ν�ӫ"y�T��N�=u�
�n)1�.�e.�"�(OgC|�N[?�P�47��{&��an���߉�iRf�!�ByǪmu^������O��W����X���Ee��1����߉��{�X1�ȥ��]U	��{�	:�g�������u��ZR�_ִ<9fK7�����^�S�-���+WyKA�ܒ�^�.��Zqe�J(�K�����|������^�D����ḘIئ׷�Ҝ�1%���"�Q[�{���穇�qF� Lʿ