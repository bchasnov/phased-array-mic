// Copyright (C) 1991-2012 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// VENDOR "Altera"
// PROGRAM "Quartus II 32-bit"
// VERSION "Version 12.0 Build 178 05/31/2012 SJ Web Edition"

// DATE "11/21/2014 14:01:54"

// 
// Device: Altera EP3C5F256C6 Package FBGA256
// 

// 
// This greybox netlist file is for third party Synthesis Tools
// for timing and resource estimation only.
// 


module fft (
	clk,
	reset_n,
	inverse,
	sink_valid,
	sink_sop,
	sink_eop,
	sink_real,
	sink_imag,
	sink_error,
	source_ready,
	sink_ready,
	source_error,
	source_sop,
	source_eop,
	source_valid,
	source_exp,
	source_real,
	source_imag)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset_n;
input 	inverse;
input 	sink_valid;
input 	sink_sop;
input 	sink_eop;
input 	[7:0] sink_real;
input 	[7:0] sink_imag;
input 	[1:0] sink_error;
input 	source_ready;
output 	sink_ready;
output 	[1:0] source_error;
output 	source_sop;
output 	source_eop;
output 	source_valid;
output 	[5:0] source_exp;
output 	[7:0] source_real;
output 	[7:0] source_imag;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_sink_1|at_sink_ready_s~q ;
wire \asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_error[0]~q ;
wire \asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_error[1]~q ;
wire \asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_sop_s~q ;
wire \asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_eop_s~q ;
wire \asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_valid_s~q ;
wire \asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[0]~q ;
wire \asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[1]~q ;
wire \asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[2]~q ;
wire \asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[3]~q ;
wire \asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[4]~q ;
wire \asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[5]~q ;
wire \asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[14]~q ;
wire \asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[15]~q ;
wire \asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[16]~q ;
wire \asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[17]~q ;
wire \asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[18]~q ;
wire \asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[19]~q ;
wire \asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[20]~q ;
wire \asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[21]~q ;
wire \asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[6]~q ;
wire \asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[7]~q ;
wire \asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[8]~q ;
wire \asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[9]~q ;
wire \asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[10]~q ;
wire \asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[11]~q ;
wire \asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[12]~q ;
wire \asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[13]~q ;
wire \~GND~combout ;
wire \clk~input_o ;
wire \reset_n~input_o ;
wire \source_ready~input_o ;
wire \sink_error[0]~input_o ;
wire \sink_error[1]~input_o ;
wire \sink_valid~input_o ;
wire \sink_sop~input_o ;
wire \sink_eop~input_o ;
wire \inverse~input_o ;
wire \sink_imag[2]~input_o ;
wire \sink_real[2]~input_o ;
wire \sink_imag[6]~input_o ;
wire \sink_real[6]~input_o ;
wire \sink_imag[4]~input_o ;
wire \sink_real[4]~input_o ;
wire \sink_imag[3]~input_o ;
wire \sink_real[3]~input_o ;
wire \sink_imag[5]~input_o ;
wire \sink_real[5]~input_o ;
wire \sink_imag[1]~input_o ;
wire \sink_real[1]~input_o ;
wire \sink_imag[0]~input_o ;
wire \sink_real[0]~input_o ;
wire \sink_imag[7]~input_o ;
wire \sink_real[7]~input_o ;


fft_asj_fft_sglstream_fft_120 asj_fft_sglstream_fft_120_inst(
	.at_sink_ready_s(\asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_sink_1|at_sink_ready_s~q ),
	.at_source_error_0(\asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_error[0]~q ),
	.at_source_error_1(\asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_error[1]~q ),
	.at_source_sop_s(\asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_sop_s~q ),
	.at_source_eop_s(\asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_eop_s~q ),
	.at_source_valid_s(\asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_valid_s~q ),
	.at_source_data_0(\asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[0]~q ),
	.at_source_data_1(\asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[1]~q ),
	.at_source_data_2(\asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[2]~q ),
	.at_source_data_3(\asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[3]~q ),
	.at_source_data_4(\asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[4]~q ),
	.at_source_data_5(\asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[5]~q ),
	.at_source_data_14(\asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[14]~q ),
	.at_source_data_15(\asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[15]~q ),
	.at_source_data_16(\asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[16]~q ),
	.at_source_data_17(\asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[17]~q ),
	.at_source_data_18(\asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[18]~q ),
	.at_source_data_19(\asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[19]~q ),
	.at_source_data_20(\asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[20]~q ),
	.at_source_data_21(\asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[21]~q ),
	.at_source_data_6(\asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[6]~q ),
	.at_source_data_7(\asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[7]~q ),
	.at_source_data_8(\asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[8]~q ),
	.at_source_data_9(\asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[9]~q ),
	.at_source_data_10(\asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[10]~q ),
	.at_source_data_11(\asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[11]~q ),
	.at_source_data_12(\asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[12]~q ),
	.at_source_data_13(\asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[13]~q ),
	.GND_port(\~GND~combout ),
	.clk(\clk~input_o ),
	.reset_n(\reset_n~input_o ),
	.source_ready(\source_ready~input_o ),
	.sink_error_0(\sink_error[0]~input_o ),
	.sink_error_1(\sink_error[1]~input_o ),
	.sink_valid(\sink_valid~input_o ),
	.sink_sop(\sink_sop~input_o ),
	.sink_eop(\sink_eop~input_o ),
	.inverse(\inverse~input_o ),
	.sink_imag({\sink_imag[7]~input_o ,\sink_imag[6]~input_o ,\sink_imag[5]~input_o ,\sink_imag[4]~input_o ,\sink_imag[3]~input_o ,\sink_imag[2]~input_o ,\sink_imag[1]~input_o ,\sink_imag[0]~input_o }),
	.sink_real({\sink_real[7]~input_o ,\sink_real[6]~input_o ,\sink_real[5]~input_o ,\sink_real[4]~input_o ,\sink_real[3]~input_o ,\sink_real[2]~input_o ,\sink_real[1]~input_o ,\sink_real[0]~input_o }));

cycloneiii_lcell_comb \~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\~GND~combout ),
	.cout());
defparam \~GND .lut_mask = 16'h0000;
defparam \~GND .sum_lutc_input = "datac";

assign \clk~input_o  = clk;

assign \reset_n~input_o  = reset_n;

assign \source_ready~input_o  = source_ready;

assign \sink_error[0]~input_o  = sink_error[0];

assign \sink_error[1]~input_o  = sink_error[1];

assign \sink_valid~input_o  = sink_valid;

assign \sink_sop~input_o  = sink_sop;

assign \sink_eop~input_o  = sink_eop;

assign \inverse~input_o  = inverse;

assign \sink_imag[2]~input_o  = sink_imag[2];

assign \sink_real[2]~input_o  = sink_real[2];

assign \sink_imag[6]~input_o  = sink_imag[6];

assign \sink_real[6]~input_o  = sink_real[6];

assign \sink_imag[4]~input_o  = sink_imag[4];

assign \sink_real[4]~input_o  = sink_real[4];

assign \sink_imag[3]~input_o  = sink_imag[3];

assign \sink_real[3]~input_o  = sink_real[3];

assign \sink_imag[5]~input_o  = sink_imag[5];

assign \sink_real[5]~input_o  = sink_real[5];

assign \sink_imag[1]~input_o  = sink_imag[1];

assign \sink_real[1]~input_o  = sink_real[1];

assign \sink_imag[0]~input_o  = sink_imag[0];

assign \sink_real[0]~input_o  = sink_real[0];

assign \sink_imag[7]~input_o  = sink_imag[7];

assign \sink_real[7]~input_o  = sink_real[7];

assign sink_ready = \asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_sink_1|at_sink_ready_s~q ;

assign source_error[0] = \asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_error[0]~q ;

assign source_error[1] = \asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_error[1]~q ;

assign source_sop = \asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_sop_s~q ;

assign source_eop = \asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_eop_s~q ;

assign source_valid = \asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_valid_s~q ;

assign source_exp[0] = \asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[0]~q ;

assign source_exp[1] = \asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[1]~q ;

assign source_exp[2] = \asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[2]~q ;

assign source_exp[3] = \asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[3]~q ;

assign source_exp[4] = \asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[4]~q ;

assign source_exp[5] = \asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[5]~q ;

assign source_real[0] = \asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[14]~q ;

assign source_real[1] = \asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[15]~q ;

assign source_real[2] = \asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[16]~q ;

assign source_real[3] = \asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[17]~q ;

assign source_real[4] = \asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[18]~q ;

assign source_real[5] = \asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[19]~q ;

assign source_real[6] = \asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[20]~q ;

assign source_real[7] = \asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[21]~q ;

assign source_imag[0] = \asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[6]~q ;

assign source_imag[1] = \asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[7]~q ;

assign source_imag[2] = \asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[8]~q ;

assign source_imag[3] = \asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[9]~q ;

assign source_imag[4] = \asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[10]~q ;

assign source_imag[5] = \asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[11]~q ;

assign source_imag[6] = \asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[12]~q ;

assign source_imag[7] = \asj_fft_sglstream_fft_120_inst|auk_dsp_atlantic_source_1|at_source_data[13]~q ;

endmodule

module fft_asj_fft_sglstream_fft_120 (
	at_sink_ready_s,
	at_source_error_0,
	at_source_error_1,
	at_source_sop_s,
	at_source_eop_s,
	at_source_valid_s,
	at_source_data_0,
	at_source_data_1,
	at_source_data_2,
	at_source_data_3,
	at_source_data_4,
	at_source_data_5,
	at_source_data_14,
	at_source_data_15,
	at_source_data_16,
	at_source_data_17,
	at_source_data_18,
	at_source_data_19,
	at_source_data_20,
	at_source_data_21,
	at_source_data_6,
	at_source_data_7,
	at_source_data_8,
	at_source_data_9,
	at_source_data_10,
	at_source_data_11,
	at_source_data_12,
	at_source_data_13,
	GND_port,
	clk,
	reset_n,
	source_ready,
	sink_error_0,
	sink_error_1,
	sink_valid,
	sink_sop,
	sink_eop,
	inverse,
	sink_imag,
	sink_real)/* synthesis synthesis_greybox=1 */;
output 	at_sink_ready_s;
output 	at_source_error_0;
output 	at_source_error_1;
output 	at_source_sop_s;
output 	at_source_eop_s;
output 	at_source_valid_s;
output 	at_source_data_0;
output 	at_source_data_1;
output 	at_source_data_2;
output 	at_source_data_3;
output 	at_source_data_4;
output 	at_source_data_5;
output 	at_source_data_14;
output 	at_source_data_15;
output 	at_source_data_16;
output 	at_source_data_17;
output 	at_source_data_18;
output 	at_source_data_19;
output 	at_source_data_20;
output 	at_source_data_21;
output 	at_source_data_6;
output 	at_source_data_7;
output 	at_source_data_8;
output 	at_source_data_9;
output 	at_source_data_10;
output 	at_source_data_11;
output 	at_source_data_12;
output 	at_source_data_13;
input 	GND_port;
input 	clk;
input 	reset_n;
input 	source_ready;
input 	sink_error_0;
input 	sink_error_1;
input 	sink_valid;
input 	sink_sop;
input 	sink_eop;
input 	inverse;
input 	[7:0] sink_imag;
input 	[7:0] sink_real;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \data_count_sig[3]~q ;
wire \data_count_sig[2]~q ;
wire \data_count_sig[1]~q ;
wire \data_count_sig[0]~q ;
wire \data_count_sig[6]~q ;
wire \data_count_sig[7]~q ;
wire \data_count_sig[4]~q ;
wire \data_count_sig[5]~q ;
wire \data_count_sig[8]~q ;
wire \data_count_sig[0]~10 ;
wire \data_count_sig[0]~9_combout ;
wire \data_count_sig[1]~12 ;
wire \data_count_sig[1]~11_combout ;
wire \data_count_sig[2]~14 ;
wire \data_count_sig[2]~13_combout ;
wire \data_count_sig[3]~16 ;
wire \data_count_sig[3]~15_combout ;
wire \data_count_sig[4]~22 ;
wire \data_count_sig[4]~21_combout ;
wire \data_count_sig[5]~24 ;
wire \data_count_sig[5]~23_combout ;
wire \data_count_sig[6]~26 ;
wire \data_count_sig[6]~25_combout ;
wire \data_count_sig[7]~28 ;
wire \data_count_sig[7]~27_combout ;
wire \data_count_sig[8]~29_combout ;
wire \fft_dirn_stream~q ;
wire \fft_s2_cur.WAIT_FOR_LPP_INPUT~q ;
wire \fft_dirn_held_o2~q ;
wire \fft_s2_cur.LPP_C_OUTPUT~q ;
wire \lpp_count_offset[0]~q ;
wire \lpp_count_offset[1]~q ;
wire \lpp_count_offset[2]~q ;
wire \lpp_count_offset[3]~q ;
wire \lpp_count_offset[4]~q ;
wire \lpp_count_offset[5]~q ;
wire \lpp_count_offset[6]~q ;
wire \lpp_count_offset[7]~q ;
wire \lpp_count_offset[8]~q ;
wire \fft_dirn_held_o~q ;
wire \gen_gt256_mk:ctrl|blk_done_int~q ;
wire \lpp_count[0]~q ;
wire \lpp_count_offset[0]~10 ;
wire \lpp_count_offset[0]~9_combout ;
wire \lpp_count[1]~q ;
wire \lpp_count_offset[1]~14 ;
wire \lpp_count_offset[1]~13_combout ;
wire \lpp_count[2]~q ;
wire \lpp_count_offset[2]~16 ;
wire \lpp_count_offset[2]~15_combout ;
wire \lpp_count[3]~q ;
wire \lpp_count_offset[3]~18 ;
wire \lpp_count_offset[3]~17_combout ;
wire \lpp_count[4]~q ;
wire \lpp_count_offset[4]~20 ;
wire \lpp_count_offset[4]~19_combout ;
wire \lpp_count[5]~q ;
wire \lpp_count_offset[5]~22 ;
wire \lpp_count_offset[5]~21_combout ;
wire \lpp_count[6]~q ;
wire \lpp_count_offset[6]~24 ;
wire \lpp_count_offset[6]~23_combout ;
wire \lpp_count[7]~q ;
wire \lpp_count_offset[7]~26 ;
wire \lpp_count_offset[7]~25_combout ;
wire \lpp_count[8]~q ;
wire \lpp_count_offset[8]~27_combout ;
wire \lpp_ram_data_out_sw[1][1]~q ;
wire \lpp_ram_data_out_sw[0][1]~q ;
wire \lpp_ram_data_out_sw[1][0]~q ;
wire \lpp_ram_data_out_sw[0][0]~q ;
wire \lpp_ram_data_out_sw[1][7]~q ;
wire \lpp_ram_data_out_sw[0][7]~q ;
wire \lpp_ram_data_out_sw[1][6]~q ;
wire \lpp_ram_data_out_sw[0][6]~q ;
wire \lpp_ram_data_out_sw[1][5]~q ;
wire \lpp_ram_data_out_sw[0][5]~q ;
wire \lpp_ram_data_out_sw[1][4]~q ;
wire \lpp_ram_data_out_sw[0][4]~q ;
wire \lpp_ram_data_out_sw[1][3]~q ;
wire \lpp_ram_data_out_sw[0][3]~q ;
wire \lpp_ram_data_out_sw[1][2]~q ;
wire \lpp_ram_data_out_sw[0][2]~q ;
wire \lpp_ram_data_out_sw[1][9]~q ;
wire \lpp_ram_data_out_sw[0][9]~q ;
wire \lpp_ram_data_out_sw[1][8]~q ;
wire \lpp_ram_data_out_sw[0][8]~q ;
wire \lpp_ram_data_out_sw[1][15]~q ;
wire \lpp_ram_data_out_sw[0][15]~q ;
wire \lpp_ram_data_out_sw[1][14]~q ;
wire \lpp_ram_data_out_sw[0][14]~q ;
wire \lpp_ram_data_out_sw[1][13]~q ;
wire \lpp_ram_data_out_sw[0][13]~q ;
wire \lpp_ram_data_out_sw[1][12]~q ;
wire \lpp_ram_data_out_sw[0][12]~q ;
wire \lpp_ram_data_out_sw[1][11]~q ;
wire \lpp_ram_data_out_sw[0][11]~q ;
wire \lpp_ram_data_out_sw[1][10]~q ;
wire \lpp_ram_data_out_sw[0][10]~q ;
wire \Add2~1 ;
wire \Add2~0_combout ;
wire \Add2~3 ;
wire \Add2~2_combout ;
wire \Add2~5 ;
wire \Add2~4_combout ;
wire \Add2~7 ;
wire \Add2~6_combout ;
wire \Add2~9 ;
wire \Add2~8_combout ;
wire \Add2~11 ;
wire \Add2~10_combout ;
wire \Add2~13 ;
wire \Add2~12_combout ;
wire \Add2~15 ;
wire \Add2~14_combout ;
wire \Add2~16_combout ;
wire \lpp_ram_data_out[2][1]~q ;
wire \lpp_ram_data_out[1][1]~q ;
wire \lpp_ram_data_out[0][1]~q ;
wire \lpp_ram_data_out[3][1]~q ;
wire \lpp_ram_data_out_sw[1][1]~2_combout ;
wire \lpp_ram_data_out_sw[0][1]~3_combout ;
wire \lpp_ram_data_out[2][0]~q ;
wire \lpp_ram_data_out[1][0]~q ;
wire \lpp_ram_data_out[0][0]~q ;
wire \lpp_ram_data_out[3][0]~q ;
wire \lpp_ram_data_out_sw[1][0]~30_combout ;
wire \lpp_ram_data_out_sw[0][0]~31_combout ;
wire \lpp_ram_data_out[2][7]~q ;
wire \lpp_ram_data_out[1][7]~q ;
wire \lpp_ram_data_out[0][7]~q ;
wire \lpp_ram_data_out[3][7]~q ;
wire \lpp_ram_data_out_sw[1][7]~26_combout ;
wire \lpp_ram_data_out_sw[0][7]~27_combout ;
wire \lpp_ram_data_out[2][6]~q ;
wire \lpp_ram_data_out[1][6]~q ;
wire \lpp_ram_data_out[0][6]~q ;
wire \lpp_ram_data_out[3][6]~q ;
wire \lpp_ram_data_out_sw[1][6]~22_combout ;
wire \lpp_ram_data_out_sw[0][6]~23_combout ;
wire \lpp_ram_data_out[2][5]~q ;
wire \lpp_ram_data_out[1][5]~q ;
wire \lpp_ram_data_out[0][5]~q ;
wire \lpp_ram_data_out[3][5]~q ;
wire \lpp_ram_data_out_sw[1][5]~18_combout ;
wire \lpp_ram_data_out_sw[0][5]~19_combout ;
wire \lpp_ram_data_out[2][4]~q ;
wire \lpp_ram_data_out[1][4]~q ;
wire \lpp_ram_data_out[0][4]~q ;
wire \lpp_ram_data_out[3][4]~q ;
wire \lpp_ram_data_out_sw[1][4]~14_combout ;
wire \lpp_ram_data_out_sw[0][4]~15_combout ;
wire \lpp_ram_data_out[2][3]~q ;
wire \lpp_ram_data_out[1][3]~q ;
wire \lpp_ram_data_out[0][3]~q ;
wire \lpp_ram_data_out[3][3]~q ;
wire \lpp_ram_data_out_sw[1][3]~10_combout ;
wire \lpp_ram_data_out_sw[0][3]~11_combout ;
wire \lpp_ram_data_out[2][2]~q ;
wire \lpp_ram_data_out[1][2]~q ;
wire \lpp_ram_data_out[0][2]~q ;
wire \lpp_ram_data_out[3][2]~q ;
wire \lpp_ram_data_out_sw[1][2]~6_combout ;
wire \lpp_ram_data_out_sw[0][2]~7_combout ;
wire \lpp_ram_data_out[2][9]~q ;
wire \lpp_ram_data_out[1][9]~q ;
wire \lpp_ram_data_out[0][9]~q ;
wire \lpp_ram_data_out[3][9]~q ;
wire \lpp_ram_data_out_sw[1][9]~0_combout ;
wire \lpp_ram_data_out_sw[0][9]~1_combout ;
wire \lpp_ram_data_out[2][8]~q ;
wire \lpp_ram_data_out[1][8]~q ;
wire \lpp_ram_data_out[0][8]~q ;
wire \lpp_ram_data_out[3][8]~q ;
wire \lpp_ram_data_out_sw[1][8]~28_combout ;
wire \lpp_ram_data_out_sw[0][8]~29_combout ;
wire \lpp_ram_data_out[2][15]~q ;
wire \lpp_ram_data_out[1][15]~q ;
wire \lpp_ram_data_out[0][15]~q ;
wire \lpp_ram_data_out[3][15]~q ;
wire \lpp_ram_data_out_sw[1][15]~24_combout ;
wire \lpp_ram_data_out_sw[0][15]~25_combout ;
wire \lpp_ram_data_out[2][14]~q ;
wire \lpp_ram_data_out[1][14]~q ;
wire \lpp_ram_data_out[0][14]~q ;
wire \lpp_ram_data_out[3][14]~q ;
wire \lpp_ram_data_out_sw[1][14]~20_combout ;
wire \lpp_ram_data_out_sw[0][14]~21_combout ;
wire \lpp_ram_data_out[2][13]~q ;
wire \lpp_ram_data_out[1][13]~q ;
wire \lpp_ram_data_out[0][13]~q ;
wire \lpp_ram_data_out[3][13]~q ;
wire \lpp_ram_data_out_sw[1][13]~16_combout ;
wire \lpp_ram_data_out_sw[0][13]~17_combout ;
wire \lpp_ram_data_out[2][12]~q ;
wire \lpp_ram_data_out[1][12]~q ;
wire \lpp_ram_data_out[0][12]~q ;
wire \lpp_ram_data_out[3][12]~q ;
wire \lpp_ram_data_out_sw[1][12]~12_combout ;
wire \lpp_ram_data_out_sw[0][12]~13_combout ;
wire \lpp_ram_data_out[2][11]~q ;
wire \lpp_ram_data_out[1][11]~q ;
wire \lpp_ram_data_out[0][11]~q ;
wire \lpp_ram_data_out[3][11]~q ;
wire \lpp_ram_data_out_sw[1][11]~8_combout ;
wire \lpp_ram_data_out_sw[0][11]~9_combout ;
wire \lpp_ram_data_out[2][10]~q ;
wire \lpp_ram_data_out[1][10]~q ;
wire \lpp_ram_data_out[0][10]~q ;
wire \lpp_ram_data_out[3][10]~q ;
wire \lpp_ram_data_out_sw[1][10]~4_combout ;
wire \lpp_ram_data_out_sw[0][10]~5_combout ;
wire \fft_dirn~q ;
wire \gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[1] ;
wire \gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[1] ;
wire \lpp_sel~q ;
wire \gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[1] ;
wire \gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[1] ;
wire \gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[1] ;
wire \gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[1] ;
wire \gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[1] ;
wire \gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[1] ;
wire \gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[0] ;
wire \gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[0] ;
wire \gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[0] ;
wire \gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[0] ;
wire \gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[0] ;
wire \gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[0] ;
wire \gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[0] ;
wire \gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[0] ;
wire \gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[7] ;
wire \gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[7] ;
wire \gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[7] ;
wire \gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[7] ;
wire \gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[7] ;
wire \gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[7] ;
wire \gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[7] ;
wire \gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[7] ;
wire \gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[6] ;
wire \gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[6] ;
wire \gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[6] ;
wire \gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[6] ;
wire \gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[6] ;
wire \gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[6] ;
wire \gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[6] ;
wire \gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[6] ;
wire \gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[5] ;
wire \gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[5] ;
wire \gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[5] ;
wire \gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[5] ;
wire \gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[5] ;
wire \gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[5] ;
wire \gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[5] ;
wire \gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[5] ;
wire \gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[4] ;
wire \gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[4] ;
wire \gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[4] ;
wire \gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[4] ;
wire \gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[4] ;
wire \gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[4] ;
wire \gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[4] ;
wire \gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[4] ;
wire \gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[3] ;
wire \gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[3] ;
wire \gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[3] ;
wire \gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[3] ;
wire \gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[3] ;
wire \gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[3] ;
wire \gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[3] ;
wire \gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[3] ;
wire \gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[2] ;
wire \gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[2] ;
wire \gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[2] ;
wire \gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[2] ;
wire \gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[2] ;
wire \gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[2] ;
wire \gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[2] ;
wire \gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[2] ;
wire \gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[9] ;
wire \gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[9] ;
wire \gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[9] ;
wire \gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[9] ;
wire \gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[9] ;
wire \gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[9] ;
wire \gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[9] ;
wire \gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[9] ;
wire \gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[8] ;
wire \gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[8] ;
wire \gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[8] ;
wire \gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[8] ;
wire \gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[8] ;
wire \gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[8] ;
wire \gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[8] ;
wire \gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[8] ;
wire \gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[15] ;
wire \gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[15] ;
wire \gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[15] ;
wire \gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[15] ;
wire \gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[15] ;
wire \gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[15] ;
wire \gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[15] ;
wire \gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[15] ;
wire \gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[14] ;
wire \gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[14] ;
wire \gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[14] ;
wire \gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[14] ;
wire \gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[14] ;
wire \gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[14] ;
wire \gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[14] ;
wire \gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[14] ;
wire \gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[13] ;
wire \gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[13] ;
wire \gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[13] ;
wire \gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[13] ;
wire \gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[13] ;
wire \gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[13] ;
wire \gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[13] ;
wire \gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[13] ;
wire \gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[12] ;
wire \gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[12] ;
wire \gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[12] ;
wire \gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[12] ;
wire \gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[12] ;
wire \gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[12] ;
wire \gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[12] ;
wire \gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[12] ;
wire \gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[11] ;
wire \gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[11] ;
wire \gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[11] ;
wire \gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[11] ;
wire \gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[11] ;
wire \gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[11] ;
wire \gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[11] ;
wire \gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[11] ;
wire \gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[10] ;
wire \gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[10] ;
wire \gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[10] ;
wire \gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[10] ;
wire \gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[10] ;
wire \gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[10] ;
wire \gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[10] ;
wire \gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[10] ;
wire \ram_cxb_wr_data|ram_in_reg[6][1]~q ;
wire \ram_cxb_wr_data|ram_in_reg[5][1]~q ;
wire \ram_cxb_wr_data|ram_in_reg[4][1]~q ;
wire \ram_cxb_wr_data|ram_in_reg[7][1]~q ;
wire \ram_cxb_wr_data|ram_in_reg[6][0]~q ;
wire \ram_cxb_wr_data|ram_in_reg[5][0]~q ;
wire \ram_cxb_wr_data|ram_in_reg[4][0]~q ;
wire \ram_cxb_wr_data|ram_in_reg[7][0]~q ;
wire \ram_cxb_wr_data|ram_in_reg[6][7]~q ;
wire \ram_cxb_wr_data|ram_in_reg[5][7]~q ;
wire \ram_cxb_wr_data|ram_in_reg[4][7]~q ;
wire \ram_cxb_wr_data|ram_in_reg[7][7]~q ;
wire \ram_cxb_wr_data|ram_in_reg[6][6]~q ;
wire \ram_cxb_wr_data|ram_in_reg[5][6]~q ;
wire \ram_cxb_wr_data|ram_in_reg[4][6]~q ;
wire \ram_cxb_wr_data|ram_in_reg[7][6]~q ;
wire \ram_cxb_wr_data|ram_in_reg[6][5]~q ;
wire \ram_cxb_wr_data|ram_in_reg[5][5]~q ;
wire \ram_cxb_wr_data|ram_in_reg[4][5]~q ;
wire \ram_cxb_wr_data|ram_in_reg[7][5]~q ;
wire \ram_cxb_wr_data|ram_in_reg[6][4]~q ;
wire \ram_cxb_wr_data|ram_in_reg[5][4]~q ;
wire \ram_cxb_wr_data|ram_in_reg[4][4]~q ;
wire \ram_cxb_wr_data|ram_in_reg[7][4]~q ;
wire \ram_cxb_wr_data|ram_in_reg[6][3]~q ;
wire \ram_cxb_wr_data|ram_in_reg[5][3]~q ;
wire \ram_cxb_wr_data|ram_in_reg[4][3]~q ;
wire \ram_cxb_wr_data|ram_in_reg[7][3]~q ;
wire \ram_cxb_wr_data|ram_in_reg[6][2]~q ;
wire \ram_cxb_wr_data|ram_in_reg[5][2]~q ;
wire \ram_cxb_wr_data|ram_in_reg[4][2]~q ;
wire \ram_cxb_wr_data|ram_in_reg[7][2]~q ;
wire \ram_cxb_wr_data|ram_in_reg[2][1]~q ;
wire \ram_cxb_wr_data|ram_in_reg[1][1]~q ;
wire \ram_cxb_wr_data|ram_in_reg[0][1]~q ;
wire \ram_cxb_wr_data|ram_in_reg[3][1]~q ;
wire \ram_cxb_wr_data|ram_in_reg[2][0]~q ;
wire \ram_cxb_wr_data|ram_in_reg[1][0]~q ;
wire \ram_cxb_wr_data|ram_in_reg[0][0]~q ;
wire \ram_cxb_wr_data|ram_in_reg[3][0]~q ;
wire \ram_cxb_wr_data|ram_in_reg[2][7]~q ;
wire \ram_cxb_wr_data|ram_in_reg[1][7]~q ;
wire \ram_cxb_wr_data|ram_in_reg[0][7]~q ;
wire \ram_cxb_wr_data|ram_in_reg[3][7]~q ;
wire \ram_cxb_wr_data|ram_in_reg[2][6]~q ;
wire \ram_cxb_wr_data|ram_in_reg[1][6]~q ;
wire \ram_cxb_wr_data|ram_in_reg[0][6]~q ;
wire \ram_cxb_wr_data|ram_in_reg[3][6]~q ;
wire \ram_cxb_wr_data|ram_in_reg[2][5]~q ;
wire \ram_cxb_wr_data|ram_in_reg[1][5]~q ;
wire \ram_cxb_wr_data|ram_in_reg[0][5]~q ;
wire \ram_cxb_wr_data|ram_in_reg[3][5]~q ;
wire \ram_cxb_wr_data|ram_in_reg[2][4]~q ;
wire \ram_cxb_wr_data|ram_in_reg[1][4]~q ;
wire \ram_cxb_wr_data|ram_in_reg[0][4]~q ;
wire \ram_cxb_wr_data|ram_in_reg[3][4]~q ;
wire \ram_cxb_wr_data|ram_in_reg[2][3]~q ;
wire \ram_cxb_wr_data|ram_in_reg[1][3]~q ;
wire \ram_cxb_wr_data|ram_in_reg[0][3]~q ;
wire \ram_cxb_wr_data|ram_in_reg[3][3]~q ;
wire \ram_cxb_wr_data|ram_in_reg[2][2]~q ;
wire \ram_cxb_wr_data|ram_in_reg[1][2]~q ;
wire \ram_cxb_wr_data|ram_in_reg[0][2]~q ;
wire \ram_cxb_wr_data|ram_in_reg[3][2]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[0][3]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[0][3]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[1][3]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[1][3]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[2][3]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[2][3]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[3][3]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[3][3]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[0][4]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[0][4]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[1][4]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[1][4]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[2][4]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[2][4]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[3][4]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[3][4]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[0][5]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[0][5]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[1][5]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[1][5]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[2][5]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[2][5]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[3][5]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[3][5]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[2][2]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[1][2]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[0][2]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[3][2]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[2][2]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[1][2]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[0][2]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[3][2]~q ;
wire \gen_radix_2_last_pass:gen_lpp_addr|sw[0]~q ;
wire \writer|data_rdy_int~q ;
wire \twrom|gen_M4K:cos_1n|gen_auto:altsyncram_component|auto_generated|q_a[0] ;
wire \twrom|gen_M4K:cos_1n|gen_auto:altsyncram_component|auto_generated|q_a[1] ;
wire \twrom|gen_M4K:cos_1n|gen_auto:altsyncram_component|auto_generated|q_a[2] ;
wire \twrom|gen_M4K:cos_1n|gen_auto:altsyncram_component|auto_generated|q_a[3] ;
wire \twrom|gen_M4K:cos_1n|gen_auto:altsyncram_component|auto_generated|q_a[4] ;
wire \twrom|gen_M4K:cos_1n|gen_auto:altsyncram_component|auto_generated|q_a[5] ;
wire \twrom|gen_M4K:cos_1n|gen_auto:altsyncram_component|auto_generated|q_a[6] ;
wire \twrom|gen_M4K:cos_1n|gen_auto:altsyncram_component|auto_generated|q_a[7] ;
wire \twrom|gen_M4K:sin_1n|gen_auto:altsyncram_component|auto_generated|q_a[0] ;
wire \twrom|gen_M4K:sin_1n|gen_auto:altsyncram_component|auto_generated|q_a[1] ;
wire \twrom|gen_M4K:sin_1n|gen_auto:altsyncram_component|auto_generated|q_a[2] ;
wire \twrom|gen_M4K:sin_1n|gen_auto:altsyncram_component|auto_generated|q_a[3] ;
wire \twrom|gen_M4K:sin_1n|gen_auto:altsyncram_component|auto_generated|q_a[4] ;
wire \twrom|gen_M4K:sin_1n|gen_auto:altsyncram_component|auto_generated|q_a[5] ;
wire \twrom|gen_M4K:sin_1n|gen_auto:altsyncram_component|auto_generated|q_a[6] ;
wire \twrom|gen_M4K:sin_1n|gen_auto:altsyncram_component|auto_generated|q_a[7] ;
wire \twrom|gen_M4K:cos_2n|gen_auto:altsyncram_component|auto_generated|q_a[0] ;
wire \twrom|gen_M4K:cos_2n|gen_auto:altsyncram_component|auto_generated|q_a[1] ;
wire \twrom|gen_M4K:cos_2n|gen_auto:altsyncram_component|auto_generated|q_a[2] ;
wire \twrom|gen_M4K:cos_2n|gen_auto:altsyncram_component|auto_generated|q_a[3] ;
wire \twrom|gen_M4K:cos_2n|gen_auto:altsyncram_component|auto_generated|q_a[4] ;
wire \twrom|gen_M4K:cos_2n|gen_auto:altsyncram_component|auto_generated|q_a[5] ;
wire \twrom|gen_M4K:cos_2n|gen_auto:altsyncram_component|auto_generated|q_a[6] ;
wire \twrom|gen_M4K:cos_2n|gen_auto:altsyncram_component|auto_generated|q_a[7] ;
wire \twrom|gen_M4K:sin_2n|gen_auto:altsyncram_component|auto_generated|q_a[0] ;
wire \twrom|gen_M4K:sin_2n|gen_auto:altsyncram_component|auto_generated|q_a[1] ;
wire \twrom|gen_M4K:sin_2n|gen_auto:altsyncram_component|auto_generated|q_a[2] ;
wire \twrom|gen_M4K:sin_2n|gen_auto:altsyncram_component|auto_generated|q_a[3] ;
wire \twrom|gen_M4K:sin_2n|gen_auto:altsyncram_component|auto_generated|q_a[4] ;
wire \twrom|gen_M4K:sin_2n|gen_auto:altsyncram_component|auto_generated|q_a[5] ;
wire \twrom|gen_M4K:sin_2n|gen_auto:altsyncram_component|auto_generated|q_a[6] ;
wire \twrom|gen_M4K:sin_2n|gen_auto:altsyncram_component|auto_generated|q_a[7] ;
wire \twrom|gen_M4K:cos_3n|gen_auto:altsyncram_component|auto_generated|q_a[0] ;
wire \twrom|gen_M4K:cos_3n|gen_auto:altsyncram_component|auto_generated|q_a[1] ;
wire \twrom|gen_M4K:cos_3n|gen_auto:altsyncram_component|auto_generated|q_a[2] ;
wire \twrom|gen_M4K:cos_3n|gen_auto:altsyncram_component|auto_generated|q_a[3] ;
wire \twrom|gen_M4K:cos_3n|gen_auto:altsyncram_component|auto_generated|q_a[4] ;
wire \twrom|gen_M4K:cos_3n|gen_auto:altsyncram_component|auto_generated|q_a[5] ;
wire \twrom|gen_M4K:cos_3n|gen_auto:altsyncram_component|auto_generated|q_a[6] ;
wire \twrom|gen_M4K:cos_3n|gen_auto:altsyncram_component|auto_generated|q_a[7] ;
wire \twrom|gen_M4K:sin_3n|gen_auto:altsyncram_component|auto_generated|q_a[0] ;
wire \twrom|gen_M4K:sin_3n|gen_auto:altsyncram_component|auto_generated|q_a[1] ;
wire \twrom|gen_M4K:sin_3n|gen_auto:altsyncram_component|auto_generated|q_a[2] ;
wire \twrom|gen_M4K:sin_3n|gen_auto:altsyncram_component|auto_generated|q_a[3] ;
wire \twrom|gen_M4K:sin_3n|gen_auto:altsyncram_component|auto_generated|q_a[4] ;
wire \twrom|gen_M4K:sin_3n|gen_auto:altsyncram_component|auto_generated|q_a[5] ;
wire \twrom|gen_M4K:sin_3n|gen_auto:altsyncram_component|auto_generated|q_a[6] ;
wire \twrom|gen_M4K:sin_3n|gen_auto:altsyncram_component|auto_generated|q_a[7] ;
wire \ram_cxb_bfp_data|ram_in_reg[0][2]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[0][6]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[0][4]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[0][3]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[0][5]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[2][2]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[2][6]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[2][4]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[2][3]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[2][5]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[0][1]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[2][1]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[0][0]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[2][0]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[1][2]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[1][6]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[1][4]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[1][3]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[1][5]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[3][2]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[3][6]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[3][4]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[3][3]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[3][5]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[1][1]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[3][1]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[1][0]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[3][0]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[0][7]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[2][7]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[1][7]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[3][7]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[4][7]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[4][3]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[4][5]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[4][4]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[4][6]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[6][7]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[6][3]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[6][5]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[6][4]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[6][6]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[4][2]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[6][2]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[4][1]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[6][1]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[4][0]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[6][0]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[5][7]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[5][3]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[5][5]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[5][4]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[5][6]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[7][3]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[7][7]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[7][5]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[7][4]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[7][6]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[5][2]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[7][2]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[5][1]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[7][1]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[5][0]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[7][0]~q ;
wire \dat_B|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[10] ;
wire \dat_A|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[10] ;
wire \dat_B|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[10] ;
wire \dat_A|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[10] ;
wire \dat_B|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[10] ;
wire \dat_A|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[10] ;
wire \dat_B|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[10] ;
wire \dat_A|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[10] ;
wire \dat_B|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[14] ;
wire \dat_A|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[14] ;
wire \dat_B|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[14] ;
wire \dat_A|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[14] ;
wire \dat_B|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[14] ;
wire \dat_A|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[14] ;
wire \dat_B|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[14] ;
wire \dat_A|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[14] ;
wire \dat_B|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[12] ;
wire \dat_A|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[12] ;
wire \dat_B|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[12] ;
wire \dat_A|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[12] ;
wire \dat_B|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[12] ;
wire \dat_A|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[12] ;
wire \dat_B|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[12] ;
wire \dat_A|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[12] ;
wire \dat_B|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[11] ;
wire \dat_A|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[11] ;
wire \dat_B|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[11] ;
wire \dat_A|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[11] ;
wire \dat_B|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[11] ;
wire \dat_A|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[11] ;
wire \dat_B|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[11] ;
wire \dat_A|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[11] ;
wire \dat_B|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[13] ;
wire \dat_A|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[13] ;
wire \dat_B|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[13] ;
wire \dat_A|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[13] ;
wire \dat_B|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[13] ;
wire \dat_A|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[13] ;
wire \dat_B|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[13] ;
wire \dat_A|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[13] ;
wire \dat_B|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[9] ;
wire \dat_A|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[9] ;
wire \dat_B|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[9] ;
wire \dat_A|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[9] ;
wire \dat_B|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[9] ;
wire \dat_A|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[9] ;
wire \dat_B|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[9] ;
wire \dat_A|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[9] ;
wire \dat_B|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[8] ;
wire \dat_A|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[8] ;
wire \dat_B|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[8] ;
wire \dat_A|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[8] ;
wire \dat_B|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[8] ;
wire \dat_A|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[8] ;
wire \dat_B|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[8] ;
wire \dat_A|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[8] ;
wire \dat_B|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[15] ;
wire \dat_A|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[15] ;
wire \dat_B|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[15] ;
wire \dat_A|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[15] ;
wire \dat_B|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[15] ;
wire \dat_A|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[15] ;
wire \dat_B|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[15] ;
wire \dat_A|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[15] ;
wire \dat_B|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[7] ;
wire \dat_A|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[7] ;
wire \dat_B|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[7] ;
wire \dat_A|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[7] ;
wire \dat_B|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[7] ;
wire \dat_A|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[7] ;
wire \dat_B|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[7] ;
wire \dat_A|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[7] ;
wire \dat_B|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[3] ;
wire \dat_A|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[3] ;
wire \dat_B|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[3] ;
wire \dat_A|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[3] ;
wire \dat_B|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[3] ;
wire \dat_A|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[3] ;
wire \dat_B|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[3] ;
wire \dat_A|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[3] ;
wire \dat_B|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[5] ;
wire \dat_A|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[5] ;
wire \dat_B|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[5] ;
wire \dat_A|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[5] ;
wire \dat_B|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[5] ;
wire \dat_A|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[5] ;
wire \dat_B|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[5] ;
wire \dat_A|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[5] ;
wire \dat_B|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[4] ;
wire \dat_A|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[4] ;
wire \dat_B|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[4] ;
wire \dat_A|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[4] ;
wire \dat_B|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[4] ;
wire \dat_A|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[4] ;
wire \dat_B|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[4] ;
wire \dat_A|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[4] ;
wire \dat_B|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[6] ;
wire \dat_A|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[6] ;
wire \dat_B|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[6] ;
wire \dat_A|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[6] ;
wire \dat_B|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[6] ;
wire \dat_A|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[6] ;
wire \dat_B|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[6] ;
wire \dat_A|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[6] ;
wire \dat_B|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[2] ;
wire \dat_A|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[2] ;
wire \dat_B|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[2] ;
wire \dat_A|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[2] ;
wire \dat_B|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[2] ;
wire \dat_A|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[2] ;
wire \dat_B|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[2] ;
wire \dat_A|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[2] ;
wire \dat_B|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[1] ;
wire \dat_A|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[1] ;
wire \dat_B|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[1] ;
wire \dat_A|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[1] ;
wire \dat_B|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[1] ;
wire \dat_A|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[1] ;
wire \dat_B|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[1] ;
wire \dat_A|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[1] ;
wire \dat_B|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[0] ;
wire \dat_A|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[0] ;
wire \dat_B|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[0] ;
wire \dat_A|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[0] ;
wire \dat_B|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[0] ;
wire \dat_A|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[0] ;
wire \dat_B|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[0] ;
wire \dat_A|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[0] ;
wire \wren_b[0]~q ;
wire \wren_a[0]~q ;
wire \wren_b[1]~q ;
wire \wren_a[1]~q ;
wire \wren_b[2]~q ;
wire \wren_a[2]~q ;
wire \wren_b[3]~q ;
wire \wren_a[3]~q ;
wire \writer|wren[0]~q ;
wire \writer|wren[1]~q ;
wire \writer|wren[2]~q ;
wire \writer|wren[3]~q ;
wire \core_real_in[2]~q ;
wire \core_real_in[6]~q ;
wire \core_real_in[4]~q ;
wire \core_real_in[3]~q ;
wire \core_real_in[5]~q ;
wire \core_real_in[1]~q ;
wire \core_real_in[0]~q ;
wire \core_real_in[7]~q ;
wire \core_imag_in[7]~q ;
wire \core_imag_in[3]~q ;
wire \core_imag_in[5]~q ;
wire \core_imag_in[4]~q ;
wire \core_imag_in[6]~q ;
wire \core_imag_in[2]~q ;
wire \core_imag_in[1]~q ;
wire \core_imag_in[0]~q ;
wire \writer|anb~q ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[2] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[10] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[14] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[4] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[12] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[3] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[11] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[13] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[1] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[9] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[0] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[8] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[15] ;
wire \auk_dsp_interface_controller_1|source_packet_error[0]~q ;
wire \auk_dsp_interface_controller_1|source_packet_error[1]~q ;
wire \auk_dsp_atlantic_source_1|valid_ctrl_int~q ;
wire \master_sink_ena~q ;
wire \auk_dsp_interface_controller_1|source_stall_reg~q ;
wire \auk_dsp_interface_controller_1|sink_stall_reg~q ;
wire \auk_dsp_interface_controller_1|sink_ready_ctrl~0_combout ;
wire \auk_dsp_atlantic_sink_1|sink_stall~combout ;
wire \auk_dsp_atlantic_sink_1|packet_error_s[0]~q ;
wire \auk_dsp_atlantic_sink_1|packet_error_s[1]~q ;
wire \master_source_ena~q ;
wire \sink_ready_ctrl_d~q ;
wire \auk_dsp_atlantic_sink_1|send_sop_s~q ;
wire \sop~q ;
wire \source_valid_ctrl_sop~0_combout ;
wire \auk_dsp_atlantic_source_1|Mux3~0_combout ;
wire \source_valid_ctrl_sop~1_combout ;
wire \auk_dsp_interface_controller_1|stall_reg~q ;
wire \auk_dsp_atlantic_source_1|source_stall_int_d~q ;
wire \exponent_out[0]~q ;
wire \exponent_out[1]~q ;
wire \exponent_out[2]~q ;
wire \exponent_out[3]~q ;
wire \exponent_out[4]~q ;
wire \exponent_out[5]~q ;
wire \fft_real_out[0]~q ;
wire \fft_real_out[1]~q ;
wire \fft_real_out[2]~q ;
wire \fft_real_out[3]~q ;
wire \fft_real_out[4]~q ;
wire \fft_real_out[5]~q ;
wire \fft_real_out[6]~q ;
wire \fft_real_out[7]~q ;
wire \fft_imag_out[0]~q ;
wire \fft_imag_out[1]~q ;
wire \fft_imag_out[2]~q ;
wire \fft_imag_out[3]~q ;
wire \fft_imag_out[4]~q ;
wire \fft_imag_out[5]~q ;
wire \fft_imag_out[6]~q ;
wire \fft_imag_out[7]~q ;
wire \global_clock_enable~0_combout ;
wire \auk_dsp_atlantic_source_1|Mux0~0_combout ;
wire \auk_dsp_atlantic_source_1|Mux0~2_combout ;
wire \oe~q ;
wire \master_source_ena~0_combout ;
wire \auk_dsp_atlantic_sink_1|send_eop_s~q ;
wire \sop~0_combout ;
wire \Equal0~0_combout ;
wire \Equal0~1_combout ;
wire \LessThan0~0_combout ;
wire \LessThan0~1_combout ;
wire \master_source_sop~q ;
wire \data_count_sig[0]~17_combout ;
wire \data_count_sig[0]~18_combout ;
wire \data_count_sig[0]~19_combout ;
wire \data_count_sig[0]~20_combout ;
wire \blk_exp_accum[0]~q ;
wire \exponent_out~0_combout ;
wire \blk_exp_accum[1]~q ;
wire \exponent_out~1_combout ;
wire \blk_exp_accum[2]~q ;
wire \exponent_out~2_combout ;
wire \blk_exp_accum[3]~q ;
wire \exponent_out~3_combout ;
wire \blk_exp_accum[4]~q ;
wire \exponent_out~4_combout ;
wire \blk_exp_accum[5]~q ;
wire \exponent_out~5_combout ;
wire \gen_radix_2_last_pass:lpp_r2|data_imag_o[0]~q ;
wire \gen_radix_2_last_pass:lpp_r2|data_real_o[0]~q ;
wire \fft_real_out~0_combout ;
wire \gen_radix_2_last_pass:lpp_r2|data_imag_o[1]~q ;
wire \gen_radix_2_last_pass:lpp_r2|data_real_o[1]~q ;
wire \fft_real_out~1_combout ;
wire \gen_radix_2_last_pass:lpp_r2|data_imag_o[2]~q ;
wire \gen_radix_2_last_pass:lpp_r2|data_real_o[2]~q ;
wire \fft_real_out~2_combout ;
wire \gen_radix_2_last_pass:lpp_r2|data_imag_o[3]~q ;
wire \gen_radix_2_last_pass:lpp_r2|data_real_o[3]~q ;
wire \fft_real_out~3_combout ;
wire \gen_radix_2_last_pass:lpp_r2|data_imag_o[4]~q ;
wire \gen_radix_2_last_pass:lpp_r2|data_real_o[4]~q ;
wire \fft_real_out~4_combout ;
wire \gen_radix_2_last_pass:lpp_r2|data_imag_o[5]~q ;
wire \gen_radix_2_last_pass:lpp_r2|data_real_o[5]~q ;
wire \fft_real_out~5_combout ;
wire \gen_radix_2_last_pass:lpp_r2|data_imag_o[6]~q ;
wire \gen_radix_2_last_pass:lpp_r2|data_real_o[6]~q ;
wire \fft_real_out~6_combout ;
wire \gen_radix_2_last_pass:lpp_r2|data_imag_o[7]~q ;
wire \gen_radix_2_last_pass:lpp_r2|data_real_o[7]~q ;
wire \fft_real_out~7_combout ;
wire \fft_imag_out~0_combout ;
wire \fft_imag_out~1_combout ;
wire \fft_imag_out~2_combout ;
wire \fft_imag_out~3_combout ;
wire \fft_imag_out~4_combout ;
wire \fft_imag_out~5_combout ;
wire \fft_imag_out~6_combout ;
wire \fft_imag_out~7_combout ;
wire \fft_s2_cur.IDLE~q ;
wire \val_out~1_combout ;
wire \sop_out~q ;
wire \master_source_sop~0_combout ;
wire \gen_dft_2:bfpc|blk_exp[0]~q ;
wire \fft_s2_cur.FIRST_LPP_C~q ;
wire \Selector5~0_combout ;
wire \gen_dft_2:bfpc|blk_exp[1]~q ;
wire \Selector4~0_combout ;
wire \gen_dft_2:bfpc|blk_exp[2]~q ;
wire \Selector3~0_combout ;
wire \gen_dft_2:bfpc|blk_exp[3]~q ;
wire \Selector2~0_combout ;
wire \gen_dft_2:bfpc|blk_exp[4]~q ;
wire \Selector1~0_combout ;
wire \gen_dft_2:bfpc|blk_exp[5]~q ;
wire \Selector0~0_combout ;
wire \fft_dirn_stream~0_combout ;
wire \fft_s2_cur.LAST_LPP_C~q ;
wire \delay_lpp_en|tdl_arr[3]~q ;
wire \Selector20~0_combout ;
wire \Equal4~0_combout ;
wire \Equal4~1_combout ;
wire \Equal4~2_combout ;
wire \fft_s2_cur.IDLE~0_combout ;
wire \sop_out~0_combout ;
wire \gen_radix_2_last_pass:gen_lpp_addr|delay_en|tdl_arr[4]~q ;
wire \fft_s2_cur~9_combout ;
wire \fft_dirn_held_o2~0_combout ;
wire \fft_s2_cur.IDLE~1_combout ;
wire \Selector22~0_combout ;
wire \lpp_count_offset[0]~11_combout ;
wire \lpp_count_offset[0]~12_combout ;
wire \gen_dft_2:bfpc|slb_last[0]~q ;
wire \gen_dft_2:bfpc|slb_last[1]~q ;
wire \gen_dft_2:bfpc|slb_last[2]~q ;
wire \fft_dirn_held~q ;
wire \writer|next_block~q ;
wire \fft_dirn_held_o~0_combout ;
wire \gen_gt256_mk:ctrl|p[2]~q ;
wire \gen_gt256_mk:ctrl|p[0]~q ;
wire \gen_gt256_mk:ctrl|p[1]~q ;
wire \Selector14~0_combout ;
wire \lpp_count~0_combout ;
wire \Selector13~0_combout ;
wire \Selector12~0_combout ;
wire \Selector11~0_combout ;
wire \Selector10~0_combout ;
wire \Selector9~0_combout ;
wire \Selector8~0_combout ;
wire \Selector7~0_combout ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_detect|slb_i[0]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_detect|slb_i[1]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_detect|slb_i[2]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_detect|slb_i[3]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_detect|Mux2~0_combout ;
wire \gen_dft_2:delay_blk_done|tdl_arr[11]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_detect|Mux1~0_combout ;
wire \gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ;
wire \Mux30~0_combout ;
wire \Mux30~1_combout ;
wire \gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ;
wire \Mux30~2_combout ;
wire \Mux30~3_combout ;
wire \gen_radix_2_last_pass:delay_mid|tdl_arr[4]~q ;
wire \Mux31~0_combout ;
wire \Mux31~1_combout ;
wire \Mux31~2_combout ;
wire \Mux31~3_combout ;
wire \Mux24~0_combout ;
wire \Mux24~1_combout ;
wire \Mux24~2_combout ;
wire \Mux24~3_combout ;
wire \Mux25~0_combout ;
wire \Mux25~1_combout ;
wire \Mux25~2_combout ;
wire \Mux25~3_combout ;
wire \Mux26~0_combout ;
wire \Mux26~1_combout ;
wire \Mux26~2_combout ;
wire \Mux26~3_combout ;
wire \Mux27~0_combout ;
wire \Mux27~1_combout ;
wire \Mux27~2_combout ;
wire \Mux27~3_combout ;
wire \Mux28~0_combout ;
wire \Mux28~1_combout ;
wire \Mux28~2_combout ;
wire \Mux28~3_combout ;
wire \Mux29~0_combout ;
wire \Mux29~1_combout ;
wire \Mux29~2_combout ;
wire \Mux29~3_combout ;
wire \Mux22~0_combout ;
wire \Mux22~1_combout ;
wire \Mux22~2_combout ;
wire \Mux22~3_combout ;
wire \Mux23~0_combout ;
wire \Mux23~1_combout ;
wire \Mux23~2_combout ;
wire \Mux23~3_combout ;
wire \Mux16~0_combout ;
wire \Mux16~1_combout ;
wire \Mux16~2_combout ;
wire \Mux16~3_combout ;
wire \Mux17~0_combout ;
wire \Mux17~1_combout ;
wire \Mux17~2_combout ;
wire \Mux17~3_combout ;
wire \Mux18~0_combout ;
wire \Mux18~1_combout ;
wire \Mux18~2_combout ;
wire \Mux18~3_combout ;
wire \Mux19~0_combout ;
wire \Mux19~1_combout ;
wire \Mux19~2_combout ;
wire \Mux19~3_combout ;
wire \Mux20~0_combout ;
wire \Mux20~1_combout ;
wire \Mux20~2_combout ;
wire \Mux20~3_combout ;
wire \Mux21~0_combout ;
wire \Mux21~1_combout ;
wire \Mux21~2_combout ;
wire \Mux21~3_combout ;
wire \fft_dirn_held~0_combout ;
wire \gen_dft_2:bfpdft|gen_cont:delay_next_blk|tdl_arr[4]~q ;
wire \data_rdy_vec[4]~q ;
wire \gen_gt256_mk:ctrl|next_pass_i~q ;
wire \gen_gt256_mk:ctrl|Equal0~0_combout ;
wire \lpp_ram_data_out~0_combout ;
wire \lpp_ram_data_out~1_combout ;
wire \lpp_ram_data_out~2_combout ;
wire \lpp_ram_data_out~3_combout ;
wire \lpp_ram_data_out~4_combout ;
wire \lpp_ram_data_out~5_combout ;
wire \lpp_ram_data_out~6_combout ;
wire \lpp_ram_data_out~7_combout ;
wire \lpp_ram_data_out~8_combout ;
wire \lpp_ram_data_out~9_combout ;
wire \lpp_ram_data_out~10_combout ;
wire \lpp_ram_data_out~11_combout ;
wire \lpp_ram_data_out~12_combout ;
wire \lpp_ram_data_out~13_combout ;
wire \lpp_ram_data_out~14_combout ;
wire \lpp_ram_data_out~15_combout ;
wire \lpp_ram_data_out~16_combout ;
wire \lpp_ram_data_out~17_combout ;
wire \lpp_ram_data_out~18_combout ;
wire \lpp_ram_data_out~19_combout ;
wire \lpp_ram_data_out~20_combout ;
wire \lpp_ram_data_out~21_combout ;
wire \lpp_ram_data_out~22_combout ;
wire \lpp_ram_data_out~23_combout ;
wire \lpp_ram_data_out~24_combout ;
wire \lpp_ram_data_out~25_combout ;
wire \lpp_ram_data_out~26_combout ;
wire \lpp_ram_data_out~27_combout ;
wire \lpp_ram_data_out~28_combout ;
wire \lpp_ram_data_out~29_combout ;
wire \lpp_ram_data_out~30_combout ;
wire \lpp_ram_data_out~31_combout ;
wire \lpp_ram_data_out~32_combout ;
wire \lpp_ram_data_out~33_combout ;
wire \lpp_ram_data_out~34_combout ;
wire \lpp_ram_data_out~35_combout ;
wire \lpp_ram_data_out~36_combout ;
wire \lpp_ram_data_out~37_combout ;
wire \lpp_ram_data_out~38_combout ;
wire \lpp_ram_data_out~39_combout ;
wire \lpp_ram_data_out~40_combout ;
wire \lpp_ram_data_out~41_combout ;
wire \lpp_ram_data_out~42_combout ;
wire \lpp_ram_data_out~43_combout ;
wire \lpp_ram_data_out~44_combout ;
wire \lpp_ram_data_out~45_combout ;
wire \lpp_ram_data_out~46_combout ;
wire \lpp_ram_data_out~47_combout ;
wire \lpp_ram_data_out~48_combout ;
wire \lpp_ram_data_out~49_combout ;
wire \lpp_ram_data_out~50_combout ;
wire \lpp_ram_data_out~51_combout ;
wire \lpp_ram_data_out~52_combout ;
wire \lpp_ram_data_out~53_combout ;
wire \lpp_ram_data_out~54_combout ;
wire \lpp_ram_data_out~55_combout ;
wire \lpp_ram_data_out~56_combout ;
wire \lpp_ram_data_out~57_combout ;
wire \lpp_ram_data_out~58_combout ;
wire \lpp_ram_data_out~59_combout ;
wire \lpp_ram_data_out~60_combout ;
wire \lpp_ram_data_out~61_combout ;
wire \lpp_ram_data_out~62_combout ;
wire \lpp_ram_data_out~63_combout ;
wire \fft_dirn~0_combout ;
wire \gen_dft_2:bfpdft|gen_cont:delay_next_blk|tdl_arr[3]~q ;
wire \data_rdy_vec[3]~q ;
wire \data_rdy_vec~0_combout ;
wire \wc_vec[6]~q ;
wire \gen_wrsw_2:ram_cxb_wr|ram_in_reg[0][0]~q ;
wire \gen_wrsw_2:ram_cxb_wr|ram_in_reg[2][1]~q ;
wire \gen_wrsw_2:ram_cxb_wr|ram_in_reg[0][2]~q ;
wire \gen_wrsw_2:ram_cxb_wr|ram_in_reg[2][3]~q ;
wire \gen_wrsw_2:ram_cxb_wr|ram_in_reg[0][4]~q ;
wire \gen_wrsw_2:ram_cxb_wr|ram_in_reg[2][5]~q ;
wire \gen_wrsw_2:ram_cxb_wr|ram_in_reg[0][6]~q ;
wire \rdaddress_c_bus[0]~q ;
wire \rdaddress_c_bus[15]~q ;
wire \rdaddress_c_bus[16]~q ;
wire \rdaddress_c_bus[10]~q ;
wire \rdaddress_c_bus[11]~q ;
wire \rdaddress_c_bus[12]~q ;
wire \rdaddress_c_bus[13]~q ;
wire \wd_vec[6]~q ;
wire \lpp_sel~0_combout ;
wire \gen_wrsw_2:ram_cxb_wr|ram_in_reg[1][0]~q ;
wire \gen_wrsw_2:ram_cxb_wr|ram_in_reg[1][1]~q ;
wire \gen_wrsw_2:ram_cxb_wr|ram_in_reg[1][2]~q ;
wire \gen_wrsw_2:ram_cxb_wr|ram_in_reg[1][3]~q ;
wire \gen_wrsw_2:ram_cxb_wr|ram_in_reg[1][4]~q ;
wire \gen_wrsw_2:ram_cxb_wr|ram_in_reg[1][5]~q ;
wire \rdaddress_c_bus[20]~q ;
wire \gen_wrsw_2:ram_cxb_wr|ram_in_reg[0][1]~q ;
wire \gen_wrsw_2:ram_cxb_wr|ram_in_reg[0][3]~q ;
wire \gen_wrsw_2:ram_cxb_wr|ram_in_reg[0][5]~q ;
wire \gen_wrsw_2:ram_cxb_wr|ram_in_reg[3][1]~q ;
wire \gen_wrsw_2:ram_cxb_wr|ram_in_reg[3][3]~q ;
wire \gen_wrsw_2:ram_cxb_wr|ram_in_reg[3][5]~q ;
wire \data_rdy_vec[2]~q ;
wire \data_rdy_vec~1_combout ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[0][7]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[0][7]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[1][7]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[1][7]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[2][7]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[2][7]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[3][7]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[3][7]~q ;
wire \gen_dft_2:bfpdft|blk_done_vec[2]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[0][6]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[0][6]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[1][6]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[1][6]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[2][6]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[2][6]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[3][6]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[3][6]~q ;
wire \wc_vec[5]~q ;
wire \wc_vec~0_combout ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[2][1]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[1][1]~q ;
wire \gen_wrsw_2:get_wr_swtiches|swa_tdl[0][0]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[0][1]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[3][1]~q ;
wire \gen_wrsw_2:get_wr_swtiches|swa_tdl[0][1]~q ;
wire \gen_radix_2_last_pass:ram_cxb_rd_lpp|ram_in_reg[0][0]~q ;
wire \rdaddress_c_bus~0_combout ;
wire \gen_radix_2_last_pass:ram_cxb_rd_lpp|ram_in_reg[0][1]~q ;
wire \rdaddress_c_bus~1_combout ;
wire \gen_radix_2_last_pass:ram_cxb_rd_lpp|ram_in_reg[0][2]~q ;
wire \rdaddress_c_bus~2_combout ;
wire \gen_radix_2_last_pass:ram_cxb_rd_lpp|ram_in_reg[0][3]~q ;
wire \rdaddress_c_bus~3_combout ;
wire \gen_radix_2_last_pass:ram_cxb_rd_lpp|ram_in_reg[0][4]~q ;
wire \rdaddress_c_bus~4_combout ;
wire \gen_radix_2_last_pass:ram_cxb_rd_lpp|ram_in_reg[0][5]~q ;
wire \rdaddress_c_bus~5_combout ;
wire \gen_radix_2_last_pass:ram_cxb_rd_lpp|ram_in_reg[1][6]~q ;
wire \rdaddress_c_bus~6_combout ;
wire \wd_vec[5]~q ;
wire \wd_vec~0_combout ;
wire \rdaddress_c_bus~7_combout ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[2][0]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[1][0]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[0][0]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[3][0]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[2][1]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[1][1]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[0][1]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[3][1]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[2][0]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[1][0]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[0][0]~q ;
wire \gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[3][0]~q ;
wire \data_rdy_vec[1]~q ;
wire \data_rdy_vec~2_combout ;
wire \gen_dft_2:delay_blk_done|tdl_arr[5]~q ;
wire \gen_dft_2:delay_blk_done2|tdl_arr[19]~q ;
wire \wc_vec[4]~q ;
wire \wc_vec~1_combout ;
wire \gen_wrsw_2:wr_adgen|rd_addr_d[0]~q ;
wire \gen_wrsw_2:wr_adgen|rd_addr_c[0]~q ;
wire \gen_wrsw_2:wr_adgen|rd_addr_d[1]~q ;
wire \gen_wrsw_2:wr_adgen|rd_addr_b[1]~q ;
wire \gen_wrsw_2:wr_adgen|rd_addr_d[2]~q ;
wire \gen_wrsw_2:wr_adgen|rd_addr_c[2]~q ;
wire \gen_wrsw_2:wr_adgen|rd_addr_d[3]~q ;
wire \gen_wrsw_2:wr_adgen|rd_addr_b[3]~q ;
wire \gen_wrsw_2:wr_adgen|rd_addr_d[4]~q ;
wire \gen_wrsw_2:wr_adgen|rd_addr_c[4]~q ;
wire \gen_wrsw_2:wr_adgen|rd_addr_d[5]~q ;
wire \gen_wrsw_2:wr_adgen|rd_addr_b[5]~q ;
wire \gen_wrsw_2:wr_adgen|rd_addr_d[6]~q ;
wire \gen_radix_2_last_pass:gen_lpp_addr|rd_addr_b[0]~q ;
wire \gen_radix_2_last_pass:gen_lpp_addr|rd_addr_b[1]~q ;
wire \gen_radix_2_last_pass:gen_lpp_addr|rd_addr_b[2]~q ;
wire \gen_radix_2_last_pass:gen_lpp_addr|rd_addr_b[3]~q ;
wire \gen_radix_2_last_pass:gen_lpp_addr|rd_addr_b[4]~q ;
wire \gen_radix_2_last_pass:gen_lpp_addr|rd_addr_b[5]~q ;
wire \gen_radix_2_last_pass:gen_lpp_addr|rd_addr_b[6]~q ;
wire \wd_vec[4]~q ;
wire \wd_vec~1_combout ;
wire \data_rdy_vec[0]~q ;
wire \data_rdy_vec~3_combout ;
wire \delay_ctrl_np|tdl_arr[5]~q ;
wire \wc_vec[3]~q ;
wire \wc_vec~2_combout ;
wire \gen_wrsw_2:k_delay|tdl_arr[20][4]~q ;
wire \gen_wrsw_2:k_delay|tdl_arr[20][6]~q ;
wire \gen_wrsw_2:k_delay|tdl_arr[20][0]~q ;
wire \gen_wrsw_2:k_delay|tdl_arr[20][2]~q ;
wire \gen_wrsw_2:p_delay|tdl_arr[1][0]~q ;
wire \gen_wrsw_2:p_delay|tdl_arr[1][2]~q ;
wire \gen_wrsw_2:p_delay|tdl_arr[1][1]~q ;
wire \gen_wrsw_2:k_delay|tdl_arr[20][1]~q ;
wire \gen_wrsw_2:k_delay|tdl_arr[20][3]~q ;
wire \gen_wrsw_2:k_delay|tdl_arr[20][5]~q ;
wire \wd_vec[3]~q ;
wire \wd_vec~2_combout ;
wire \data_rdy_vec~4_combout ;
wire \wc_vec[2]~q ;
wire \wc_vec~3_combout ;
wire \wd_vec[2]~q ;
wire \wd_vec~3_combout ;
wire \wc_vec[1]~q ;
wire \wc_vec~4_combout ;
wire \p_tdl[18][0]~q ;
wire \p_tdl[18][2]~q ;
wire \p_tdl[18][1]~q ;
wire \wd_vec[1]~q ;
wire \wd_vec~4_combout ;
wire \wc_vec[0]~q ;
wire \wc_vec~5_combout ;
wire \p_tdl[17][0]~q ;
wire \p_tdl[17][2]~q ;
wire \p_tdl[17][1]~q ;
wire \wd_vec[0]~q ;
wire \wd_vec~5_combout ;
wire \twiddle_data[0][0][0]~q ;
wire \twiddle_data[0][0][1]~q ;
wire \twiddle_data[0][0][2]~q ;
wire \twiddle_data[0][0][3]~q ;
wire \twiddle_data[0][0][4]~q ;
wire \twiddle_data[0][0][5]~q ;
wire \twiddle_data[0][0][6]~q ;
wire \twiddle_data[0][0][7]~q ;
wire \twiddle_data[0][1][0]~q ;
wire \twiddle_data[0][1][1]~q ;
wire \twiddle_data[0][1][2]~q ;
wire \twiddle_data[0][1][3]~q ;
wire \twiddle_data[0][1][4]~q ;
wire \twiddle_data[0][1][5]~q ;
wire \twiddle_data[0][1][6]~q ;
wire \twiddle_data[0][1][7]~q ;
wire \twiddle_data[1][0][0]~q ;
wire \twiddle_data[1][0][1]~q ;
wire \twiddle_data[1][0][2]~q ;
wire \twiddle_data[1][0][3]~q ;
wire \twiddle_data[1][0][4]~q ;
wire \twiddle_data[1][0][5]~q ;
wire \twiddle_data[1][0][6]~q ;
wire \twiddle_data[1][0][7]~q ;
wire \twiddle_data[1][1][0]~q ;
wire \twiddle_data[1][1][1]~q ;
wire \twiddle_data[1][1][2]~q ;
wire \twiddle_data[1][1][3]~q ;
wire \twiddle_data[1][1][4]~q ;
wire \twiddle_data[1][1][5]~q ;
wire \twiddle_data[1][1][6]~q ;
wire \twiddle_data[1][1][7]~q ;
wire \twiddle_data[2][0][0]~q ;
wire \twiddle_data[2][0][1]~q ;
wire \twiddle_data[2][0][2]~q ;
wire \twiddle_data[2][0][3]~q ;
wire \twiddle_data[2][0][4]~q ;
wire \twiddle_data[2][0][5]~q ;
wire \twiddle_data[2][0][6]~q ;
wire \twiddle_data[2][0][7]~q ;
wire \twiddle_data[2][1][0]~q ;
wire \twiddle_data[2][1][1]~q ;
wire \twiddle_data[2][1][2]~q ;
wire \twiddle_data[2][1][3]~q ;
wire \twiddle_data[2][1][4]~q ;
wire \twiddle_data[2][1][5]~q ;
wire \twiddle_data[2][1][6]~q ;
wire \twiddle_data[2][1][7]~q ;
wire \sel_we|wc_i~q ;
wire \wc_vec~6_combout ;
wire \p_tdl[16][0]~q ;
wire \p_tdl[16][2]~q ;
wire \p_tdl[16][1]~q ;
wire \sel_we|wd_i~q ;
wire \wd_vec~6_combout ;
wire \twiddle_data~0_combout ;
wire \twiddle_data~1_combout ;
wire \twiddle_data~2_combout ;
wire \twiddle_data~3_combout ;
wire \twiddle_data~4_combout ;
wire \twiddle_data~5_combout ;
wire \twiddle_data~6_combout ;
wire \twiddle_data~7_combout ;
wire \twiddle_data~8_combout ;
wire \twiddle_data~9_combout ;
wire \twiddle_data~10_combout ;
wire \twiddle_data~11_combout ;
wire \twiddle_data~12_combout ;
wire \twiddle_data~13_combout ;
wire \twiddle_data~14_combout ;
wire \twiddle_data~15_combout ;
wire \twiddle_data~16_combout ;
wire \twiddle_data~17_combout ;
wire \twiddle_data~18_combout ;
wire \twiddle_data~19_combout ;
wire \twiddle_data~20_combout ;
wire \twiddle_data~21_combout ;
wire \twiddle_data~22_combout ;
wire \twiddle_data~23_combout ;
wire \twiddle_data~24_combout ;
wire \twiddle_data~25_combout ;
wire \twiddle_data~26_combout ;
wire \twiddle_data~27_combout ;
wire \twiddle_data~28_combout ;
wire \twiddle_data~29_combout ;
wire \twiddle_data~30_combout ;
wire \twiddle_data~31_combout ;
wire \twiddle_data~32_combout ;
wire \twiddle_data~33_combout ;
wire \twiddle_data~34_combout ;
wire \twiddle_data~35_combout ;
wire \twiddle_data~36_combout ;
wire \twiddle_data~37_combout ;
wire \twiddle_data~38_combout ;
wire \twiddle_data~39_combout ;
wire \twiddle_data~40_combout ;
wire \twiddle_data~41_combout ;
wire \twiddle_data~42_combout ;
wire \twiddle_data~43_combout ;
wire \twiddle_data~44_combout ;
wire \twiddle_data~45_combout ;
wire \twiddle_data~46_combout ;
wire \twiddle_data~47_combout ;
wire \en_slb~q ;
wire \ram_a_not_b_vec[26]~q ;
wire \p_cd_en[2]~q ;
wire \p_cd_en[0]~q ;
wire \p_cd_en[1]~q ;
wire \twid_factors|twad_tdl[6][0]~q ;
wire \twid_factors|twad_tdl[6][1]~q ;
wire \twid_factors|twad_tdl[6][2]~q ;
wire \twid_factors|twad_tdl[6][3]~q ;
wire \twid_factors|twad_tdl[6][4]~q ;
wire \twid_factors|twad_tdl[6][5]~q ;
wire \twid_factors|twad_tdl[6][6]~q ;
wire \gen_dft_2:bfpdft|next_pass_vec[2]~q ;
wire \delay_ctrl_np|tdl_arr[9]~q ;
wire \en_slb~0_combout ;
wire \ram_a_not_b_vec[25]~q ;
wire \ram_a_not_b_vec~0_combout ;
wire \p_tdl[14][2]~q ;
wire \p_tdl[14][0]~q ;
wire \p_tdl[14][1]~q ;
wire \ram_a_not_b_vec[24]~q ;
wire \ram_a_not_b_vec~1_combout ;
wire \p_tdl[13][2]~q ;
wire \p_tdl[13][0]~q ;
wire \p_tdl[13][1]~q ;
wire \ram_a_not_b_vec[23]~q ;
wire \ram_a_not_b_vec~2_combout ;
wire \p_tdl[12][2]~q ;
wire \p_tdl[12][0]~q ;
wire \p_tdl[12][1]~q ;
wire \ccc|ram_data_out0[10]~q ;
wire \ccc|ram_data_out1[10]~q ;
wire \sw_r_tdl[4][0]~q ;
wire \ccc|ram_data_out2[10]~q ;
wire \ccc|ram_data_out3[10]~q ;
wire \sw_r_tdl[4][1]~q ;
wire \ccc|ram_data_out0[14]~q ;
wire \ccc|ram_data_out1[14]~q ;
wire \ccc|ram_data_out2[14]~q ;
wire \ccc|ram_data_out3[14]~q ;
wire \ccc|ram_data_out0[12]~q ;
wire \ccc|ram_data_out1[12]~q ;
wire \ccc|ram_data_out2[12]~q ;
wire \ccc|ram_data_out3[12]~q ;
wire \ccc|ram_data_out0[11]~q ;
wire \ccc|ram_data_out1[11]~q ;
wire \ccc|ram_data_out2[11]~q ;
wire \ccc|ram_data_out3[11]~q ;
wire \ccc|ram_data_out0[13]~q ;
wire \ccc|ram_data_out1[13]~q ;
wire \ccc|ram_data_out2[13]~q ;
wire \ccc|ram_data_out3[13]~q ;
wire \ccc|ram_data_out0[9]~q ;
wire \ccc|ram_data_out1[9]~q ;
wire \ccc|ram_data_out2[9]~q ;
wire \ccc|ram_data_out3[9]~q ;
wire \ccc|ram_data_out0[8]~q ;
wire \ccc|ram_data_out1[8]~q ;
wire \ccc|ram_data_out2[8]~q ;
wire \ccc|ram_data_out3[8]~q ;
wire \ccc|ram_data_out0[15]~q ;
wire \ccc|ram_data_out1[15]~q ;
wire \ccc|ram_data_out2[15]~q ;
wire \ccc|ram_data_out3[15]~q ;
wire \ccc|ram_data_out0[7]~q ;
wire \ccc|ram_data_out1[7]~q ;
wire \ccc|ram_data_out2[7]~q ;
wire \ccc|ram_data_out3[7]~q ;
wire \ccc|ram_data_out0[3]~q ;
wire \ccc|ram_data_out1[3]~q ;
wire \ccc|ram_data_out2[3]~q ;
wire \ccc|ram_data_out3[3]~q ;
wire \ccc|ram_data_out0[5]~q ;
wire \ccc|ram_data_out1[5]~q ;
wire \ccc|ram_data_out2[5]~q ;
wire \ccc|ram_data_out3[5]~q ;
wire \ccc|ram_data_out0[4]~q ;
wire \ccc|ram_data_out1[4]~q ;
wire \ccc|ram_data_out2[4]~q ;
wire \ccc|ram_data_out3[4]~q ;
wire \ccc|ram_data_out0[6]~q ;
wire \ccc|ram_data_out1[6]~q ;
wire \ccc|ram_data_out2[6]~q ;
wire \ccc|ram_data_out3[6]~q ;
wire \ccc|ram_data_out0[2]~q ;
wire \ccc|ram_data_out1[2]~q ;
wire \ccc|ram_data_out2[2]~q ;
wire \ccc|ram_data_out3[2]~q ;
wire \ccc|ram_data_out0[1]~q ;
wire \ccc|ram_data_out1[1]~q ;
wire \ccc|ram_data_out2[1]~q ;
wire \ccc|ram_data_out3[1]~q ;
wire \ccc|ram_data_out0[0]~q ;
wire \ccc|ram_data_out1[0]~q ;
wire \ccc|ram_data_out2[0]~q ;
wire \ccc|ram_data_out3[0]~q ;
wire \ram_a_not_b_vec[22]~q ;
wire \ram_a_not_b_vec~3_combout ;
wire \p_tdl[11][2]~q ;
wire \p_tdl[11][0]~q ;
wire \p_tdl[11][1]~q ;
wire \data_rdy_vec[10]~q ;
wire \ram_a_not_b_vec[10]~q ;
wire \sw_r_tdl[3][0]~q ;
wire \sw_r_tdl[3][1]~q ;
wire \ram_a_not_b_vec[21]~q ;
wire \ram_a_not_b_vec~4_combout ;
wire \p_tdl[10][2]~q ;
wire \p_tdl[10][0]~q ;
wire \p_tdl[10][1]~q ;
wire \ccc|b_ram_data_in_bus[58]~q ;
wire \ccc|wraddress_b_bus[21]~q ;
wire \ccc|wraddress_b_bus[22]~q ;
wire \ccc|wraddress_b_bus[23]~q ;
wire \ccc|wraddress_b_bus[24]~q ;
wire \ccc|wraddress_b_bus[11]~q ;
wire \ccc|wraddress_b_bus[26]~q ;
wire \ccc|wraddress_b_bus[13]~q ;
wire \ccc|rdaddress_b_bus[21]~q ;
wire \ccc|rdaddress_b_bus[22]~q ;
wire \ccc|rdaddress_b_bus[23]~q ;
wire \ccc|rdaddress_b_bus[24]~q ;
wire \ccc|rdaddress_b_bus[11]~q ;
wire \ccc|rdaddress_b_bus[26]~q ;
wire \ccc|rdaddress_b_bus[13]~q ;
wire \ccc|a_ram_data_in_bus[58]~q ;
wire \ccc|wraddress_a_bus[21]~q ;
wire \ccc|wraddress_a_bus[22]~q ;
wire \ccc|wraddress_a_bus[23]~q ;
wire \ccc|wraddress_a_bus[24]~q ;
wire \ccc|wraddress_a_bus[11]~q ;
wire \ccc|wraddress_a_bus[26]~q ;
wire \ccc|wraddress_a_bus[13]~q ;
wire \ccc|rdaddress_a_bus[21]~q ;
wire \ccc|rdaddress_a_bus[22]~q ;
wire \ccc|rdaddress_a_bus[23]~q ;
wire \ccc|rdaddress_a_bus[24]~q ;
wire \ccc|rdaddress_a_bus[11]~q ;
wire \ccc|rdaddress_a_bus[26]~q ;
wire \ccc|rdaddress_a_bus[13]~q ;
wire \data_rdy_vec[9]~q ;
wire \data_rdy_vec~5_combout ;
wire \ram_a_not_b_vec[9]~q ;
wire \ram_a_not_b_vec~5_combout ;
wire \ccc|b_ram_data_in_bus[42]~q ;
wire \ccc|wraddress_b_bus[0]~q ;
wire \ccc|wraddress_b_bus[15]~q ;
wire \ccc|wraddress_b_bus[16]~q ;
wire \ccc|wraddress_b_bus[17]~q ;
wire \ccc|wraddress_b_bus[18]~q ;
wire \ccc|wraddress_b_bus[19]~q ;
wire \ccc|rdaddress_b_bus[0]~q ;
wire \ccc|rdaddress_b_bus[15]~q ;
wire \ccc|rdaddress_b_bus[16]~q ;
wire \ccc|rdaddress_b_bus[17]~q ;
wire \ccc|rdaddress_b_bus[18]~q ;
wire \ccc|rdaddress_b_bus[19]~q ;
wire \ccc|a_ram_data_in_bus[42]~q ;
wire \ccc|wraddress_a_bus[0]~q ;
wire \ccc|wraddress_a_bus[15]~q ;
wire \ccc|wraddress_a_bus[16]~q ;
wire \ccc|wraddress_a_bus[17]~q ;
wire \ccc|wraddress_a_bus[18]~q ;
wire \ccc|wraddress_a_bus[19]~q ;
wire \ccc|rdaddress_a_bus[0]~q ;
wire \ccc|rdaddress_a_bus[15]~q ;
wire \ccc|rdaddress_a_bus[16]~q ;
wire \ccc|rdaddress_a_bus[17]~q ;
wire \ccc|rdaddress_a_bus[18]~q ;
wire \ccc|rdaddress_a_bus[19]~q ;
wire \sw_r_tdl[2][0]~q ;
wire \ccc|b_ram_data_in_bus[26]~q ;
wire \ccc|wraddress_b_bus[8]~q ;
wire \ccc|wraddress_b_bus[10]~q ;
wire \ccc|wraddress_b_bus[12]~q ;
wire \ccc|rdaddress_b_bus[8]~q ;
wire \ccc|rdaddress_b_bus[10]~q ;
wire \ccc|rdaddress_b_bus[12]~q ;
wire \ccc|a_ram_data_in_bus[26]~q ;
wire \ccc|wraddress_a_bus[8]~q ;
wire \ccc|wraddress_a_bus[10]~q ;
wire \ccc|wraddress_a_bus[12]~q ;
wire \ccc|rdaddress_a_bus[8]~q ;
wire \ccc|rdaddress_a_bus[10]~q ;
wire \ccc|rdaddress_a_bus[12]~q ;
wire \ccc|b_ram_data_in_bus[10]~q ;
wire \ccc|wraddress_b_bus[1]~q ;
wire \ccc|wraddress_b_bus[3]~q ;
wire \ccc|wraddress_b_bus[5]~q ;
wire \ccc|rdaddress_b_bus[1]~q ;
wire \ccc|rdaddress_b_bus[3]~q ;
wire \ccc|rdaddress_b_bus[5]~q ;
wire \ccc|a_ram_data_in_bus[10]~q ;
wire \ccc|wraddress_a_bus[1]~q ;
wire \ccc|wraddress_a_bus[3]~q ;
wire \ccc|wraddress_a_bus[5]~q ;
wire \ccc|rdaddress_a_bus[1]~q ;
wire \ccc|rdaddress_a_bus[3]~q ;
wire \ccc|rdaddress_a_bus[5]~q ;
wire \sw_r_tdl[2][1]~q ;
wire \ccc|b_ram_data_in_bus[62]~q ;
wire \ccc|a_ram_data_in_bus[62]~q ;
wire \ccc|b_ram_data_in_bus[46]~q ;
wire \ccc|a_ram_data_in_bus[46]~q ;
wire \ccc|b_ram_data_in_bus[30]~q ;
wire \ccc|a_ram_data_in_bus[30]~q ;
wire \ccc|b_ram_data_in_bus[14]~q ;
wire \ccc|a_ram_data_in_bus[14]~q ;
wire \ccc|b_ram_data_in_bus[60]~q ;
wire \ccc|a_ram_data_in_bus[60]~q ;
wire \ccc|b_ram_data_in_bus[44]~q ;
wire \ccc|a_ram_data_in_bus[44]~q ;
wire \ccc|b_ram_data_in_bus[28]~q ;
wire \ccc|a_ram_data_in_bus[28]~q ;
wire \ccc|b_ram_data_in_bus[12]~q ;
wire \ccc|a_ram_data_in_bus[12]~q ;
wire \ccc|b_ram_data_in_bus[59]~q ;
wire \ccc|a_ram_data_in_bus[59]~q ;
wire \ccc|b_ram_data_in_bus[43]~q ;
wire \ccc|a_ram_data_in_bus[43]~q ;
wire \ccc|b_ram_data_in_bus[27]~q ;
wire \ccc|a_ram_data_in_bus[27]~q ;
wire \ccc|b_ram_data_in_bus[11]~q ;
wire \ccc|a_ram_data_in_bus[11]~q ;
wire \ccc|b_ram_data_in_bus[61]~q ;
wire \ccc|a_ram_data_in_bus[61]~q ;
wire \ccc|b_ram_data_in_bus[45]~q ;
wire \ccc|a_ram_data_in_bus[45]~q ;
wire \ccc|b_ram_data_in_bus[29]~q ;
wire \ccc|a_ram_data_in_bus[29]~q ;
wire \ccc|b_ram_data_in_bus[13]~q ;
wire \ccc|a_ram_data_in_bus[13]~q ;
wire \ccc|b_ram_data_in_bus[57]~q ;
wire \ccc|a_ram_data_in_bus[57]~q ;
wire \ccc|b_ram_data_in_bus[41]~q ;
wire \ccc|a_ram_data_in_bus[41]~q ;
wire \ccc|b_ram_data_in_bus[25]~q ;
wire \ccc|a_ram_data_in_bus[25]~q ;
wire \ccc|b_ram_data_in_bus[9]~q ;
wire \ccc|a_ram_data_in_bus[9]~q ;
wire \ccc|b_ram_data_in_bus[56]~q ;
wire \ccc|a_ram_data_in_bus[56]~q ;
wire \ccc|b_ram_data_in_bus[40]~q ;
wire \ccc|a_ram_data_in_bus[40]~q ;
wire \ccc|b_ram_data_in_bus[24]~q ;
wire \ccc|a_ram_data_in_bus[24]~q ;
wire \ccc|b_ram_data_in_bus[8]~q ;
wire \ccc|a_ram_data_in_bus[8]~q ;
wire \ccc|b_ram_data_in_bus[63]~q ;
wire \ccc|a_ram_data_in_bus[63]~q ;
wire \ccc|b_ram_data_in_bus[47]~q ;
wire \ccc|a_ram_data_in_bus[47]~q ;
wire \ccc|b_ram_data_in_bus[31]~q ;
wire \ccc|a_ram_data_in_bus[31]~q ;
wire \ccc|b_ram_data_in_bus[15]~q ;
wire \ccc|a_ram_data_in_bus[15]~q ;
wire \ccc|b_ram_data_in_bus[55]~q ;
wire \ccc|a_ram_data_in_bus[55]~q ;
wire \ccc|b_ram_data_in_bus[39]~q ;
wire \ccc|a_ram_data_in_bus[39]~q ;
wire \ccc|b_ram_data_in_bus[23]~q ;
wire \ccc|a_ram_data_in_bus[23]~q ;
wire \ccc|b_ram_data_in_bus[7]~q ;
wire \ccc|a_ram_data_in_bus[7]~q ;
wire \ccc|b_ram_data_in_bus[51]~q ;
wire \ccc|a_ram_data_in_bus[51]~q ;
wire \ccc|b_ram_data_in_bus[35]~q ;
wire \ccc|a_ram_data_in_bus[35]~q ;
wire \ccc|b_ram_data_in_bus[19]~q ;
wire \ccc|a_ram_data_in_bus[19]~q ;
wire \ccc|b_ram_data_in_bus[3]~q ;
wire \ccc|a_ram_data_in_bus[3]~q ;
wire \ccc|b_ram_data_in_bus[53]~q ;
wire \ccc|a_ram_data_in_bus[53]~q ;
wire \ccc|b_ram_data_in_bus[37]~q ;
wire \ccc|a_ram_data_in_bus[37]~q ;
wire \ccc|b_ram_data_in_bus[21]~q ;
wire \ccc|a_ram_data_in_bus[21]~q ;
wire \ccc|b_ram_data_in_bus[5]~q ;
wire \ccc|a_ram_data_in_bus[5]~q ;
wire \ccc|b_ram_data_in_bus[52]~q ;
wire \ccc|a_ram_data_in_bus[52]~q ;
wire \ccc|b_ram_data_in_bus[36]~q ;
wire \ccc|a_ram_data_in_bus[36]~q ;
wire \ccc|b_ram_data_in_bus[20]~q ;
wire \ccc|a_ram_data_in_bus[20]~q ;
wire \ccc|b_ram_data_in_bus[4]~q ;
wire \ccc|a_ram_data_in_bus[4]~q ;
wire \ccc|b_ram_data_in_bus[54]~q ;
wire \ccc|a_ram_data_in_bus[54]~q ;
wire \ccc|b_ram_data_in_bus[38]~q ;
wire \ccc|a_ram_data_in_bus[38]~q ;
wire \ccc|b_ram_data_in_bus[22]~q ;
wire \ccc|a_ram_data_in_bus[22]~q ;
wire \ccc|b_ram_data_in_bus[6]~q ;
wire \ccc|a_ram_data_in_bus[6]~q ;
wire \ccc|b_ram_data_in_bus[50]~q ;
wire \ccc|a_ram_data_in_bus[50]~q ;
wire \ccc|b_ram_data_in_bus[34]~q ;
wire \ccc|a_ram_data_in_bus[34]~q ;
wire \ccc|b_ram_data_in_bus[18]~q ;
wire \ccc|a_ram_data_in_bus[18]~q ;
wire \ccc|b_ram_data_in_bus[2]~q ;
wire \ccc|a_ram_data_in_bus[2]~q ;
wire \ccc|b_ram_data_in_bus[49]~q ;
wire \ccc|a_ram_data_in_bus[49]~q ;
wire \ccc|b_ram_data_in_bus[33]~q ;
wire \ccc|a_ram_data_in_bus[33]~q ;
wire \ccc|b_ram_data_in_bus[17]~q ;
wire \ccc|a_ram_data_in_bus[17]~q ;
wire \ccc|b_ram_data_in_bus[1]~q ;
wire \ccc|a_ram_data_in_bus[1]~q ;
wire \ccc|b_ram_data_in_bus[48]~q ;
wire \ccc|a_ram_data_in_bus[48]~q ;
wire \ccc|b_ram_data_in_bus[32]~q ;
wire \ccc|a_ram_data_in_bus[32]~q ;
wire \ccc|b_ram_data_in_bus[16]~q ;
wire \ccc|a_ram_data_in_bus[16]~q ;
wire \ccc|b_ram_data_in_bus[0]~q ;
wire \ccc|a_ram_data_in_bus[0]~q ;
wire \ram_a_not_b_vec[20]~q ;
wire \ram_a_not_b_vec~6_combout ;
wire \p_tdl[9][2]~q ;
wire \p_tdl[9][0]~q ;
wire \p_tdl[9][1]~q ;
wire \ram_a_not_b_vec[29]~q ;
wire \ram_a_not_b_vec[1]~q ;
wire \wren_b~0_combout ;
wire \writer|data_in_r[2]~q ;
wire \writer|wr_address_i_int[0]~q ;
wire \writer|wr_address_i_int[1]~q ;
wire \writer|wr_address_i_int[2]~q ;
wire \writer|wr_address_i_int[3]~q ;
wire \writer|wr_address_i_int[4]~q ;
wire \writer|wr_address_i_int[5]~q ;
wire \writer|wr_address_i_int[6]~q ;
wire \ram_a_not_b_vec[7]~q ;
wire \ram_cxb_rd|ram_in_reg[0][0]~q ;
wire \ram_cxb_rd|ram_in_reg[0][1]~q ;
wire \ram_cxb_rd|ram_in_reg[0][2]~q ;
wire \ram_cxb_rd|ram_in_reg[0][3]~q ;
wire \ram_cxb_rd|ram_in_reg[0][4]~q ;
wire \ram_cxb_rd|ram_in_reg[0][5]~q ;
wire \gen_wrsw_2:k_delay|tdl_arr[1][6]~q ;
wire \wren_a~0_combout ;
wire \data_rdy_vec[8]~q ;
wire \data_rdy_vec~6_combout ;
wire \ram_a_not_b_vec[8]~q ;
wire \ram_a_not_b_vec~7_combout ;
wire \wren_b~1_combout ;
wire \ram_cxb_rd|ram_in_reg[1][0]~q ;
wire \ram_cxb_rd|ram_in_reg[1][1]~q ;
wire \ram_cxb_rd|ram_in_reg[1][2]~q ;
wire \ram_cxb_rd|ram_in_reg[1][3]~q ;
wire \ram_cxb_rd|ram_in_reg[1][4]~q ;
wire \ram_cxb_rd|ram_in_reg[1][5]~q ;
wire \wren_a~1_combout ;
wire \sw_r_tdl[1][0]~q ;
wire \wren_b~2_combout ;
wire \ram_cxb_rd|ram_in_reg[2][1]~q ;
wire \ram_cxb_rd|ram_in_reg[2][3]~q ;
wire \ram_cxb_rd|ram_in_reg[2][5]~q ;
wire \wren_a~2_combout ;
wire \wren_b~3_combout ;
wire \ram_cxb_rd|ram_in_reg[3][1]~q ;
wire \ram_cxb_rd|ram_in_reg[3][3]~q ;
wire \ram_cxb_rd|ram_in_reg[3][5]~q ;
wire \wren_a~3_combout ;
wire \sw_r_tdl[1][1]~q ;
wire \writer|data_in_r[6]~q ;
wire \writer|data_in_r[4]~q ;
wire \writer|data_in_r[3]~q ;
wire \writer|data_in_r[5]~q ;
wire \writer|data_in_r[1]~q ;
wire \writer|data_in_r[0]~q ;
wire \writer|data_in_r[7]~q ;
wire \writer|data_in_i[7]~q ;
wire \writer|data_in_i[3]~q ;
wire \writer|data_in_i[5]~q ;
wire \writer|data_in_i[4]~q ;
wire \writer|data_in_i[6]~q ;
wire \writer|data_in_i[2]~q ;
wire \writer|data_in_i[1]~q ;
wire \writer|data_in_i[0]~q ;
wire \ram_a_not_b_vec[19]~q ;
wire \ram_a_not_b_vec~8_combout ;
wire \p_tdl[8][2]~q ;
wire \p_tdl[8][0]~q ;
wire \p_tdl[8][1]~q ;
wire \ram_a_not_b_vec[28]~q ;
wire \ram_a_not_b_vec~9_combout ;
wire \ram_a_not_b_vec[0]~q ;
wire \ram_a_not_b_vec~10_combout ;
wire \ram_a_not_b_vec[6]~q ;
wire \ram_a_not_b_vec~11_combout ;
wire \rd_adgen|rd_addr_d[0]~q ;
wire \rd_adgen|rd_addr_c[0]~q ;
wire \rd_adgen|sw[0]~q ;
wire \rd_adgen|rd_addr_b[1]~q ;
wire \rd_adgen|rd_addr_d[1]~q ;
wire \rd_adgen|sw[1]~q ;
wire \rd_adgen|rd_addr_d[2]~q ;
wire \rd_adgen|rd_addr_c[2]~q ;
wire \rd_adgen|rd_addr_b[3]~q ;
wire \rd_adgen|rd_addr_d[3]~q ;
wire \rd_adgen|rd_addr_d[4]~q ;
wire \rd_adgen|rd_addr_c[4]~q ;
wire \rd_adgen|rd_addr_b[5]~q ;
wire \rd_adgen|rd_addr_d[5]~q ;
wire \data_rdy_vec[7]~q ;
wire \data_rdy_vec~7_combout ;
wire \ram_a_not_b_vec~12_combout ;
wire \sw_r_tdl[0][0]~q ;
wire \sw_r_tdl[0][1]~q ;
wire \ram_a_not_b_vec[18]~q ;
wire \ram_a_not_b_vec~13_combout ;
wire \p_tdl[7][2]~q ;
wire \p_tdl[7][0]~q ;
wire \p_tdl[7][1]~q ;
wire \ram_a_not_b_vec[27]~q ;
wire \ram_a_not_b_vec~14_combout ;
wire \ram_a_not_b_vec~15_combout ;
wire \data_imag_in_reg[2]~q ;
wire \data_real_in_reg[2]~q ;
wire \core_real_in~0_combout ;
wire \ram_a_not_b_vec[5]~q ;
wire \ram_a_not_b_vec~16_combout ;
wire \gen_gt256_mk:ctrl|k_count[0]~q ;
wire \gen_gt256_mk:ctrl|k_count[2]~q ;
wire \rd_adgen|Mux7~1_combout ;
wire \rd_adgen|Mux1~0_combout ;
wire \gen_gt256_mk:ctrl|k_count[4]~q ;
wire \rd_adgen|Mux1~1_combout ;
wire \gen_gt256_mk:ctrl|k_count[1]~q ;
wire \gen_gt256_mk:ctrl|k_count[3]~q ;
wire \gen_gt256_mk:ctrl|k_count[5]~q ;
wire \gen_gt256_mk:ctrl|k_count[6]~q ;
wire \data_rdy_vec[6]~q ;
wire \data_rdy_vec~8_combout ;
wire \data_imag_in_reg[6]~q ;
wire \data_real_in_reg[6]~q ;
wire \core_real_in~1_combout ;
wire \data_imag_in_reg[4]~q ;
wire \data_real_in_reg[4]~q ;
wire \core_real_in~2_combout ;
wire \data_imag_in_reg[3]~q ;
wire \data_real_in_reg[3]~q ;
wire \core_real_in~3_combout ;
wire \data_imag_in_reg[5]~q ;
wire \data_real_in_reg[5]~q ;
wire \core_real_in~4_combout ;
wire \data_imag_in_reg[1]~q ;
wire \data_real_in_reg[1]~q ;
wire \core_real_in~5_combout ;
wire \data_imag_in_reg[0]~q ;
wire \data_real_in_reg[0]~q ;
wire \core_real_in~6_combout ;
wire \data_imag_in_reg[7]~q ;
wire \data_real_in_reg[7]~q ;
wire \core_real_in~7_combout ;
wire \core_imag_in~0_combout ;
wire \core_imag_in~1_combout ;
wire \core_imag_in~2_combout ;
wire \core_imag_in~3_combout ;
wire \core_imag_in~4_combout ;
wire \core_imag_in~5_combout ;
wire \core_imag_in~6_combout ;
wire \core_imag_in~7_combout ;
wire \ram_a_not_b_vec[17]~q ;
wire \ram_a_not_b_vec~17_combout ;
wire \p_tdl[6][2]~q ;
wire \p_tdl[6][0]~q ;
wire \p_tdl[6][1]~q ;
wire \ram_a_not_b_vec~18_combout ;
wire \data_imag_in_reg~0_combout ;
wire \data_real_in_reg~0_combout ;
wire \ram_a_not_b_vec[4]~q ;
wire \ram_a_not_b_vec~19_combout ;
wire \data_rdy_vec[5]~q ;
wire \data_rdy_vec~9_combout ;
wire \data_imag_in_reg~1_combout ;
wire \data_real_in_reg~1_combout ;
wire \data_imag_in_reg~2_combout ;
wire \data_real_in_reg~2_combout ;
wire \data_imag_in_reg~3_combout ;
wire \data_real_in_reg~3_combout ;
wire \data_imag_in_reg~4_combout ;
wire \data_real_in_reg~4_combout ;
wire \data_imag_in_reg~5_combout ;
wire \data_real_in_reg~5_combout ;
wire \data_imag_in_reg~6_combout ;
wire \data_real_in_reg~6_combout ;
wire \data_imag_in_reg~7_combout ;
wire \data_real_in_reg~7_combout ;
wire \ram_a_not_b_vec[16]~q ;
wire \ram_a_not_b_vec~20_combout ;
wire \p_tdl[5][2]~q ;
wire \p_tdl[5][0]~q ;
wire \p_tdl[5][1]~q ;
wire \ram_a_not_b_vec[3]~q ;
wire \ram_a_not_b_vec~21_combout ;
wire \data_rdy_vec~10_combout ;
wire \ram_a_not_b_vec[15]~q ;
wire \ram_a_not_b_vec~22_combout ;
wire \p_tdl[4][2]~q ;
wire \p_tdl[4][0]~q ;
wire \p_tdl[4][1]~q ;
wire \ram_a_not_b_vec[2]~q ;
wire \ram_a_not_b_vec~23_combout ;
wire \ram_a_not_b_vec[14]~q ;
wire \ram_a_not_b_vec~24_combout ;
wire \p_tdl[3][2]~q ;
wire \p_tdl[3][0]~q ;
wire \p_tdl[3][1]~q ;
wire \ram_a_not_b_vec~25_combout ;
wire \ram_a_not_b_vec[13]~q ;
wire \ram_a_not_b_vec~26_combout ;
wire \p_tdl[2][2]~q ;
wire \p_tdl[2][0]~q ;
wire \p_tdl[2][1]~q ;
wire \ram_a_not_b_vec[12]~q ;
wire \ram_a_not_b_vec~27_combout ;
wire \p_tdl[1][2]~q ;
wire \p_tdl[1][0]~q ;
wire \p_tdl[1][1]~q ;
wire \ram_a_not_b_vec[11]~q ;
wire \ram_a_not_b_vec~28_combout ;
wire \p_tdl[0][2]~q ;
wire \p_tdl[0][0]~q ;
wire \p_tdl[0][1]~q ;
wire \ram_a_not_b_vec~29_combout ;


fft_asj_fft_tdl_bit_rst_fft_120_7 delay_lpp_en(
	.global_clock_enable(\global_clock_enable~0_combout ),
	.tdl_arr_3(\delay_lpp_en|tdl_arr[3]~q ),
	.tdl_arr_4(\gen_radix_2_last_pass:gen_lpp_addr|delay_en|tdl_arr[4]~q ),
	.clk(clk),
	.reset_n(reset_n));

fft_asj_fft_lpp_serial_r2_fft_120 \gen_radix_2_last_pass:lpp_r2 (
	.lpp_ram_data_out_sw_1_1(\lpp_ram_data_out_sw[1][1]~q ),
	.lpp_ram_data_out_sw_1_0(\lpp_ram_data_out_sw[0][1]~q ),
	.lpp_ram_data_out_sw_0_1(\lpp_ram_data_out_sw[1][0]~q ),
	.lpp_ram_data_out_sw_0_0(\lpp_ram_data_out_sw[0][0]~q ),
	.lpp_ram_data_out_sw_7_1(\lpp_ram_data_out_sw[1][7]~q ),
	.lpp_ram_data_out_sw_7_0(\lpp_ram_data_out_sw[0][7]~q ),
	.lpp_ram_data_out_sw_6_1(\lpp_ram_data_out_sw[1][6]~q ),
	.lpp_ram_data_out_sw_6_0(\lpp_ram_data_out_sw[0][6]~q ),
	.lpp_ram_data_out_sw_5_1(\lpp_ram_data_out_sw[1][5]~q ),
	.lpp_ram_data_out_sw_5_0(\lpp_ram_data_out_sw[0][5]~q ),
	.lpp_ram_data_out_sw_4_1(\lpp_ram_data_out_sw[1][4]~q ),
	.lpp_ram_data_out_sw_4_0(\lpp_ram_data_out_sw[0][4]~q ),
	.lpp_ram_data_out_sw_3_1(\lpp_ram_data_out_sw[1][3]~q ),
	.lpp_ram_data_out_sw_3_0(\lpp_ram_data_out_sw[0][3]~q ),
	.lpp_ram_data_out_sw_2_1(\lpp_ram_data_out_sw[1][2]~q ),
	.lpp_ram_data_out_sw_2_0(\lpp_ram_data_out_sw[0][2]~q ),
	.lpp_ram_data_out_sw_9_1(\lpp_ram_data_out_sw[1][9]~q ),
	.lpp_ram_data_out_sw_9_0(\lpp_ram_data_out_sw[0][9]~q ),
	.lpp_ram_data_out_sw_8_1(\lpp_ram_data_out_sw[1][8]~q ),
	.lpp_ram_data_out_sw_8_0(\lpp_ram_data_out_sw[0][8]~q ),
	.lpp_ram_data_out_sw_15_1(\lpp_ram_data_out_sw[1][15]~q ),
	.lpp_ram_data_out_sw_15_0(\lpp_ram_data_out_sw[0][15]~q ),
	.lpp_ram_data_out_sw_14_1(\lpp_ram_data_out_sw[1][14]~q ),
	.lpp_ram_data_out_sw_14_0(\lpp_ram_data_out_sw[0][14]~q ),
	.lpp_ram_data_out_sw_13_1(\lpp_ram_data_out_sw[1][13]~q ),
	.lpp_ram_data_out_sw_13_0(\lpp_ram_data_out_sw[0][13]~q ),
	.lpp_ram_data_out_sw_12_1(\lpp_ram_data_out_sw[1][12]~q ),
	.lpp_ram_data_out_sw_12_0(\lpp_ram_data_out_sw[0][12]~q ),
	.lpp_ram_data_out_sw_11_1(\lpp_ram_data_out_sw[1][11]~q ),
	.lpp_ram_data_out_sw_11_0(\lpp_ram_data_out_sw[0][11]~q ),
	.lpp_ram_data_out_sw_10_1(\lpp_ram_data_out_sw[1][10]~q ),
	.lpp_ram_data_out_sw_10_0(\lpp_ram_data_out_sw[0][10]~q ),
	.source_valid_ctrl_sop(\source_valid_ctrl_sop~1_combout ),
	.stall_reg(\auk_dsp_interface_controller_1|stall_reg~q ),
	.source_stall_int_d(\auk_dsp_atlantic_source_1|source_stall_int_d~q ),
	.global_clock_enable(\global_clock_enable~0_combout ),
	.data_imag_o_0(\gen_radix_2_last_pass:lpp_r2|data_imag_o[0]~q ),
	.data_real_o_0(\gen_radix_2_last_pass:lpp_r2|data_real_o[0]~q ),
	.data_imag_o_1(\gen_radix_2_last_pass:lpp_r2|data_imag_o[1]~q ),
	.data_real_o_1(\gen_radix_2_last_pass:lpp_r2|data_real_o[1]~q ),
	.data_imag_o_2(\gen_radix_2_last_pass:lpp_r2|data_imag_o[2]~q ),
	.data_real_o_2(\gen_radix_2_last_pass:lpp_r2|data_real_o[2]~q ),
	.data_imag_o_3(\gen_radix_2_last_pass:lpp_r2|data_imag_o[3]~q ),
	.data_real_o_3(\gen_radix_2_last_pass:lpp_r2|data_real_o[3]~q ),
	.data_imag_o_4(\gen_radix_2_last_pass:lpp_r2|data_imag_o[4]~q ),
	.data_real_o_4(\gen_radix_2_last_pass:lpp_r2|data_real_o[4]~q ),
	.data_imag_o_5(\gen_radix_2_last_pass:lpp_r2|data_imag_o[5]~q ),
	.data_real_o_5(\gen_radix_2_last_pass:lpp_r2|data_real_o[5]~q ),
	.data_imag_o_6(\gen_radix_2_last_pass:lpp_r2|data_imag_o[6]~q ),
	.data_real_o_6(\gen_radix_2_last_pass:lpp_r2|data_real_o[6]~q ),
	.data_imag_o_7(\gen_radix_2_last_pass:lpp_r2|data_imag_o[7]~q ),
	.data_real_o_7(\gen_radix_2_last_pass:lpp_r2|data_real_o[7]~q ),
	.tdl_arr_4(\gen_radix_2_last_pass:gen_lpp_addr|delay_en|tdl_arr[4]~q ),
	.clk(clk),
	.reset_n(reset_n));

fft_asj_fft_tdl_bit_fft_120_4 \gen_radix_2_last_pass:delay_mid (
	.global_clock_enable(\global_clock_enable~0_combout ),
	.tdl_arr_4(\gen_radix_2_last_pass:delay_mid|tdl_arr[4]~q ),
	.rd_addr_b_6(\gen_radix_2_last_pass:gen_lpp_addr|rd_addr_b[6]~q ),
	.clk(clk));

fft_asj_fft_cxb_addr_fft_120 \gen_radix_2_last_pass:ram_cxb_rd_lpp (
	.sw_0(\gen_radix_2_last_pass:gen_lpp_addr|sw[0]~q ),
	.global_clock_enable(\global_clock_enable~0_combout ),
	.ram_in_reg_0_0(\gen_radix_2_last_pass:ram_cxb_rd_lpp|ram_in_reg[0][0]~q ),
	.ram_in_reg_1_0(\gen_radix_2_last_pass:ram_cxb_rd_lpp|ram_in_reg[0][1]~q ),
	.ram_in_reg_2_0(\gen_radix_2_last_pass:ram_cxb_rd_lpp|ram_in_reg[0][2]~q ),
	.ram_in_reg_3_0(\gen_radix_2_last_pass:ram_cxb_rd_lpp|ram_in_reg[0][3]~q ),
	.ram_in_reg_4_0(\gen_radix_2_last_pass:ram_cxb_rd_lpp|ram_in_reg[0][4]~q ),
	.ram_in_reg_5_0(\gen_radix_2_last_pass:ram_cxb_rd_lpp|ram_in_reg[0][5]~q ),
	.ram_in_reg_6_1(\gen_radix_2_last_pass:ram_cxb_rd_lpp|ram_in_reg[1][6]~q ),
	.rd_addr_b_0(\gen_radix_2_last_pass:gen_lpp_addr|rd_addr_b[0]~q ),
	.rd_addr_b_1(\gen_radix_2_last_pass:gen_lpp_addr|rd_addr_b[1]~q ),
	.rd_addr_b_2(\gen_radix_2_last_pass:gen_lpp_addr|rd_addr_b[2]~q ),
	.rd_addr_b_3(\gen_radix_2_last_pass:gen_lpp_addr|rd_addr_b[3]~q ),
	.rd_addr_b_4(\gen_radix_2_last_pass:gen_lpp_addr|rd_addr_b[4]~q ),
	.rd_addr_b_5(\gen_radix_2_last_pass:gen_lpp_addr|rd_addr_b[5]~q ),
	.rd_addr_b_6(\gen_radix_2_last_pass:gen_lpp_addr|rd_addr_b[6]~q ),
	.clk(clk));

fft_asj_fft_lpprdadr2gen_fft_120 \gen_radix_2_last_pass:gen_lpp_addr (
	.sw_0(\gen_radix_2_last_pass:gen_lpp_addr|sw[0]~q ),
	.global_clock_enable(\global_clock_enable~0_combout ),
	.tdl_arr_4(\gen_radix_2_last_pass:gen_lpp_addr|delay_en|tdl_arr[4]~q ),
	.tdl_arr_0_4(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.tdl_arr_1_4(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.tdl_arr_19(\gen_dft_2:delay_blk_done2|tdl_arr[19]~q ),
	.rd_addr_b_0(\gen_radix_2_last_pass:gen_lpp_addr|rd_addr_b[0]~q ),
	.rd_addr_b_1(\gen_radix_2_last_pass:gen_lpp_addr|rd_addr_b[1]~q ),
	.rd_addr_b_2(\gen_radix_2_last_pass:gen_lpp_addr|rd_addr_b[2]~q ),
	.rd_addr_b_3(\gen_radix_2_last_pass:gen_lpp_addr|rd_addr_b[3]~q ),
	.rd_addr_b_4(\gen_radix_2_last_pass:gen_lpp_addr|rd_addr_b[4]~q ),
	.rd_addr_b_5(\gen_radix_2_last_pass:gen_lpp_addr|rd_addr_b[5]~q ),
	.rd_addr_b_6(\gen_radix_2_last_pass:gen_lpp_addr|rd_addr_b[6]~q ),
	.clk(clk),
	.reset_n(reset_n));

fft_asj_fft_3dp_rom_fft_120 twrom(
	.q_a_0(\twrom|gen_M4K:cos_1n|gen_auto:altsyncram_component|auto_generated|q_a[0] ),
	.q_a_1(\twrom|gen_M4K:cos_1n|gen_auto:altsyncram_component|auto_generated|q_a[1] ),
	.q_a_2(\twrom|gen_M4K:cos_1n|gen_auto:altsyncram_component|auto_generated|q_a[2] ),
	.q_a_3(\twrom|gen_M4K:cos_1n|gen_auto:altsyncram_component|auto_generated|q_a[3] ),
	.q_a_4(\twrom|gen_M4K:cos_1n|gen_auto:altsyncram_component|auto_generated|q_a[4] ),
	.q_a_5(\twrom|gen_M4K:cos_1n|gen_auto:altsyncram_component|auto_generated|q_a[5] ),
	.q_a_6(\twrom|gen_M4K:cos_1n|gen_auto:altsyncram_component|auto_generated|q_a[6] ),
	.q_a_7(\twrom|gen_M4K:cos_1n|gen_auto:altsyncram_component|auto_generated|q_a[7] ),
	.q_a_01(\twrom|gen_M4K:sin_1n|gen_auto:altsyncram_component|auto_generated|q_a[0] ),
	.q_a_11(\twrom|gen_M4K:sin_1n|gen_auto:altsyncram_component|auto_generated|q_a[1] ),
	.q_a_21(\twrom|gen_M4K:sin_1n|gen_auto:altsyncram_component|auto_generated|q_a[2] ),
	.q_a_31(\twrom|gen_M4K:sin_1n|gen_auto:altsyncram_component|auto_generated|q_a[3] ),
	.q_a_41(\twrom|gen_M4K:sin_1n|gen_auto:altsyncram_component|auto_generated|q_a[4] ),
	.q_a_51(\twrom|gen_M4K:sin_1n|gen_auto:altsyncram_component|auto_generated|q_a[5] ),
	.q_a_61(\twrom|gen_M4K:sin_1n|gen_auto:altsyncram_component|auto_generated|q_a[6] ),
	.q_a_71(\twrom|gen_M4K:sin_1n|gen_auto:altsyncram_component|auto_generated|q_a[7] ),
	.q_a_02(\twrom|gen_M4K:cos_2n|gen_auto:altsyncram_component|auto_generated|q_a[0] ),
	.q_a_12(\twrom|gen_M4K:cos_2n|gen_auto:altsyncram_component|auto_generated|q_a[1] ),
	.q_a_22(\twrom|gen_M4K:cos_2n|gen_auto:altsyncram_component|auto_generated|q_a[2] ),
	.q_a_32(\twrom|gen_M4K:cos_2n|gen_auto:altsyncram_component|auto_generated|q_a[3] ),
	.q_a_42(\twrom|gen_M4K:cos_2n|gen_auto:altsyncram_component|auto_generated|q_a[4] ),
	.q_a_52(\twrom|gen_M4K:cos_2n|gen_auto:altsyncram_component|auto_generated|q_a[5] ),
	.q_a_62(\twrom|gen_M4K:cos_2n|gen_auto:altsyncram_component|auto_generated|q_a[6] ),
	.q_a_72(\twrom|gen_M4K:cos_2n|gen_auto:altsyncram_component|auto_generated|q_a[7] ),
	.q_a_03(\twrom|gen_M4K:sin_2n|gen_auto:altsyncram_component|auto_generated|q_a[0] ),
	.q_a_13(\twrom|gen_M4K:sin_2n|gen_auto:altsyncram_component|auto_generated|q_a[1] ),
	.q_a_23(\twrom|gen_M4K:sin_2n|gen_auto:altsyncram_component|auto_generated|q_a[2] ),
	.q_a_33(\twrom|gen_M4K:sin_2n|gen_auto:altsyncram_component|auto_generated|q_a[3] ),
	.q_a_43(\twrom|gen_M4K:sin_2n|gen_auto:altsyncram_component|auto_generated|q_a[4] ),
	.q_a_53(\twrom|gen_M4K:sin_2n|gen_auto:altsyncram_component|auto_generated|q_a[5] ),
	.q_a_63(\twrom|gen_M4K:sin_2n|gen_auto:altsyncram_component|auto_generated|q_a[6] ),
	.q_a_73(\twrom|gen_M4K:sin_2n|gen_auto:altsyncram_component|auto_generated|q_a[7] ),
	.q_a_04(\twrom|gen_M4K:cos_3n|gen_auto:altsyncram_component|auto_generated|q_a[0] ),
	.q_a_14(\twrom|gen_M4K:cos_3n|gen_auto:altsyncram_component|auto_generated|q_a[1] ),
	.q_a_24(\twrom|gen_M4K:cos_3n|gen_auto:altsyncram_component|auto_generated|q_a[2] ),
	.q_a_34(\twrom|gen_M4K:cos_3n|gen_auto:altsyncram_component|auto_generated|q_a[3] ),
	.q_a_44(\twrom|gen_M4K:cos_3n|gen_auto:altsyncram_component|auto_generated|q_a[4] ),
	.q_a_54(\twrom|gen_M4K:cos_3n|gen_auto:altsyncram_component|auto_generated|q_a[5] ),
	.q_a_64(\twrom|gen_M4K:cos_3n|gen_auto:altsyncram_component|auto_generated|q_a[6] ),
	.q_a_74(\twrom|gen_M4K:cos_3n|gen_auto:altsyncram_component|auto_generated|q_a[7] ),
	.q_a_05(\twrom|gen_M4K:sin_3n|gen_auto:altsyncram_component|auto_generated|q_a[0] ),
	.q_a_15(\twrom|gen_M4K:sin_3n|gen_auto:altsyncram_component|auto_generated|q_a[1] ),
	.q_a_25(\twrom|gen_M4K:sin_3n|gen_auto:altsyncram_component|auto_generated|q_a[2] ),
	.q_a_35(\twrom|gen_M4K:sin_3n|gen_auto:altsyncram_component|auto_generated|q_a[3] ),
	.q_a_45(\twrom|gen_M4K:sin_3n|gen_auto:altsyncram_component|auto_generated|q_a[4] ),
	.q_a_55(\twrom|gen_M4K:sin_3n|gen_auto:altsyncram_component|auto_generated|q_a[5] ),
	.q_a_65(\twrom|gen_M4K:sin_3n|gen_auto:altsyncram_component|auto_generated|q_a[6] ),
	.q_a_75(\twrom|gen_M4K:sin_3n|gen_auto:altsyncram_component|auto_generated|q_a[7] ),
	.global_clock_enable(\global_clock_enable~0_combout ),
	.twad_tdl_0_6(\twid_factors|twad_tdl[6][0]~q ),
	.twad_tdl_1_6(\twid_factors|twad_tdl[6][1]~q ),
	.twad_tdl_2_6(\twid_factors|twad_tdl[6][2]~q ),
	.twad_tdl_3_6(\twid_factors|twad_tdl[6][3]~q ),
	.twad_tdl_4_6(\twid_factors|twad_tdl[6][4]~q ),
	.twad_tdl_5_6(\twid_factors|twad_tdl[6][5]~q ),
	.twad_tdl_6_6(\twid_factors|twad_tdl[6][6]~q ),
	.clk(clk));

fft_asj_fft_twadgen_fft_120 twid_factors(
	.global_clock_enable(\global_clock_enable~0_combout ),
	.p_2(\gen_gt256_mk:ctrl|p[2]~q ),
	.p_0(\gen_gt256_mk:ctrl|p[0]~q ),
	.p_1(\gen_gt256_mk:ctrl|p[1]~q ),
	.twad_tdl_0_6(\twid_factors|twad_tdl[6][0]~q ),
	.twad_tdl_1_6(\twid_factors|twad_tdl[6][1]~q ),
	.twad_tdl_2_6(\twid_factors|twad_tdl[6][2]~q ),
	.twad_tdl_3_6(\twid_factors|twad_tdl[6][3]~q ),
	.twad_tdl_4_6(\twid_factors|twad_tdl[6][4]~q ),
	.twad_tdl_5_6(\twid_factors|twad_tdl[6][5]~q ),
	.twad_tdl_6_6(\twid_factors|twad_tdl[6][6]~q ),
	.k_count_2(\gen_gt256_mk:ctrl|k_count[2]~q ),
	.Mux7(\rd_adgen|Mux7~1_combout ),
	.Mux1(\rd_adgen|Mux1~0_combout ),
	.k_count_4(\gen_gt256_mk:ctrl|k_count[4]~q ),
	.Mux11(\rd_adgen|Mux1~1_combout ),
	.k_count_1(\gen_gt256_mk:ctrl|k_count[1]~q ),
	.k_count_3(\gen_gt256_mk:ctrl|k_count[3]~q ),
	.k_count_5(\gen_gt256_mk:ctrl|k_count[5]~q ),
	.k_count_6(\gen_gt256_mk:ctrl|k_count[6]~q ),
	.clk(clk));

fft_asj_fft_tdl_bit_rst_fft_120_4 \gen_dft_2:delay_blk_done2 (
	.global_clock_enable(\global_clock_enable~0_combout ),
	.tdl_arr_11(\gen_dft_2:delay_blk_done|tdl_arr[11]~q ),
	.tdl_arr_19(\gen_dft_2:delay_blk_done2|tdl_arr[19]~q ),
	.clk(clk),
	.reset_n(reset_n));

fft_asj_fft_bfp_ctrl_fft_120 \gen_dft_2:bfpc (
	.source_valid_ctrl_sop(\source_valid_ctrl_sop~1_combout ),
	.stall_reg(\auk_dsp_interface_controller_1|stall_reg~q ),
	.source_stall_int_d(\auk_dsp_atlantic_source_1|source_stall_int_d~q ),
	.global_clock_enable(\global_clock_enable~0_combout ),
	.blk_exp_0(\gen_dft_2:bfpc|blk_exp[0]~q ),
	.blk_exp_1(\gen_dft_2:bfpc|blk_exp[1]~q ),
	.blk_exp_2(\gen_dft_2:bfpc|blk_exp[2]~q ),
	.blk_exp_3(\gen_dft_2:bfpc|blk_exp[3]~q ),
	.blk_exp_4(\gen_dft_2:bfpc|blk_exp[4]~q ),
	.blk_exp_5(\gen_dft_2:bfpc|blk_exp[5]~q ),
	.tdl_arr_4(\gen_radix_2_last_pass:gen_lpp_addr|delay_en|tdl_arr[4]~q ),
	.slb_last_0(\gen_dft_2:bfpc|slb_last[0]~q ),
	.slb_last_1(\gen_dft_2:bfpc|slb_last[1]~q ),
	.slb_last_2(\gen_dft_2:bfpc|slb_last[2]~q ),
	.slb_i_0(\gen_dft_2:bfpdft|gen_cont:bfp_detect|slb_i[0]~q ),
	.slb_i_1(\gen_dft_2:bfpdft|gen_cont:bfp_detect|slb_i[1]~q ),
	.slb_i_2(\gen_dft_2:bfpdft|gen_cont:bfp_detect|slb_i[2]~q ),
	.slb_i_3(\gen_dft_2:bfpdft|gen_cont:bfp_detect|slb_i[3]~q ),
	.Mux2(\gen_dft_2:bfpdft|gen_cont:bfp_detect|Mux2~0_combout ),
	.tdl_arr_11(\gen_dft_2:delay_blk_done|tdl_arr[11]~q ),
	.Mux1(\gen_dft_2:bfpdft|gen_cont:bfp_detect|Mux1~0_combout ),
	.en_slb(\en_slb~q ),
	.GND_port(GND_port),
	.clk(clk),
	.reset_n(reset_n));

fft_asj_fft_tdl_bit_rst_fft_120_3 \gen_dft_2:delay_blk_done (
	.blk_done_int(\gen_gt256_mk:ctrl|blk_done_int~q ),
	.global_clock_enable(\global_clock_enable~0_combout ),
	.tdl_arr_11(\gen_dft_2:delay_blk_done|tdl_arr[11]~q ),
	.blk_done_vec_2(\gen_dft_2:bfpdft|blk_done_vec[2]~q ),
	.tdl_arr_5(\gen_dft_2:delay_blk_done|tdl_arr[5]~q ),
	.clk(clk),
	.reset_n(reset_n));

fft_asj_fft_dft_bfp_fft_120 \gen_dft_2:bfpdft (
	.r_array_out_3_0(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[0][3]~q ),
	.i_array_out_3_0(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[0][3]~q ),
	.r_array_out_3_1(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[1][3]~q ),
	.i_array_out_3_1(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[1][3]~q ),
	.r_array_out_3_2(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[2][3]~q ),
	.i_array_out_3_2(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[2][3]~q ),
	.r_array_out_3_3(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[3][3]~q ),
	.i_array_out_3_3(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[3][3]~q ),
	.r_array_out_4_0(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[0][4]~q ),
	.i_array_out_4_0(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[0][4]~q ),
	.r_array_out_4_1(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[1][4]~q ),
	.i_array_out_4_1(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[1][4]~q ),
	.r_array_out_4_2(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[2][4]~q ),
	.i_array_out_4_2(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[2][4]~q ),
	.r_array_out_4_3(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[3][4]~q ),
	.i_array_out_4_3(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[3][4]~q ),
	.r_array_out_5_0(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[0][5]~q ),
	.i_array_out_5_0(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[0][5]~q ),
	.r_array_out_5_1(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[1][5]~q ),
	.i_array_out_5_1(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[1][5]~q ),
	.r_array_out_5_2(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[2][5]~q ),
	.i_array_out_5_2(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[2][5]~q ),
	.r_array_out_5_3(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[3][5]~q ),
	.i_array_out_5_3(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[3][5]~q ),
	.i_array_out_2_2(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[2][2]~q ),
	.i_array_out_2_1(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[1][2]~q ),
	.i_array_out_2_0(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[0][2]~q ),
	.i_array_out_2_3(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[3][2]~q ),
	.r_array_out_2_2(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[2][2]~q ),
	.r_array_out_2_1(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[1][2]~q ),
	.r_array_out_2_0(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[0][2]~q ),
	.r_array_out_2_3(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[3][2]~q ),
	.ram_in_reg_2_0(\ram_cxb_bfp_data|ram_in_reg[0][2]~q ),
	.ram_in_reg_6_0(\ram_cxb_bfp_data|ram_in_reg[0][6]~q ),
	.ram_in_reg_4_0(\ram_cxb_bfp_data|ram_in_reg[0][4]~q ),
	.ram_in_reg_3_0(\ram_cxb_bfp_data|ram_in_reg[0][3]~q ),
	.ram_in_reg_5_0(\ram_cxb_bfp_data|ram_in_reg[0][5]~q ),
	.ram_in_reg_2_2(\ram_cxb_bfp_data|ram_in_reg[2][2]~q ),
	.ram_in_reg_6_2(\ram_cxb_bfp_data|ram_in_reg[2][6]~q ),
	.ram_in_reg_4_2(\ram_cxb_bfp_data|ram_in_reg[2][4]~q ),
	.ram_in_reg_3_2(\ram_cxb_bfp_data|ram_in_reg[2][3]~q ),
	.ram_in_reg_5_2(\ram_cxb_bfp_data|ram_in_reg[2][5]~q ),
	.ram_in_reg_1_0(\ram_cxb_bfp_data|ram_in_reg[0][1]~q ),
	.ram_in_reg_1_2(\ram_cxb_bfp_data|ram_in_reg[2][1]~q ),
	.ram_in_reg_0_0(\ram_cxb_bfp_data|ram_in_reg[0][0]~q ),
	.ram_in_reg_0_2(\ram_cxb_bfp_data|ram_in_reg[2][0]~q ),
	.ram_in_reg_2_1(\ram_cxb_bfp_data|ram_in_reg[1][2]~q ),
	.ram_in_reg_6_1(\ram_cxb_bfp_data|ram_in_reg[1][6]~q ),
	.ram_in_reg_4_1(\ram_cxb_bfp_data|ram_in_reg[1][4]~q ),
	.ram_in_reg_3_1(\ram_cxb_bfp_data|ram_in_reg[1][3]~q ),
	.ram_in_reg_5_1(\ram_cxb_bfp_data|ram_in_reg[1][5]~q ),
	.ram_in_reg_2_3(\ram_cxb_bfp_data|ram_in_reg[3][2]~q ),
	.ram_in_reg_6_3(\ram_cxb_bfp_data|ram_in_reg[3][6]~q ),
	.ram_in_reg_4_3(\ram_cxb_bfp_data|ram_in_reg[3][4]~q ),
	.ram_in_reg_3_3(\ram_cxb_bfp_data|ram_in_reg[3][3]~q ),
	.ram_in_reg_5_3(\ram_cxb_bfp_data|ram_in_reg[3][5]~q ),
	.ram_in_reg_1_1(\ram_cxb_bfp_data|ram_in_reg[1][1]~q ),
	.ram_in_reg_1_3(\ram_cxb_bfp_data|ram_in_reg[3][1]~q ),
	.ram_in_reg_0_1(\ram_cxb_bfp_data|ram_in_reg[1][0]~q ),
	.ram_in_reg_0_3(\ram_cxb_bfp_data|ram_in_reg[3][0]~q ),
	.ram_in_reg_7_0(\ram_cxb_bfp_data|ram_in_reg[0][7]~q ),
	.ram_in_reg_7_2(\ram_cxb_bfp_data|ram_in_reg[2][7]~q ),
	.ram_in_reg_7_1(\ram_cxb_bfp_data|ram_in_reg[1][7]~q ),
	.ram_in_reg_7_3(\ram_cxb_bfp_data|ram_in_reg[3][7]~q ),
	.ram_in_reg_7_4(\ram_cxb_bfp_data|ram_in_reg[4][7]~q ),
	.ram_in_reg_3_4(\ram_cxb_bfp_data|ram_in_reg[4][3]~q ),
	.ram_in_reg_5_4(\ram_cxb_bfp_data|ram_in_reg[4][5]~q ),
	.ram_in_reg_4_4(\ram_cxb_bfp_data|ram_in_reg[4][4]~q ),
	.ram_in_reg_6_4(\ram_cxb_bfp_data|ram_in_reg[4][6]~q ),
	.ram_in_reg_7_6(\ram_cxb_bfp_data|ram_in_reg[6][7]~q ),
	.ram_in_reg_3_6(\ram_cxb_bfp_data|ram_in_reg[6][3]~q ),
	.ram_in_reg_5_6(\ram_cxb_bfp_data|ram_in_reg[6][5]~q ),
	.ram_in_reg_4_6(\ram_cxb_bfp_data|ram_in_reg[6][4]~q ),
	.ram_in_reg_6_6(\ram_cxb_bfp_data|ram_in_reg[6][6]~q ),
	.ram_in_reg_2_4(\ram_cxb_bfp_data|ram_in_reg[4][2]~q ),
	.ram_in_reg_2_6(\ram_cxb_bfp_data|ram_in_reg[6][2]~q ),
	.ram_in_reg_1_4(\ram_cxb_bfp_data|ram_in_reg[4][1]~q ),
	.ram_in_reg_1_6(\ram_cxb_bfp_data|ram_in_reg[6][1]~q ),
	.ram_in_reg_0_4(\ram_cxb_bfp_data|ram_in_reg[4][0]~q ),
	.ram_in_reg_0_6(\ram_cxb_bfp_data|ram_in_reg[6][0]~q ),
	.ram_in_reg_7_5(\ram_cxb_bfp_data|ram_in_reg[5][7]~q ),
	.ram_in_reg_3_5(\ram_cxb_bfp_data|ram_in_reg[5][3]~q ),
	.ram_in_reg_5_5(\ram_cxb_bfp_data|ram_in_reg[5][5]~q ),
	.ram_in_reg_4_5(\ram_cxb_bfp_data|ram_in_reg[5][4]~q ),
	.ram_in_reg_6_5(\ram_cxb_bfp_data|ram_in_reg[5][6]~q ),
	.ram_in_reg_3_7(\ram_cxb_bfp_data|ram_in_reg[7][3]~q ),
	.ram_in_reg_7_7(\ram_cxb_bfp_data|ram_in_reg[7][7]~q ),
	.ram_in_reg_5_7(\ram_cxb_bfp_data|ram_in_reg[7][5]~q ),
	.ram_in_reg_4_7(\ram_cxb_bfp_data|ram_in_reg[7][4]~q ),
	.ram_in_reg_6_7(\ram_cxb_bfp_data|ram_in_reg[7][6]~q ),
	.ram_in_reg_2_5(\ram_cxb_bfp_data|ram_in_reg[5][2]~q ),
	.ram_in_reg_2_7(\ram_cxb_bfp_data|ram_in_reg[7][2]~q ),
	.ram_in_reg_1_5(\ram_cxb_bfp_data|ram_in_reg[5][1]~q ),
	.ram_in_reg_1_7(\ram_cxb_bfp_data|ram_in_reg[7][1]~q ),
	.ram_in_reg_0_5(\ram_cxb_bfp_data|ram_in_reg[5][0]~q ),
	.ram_in_reg_0_7(\ram_cxb_bfp_data|ram_in_reg[7][0]~q ),
	.global_clock_enable(\global_clock_enable~0_combout ),
	.slb_last_0(\gen_dft_2:bfpc|slb_last[0]~q ),
	.slb_last_1(\gen_dft_2:bfpc|slb_last[1]~q ),
	.slb_last_2(\gen_dft_2:bfpc|slb_last[2]~q ),
	.next_block(\writer|next_block~q ),
	.slb_i_0(\gen_dft_2:bfpdft|gen_cont:bfp_detect|slb_i[0]~q ),
	.slb_i_1(\gen_dft_2:bfpdft|gen_cont:bfp_detect|slb_i[1]~q ),
	.slb_i_2(\gen_dft_2:bfpdft|gen_cont:bfp_detect|slb_i[2]~q ),
	.slb_i_3(\gen_dft_2:bfpdft|gen_cont:bfp_detect|slb_i[3]~q ),
	.Mux2(\gen_dft_2:bfpdft|gen_cont:bfp_detect|Mux2~0_combout ),
	.Mux1(\gen_dft_2:bfpdft|gen_cont:bfp_detect|Mux1~0_combout ),
	.tdl_arr_4(\gen_dft_2:bfpdft|gen_cont:delay_next_blk|tdl_arr[4]~q ),
	.tdl_arr_3(\gen_dft_2:bfpdft|gen_cont:delay_next_blk|tdl_arr[3]~q ),
	.r_array_out_7_0(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[0][7]~q ),
	.i_array_out_7_0(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[0][7]~q ),
	.r_array_out_7_1(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[1][7]~q ),
	.i_array_out_7_1(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[1][7]~q ),
	.r_array_out_7_2(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[2][7]~q ),
	.i_array_out_7_2(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[2][7]~q ),
	.r_array_out_7_3(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[3][7]~q ),
	.i_array_out_7_3(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[3][7]~q ),
	.blk_done_vec_2(\gen_dft_2:bfpdft|blk_done_vec[2]~q ),
	.r_array_out_6_0(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[0][6]~q ),
	.i_array_out_6_0(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[0][6]~q ),
	.r_array_out_6_1(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[1][6]~q ),
	.i_array_out_6_1(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[1][6]~q ),
	.r_array_out_6_2(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[2][6]~q ),
	.i_array_out_6_2(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[2][6]~q ),
	.r_array_out_6_3(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[3][6]~q ),
	.i_array_out_6_3(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[3][6]~q ),
	.i_array_out_1_2(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[2][1]~q ),
	.i_array_out_1_1(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[1][1]~q ),
	.i_array_out_1_0(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[0][1]~q ),
	.i_array_out_1_3(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[3][1]~q ),
	.i_array_out_0_2(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[2][0]~q ),
	.i_array_out_0_1(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[1][0]~q ),
	.i_array_out_0_0(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[0][0]~q ),
	.i_array_out_0_3(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[3][0]~q ),
	.r_array_out_1_2(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[2][1]~q ),
	.r_array_out_1_1(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[1][1]~q ),
	.r_array_out_1_0(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[0][1]~q ),
	.r_array_out_1_3(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[3][1]~q ),
	.r_array_out_0_2(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[2][0]~q ),
	.r_array_out_0_1(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[1][0]~q ),
	.r_array_out_0_0(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[0][0]~q ),
	.r_array_out_0_3(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[3][0]~q ),
	.tdl_arr_5(\gen_dft_2:delay_blk_done|tdl_arr[5]~q ),
	.tdl_arr_51(\delay_ctrl_np|tdl_arr[5]~q ),
	.twiddle_data000(\twiddle_data[0][0][0]~q ),
	.twiddle_data001(\twiddle_data[0][0][1]~q ),
	.twiddle_data002(\twiddle_data[0][0][2]~q ),
	.twiddle_data003(\twiddle_data[0][0][3]~q ),
	.twiddle_data004(\twiddle_data[0][0][4]~q ),
	.twiddle_data005(\twiddle_data[0][0][5]~q ),
	.twiddle_data006(\twiddle_data[0][0][6]~q ),
	.twiddle_data007(\twiddle_data[0][0][7]~q ),
	.twiddle_data010(\twiddle_data[0][1][0]~q ),
	.twiddle_data011(\twiddle_data[0][1][1]~q ),
	.twiddle_data012(\twiddle_data[0][1][2]~q ),
	.twiddle_data013(\twiddle_data[0][1][3]~q ),
	.twiddle_data014(\twiddle_data[0][1][4]~q ),
	.twiddle_data015(\twiddle_data[0][1][5]~q ),
	.twiddle_data016(\twiddle_data[0][1][6]~q ),
	.twiddle_data017(\twiddle_data[0][1][7]~q ),
	.twiddle_data100(\twiddle_data[1][0][0]~q ),
	.twiddle_data101(\twiddle_data[1][0][1]~q ),
	.twiddle_data102(\twiddle_data[1][0][2]~q ),
	.twiddle_data103(\twiddle_data[1][0][3]~q ),
	.twiddle_data104(\twiddle_data[1][0][4]~q ),
	.twiddle_data105(\twiddle_data[1][0][5]~q ),
	.twiddle_data106(\twiddle_data[1][0][6]~q ),
	.twiddle_data107(\twiddle_data[1][0][7]~q ),
	.twiddle_data110(\twiddle_data[1][1][0]~q ),
	.twiddle_data111(\twiddle_data[1][1][1]~q ),
	.twiddle_data112(\twiddle_data[1][1][2]~q ),
	.twiddle_data113(\twiddle_data[1][1][3]~q ),
	.twiddle_data114(\twiddle_data[1][1][4]~q ),
	.twiddle_data115(\twiddle_data[1][1][5]~q ),
	.twiddle_data116(\twiddle_data[1][1][6]~q ),
	.twiddle_data117(\twiddle_data[1][1][7]~q ),
	.twiddle_data200(\twiddle_data[2][0][0]~q ),
	.twiddle_data201(\twiddle_data[2][0][1]~q ),
	.twiddle_data202(\twiddle_data[2][0][2]~q ),
	.twiddle_data203(\twiddle_data[2][0][3]~q ),
	.twiddle_data204(\twiddle_data[2][0][4]~q ),
	.twiddle_data205(\twiddle_data[2][0][5]~q ),
	.twiddle_data206(\twiddle_data[2][0][6]~q ),
	.twiddle_data207(\twiddle_data[2][0][7]~q ),
	.twiddle_data210(\twiddle_data[2][1][0]~q ),
	.twiddle_data211(\twiddle_data[2][1][1]~q ),
	.twiddle_data212(\twiddle_data[2][1][2]~q ),
	.twiddle_data213(\twiddle_data[2][1][3]~q ),
	.twiddle_data214(\twiddle_data[2][1][4]~q ),
	.twiddle_data215(\twiddle_data[2][1][5]~q ),
	.twiddle_data216(\twiddle_data[2][1][6]~q ),
	.twiddle_data217(\twiddle_data[2][1][7]~q ),
	.next_pass_vec_2(\gen_dft_2:bfpdft|next_pass_vec[2]~q ),
	.clk(clk),
	.reset_n(reset_n));

fft_asj_fft_cxb_data_r_fft_120 ram_cxb_bfp_data(
	.ram_in_reg_2_0(\ram_cxb_bfp_data|ram_in_reg[0][2]~q ),
	.ram_in_reg_6_0(\ram_cxb_bfp_data|ram_in_reg[0][6]~q ),
	.ram_in_reg_4_0(\ram_cxb_bfp_data|ram_in_reg[0][4]~q ),
	.ram_in_reg_3_0(\ram_cxb_bfp_data|ram_in_reg[0][3]~q ),
	.ram_in_reg_5_0(\ram_cxb_bfp_data|ram_in_reg[0][5]~q ),
	.ram_in_reg_2_2(\ram_cxb_bfp_data|ram_in_reg[2][2]~q ),
	.ram_in_reg_6_2(\ram_cxb_bfp_data|ram_in_reg[2][6]~q ),
	.ram_in_reg_4_2(\ram_cxb_bfp_data|ram_in_reg[2][4]~q ),
	.ram_in_reg_3_2(\ram_cxb_bfp_data|ram_in_reg[2][3]~q ),
	.ram_in_reg_5_2(\ram_cxb_bfp_data|ram_in_reg[2][5]~q ),
	.ram_in_reg_1_0(\ram_cxb_bfp_data|ram_in_reg[0][1]~q ),
	.ram_in_reg_1_2(\ram_cxb_bfp_data|ram_in_reg[2][1]~q ),
	.ram_in_reg_0_0(\ram_cxb_bfp_data|ram_in_reg[0][0]~q ),
	.ram_in_reg_0_2(\ram_cxb_bfp_data|ram_in_reg[2][0]~q ),
	.ram_in_reg_2_1(\ram_cxb_bfp_data|ram_in_reg[1][2]~q ),
	.ram_in_reg_6_1(\ram_cxb_bfp_data|ram_in_reg[1][6]~q ),
	.ram_in_reg_4_1(\ram_cxb_bfp_data|ram_in_reg[1][4]~q ),
	.ram_in_reg_3_1(\ram_cxb_bfp_data|ram_in_reg[1][3]~q ),
	.ram_in_reg_5_1(\ram_cxb_bfp_data|ram_in_reg[1][5]~q ),
	.ram_in_reg_2_3(\ram_cxb_bfp_data|ram_in_reg[3][2]~q ),
	.ram_in_reg_6_3(\ram_cxb_bfp_data|ram_in_reg[3][6]~q ),
	.ram_in_reg_4_3(\ram_cxb_bfp_data|ram_in_reg[3][4]~q ),
	.ram_in_reg_3_3(\ram_cxb_bfp_data|ram_in_reg[3][3]~q ),
	.ram_in_reg_5_3(\ram_cxb_bfp_data|ram_in_reg[3][5]~q ),
	.ram_in_reg_1_1(\ram_cxb_bfp_data|ram_in_reg[1][1]~q ),
	.ram_in_reg_1_3(\ram_cxb_bfp_data|ram_in_reg[3][1]~q ),
	.ram_in_reg_0_1(\ram_cxb_bfp_data|ram_in_reg[1][0]~q ),
	.ram_in_reg_0_3(\ram_cxb_bfp_data|ram_in_reg[3][0]~q ),
	.ram_in_reg_7_0(\ram_cxb_bfp_data|ram_in_reg[0][7]~q ),
	.ram_in_reg_7_2(\ram_cxb_bfp_data|ram_in_reg[2][7]~q ),
	.ram_in_reg_7_1(\ram_cxb_bfp_data|ram_in_reg[1][7]~q ),
	.ram_in_reg_7_3(\ram_cxb_bfp_data|ram_in_reg[3][7]~q ),
	.ram_in_reg_7_4(\ram_cxb_bfp_data|ram_in_reg[4][7]~q ),
	.ram_in_reg_3_4(\ram_cxb_bfp_data|ram_in_reg[4][3]~q ),
	.ram_in_reg_5_4(\ram_cxb_bfp_data|ram_in_reg[4][5]~q ),
	.ram_in_reg_4_4(\ram_cxb_bfp_data|ram_in_reg[4][4]~q ),
	.ram_in_reg_6_4(\ram_cxb_bfp_data|ram_in_reg[4][6]~q ),
	.ram_in_reg_7_6(\ram_cxb_bfp_data|ram_in_reg[6][7]~q ),
	.ram_in_reg_3_6(\ram_cxb_bfp_data|ram_in_reg[6][3]~q ),
	.ram_in_reg_5_6(\ram_cxb_bfp_data|ram_in_reg[6][5]~q ),
	.ram_in_reg_4_6(\ram_cxb_bfp_data|ram_in_reg[6][4]~q ),
	.ram_in_reg_6_6(\ram_cxb_bfp_data|ram_in_reg[6][6]~q ),
	.ram_in_reg_2_4(\ram_cxb_bfp_data|ram_in_reg[4][2]~q ),
	.ram_in_reg_2_6(\ram_cxb_bfp_data|ram_in_reg[6][2]~q ),
	.ram_in_reg_1_4(\ram_cxb_bfp_data|ram_in_reg[4][1]~q ),
	.ram_in_reg_1_6(\ram_cxb_bfp_data|ram_in_reg[6][1]~q ),
	.ram_in_reg_0_4(\ram_cxb_bfp_data|ram_in_reg[4][0]~q ),
	.ram_in_reg_0_6(\ram_cxb_bfp_data|ram_in_reg[6][0]~q ),
	.ram_in_reg_7_5(\ram_cxb_bfp_data|ram_in_reg[5][7]~q ),
	.ram_in_reg_3_5(\ram_cxb_bfp_data|ram_in_reg[5][3]~q ),
	.ram_in_reg_5_5(\ram_cxb_bfp_data|ram_in_reg[5][5]~q ),
	.ram_in_reg_4_5(\ram_cxb_bfp_data|ram_in_reg[5][4]~q ),
	.ram_in_reg_6_5(\ram_cxb_bfp_data|ram_in_reg[5][6]~q ),
	.ram_in_reg_3_7(\ram_cxb_bfp_data|ram_in_reg[7][3]~q ),
	.ram_in_reg_7_7(\ram_cxb_bfp_data|ram_in_reg[7][7]~q ),
	.ram_in_reg_5_7(\ram_cxb_bfp_data|ram_in_reg[7][5]~q ),
	.ram_in_reg_4_7(\ram_cxb_bfp_data|ram_in_reg[7][4]~q ),
	.ram_in_reg_6_7(\ram_cxb_bfp_data|ram_in_reg[7][6]~q ),
	.ram_in_reg_2_5(\ram_cxb_bfp_data|ram_in_reg[5][2]~q ),
	.ram_in_reg_2_7(\ram_cxb_bfp_data|ram_in_reg[7][2]~q ),
	.ram_in_reg_1_5(\ram_cxb_bfp_data|ram_in_reg[5][1]~q ),
	.ram_in_reg_1_7(\ram_cxb_bfp_data|ram_in_reg[7][1]~q ),
	.ram_in_reg_0_5(\ram_cxb_bfp_data|ram_in_reg[5][0]~q ),
	.ram_in_reg_0_7(\ram_cxb_bfp_data|ram_in_reg[7][0]~q ),
	.global_clock_enable(\global_clock_enable~0_combout ),
	.ram_data_out0_10(\ccc|ram_data_out0[10]~q ),
	.ram_data_out1_10(\ccc|ram_data_out1[10]~q ),
	.sw_r_tdl_0_4(\sw_r_tdl[4][0]~q ),
	.ram_data_out2_10(\ccc|ram_data_out2[10]~q ),
	.ram_data_out3_10(\ccc|ram_data_out3[10]~q ),
	.sw_r_tdl_1_4(\sw_r_tdl[4][1]~q ),
	.ram_data_out0_14(\ccc|ram_data_out0[14]~q ),
	.ram_data_out1_14(\ccc|ram_data_out1[14]~q ),
	.ram_data_out2_14(\ccc|ram_data_out2[14]~q ),
	.ram_data_out3_14(\ccc|ram_data_out3[14]~q ),
	.ram_data_out0_12(\ccc|ram_data_out0[12]~q ),
	.ram_data_out1_12(\ccc|ram_data_out1[12]~q ),
	.ram_data_out2_12(\ccc|ram_data_out2[12]~q ),
	.ram_data_out3_12(\ccc|ram_data_out3[12]~q ),
	.ram_data_out0_11(\ccc|ram_data_out0[11]~q ),
	.ram_data_out1_11(\ccc|ram_data_out1[11]~q ),
	.ram_data_out2_11(\ccc|ram_data_out2[11]~q ),
	.ram_data_out3_11(\ccc|ram_data_out3[11]~q ),
	.ram_data_out0_13(\ccc|ram_data_out0[13]~q ),
	.ram_data_out1_13(\ccc|ram_data_out1[13]~q ),
	.ram_data_out2_13(\ccc|ram_data_out2[13]~q ),
	.ram_data_out3_13(\ccc|ram_data_out3[13]~q ),
	.ram_data_out0_9(\ccc|ram_data_out0[9]~q ),
	.ram_data_out1_9(\ccc|ram_data_out1[9]~q ),
	.ram_data_out2_9(\ccc|ram_data_out2[9]~q ),
	.ram_data_out3_9(\ccc|ram_data_out3[9]~q ),
	.ram_data_out0_8(\ccc|ram_data_out0[8]~q ),
	.ram_data_out1_8(\ccc|ram_data_out1[8]~q ),
	.ram_data_out2_8(\ccc|ram_data_out2[8]~q ),
	.ram_data_out3_8(\ccc|ram_data_out3[8]~q ),
	.ram_data_out0_15(\ccc|ram_data_out0[15]~q ),
	.ram_data_out1_15(\ccc|ram_data_out1[15]~q ),
	.ram_data_out2_15(\ccc|ram_data_out2[15]~q ),
	.ram_data_out3_15(\ccc|ram_data_out3[15]~q ),
	.ram_data_out0_7(\ccc|ram_data_out0[7]~q ),
	.ram_data_out1_7(\ccc|ram_data_out1[7]~q ),
	.ram_data_out2_7(\ccc|ram_data_out2[7]~q ),
	.ram_data_out3_7(\ccc|ram_data_out3[7]~q ),
	.ram_data_out0_3(\ccc|ram_data_out0[3]~q ),
	.ram_data_out1_3(\ccc|ram_data_out1[3]~q ),
	.ram_data_out2_3(\ccc|ram_data_out2[3]~q ),
	.ram_data_out3_3(\ccc|ram_data_out3[3]~q ),
	.ram_data_out0_5(\ccc|ram_data_out0[5]~q ),
	.ram_data_out1_5(\ccc|ram_data_out1[5]~q ),
	.ram_data_out2_5(\ccc|ram_data_out2[5]~q ),
	.ram_data_out3_5(\ccc|ram_data_out3[5]~q ),
	.ram_data_out0_4(\ccc|ram_data_out0[4]~q ),
	.ram_data_out1_4(\ccc|ram_data_out1[4]~q ),
	.ram_data_out2_4(\ccc|ram_data_out2[4]~q ),
	.ram_data_out3_4(\ccc|ram_data_out3[4]~q ),
	.ram_data_out0_6(\ccc|ram_data_out0[6]~q ),
	.ram_data_out1_6(\ccc|ram_data_out1[6]~q ),
	.ram_data_out2_6(\ccc|ram_data_out2[6]~q ),
	.ram_data_out3_6(\ccc|ram_data_out3[6]~q ),
	.ram_data_out0_2(\ccc|ram_data_out0[2]~q ),
	.ram_data_out1_2(\ccc|ram_data_out1[2]~q ),
	.ram_data_out2_2(\ccc|ram_data_out2[2]~q ),
	.ram_data_out3_2(\ccc|ram_data_out3[2]~q ),
	.ram_data_out0_1(\ccc|ram_data_out0[1]~q ),
	.ram_data_out1_1(\ccc|ram_data_out1[1]~q ),
	.ram_data_out2_1(\ccc|ram_data_out2[1]~q ),
	.ram_data_out3_1(\ccc|ram_data_out3[1]~q ),
	.ram_data_out0_0(\ccc|ram_data_out0[0]~q ),
	.ram_data_out1_0(\ccc|ram_data_out1[0]~q ),
	.ram_data_out2_0(\ccc|ram_data_out2[0]~q ),
	.ram_data_out3_0(\ccc|ram_data_out3[0]~q ),
	.clk(clk));

fft_asj_fft_cxb_data_fft_120 ram_cxb_wr_data(
	.ram_in_reg_1_6(\ram_cxb_wr_data|ram_in_reg[6][1]~q ),
	.ram_in_reg_1_5(\ram_cxb_wr_data|ram_in_reg[5][1]~q ),
	.ram_in_reg_1_4(\ram_cxb_wr_data|ram_in_reg[4][1]~q ),
	.ram_in_reg_1_7(\ram_cxb_wr_data|ram_in_reg[7][1]~q ),
	.ram_in_reg_0_6(\ram_cxb_wr_data|ram_in_reg[6][0]~q ),
	.ram_in_reg_0_5(\ram_cxb_wr_data|ram_in_reg[5][0]~q ),
	.ram_in_reg_0_4(\ram_cxb_wr_data|ram_in_reg[4][0]~q ),
	.ram_in_reg_0_7(\ram_cxb_wr_data|ram_in_reg[7][0]~q ),
	.ram_in_reg_7_6(\ram_cxb_wr_data|ram_in_reg[6][7]~q ),
	.ram_in_reg_7_5(\ram_cxb_wr_data|ram_in_reg[5][7]~q ),
	.ram_in_reg_7_4(\ram_cxb_wr_data|ram_in_reg[4][7]~q ),
	.ram_in_reg_7_7(\ram_cxb_wr_data|ram_in_reg[7][7]~q ),
	.ram_in_reg_6_6(\ram_cxb_wr_data|ram_in_reg[6][6]~q ),
	.ram_in_reg_6_5(\ram_cxb_wr_data|ram_in_reg[5][6]~q ),
	.ram_in_reg_6_4(\ram_cxb_wr_data|ram_in_reg[4][6]~q ),
	.ram_in_reg_6_7(\ram_cxb_wr_data|ram_in_reg[7][6]~q ),
	.ram_in_reg_5_6(\ram_cxb_wr_data|ram_in_reg[6][5]~q ),
	.ram_in_reg_5_5(\ram_cxb_wr_data|ram_in_reg[5][5]~q ),
	.ram_in_reg_5_4(\ram_cxb_wr_data|ram_in_reg[4][5]~q ),
	.ram_in_reg_5_7(\ram_cxb_wr_data|ram_in_reg[7][5]~q ),
	.ram_in_reg_4_6(\ram_cxb_wr_data|ram_in_reg[6][4]~q ),
	.ram_in_reg_4_5(\ram_cxb_wr_data|ram_in_reg[5][4]~q ),
	.ram_in_reg_4_4(\ram_cxb_wr_data|ram_in_reg[4][4]~q ),
	.ram_in_reg_4_7(\ram_cxb_wr_data|ram_in_reg[7][4]~q ),
	.ram_in_reg_3_6(\ram_cxb_wr_data|ram_in_reg[6][3]~q ),
	.ram_in_reg_3_5(\ram_cxb_wr_data|ram_in_reg[5][3]~q ),
	.ram_in_reg_3_4(\ram_cxb_wr_data|ram_in_reg[4][3]~q ),
	.ram_in_reg_3_7(\ram_cxb_wr_data|ram_in_reg[7][3]~q ),
	.ram_in_reg_2_6(\ram_cxb_wr_data|ram_in_reg[6][2]~q ),
	.ram_in_reg_2_5(\ram_cxb_wr_data|ram_in_reg[5][2]~q ),
	.ram_in_reg_2_4(\ram_cxb_wr_data|ram_in_reg[4][2]~q ),
	.ram_in_reg_2_7(\ram_cxb_wr_data|ram_in_reg[7][2]~q ),
	.ram_in_reg_1_2(\ram_cxb_wr_data|ram_in_reg[2][1]~q ),
	.ram_in_reg_1_1(\ram_cxb_wr_data|ram_in_reg[1][1]~q ),
	.ram_in_reg_1_0(\ram_cxb_wr_data|ram_in_reg[0][1]~q ),
	.ram_in_reg_1_3(\ram_cxb_wr_data|ram_in_reg[3][1]~q ),
	.ram_in_reg_0_2(\ram_cxb_wr_data|ram_in_reg[2][0]~q ),
	.ram_in_reg_0_1(\ram_cxb_wr_data|ram_in_reg[1][0]~q ),
	.ram_in_reg_0_0(\ram_cxb_wr_data|ram_in_reg[0][0]~q ),
	.ram_in_reg_0_3(\ram_cxb_wr_data|ram_in_reg[3][0]~q ),
	.ram_in_reg_7_2(\ram_cxb_wr_data|ram_in_reg[2][7]~q ),
	.ram_in_reg_7_1(\ram_cxb_wr_data|ram_in_reg[1][7]~q ),
	.ram_in_reg_7_0(\ram_cxb_wr_data|ram_in_reg[0][7]~q ),
	.ram_in_reg_7_3(\ram_cxb_wr_data|ram_in_reg[3][7]~q ),
	.ram_in_reg_6_2(\ram_cxb_wr_data|ram_in_reg[2][6]~q ),
	.ram_in_reg_6_1(\ram_cxb_wr_data|ram_in_reg[1][6]~q ),
	.ram_in_reg_6_0(\ram_cxb_wr_data|ram_in_reg[0][6]~q ),
	.ram_in_reg_6_3(\ram_cxb_wr_data|ram_in_reg[3][6]~q ),
	.ram_in_reg_5_2(\ram_cxb_wr_data|ram_in_reg[2][5]~q ),
	.ram_in_reg_5_1(\ram_cxb_wr_data|ram_in_reg[1][5]~q ),
	.ram_in_reg_5_0(\ram_cxb_wr_data|ram_in_reg[0][5]~q ),
	.ram_in_reg_5_3(\ram_cxb_wr_data|ram_in_reg[3][5]~q ),
	.ram_in_reg_4_2(\ram_cxb_wr_data|ram_in_reg[2][4]~q ),
	.ram_in_reg_4_1(\ram_cxb_wr_data|ram_in_reg[1][4]~q ),
	.ram_in_reg_4_0(\ram_cxb_wr_data|ram_in_reg[0][4]~q ),
	.ram_in_reg_4_3(\ram_cxb_wr_data|ram_in_reg[3][4]~q ),
	.ram_in_reg_3_2(\ram_cxb_wr_data|ram_in_reg[2][3]~q ),
	.ram_in_reg_3_1(\ram_cxb_wr_data|ram_in_reg[1][3]~q ),
	.ram_in_reg_3_0(\ram_cxb_wr_data|ram_in_reg[0][3]~q ),
	.ram_in_reg_3_3(\ram_cxb_wr_data|ram_in_reg[3][3]~q ),
	.ram_in_reg_2_2(\ram_cxb_wr_data|ram_in_reg[2][2]~q ),
	.ram_in_reg_2_1(\ram_cxb_wr_data|ram_in_reg[1][2]~q ),
	.ram_in_reg_2_0(\ram_cxb_wr_data|ram_in_reg[0][2]~q ),
	.ram_in_reg_2_3(\ram_cxb_wr_data|ram_in_reg[3][2]~q ),
	.r_array_out_3_0(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[0][3]~q ),
	.i_array_out_3_0(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[0][3]~q ),
	.r_array_out_3_1(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[1][3]~q ),
	.i_array_out_3_1(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[1][3]~q ),
	.r_array_out_3_2(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[2][3]~q ),
	.i_array_out_3_2(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[2][3]~q ),
	.r_array_out_3_3(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[3][3]~q ),
	.i_array_out_3_3(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[3][3]~q ),
	.r_array_out_4_0(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[0][4]~q ),
	.i_array_out_4_0(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[0][4]~q ),
	.r_array_out_4_1(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[1][4]~q ),
	.i_array_out_4_1(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[1][4]~q ),
	.r_array_out_4_2(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[2][4]~q ),
	.i_array_out_4_2(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[2][4]~q ),
	.r_array_out_4_3(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[3][4]~q ),
	.i_array_out_4_3(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[3][4]~q ),
	.r_array_out_5_0(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[0][5]~q ),
	.i_array_out_5_0(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[0][5]~q ),
	.r_array_out_5_1(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[1][5]~q ),
	.i_array_out_5_1(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[1][5]~q ),
	.r_array_out_5_2(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[2][5]~q ),
	.i_array_out_5_2(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[2][5]~q ),
	.r_array_out_5_3(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[3][5]~q ),
	.i_array_out_5_3(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[3][5]~q ),
	.i_array_out_2_2(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[2][2]~q ),
	.i_array_out_2_1(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[1][2]~q ),
	.i_array_out_2_0(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[0][2]~q ),
	.i_array_out_2_3(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[3][2]~q ),
	.r_array_out_2_2(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[2][2]~q ),
	.r_array_out_2_1(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[1][2]~q ),
	.r_array_out_2_0(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[0][2]~q ),
	.r_array_out_2_3(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[3][2]~q ),
	.global_clock_enable(\global_clock_enable~0_combout ),
	.r_array_out_7_0(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[0][7]~q ),
	.i_array_out_7_0(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[0][7]~q ),
	.r_array_out_7_1(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[1][7]~q ),
	.i_array_out_7_1(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[1][7]~q ),
	.r_array_out_7_2(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[2][7]~q ),
	.i_array_out_7_2(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[2][7]~q ),
	.r_array_out_7_3(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[3][7]~q ),
	.i_array_out_7_3(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[3][7]~q ),
	.r_array_out_6_0(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[0][6]~q ),
	.i_array_out_6_0(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[0][6]~q ),
	.r_array_out_6_1(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[1][6]~q ),
	.i_array_out_6_1(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[1][6]~q ),
	.r_array_out_6_2(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[2][6]~q ),
	.i_array_out_6_2(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[2][6]~q ),
	.r_array_out_6_3(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[3][6]~q ),
	.i_array_out_6_3(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[3][6]~q ),
	.i_array_out_1_2(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[2][1]~q ),
	.i_array_out_1_1(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[1][1]~q ),
	.swa_tdl_0_0(\gen_wrsw_2:get_wr_swtiches|swa_tdl[0][0]~q ),
	.i_array_out_1_0(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[0][1]~q ),
	.i_array_out_1_3(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[3][1]~q ),
	.swa_tdl_1_0(\gen_wrsw_2:get_wr_swtiches|swa_tdl[0][1]~q ),
	.i_array_out_0_2(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[2][0]~q ),
	.i_array_out_0_1(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[1][0]~q ),
	.i_array_out_0_0(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[0][0]~q ),
	.i_array_out_0_3(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|i_array_out[3][0]~q ),
	.r_array_out_1_2(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[2][1]~q ),
	.r_array_out_1_1(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[1][1]~q ),
	.r_array_out_1_0(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[0][1]~q ),
	.r_array_out_1_3(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[3][1]~q ),
	.r_array_out_0_2(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[2][0]~q ),
	.r_array_out_0_1(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[1][0]~q ),
	.r_array_out_0_0(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[0][0]~q ),
	.r_array_out_0_3(\gen_dft_2:bfpdft|gen_cont:bfp_scale_1pt|r_array_out[3][0]~q ),
	.clk(clk));

fft_asj_fft_cxb_addr_fft_120_1 \gen_wrsw_2:ram_cxb_wr (
	.global_clock_enable(\global_clock_enable~0_combout ),
	.ram_in_reg_0_0(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[0][0]~q ),
	.ram_in_reg_1_2(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[2][1]~q ),
	.ram_in_reg_2_0(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[0][2]~q ),
	.ram_in_reg_3_2(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[2][3]~q ),
	.ram_in_reg_4_0(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[0][4]~q ),
	.ram_in_reg_5_2(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[2][5]~q ),
	.ram_in_reg_6_0(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[0][6]~q ),
	.ram_in_reg_0_1(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[1][0]~q ),
	.ram_in_reg_1_1(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[1][1]~q ),
	.ram_in_reg_2_1(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[1][2]~q ),
	.ram_in_reg_3_1(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[1][3]~q ),
	.ram_in_reg_4_1(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[1][4]~q ),
	.ram_in_reg_5_1(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[1][5]~q ),
	.ram_in_reg_1_0(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[0][1]~q ),
	.ram_in_reg_3_0(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[0][3]~q ),
	.ram_in_reg_5_0(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[0][5]~q ),
	.ram_in_reg_1_3(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[3][1]~q ),
	.ram_in_reg_3_3(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[3][3]~q ),
	.ram_in_reg_5_3(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[3][5]~q ),
	.swa_tdl_0_0(\gen_wrsw_2:get_wr_swtiches|swa_tdl[0][0]~q ),
	.swa_tdl_1_0(\gen_wrsw_2:get_wr_swtiches|swa_tdl[0][1]~q ),
	.sw_3_in({\gen_wrsw_2:wr_adgen|rd_addr_d[6]~q ,\gen_wrsw_2:wr_adgen|rd_addr_d[5]~q ,\gen_wrsw_2:wr_adgen|rd_addr_d[4]~q ,\gen_wrsw_2:wr_adgen|rd_addr_d[3]~q ,\gen_wrsw_2:wr_adgen|rd_addr_d[2]~q ,\gen_wrsw_2:wr_adgen|rd_addr_d[1]~q ,\gen_wrsw_2:wr_adgen|rd_addr_d[0]~q }),
	.sw_2_in({gnd,gnd,\gen_wrsw_2:wr_adgen|rd_addr_c[4]~q ,gnd,\gen_wrsw_2:wr_adgen|rd_addr_c[2]~q ,gnd,\gen_wrsw_2:wr_adgen|rd_addr_c[0]~q }),
	.sw_1_in({gnd,\gen_wrsw_2:wr_adgen|rd_addr_b[5]~q ,gnd,\gen_wrsw_2:wr_adgen|rd_addr_b[3]~q ,gnd,\gen_wrsw_2:wr_adgen|rd_addr_b[1]~q ,gnd}),
	.clk(clk));

fft_asj_fft_dataadgen_fft_120 \gen_wrsw_2:wr_adgen (
	.global_clock_enable(\global_clock_enable~0_combout ),
	.rd_addr_d_0(\gen_wrsw_2:wr_adgen|rd_addr_d[0]~q ),
	.rd_addr_c_0(\gen_wrsw_2:wr_adgen|rd_addr_c[0]~q ),
	.rd_addr_d_1(\gen_wrsw_2:wr_adgen|rd_addr_d[1]~q ),
	.rd_addr_b_1(\gen_wrsw_2:wr_adgen|rd_addr_b[1]~q ),
	.rd_addr_d_2(\gen_wrsw_2:wr_adgen|rd_addr_d[2]~q ),
	.rd_addr_c_2(\gen_wrsw_2:wr_adgen|rd_addr_c[2]~q ),
	.rd_addr_d_3(\gen_wrsw_2:wr_adgen|rd_addr_d[3]~q ),
	.rd_addr_b_3(\gen_wrsw_2:wr_adgen|rd_addr_b[3]~q ),
	.rd_addr_d_4(\gen_wrsw_2:wr_adgen|rd_addr_d[4]~q ),
	.rd_addr_c_4(\gen_wrsw_2:wr_adgen|rd_addr_c[4]~q ),
	.rd_addr_d_5(\gen_wrsw_2:wr_adgen|rd_addr_d[5]~q ),
	.rd_addr_b_5(\gen_wrsw_2:wr_adgen|rd_addr_b[5]~q ),
	.rd_addr_d_6(\gen_wrsw_2:wr_adgen|rd_addr_d[6]~q ),
	.tdl_arr_4_20(\gen_wrsw_2:k_delay|tdl_arr[20][4]~q ),
	.tdl_arr_6_20(\gen_wrsw_2:k_delay|tdl_arr[20][6]~q ),
	.tdl_arr_0_20(\gen_wrsw_2:k_delay|tdl_arr[20][0]~q ),
	.tdl_arr_2_20(\gen_wrsw_2:k_delay|tdl_arr[20][2]~q ),
	.tdl_arr_0_1(\gen_wrsw_2:p_delay|tdl_arr[1][0]~q ),
	.tdl_arr_2_1(\gen_wrsw_2:p_delay|tdl_arr[1][2]~q ),
	.tdl_arr_1_1(\gen_wrsw_2:p_delay|tdl_arr[1][1]~q ),
	.tdl_arr_1_20(\gen_wrsw_2:k_delay|tdl_arr[20][1]~q ),
	.tdl_arr_3_20(\gen_wrsw_2:k_delay|tdl_arr[20][3]~q ),
	.tdl_arr_5_20(\gen_wrsw_2:k_delay|tdl_arr[20][5]~q ),
	.clk(clk));

fft_asj_fft_wrswgen_fft_120 \gen_wrsw_2:get_wr_swtiches (
	.global_clock_enable(\global_clock_enable~0_combout ),
	.swa_tdl_0_0(\gen_wrsw_2:get_wr_swtiches|swa_tdl[0][0]~q ),
	.swa_tdl_1_0(\gen_wrsw_2:get_wr_swtiches|swa_tdl[0][1]~q ),
	.tdl_arr_4_20(\gen_wrsw_2:k_delay|tdl_arr[20][4]~q ),
	.tdl_arr_6_20(\gen_wrsw_2:k_delay|tdl_arr[20][6]~q ),
	.tdl_arr_0_20(\gen_wrsw_2:k_delay|tdl_arr[20][0]~q ),
	.tdl_arr_2_20(\gen_wrsw_2:k_delay|tdl_arr[20][2]~q ),
	.tdl_arr_0_1(\gen_wrsw_2:p_delay|tdl_arr[1][0]~q ),
	.tdl_arr_2_1(\gen_wrsw_2:p_delay|tdl_arr[1][2]~q ),
	.tdl_arr_1_1(\gen_wrsw_2:p_delay|tdl_arr[1][1]~q ),
	.tdl_arr_1_20(\gen_wrsw_2:k_delay|tdl_arr[20][1]~q ),
	.tdl_arr_3_20(\gen_wrsw_2:k_delay|tdl_arr[20][3]~q ),
	.tdl_arr_5_20(\gen_wrsw_2:k_delay|tdl_arr[20][5]~q ),
	.clk(clk));

fft_asj_fft_tdl_fft_120_1 \gen_wrsw_2:p_delay (
	.global_clock_enable(\global_clock_enable~0_combout ),
	.tdl_arr_0_1(\gen_wrsw_2:p_delay|tdl_arr[1][0]~q ),
	.tdl_arr_2_1(\gen_wrsw_2:p_delay|tdl_arr[1][2]~q ),
	.tdl_arr_1_1(\gen_wrsw_2:p_delay|tdl_arr[1][1]~q ),
	.data_in({gnd,gnd,gnd,gnd,\p_tdl[18][2]~q ,\p_tdl[18][1]~q ,\p_tdl[18][0]~q }),
	.clk(clk));

fft_asj_fft_tdl_fft_120 \gen_wrsw_2:k_delay (
	.global_clock_enable(\global_clock_enable~0_combout ),
	.tdl_arr_4_20(\gen_wrsw_2:k_delay|tdl_arr[20][4]~q ),
	.tdl_arr_6_20(\gen_wrsw_2:k_delay|tdl_arr[20][6]~q ),
	.tdl_arr_0_20(\gen_wrsw_2:k_delay|tdl_arr[20][0]~q ),
	.tdl_arr_2_20(\gen_wrsw_2:k_delay|tdl_arr[20][2]~q ),
	.tdl_arr_1_20(\gen_wrsw_2:k_delay|tdl_arr[20][1]~q ),
	.tdl_arr_3_20(\gen_wrsw_2:k_delay|tdl_arr[20][3]~q ),
	.tdl_arr_5_20(\gen_wrsw_2:k_delay|tdl_arr[20][5]~q ),
	.tdl_arr_6_1(\gen_wrsw_2:k_delay|tdl_arr[1][6]~q ),
	.data_in({\gen_gt256_mk:ctrl|k_count[6]~q ,\gen_gt256_mk:ctrl|k_count[5]~q ,\gen_gt256_mk:ctrl|k_count[4]~q ,\gen_gt256_mk:ctrl|k_count[3]~q ,\gen_gt256_mk:ctrl|k_count[2]~q ,\gen_gt256_mk:ctrl|k_count[1]~q ,\gen_gt256_mk:ctrl|k_count[0]~q }),
	.clk(clk));

fft_asj_fft_cxb_addr_fft_120_2 ram_cxb_rd(
	.global_clock_enable(\global_clock_enable~0_combout ),
	.ram_in_reg_0_0(\ram_cxb_rd|ram_in_reg[0][0]~q ),
	.ram_in_reg_1_0(\ram_cxb_rd|ram_in_reg[0][1]~q ),
	.ram_in_reg_2_0(\ram_cxb_rd|ram_in_reg[0][2]~q ),
	.ram_in_reg_3_0(\ram_cxb_rd|ram_in_reg[0][3]~q ),
	.ram_in_reg_4_0(\ram_cxb_rd|ram_in_reg[0][4]~q ),
	.ram_in_reg_5_0(\ram_cxb_rd|ram_in_reg[0][5]~q ),
	.ram_in_reg_0_1(\ram_cxb_rd|ram_in_reg[1][0]~q ),
	.ram_in_reg_1_1(\ram_cxb_rd|ram_in_reg[1][1]~q ),
	.ram_in_reg_2_1(\ram_cxb_rd|ram_in_reg[1][2]~q ),
	.ram_in_reg_3_1(\ram_cxb_rd|ram_in_reg[1][3]~q ),
	.ram_in_reg_4_1(\ram_cxb_rd|ram_in_reg[1][4]~q ),
	.ram_in_reg_5_1(\ram_cxb_rd|ram_in_reg[1][5]~q ),
	.ram_in_reg_1_2(\ram_cxb_rd|ram_in_reg[2][1]~q ),
	.ram_in_reg_3_2(\ram_cxb_rd|ram_in_reg[2][3]~q ),
	.ram_in_reg_5_2(\ram_cxb_rd|ram_in_reg[2][5]~q ),
	.ram_in_reg_1_3(\ram_cxb_rd|ram_in_reg[3][1]~q ),
	.ram_in_reg_3_3(\ram_cxb_rd|ram_in_reg[3][3]~q ),
	.ram_in_reg_5_3(\ram_cxb_rd|ram_in_reg[3][5]~q ),
	.rd_addr_d_0(\rd_adgen|rd_addr_d[0]~q ),
	.rd_addr_c_0(\rd_adgen|rd_addr_c[0]~q ),
	.sw_0(\rd_adgen|sw[0]~q ),
	.rd_addr_b_1(\rd_adgen|rd_addr_b[1]~q ),
	.rd_addr_d_1(\rd_adgen|rd_addr_d[1]~q ),
	.sw_1(\rd_adgen|sw[1]~q ),
	.rd_addr_d_2(\rd_adgen|rd_addr_d[2]~q ),
	.rd_addr_c_2(\rd_adgen|rd_addr_c[2]~q ),
	.rd_addr_b_3(\rd_adgen|rd_addr_b[3]~q ),
	.rd_addr_d_3(\rd_adgen|rd_addr_d[3]~q ),
	.rd_addr_d_4(\rd_adgen|rd_addr_d[4]~q ),
	.rd_addr_c_4(\rd_adgen|rd_addr_c[4]~q ),
	.rd_addr_b_5(\rd_adgen|rd_addr_b[5]~q ),
	.rd_addr_d_5(\rd_adgen|rd_addr_d[5]~q ),
	.clk(clk));

fft_asj_fft_dataadgen_fft_120_1 rd_adgen(
	.global_clock_enable(\global_clock_enable~0_combout ),
	.p_2(\gen_gt256_mk:ctrl|p[2]~q ),
	.p_0(\gen_gt256_mk:ctrl|p[0]~q ),
	.p_1(\gen_gt256_mk:ctrl|p[1]~q ),
	.Equal0(\gen_gt256_mk:ctrl|Equal0~0_combout ),
	.rd_addr_d_0(\rd_adgen|rd_addr_d[0]~q ),
	.rd_addr_c_0(\rd_adgen|rd_addr_c[0]~q ),
	.sw_0(\rd_adgen|sw[0]~q ),
	.rd_addr_b_1(\rd_adgen|rd_addr_b[1]~q ),
	.rd_addr_d_1(\rd_adgen|rd_addr_d[1]~q ),
	.sw_1(\rd_adgen|sw[1]~q ),
	.rd_addr_d_2(\rd_adgen|rd_addr_d[2]~q ),
	.rd_addr_c_2(\rd_adgen|rd_addr_c[2]~q ),
	.rd_addr_b_3(\rd_adgen|rd_addr_b[3]~q ),
	.rd_addr_d_3(\rd_adgen|rd_addr_d[3]~q ),
	.rd_addr_d_4(\rd_adgen|rd_addr_d[4]~q ),
	.rd_addr_c_4(\rd_adgen|rd_addr_c[4]~q ),
	.rd_addr_b_5(\rd_adgen|rd_addr_b[5]~q ),
	.rd_addr_d_5(\rd_adgen|rd_addr_d[5]~q ),
	.k_count_0(\gen_gt256_mk:ctrl|k_count[0]~q ),
	.k_count_2(\gen_gt256_mk:ctrl|k_count[2]~q ),
	.Mux7(\rd_adgen|Mux7~1_combout ),
	.Mux1(\rd_adgen|Mux1~0_combout ),
	.k_count_4(\gen_gt256_mk:ctrl|k_count[4]~q ),
	.Mux11(\rd_adgen|Mux1~1_combout ),
	.k_count_1(\gen_gt256_mk:ctrl|k_count[1]~q ),
	.k_count_3(\gen_gt256_mk:ctrl|k_count[3]~q ),
	.k_count_5(\gen_gt256_mk:ctrl|k_count[5]~q ),
	.k_count_6(\gen_gt256_mk:ctrl|k_count[6]~q ),
	.clk(clk));

fft_asj_fft_4dp_ram_fft_120_1 \gen_M4K_Output:dat_D (
	.q_b_1(\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[1] ),
	.q_b_11(\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[1] ),
	.q_b_12(\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[1] ),
	.q_b_13(\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[1] ),
	.q_b_0(\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[0] ),
	.q_b_01(\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[0] ),
	.q_b_02(\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[0] ),
	.q_b_03(\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[0] ),
	.q_b_7(\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[7] ),
	.q_b_71(\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[7] ),
	.q_b_72(\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[7] ),
	.q_b_73(\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[7] ),
	.q_b_6(\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[6] ),
	.q_b_61(\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[6] ),
	.q_b_62(\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[6] ),
	.q_b_63(\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[6] ),
	.q_b_5(\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[5] ),
	.q_b_51(\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[5] ),
	.q_b_52(\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[5] ),
	.q_b_53(\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[5] ),
	.q_b_4(\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[4] ),
	.q_b_41(\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[4] ),
	.q_b_42(\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[4] ),
	.q_b_43(\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[4] ),
	.q_b_3(\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[3] ),
	.q_b_31(\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[3] ),
	.q_b_32(\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[3] ),
	.q_b_33(\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[3] ),
	.q_b_2(\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[2] ),
	.q_b_21(\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[2] ),
	.q_b_22(\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[2] ),
	.q_b_23(\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[2] ),
	.q_b_9(\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[9] ),
	.q_b_91(\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[9] ),
	.q_b_92(\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[9] ),
	.q_b_93(\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[9] ),
	.q_b_8(\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[8] ),
	.q_b_81(\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[8] ),
	.q_b_82(\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[8] ),
	.q_b_83(\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[8] ),
	.q_b_15(\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[15] ),
	.q_b_151(\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[15] ),
	.q_b_152(\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[15] ),
	.q_b_153(\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[15] ),
	.q_b_14(\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[14] ),
	.q_b_141(\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[14] ),
	.q_b_142(\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[14] ),
	.q_b_143(\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[14] ),
	.q_b_131(\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[13] ),
	.q_b_132(\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[13] ),
	.q_b_133(\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[13] ),
	.q_b_134(\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[13] ),
	.q_b_121(\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[12] ),
	.q_b_122(\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[12] ),
	.q_b_123(\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[12] ),
	.q_b_124(\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[12] ),
	.q_b_111(\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[11] ),
	.q_b_112(\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[11] ),
	.q_b_113(\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[11] ),
	.q_b_114(\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[11] ),
	.q_b_10(\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[10] ),
	.q_b_101(\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[10] ),
	.q_b_102(\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[10] ),
	.q_b_103(\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[10] ),
	.ram_in_reg_1_6(\ram_cxb_wr_data|ram_in_reg[6][1]~q ),
	.ram_in_reg_1_5(\ram_cxb_wr_data|ram_in_reg[5][1]~q ),
	.ram_in_reg_1_4(\ram_cxb_wr_data|ram_in_reg[4][1]~q ),
	.ram_in_reg_1_7(\ram_cxb_wr_data|ram_in_reg[7][1]~q ),
	.ram_in_reg_0_6(\ram_cxb_wr_data|ram_in_reg[6][0]~q ),
	.ram_in_reg_0_5(\ram_cxb_wr_data|ram_in_reg[5][0]~q ),
	.ram_in_reg_0_4(\ram_cxb_wr_data|ram_in_reg[4][0]~q ),
	.ram_in_reg_0_7(\ram_cxb_wr_data|ram_in_reg[7][0]~q ),
	.ram_in_reg_7_6(\ram_cxb_wr_data|ram_in_reg[6][7]~q ),
	.ram_in_reg_7_5(\ram_cxb_wr_data|ram_in_reg[5][7]~q ),
	.ram_in_reg_7_4(\ram_cxb_wr_data|ram_in_reg[4][7]~q ),
	.ram_in_reg_7_7(\ram_cxb_wr_data|ram_in_reg[7][7]~q ),
	.ram_in_reg_6_6(\ram_cxb_wr_data|ram_in_reg[6][6]~q ),
	.ram_in_reg_6_5(\ram_cxb_wr_data|ram_in_reg[5][6]~q ),
	.ram_in_reg_6_4(\ram_cxb_wr_data|ram_in_reg[4][6]~q ),
	.ram_in_reg_6_7(\ram_cxb_wr_data|ram_in_reg[7][6]~q ),
	.ram_in_reg_5_6(\ram_cxb_wr_data|ram_in_reg[6][5]~q ),
	.ram_in_reg_5_5(\ram_cxb_wr_data|ram_in_reg[5][5]~q ),
	.ram_in_reg_5_4(\ram_cxb_wr_data|ram_in_reg[4][5]~q ),
	.ram_in_reg_5_7(\ram_cxb_wr_data|ram_in_reg[7][5]~q ),
	.ram_in_reg_4_6(\ram_cxb_wr_data|ram_in_reg[6][4]~q ),
	.ram_in_reg_4_5(\ram_cxb_wr_data|ram_in_reg[5][4]~q ),
	.ram_in_reg_4_4(\ram_cxb_wr_data|ram_in_reg[4][4]~q ),
	.ram_in_reg_4_7(\ram_cxb_wr_data|ram_in_reg[7][4]~q ),
	.ram_in_reg_3_6(\ram_cxb_wr_data|ram_in_reg[6][3]~q ),
	.ram_in_reg_3_5(\ram_cxb_wr_data|ram_in_reg[5][3]~q ),
	.ram_in_reg_3_4(\ram_cxb_wr_data|ram_in_reg[4][3]~q ),
	.ram_in_reg_3_7(\ram_cxb_wr_data|ram_in_reg[7][3]~q ),
	.ram_in_reg_2_6(\ram_cxb_wr_data|ram_in_reg[6][2]~q ),
	.ram_in_reg_2_5(\ram_cxb_wr_data|ram_in_reg[5][2]~q ),
	.ram_in_reg_2_4(\ram_cxb_wr_data|ram_in_reg[4][2]~q ),
	.ram_in_reg_2_7(\ram_cxb_wr_data|ram_in_reg[7][2]~q ),
	.ram_in_reg_1_2(\ram_cxb_wr_data|ram_in_reg[2][1]~q ),
	.ram_in_reg_1_1(\ram_cxb_wr_data|ram_in_reg[1][1]~q ),
	.ram_in_reg_1_0(\ram_cxb_wr_data|ram_in_reg[0][1]~q ),
	.ram_in_reg_1_3(\ram_cxb_wr_data|ram_in_reg[3][1]~q ),
	.ram_in_reg_0_2(\ram_cxb_wr_data|ram_in_reg[2][0]~q ),
	.ram_in_reg_0_1(\ram_cxb_wr_data|ram_in_reg[1][0]~q ),
	.ram_in_reg_0_0(\ram_cxb_wr_data|ram_in_reg[0][0]~q ),
	.ram_in_reg_0_3(\ram_cxb_wr_data|ram_in_reg[3][0]~q ),
	.ram_in_reg_7_2(\ram_cxb_wr_data|ram_in_reg[2][7]~q ),
	.ram_in_reg_7_1(\ram_cxb_wr_data|ram_in_reg[1][7]~q ),
	.ram_in_reg_7_0(\ram_cxb_wr_data|ram_in_reg[0][7]~q ),
	.ram_in_reg_7_3(\ram_cxb_wr_data|ram_in_reg[3][7]~q ),
	.ram_in_reg_6_2(\ram_cxb_wr_data|ram_in_reg[2][6]~q ),
	.ram_in_reg_6_1(\ram_cxb_wr_data|ram_in_reg[1][6]~q ),
	.ram_in_reg_6_0(\ram_cxb_wr_data|ram_in_reg[0][6]~q ),
	.ram_in_reg_6_3(\ram_cxb_wr_data|ram_in_reg[3][6]~q ),
	.ram_in_reg_5_2(\ram_cxb_wr_data|ram_in_reg[2][5]~q ),
	.ram_in_reg_5_1(\ram_cxb_wr_data|ram_in_reg[1][5]~q ),
	.ram_in_reg_5_0(\ram_cxb_wr_data|ram_in_reg[0][5]~q ),
	.ram_in_reg_5_3(\ram_cxb_wr_data|ram_in_reg[3][5]~q ),
	.ram_in_reg_4_2(\ram_cxb_wr_data|ram_in_reg[2][4]~q ),
	.ram_in_reg_4_1(\ram_cxb_wr_data|ram_in_reg[1][4]~q ),
	.ram_in_reg_4_0(\ram_cxb_wr_data|ram_in_reg[0][4]~q ),
	.ram_in_reg_4_3(\ram_cxb_wr_data|ram_in_reg[3][4]~q ),
	.ram_in_reg_3_2(\ram_cxb_wr_data|ram_in_reg[2][3]~q ),
	.ram_in_reg_3_1(\ram_cxb_wr_data|ram_in_reg[1][3]~q ),
	.ram_in_reg_3_0(\ram_cxb_wr_data|ram_in_reg[0][3]~q ),
	.ram_in_reg_3_3(\ram_cxb_wr_data|ram_in_reg[3][3]~q ),
	.ram_in_reg_2_2(\ram_cxb_wr_data|ram_in_reg[2][2]~q ),
	.ram_in_reg_2_1(\ram_cxb_wr_data|ram_in_reg[1][2]~q ),
	.ram_in_reg_2_0(\ram_cxb_wr_data|ram_in_reg[0][2]~q ),
	.ram_in_reg_2_3(\ram_cxb_wr_data|ram_in_reg[3][2]~q ),
	.global_clock_enable(\global_clock_enable~0_combout ),
	.ram_in_reg_0_01(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[0][0]~q ),
	.ram_in_reg_1_21(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[2][1]~q ),
	.ram_in_reg_2_01(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[0][2]~q ),
	.ram_in_reg_3_21(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[2][3]~q ),
	.ram_in_reg_4_01(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[0][4]~q ),
	.ram_in_reg_5_21(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[2][5]~q ),
	.ram_in_reg_6_01(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[0][6]~q ),
	.rdaddress_c_bus_0(\rdaddress_c_bus[0]~q ),
	.rdaddress_c_bus_15(\rdaddress_c_bus[15]~q ),
	.rdaddress_c_bus_16(\rdaddress_c_bus[16]~q ),
	.rdaddress_c_bus_10(\rdaddress_c_bus[10]~q ),
	.rdaddress_c_bus_11(\rdaddress_c_bus[11]~q ),
	.rdaddress_c_bus_12(\rdaddress_c_bus[12]~q ),
	.rdaddress_c_bus_13(\rdaddress_c_bus[13]~q ),
	.wd_vec_6(\wd_vec[6]~q ),
	.ram_in_reg_0_11(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[1][0]~q ),
	.ram_in_reg_1_11(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[1][1]~q ),
	.ram_in_reg_2_11(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[1][2]~q ),
	.ram_in_reg_3_11(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[1][3]~q ),
	.ram_in_reg_4_11(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[1][4]~q ),
	.ram_in_reg_5_11(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[1][5]~q ),
	.rdaddress_c_bus_20(\rdaddress_c_bus[20]~q ),
	.ram_in_reg_1_01(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[0][1]~q ),
	.ram_in_reg_3_01(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[0][3]~q ),
	.ram_in_reg_5_01(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[0][5]~q ),
	.ram_in_reg_1_31(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[3][1]~q ),
	.ram_in_reg_3_31(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[3][3]~q ),
	.ram_in_reg_5_31(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[3][5]~q ),
	.clk(clk));

fft_asj_fft_4dp_ram_fft_120 \gen_M4K_Output:dat_C (
	.q_b_1(\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[1] ),
	.q_b_11(\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[1] ),
	.q_b_12(\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[1] ),
	.q_b_13(\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[1] ),
	.q_b_0(\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[0] ),
	.q_b_01(\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[0] ),
	.q_b_02(\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[0] ),
	.q_b_03(\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[0] ),
	.q_b_7(\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[7] ),
	.q_b_71(\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[7] ),
	.q_b_72(\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[7] ),
	.q_b_73(\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[7] ),
	.q_b_6(\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[6] ),
	.q_b_61(\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[6] ),
	.q_b_62(\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[6] ),
	.q_b_63(\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[6] ),
	.q_b_5(\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[5] ),
	.q_b_51(\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[5] ),
	.q_b_52(\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[5] ),
	.q_b_53(\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[5] ),
	.q_b_4(\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[4] ),
	.q_b_41(\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[4] ),
	.q_b_42(\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[4] ),
	.q_b_43(\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[4] ),
	.q_b_3(\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[3] ),
	.q_b_31(\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[3] ),
	.q_b_32(\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[3] ),
	.q_b_33(\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[3] ),
	.q_b_2(\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[2] ),
	.q_b_21(\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[2] ),
	.q_b_22(\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[2] ),
	.q_b_23(\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[2] ),
	.q_b_9(\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[9] ),
	.q_b_91(\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[9] ),
	.q_b_92(\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[9] ),
	.q_b_93(\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[9] ),
	.q_b_8(\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[8] ),
	.q_b_81(\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[8] ),
	.q_b_82(\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[8] ),
	.q_b_83(\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[8] ),
	.q_b_15(\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[15] ),
	.q_b_151(\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[15] ),
	.q_b_152(\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[15] ),
	.q_b_153(\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[15] ),
	.q_b_14(\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[14] ),
	.q_b_141(\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[14] ),
	.q_b_142(\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[14] ),
	.q_b_143(\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[14] ),
	.q_b_131(\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[13] ),
	.q_b_132(\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[13] ),
	.q_b_133(\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[13] ),
	.q_b_134(\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[13] ),
	.q_b_121(\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[12] ),
	.q_b_122(\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[12] ),
	.q_b_123(\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[12] ),
	.q_b_124(\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[12] ),
	.q_b_111(\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[11] ),
	.q_b_112(\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[11] ),
	.q_b_113(\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[11] ),
	.q_b_114(\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[11] ),
	.q_b_10(\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[10] ),
	.q_b_101(\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[10] ),
	.q_b_102(\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[10] ),
	.q_b_103(\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[10] ),
	.ram_in_reg_1_6(\ram_cxb_wr_data|ram_in_reg[6][1]~q ),
	.ram_in_reg_1_5(\ram_cxb_wr_data|ram_in_reg[5][1]~q ),
	.ram_in_reg_1_4(\ram_cxb_wr_data|ram_in_reg[4][1]~q ),
	.ram_in_reg_1_7(\ram_cxb_wr_data|ram_in_reg[7][1]~q ),
	.ram_in_reg_0_6(\ram_cxb_wr_data|ram_in_reg[6][0]~q ),
	.ram_in_reg_0_5(\ram_cxb_wr_data|ram_in_reg[5][0]~q ),
	.ram_in_reg_0_4(\ram_cxb_wr_data|ram_in_reg[4][0]~q ),
	.ram_in_reg_0_7(\ram_cxb_wr_data|ram_in_reg[7][0]~q ),
	.ram_in_reg_7_6(\ram_cxb_wr_data|ram_in_reg[6][7]~q ),
	.ram_in_reg_7_5(\ram_cxb_wr_data|ram_in_reg[5][7]~q ),
	.ram_in_reg_7_4(\ram_cxb_wr_data|ram_in_reg[4][7]~q ),
	.ram_in_reg_7_7(\ram_cxb_wr_data|ram_in_reg[7][7]~q ),
	.ram_in_reg_6_6(\ram_cxb_wr_data|ram_in_reg[6][6]~q ),
	.ram_in_reg_6_5(\ram_cxb_wr_data|ram_in_reg[5][6]~q ),
	.ram_in_reg_6_4(\ram_cxb_wr_data|ram_in_reg[4][6]~q ),
	.ram_in_reg_6_7(\ram_cxb_wr_data|ram_in_reg[7][6]~q ),
	.ram_in_reg_5_6(\ram_cxb_wr_data|ram_in_reg[6][5]~q ),
	.ram_in_reg_5_5(\ram_cxb_wr_data|ram_in_reg[5][5]~q ),
	.ram_in_reg_5_4(\ram_cxb_wr_data|ram_in_reg[4][5]~q ),
	.ram_in_reg_5_7(\ram_cxb_wr_data|ram_in_reg[7][5]~q ),
	.ram_in_reg_4_6(\ram_cxb_wr_data|ram_in_reg[6][4]~q ),
	.ram_in_reg_4_5(\ram_cxb_wr_data|ram_in_reg[5][4]~q ),
	.ram_in_reg_4_4(\ram_cxb_wr_data|ram_in_reg[4][4]~q ),
	.ram_in_reg_4_7(\ram_cxb_wr_data|ram_in_reg[7][4]~q ),
	.ram_in_reg_3_6(\ram_cxb_wr_data|ram_in_reg[6][3]~q ),
	.ram_in_reg_3_5(\ram_cxb_wr_data|ram_in_reg[5][3]~q ),
	.ram_in_reg_3_4(\ram_cxb_wr_data|ram_in_reg[4][3]~q ),
	.ram_in_reg_3_7(\ram_cxb_wr_data|ram_in_reg[7][3]~q ),
	.ram_in_reg_2_6(\ram_cxb_wr_data|ram_in_reg[6][2]~q ),
	.ram_in_reg_2_5(\ram_cxb_wr_data|ram_in_reg[5][2]~q ),
	.ram_in_reg_2_4(\ram_cxb_wr_data|ram_in_reg[4][2]~q ),
	.ram_in_reg_2_7(\ram_cxb_wr_data|ram_in_reg[7][2]~q ),
	.ram_in_reg_1_2(\ram_cxb_wr_data|ram_in_reg[2][1]~q ),
	.ram_in_reg_1_1(\ram_cxb_wr_data|ram_in_reg[1][1]~q ),
	.ram_in_reg_1_0(\ram_cxb_wr_data|ram_in_reg[0][1]~q ),
	.ram_in_reg_1_3(\ram_cxb_wr_data|ram_in_reg[3][1]~q ),
	.ram_in_reg_0_2(\ram_cxb_wr_data|ram_in_reg[2][0]~q ),
	.ram_in_reg_0_1(\ram_cxb_wr_data|ram_in_reg[1][0]~q ),
	.ram_in_reg_0_0(\ram_cxb_wr_data|ram_in_reg[0][0]~q ),
	.ram_in_reg_0_3(\ram_cxb_wr_data|ram_in_reg[3][0]~q ),
	.ram_in_reg_7_2(\ram_cxb_wr_data|ram_in_reg[2][7]~q ),
	.ram_in_reg_7_1(\ram_cxb_wr_data|ram_in_reg[1][7]~q ),
	.ram_in_reg_7_0(\ram_cxb_wr_data|ram_in_reg[0][7]~q ),
	.ram_in_reg_7_3(\ram_cxb_wr_data|ram_in_reg[3][7]~q ),
	.ram_in_reg_6_2(\ram_cxb_wr_data|ram_in_reg[2][6]~q ),
	.ram_in_reg_6_1(\ram_cxb_wr_data|ram_in_reg[1][6]~q ),
	.ram_in_reg_6_0(\ram_cxb_wr_data|ram_in_reg[0][6]~q ),
	.ram_in_reg_6_3(\ram_cxb_wr_data|ram_in_reg[3][6]~q ),
	.ram_in_reg_5_2(\ram_cxb_wr_data|ram_in_reg[2][5]~q ),
	.ram_in_reg_5_1(\ram_cxb_wr_data|ram_in_reg[1][5]~q ),
	.ram_in_reg_5_0(\ram_cxb_wr_data|ram_in_reg[0][5]~q ),
	.ram_in_reg_5_3(\ram_cxb_wr_data|ram_in_reg[3][5]~q ),
	.ram_in_reg_4_2(\ram_cxb_wr_data|ram_in_reg[2][4]~q ),
	.ram_in_reg_4_1(\ram_cxb_wr_data|ram_in_reg[1][4]~q ),
	.ram_in_reg_4_0(\ram_cxb_wr_data|ram_in_reg[0][4]~q ),
	.ram_in_reg_4_3(\ram_cxb_wr_data|ram_in_reg[3][4]~q ),
	.ram_in_reg_3_2(\ram_cxb_wr_data|ram_in_reg[2][3]~q ),
	.ram_in_reg_3_1(\ram_cxb_wr_data|ram_in_reg[1][3]~q ),
	.ram_in_reg_3_0(\ram_cxb_wr_data|ram_in_reg[0][3]~q ),
	.ram_in_reg_3_3(\ram_cxb_wr_data|ram_in_reg[3][3]~q ),
	.ram_in_reg_2_2(\ram_cxb_wr_data|ram_in_reg[2][2]~q ),
	.ram_in_reg_2_1(\ram_cxb_wr_data|ram_in_reg[1][2]~q ),
	.ram_in_reg_2_0(\ram_cxb_wr_data|ram_in_reg[0][2]~q ),
	.ram_in_reg_2_3(\ram_cxb_wr_data|ram_in_reg[3][2]~q ),
	.global_clock_enable(\global_clock_enable~0_combout ),
	.wc_vec_6(\wc_vec[6]~q ),
	.ram_in_reg_0_01(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[0][0]~q ),
	.ram_in_reg_1_21(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[2][1]~q ),
	.ram_in_reg_2_01(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[0][2]~q ),
	.ram_in_reg_3_21(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[2][3]~q ),
	.ram_in_reg_4_01(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[0][4]~q ),
	.ram_in_reg_5_21(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[2][5]~q ),
	.ram_in_reg_6_01(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[0][6]~q ),
	.rdaddress_c_bus_0(\rdaddress_c_bus[0]~q ),
	.rdaddress_c_bus_15(\rdaddress_c_bus[15]~q ),
	.rdaddress_c_bus_16(\rdaddress_c_bus[16]~q ),
	.rdaddress_c_bus_10(\rdaddress_c_bus[10]~q ),
	.rdaddress_c_bus_11(\rdaddress_c_bus[11]~q ),
	.rdaddress_c_bus_12(\rdaddress_c_bus[12]~q ),
	.rdaddress_c_bus_13(\rdaddress_c_bus[13]~q ),
	.ram_in_reg_0_11(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[1][0]~q ),
	.ram_in_reg_1_11(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[1][1]~q ),
	.ram_in_reg_2_11(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[1][2]~q ),
	.ram_in_reg_3_11(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[1][3]~q ),
	.ram_in_reg_4_11(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[1][4]~q ),
	.ram_in_reg_5_11(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[1][5]~q ),
	.rdaddress_c_bus_20(\rdaddress_c_bus[20]~q ),
	.ram_in_reg_1_01(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[0][1]~q ),
	.ram_in_reg_3_01(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[0][3]~q ),
	.ram_in_reg_5_01(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[0][5]~q ),
	.ram_in_reg_1_31(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[3][1]~q ),
	.ram_in_reg_3_31(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[3][3]~q ),
	.ram_in_reg_5_31(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[3][5]~q ),
	.clk(clk));

fft_asj_fft_4dp_ram_fft_120_3 dat_B(
	.q_b_10(\dat_B|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[10] ),
	.q_b_101(\dat_B|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[10] ),
	.q_b_102(\dat_B|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[10] ),
	.q_b_103(\dat_B|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[10] ),
	.q_b_14(\dat_B|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[14] ),
	.q_b_141(\dat_B|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[14] ),
	.q_b_142(\dat_B|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[14] ),
	.q_b_143(\dat_B|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[14] ),
	.q_b_12(\dat_B|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[12] ),
	.q_b_121(\dat_B|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[12] ),
	.q_b_122(\dat_B|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[12] ),
	.q_b_123(\dat_B|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[12] ),
	.q_b_11(\dat_B|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[11] ),
	.q_b_111(\dat_B|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[11] ),
	.q_b_112(\dat_B|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[11] ),
	.q_b_113(\dat_B|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[11] ),
	.q_b_13(\dat_B|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[13] ),
	.q_b_131(\dat_B|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[13] ),
	.q_b_132(\dat_B|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[13] ),
	.q_b_133(\dat_B|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[13] ),
	.q_b_9(\dat_B|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[9] ),
	.q_b_91(\dat_B|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[9] ),
	.q_b_92(\dat_B|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[9] ),
	.q_b_93(\dat_B|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[9] ),
	.q_b_8(\dat_B|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[8] ),
	.q_b_81(\dat_B|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[8] ),
	.q_b_82(\dat_B|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[8] ),
	.q_b_83(\dat_B|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[8] ),
	.q_b_15(\dat_B|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[15] ),
	.q_b_151(\dat_B|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[15] ),
	.q_b_152(\dat_B|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[15] ),
	.q_b_153(\dat_B|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[15] ),
	.q_b_7(\dat_B|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[7] ),
	.q_b_71(\dat_B|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[7] ),
	.q_b_72(\dat_B|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[7] ),
	.q_b_73(\dat_B|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[7] ),
	.q_b_3(\dat_B|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[3] ),
	.q_b_31(\dat_B|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[3] ),
	.q_b_32(\dat_B|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[3] ),
	.q_b_33(\dat_B|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[3] ),
	.q_b_5(\dat_B|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[5] ),
	.q_b_51(\dat_B|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[5] ),
	.q_b_52(\dat_B|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[5] ),
	.q_b_53(\dat_B|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[5] ),
	.q_b_4(\dat_B|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[4] ),
	.q_b_41(\dat_B|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[4] ),
	.q_b_42(\dat_B|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[4] ),
	.q_b_43(\dat_B|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[4] ),
	.q_b_6(\dat_B|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[6] ),
	.q_b_61(\dat_B|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[6] ),
	.q_b_62(\dat_B|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[6] ),
	.q_b_63(\dat_B|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[6] ),
	.q_b_2(\dat_B|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[2] ),
	.q_b_21(\dat_B|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[2] ),
	.q_b_22(\dat_B|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[2] ),
	.q_b_23(\dat_B|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[2] ),
	.q_b_1(\dat_B|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[1] ),
	.q_b_16(\dat_B|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[1] ),
	.q_b_17(\dat_B|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[1] ),
	.q_b_18(\dat_B|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[1] ),
	.q_b_0(\dat_B|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[0] ),
	.q_b_01(\dat_B|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[0] ),
	.q_b_02(\dat_B|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[0] ),
	.q_b_03(\dat_B|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[0] ),
	.wren_b_0(\wren_b[0]~q ),
	.wren_b_1(\wren_b[1]~q ),
	.wren_b_2(\wren_b[2]~q ),
	.wren_b_3(\wren_b[3]~q ),
	.global_clock_enable(\global_clock_enable~0_combout ),
	.b_ram_data_in_bus_58(\ccc|b_ram_data_in_bus[58]~q ),
	.wraddress_b_bus_21(\ccc|wraddress_b_bus[21]~q ),
	.wraddress_b_bus_22(\ccc|wraddress_b_bus[22]~q ),
	.wraddress_b_bus_23(\ccc|wraddress_b_bus[23]~q ),
	.wraddress_b_bus_24(\ccc|wraddress_b_bus[24]~q ),
	.wraddress_b_bus_11(\ccc|wraddress_b_bus[11]~q ),
	.wraddress_b_bus_26(\ccc|wraddress_b_bus[26]~q ),
	.wraddress_b_bus_13(\ccc|wraddress_b_bus[13]~q ),
	.rdaddress_b_bus_21(\ccc|rdaddress_b_bus[21]~q ),
	.rdaddress_b_bus_22(\ccc|rdaddress_b_bus[22]~q ),
	.rdaddress_b_bus_23(\ccc|rdaddress_b_bus[23]~q ),
	.rdaddress_b_bus_24(\ccc|rdaddress_b_bus[24]~q ),
	.rdaddress_b_bus_11(\ccc|rdaddress_b_bus[11]~q ),
	.rdaddress_b_bus_26(\ccc|rdaddress_b_bus[26]~q ),
	.rdaddress_b_bus_13(\ccc|rdaddress_b_bus[13]~q ),
	.b_ram_data_in_bus_42(\ccc|b_ram_data_in_bus[42]~q ),
	.wraddress_b_bus_0(\ccc|wraddress_b_bus[0]~q ),
	.wraddress_b_bus_15(\ccc|wraddress_b_bus[15]~q ),
	.wraddress_b_bus_16(\ccc|wraddress_b_bus[16]~q ),
	.wraddress_b_bus_17(\ccc|wraddress_b_bus[17]~q ),
	.wraddress_b_bus_18(\ccc|wraddress_b_bus[18]~q ),
	.wraddress_b_bus_19(\ccc|wraddress_b_bus[19]~q ),
	.rdaddress_b_bus_0(\ccc|rdaddress_b_bus[0]~q ),
	.rdaddress_b_bus_15(\ccc|rdaddress_b_bus[15]~q ),
	.rdaddress_b_bus_16(\ccc|rdaddress_b_bus[16]~q ),
	.rdaddress_b_bus_17(\ccc|rdaddress_b_bus[17]~q ),
	.rdaddress_b_bus_18(\ccc|rdaddress_b_bus[18]~q ),
	.rdaddress_b_bus_19(\ccc|rdaddress_b_bus[19]~q ),
	.b_ram_data_in_bus_26(\ccc|b_ram_data_in_bus[26]~q ),
	.wraddress_b_bus_8(\ccc|wraddress_b_bus[8]~q ),
	.wraddress_b_bus_10(\ccc|wraddress_b_bus[10]~q ),
	.wraddress_b_bus_12(\ccc|wraddress_b_bus[12]~q ),
	.rdaddress_b_bus_8(\ccc|rdaddress_b_bus[8]~q ),
	.rdaddress_b_bus_10(\ccc|rdaddress_b_bus[10]~q ),
	.rdaddress_b_bus_12(\ccc|rdaddress_b_bus[12]~q ),
	.b_ram_data_in_bus_10(\ccc|b_ram_data_in_bus[10]~q ),
	.wraddress_b_bus_1(\ccc|wraddress_b_bus[1]~q ),
	.wraddress_b_bus_3(\ccc|wraddress_b_bus[3]~q ),
	.wraddress_b_bus_5(\ccc|wraddress_b_bus[5]~q ),
	.rdaddress_b_bus_1(\ccc|rdaddress_b_bus[1]~q ),
	.rdaddress_b_bus_3(\ccc|rdaddress_b_bus[3]~q ),
	.rdaddress_b_bus_5(\ccc|rdaddress_b_bus[5]~q ),
	.b_ram_data_in_bus_62(\ccc|b_ram_data_in_bus[62]~q ),
	.b_ram_data_in_bus_46(\ccc|b_ram_data_in_bus[46]~q ),
	.b_ram_data_in_bus_30(\ccc|b_ram_data_in_bus[30]~q ),
	.b_ram_data_in_bus_14(\ccc|b_ram_data_in_bus[14]~q ),
	.b_ram_data_in_bus_60(\ccc|b_ram_data_in_bus[60]~q ),
	.b_ram_data_in_bus_44(\ccc|b_ram_data_in_bus[44]~q ),
	.b_ram_data_in_bus_28(\ccc|b_ram_data_in_bus[28]~q ),
	.b_ram_data_in_bus_12(\ccc|b_ram_data_in_bus[12]~q ),
	.b_ram_data_in_bus_59(\ccc|b_ram_data_in_bus[59]~q ),
	.b_ram_data_in_bus_43(\ccc|b_ram_data_in_bus[43]~q ),
	.b_ram_data_in_bus_27(\ccc|b_ram_data_in_bus[27]~q ),
	.b_ram_data_in_bus_11(\ccc|b_ram_data_in_bus[11]~q ),
	.b_ram_data_in_bus_61(\ccc|b_ram_data_in_bus[61]~q ),
	.b_ram_data_in_bus_45(\ccc|b_ram_data_in_bus[45]~q ),
	.b_ram_data_in_bus_29(\ccc|b_ram_data_in_bus[29]~q ),
	.b_ram_data_in_bus_13(\ccc|b_ram_data_in_bus[13]~q ),
	.b_ram_data_in_bus_57(\ccc|b_ram_data_in_bus[57]~q ),
	.b_ram_data_in_bus_41(\ccc|b_ram_data_in_bus[41]~q ),
	.b_ram_data_in_bus_25(\ccc|b_ram_data_in_bus[25]~q ),
	.b_ram_data_in_bus_9(\ccc|b_ram_data_in_bus[9]~q ),
	.b_ram_data_in_bus_56(\ccc|b_ram_data_in_bus[56]~q ),
	.b_ram_data_in_bus_40(\ccc|b_ram_data_in_bus[40]~q ),
	.b_ram_data_in_bus_24(\ccc|b_ram_data_in_bus[24]~q ),
	.b_ram_data_in_bus_8(\ccc|b_ram_data_in_bus[8]~q ),
	.b_ram_data_in_bus_63(\ccc|b_ram_data_in_bus[63]~q ),
	.b_ram_data_in_bus_47(\ccc|b_ram_data_in_bus[47]~q ),
	.b_ram_data_in_bus_31(\ccc|b_ram_data_in_bus[31]~q ),
	.b_ram_data_in_bus_15(\ccc|b_ram_data_in_bus[15]~q ),
	.b_ram_data_in_bus_55(\ccc|b_ram_data_in_bus[55]~q ),
	.b_ram_data_in_bus_39(\ccc|b_ram_data_in_bus[39]~q ),
	.b_ram_data_in_bus_23(\ccc|b_ram_data_in_bus[23]~q ),
	.b_ram_data_in_bus_7(\ccc|b_ram_data_in_bus[7]~q ),
	.b_ram_data_in_bus_51(\ccc|b_ram_data_in_bus[51]~q ),
	.b_ram_data_in_bus_35(\ccc|b_ram_data_in_bus[35]~q ),
	.b_ram_data_in_bus_19(\ccc|b_ram_data_in_bus[19]~q ),
	.b_ram_data_in_bus_3(\ccc|b_ram_data_in_bus[3]~q ),
	.b_ram_data_in_bus_53(\ccc|b_ram_data_in_bus[53]~q ),
	.b_ram_data_in_bus_37(\ccc|b_ram_data_in_bus[37]~q ),
	.b_ram_data_in_bus_21(\ccc|b_ram_data_in_bus[21]~q ),
	.b_ram_data_in_bus_5(\ccc|b_ram_data_in_bus[5]~q ),
	.b_ram_data_in_bus_52(\ccc|b_ram_data_in_bus[52]~q ),
	.b_ram_data_in_bus_36(\ccc|b_ram_data_in_bus[36]~q ),
	.b_ram_data_in_bus_20(\ccc|b_ram_data_in_bus[20]~q ),
	.b_ram_data_in_bus_4(\ccc|b_ram_data_in_bus[4]~q ),
	.b_ram_data_in_bus_54(\ccc|b_ram_data_in_bus[54]~q ),
	.b_ram_data_in_bus_38(\ccc|b_ram_data_in_bus[38]~q ),
	.b_ram_data_in_bus_22(\ccc|b_ram_data_in_bus[22]~q ),
	.b_ram_data_in_bus_6(\ccc|b_ram_data_in_bus[6]~q ),
	.b_ram_data_in_bus_50(\ccc|b_ram_data_in_bus[50]~q ),
	.b_ram_data_in_bus_34(\ccc|b_ram_data_in_bus[34]~q ),
	.b_ram_data_in_bus_18(\ccc|b_ram_data_in_bus[18]~q ),
	.b_ram_data_in_bus_2(\ccc|b_ram_data_in_bus[2]~q ),
	.b_ram_data_in_bus_49(\ccc|b_ram_data_in_bus[49]~q ),
	.b_ram_data_in_bus_33(\ccc|b_ram_data_in_bus[33]~q ),
	.b_ram_data_in_bus_17(\ccc|b_ram_data_in_bus[17]~q ),
	.b_ram_data_in_bus_1(\ccc|b_ram_data_in_bus[1]~q ),
	.b_ram_data_in_bus_48(\ccc|b_ram_data_in_bus[48]~q ),
	.b_ram_data_in_bus_32(\ccc|b_ram_data_in_bus[32]~q ),
	.b_ram_data_in_bus_16(\ccc|b_ram_data_in_bus[16]~q ),
	.b_ram_data_in_bus_0(\ccc|b_ram_data_in_bus[0]~q ),
	.clk(clk));

fft_asj_fft_4dp_ram_fft_120_2 dat_A(
	.q_b_10(\dat_A|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[10] ),
	.q_b_101(\dat_A|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[10] ),
	.q_b_102(\dat_A|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[10] ),
	.q_b_103(\dat_A|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[10] ),
	.q_b_14(\dat_A|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[14] ),
	.q_b_141(\dat_A|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[14] ),
	.q_b_142(\dat_A|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[14] ),
	.q_b_143(\dat_A|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[14] ),
	.q_b_12(\dat_A|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[12] ),
	.q_b_121(\dat_A|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[12] ),
	.q_b_122(\dat_A|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[12] ),
	.q_b_123(\dat_A|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[12] ),
	.q_b_11(\dat_A|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[11] ),
	.q_b_111(\dat_A|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[11] ),
	.q_b_112(\dat_A|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[11] ),
	.q_b_113(\dat_A|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[11] ),
	.q_b_13(\dat_A|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[13] ),
	.q_b_131(\dat_A|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[13] ),
	.q_b_132(\dat_A|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[13] ),
	.q_b_133(\dat_A|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[13] ),
	.q_b_9(\dat_A|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[9] ),
	.q_b_91(\dat_A|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[9] ),
	.q_b_92(\dat_A|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[9] ),
	.q_b_93(\dat_A|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[9] ),
	.q_b_8(\dat_A|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[8] ),
	.q_b_81(\dat_A|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[8] ),
	.q_b_82(\dat_A|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[8] ),
	.q_b_83(\dat_A|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[8] ),
	.q_b_15(\dat_A|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[15] ),
	.q_b_151(\dat_A|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[15] ),
	.q_b_152(\dat_A|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[15] ),
	.q_b_153(\dat_A|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[15] ),
	.q_b_7(\dat_A|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[7] ),
	.q_b_71(\dat_A|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[7] ),
	.q_b_72(\dat_A|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[7] ),
	.q_b_73(\dat_A|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[7] ),
	.q_b_3(\dat_A|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[3] ),
	.q_b_31(\dat_A|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[3] ),
	.q_b_32(\dat_A|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[3] ),
	.q_b_33(\dat_A|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[3] ),
	.q_b_5(\dat_A|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[5] ),
	.q_b_51(\dat_A|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[5] ),
	.q_b_52(\dat_A|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[5] ),
	.q_b_53(\dat_A|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[5] ),
	.q_b_4(\dat_A|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[4] ),
	.q_b_41(\dat_A|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[4] ),
	.q_b_42(\dat_A|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[4] ),
	.q_b_43(\dat_A|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[4] ),
	.q_b_6(\dat_A|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[6] ),
	.q_b_61(\dat_A|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[6] ),
	.q_b_62(\dat_A|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[6] ),
	.q_b_63(\dat_A|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[6] ),
	.q_b_2(\dat_A|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[2] ),
	.q_b_21(\dat_A|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[2] ),
	.q_b_22(\dat_A|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[2] ),
	.q_b_23(\dat_A|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[2] ),
	.q_b_1(\dat_A|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[1] ),
	.q_b_16(\dat_A|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[1] ),
	.q_b_17(\dat_A|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[1] ),
	.q_b_18(\dat_A|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[1] ),
	.q_b_0(\dat_A|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[0] ),
	.q_b_01(\dat_A|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[0] ),
	.q_b_02(\dat_A|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[0] ),
	.q_b_03(\dat_A|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[0] ),
	.wren_a_0(\wren_a[0]~q ),
	.wren_a_1(\wren_a[1]~q ),
	.wren_a_2(\wren_a[2]~q ),
	.wren_a_3(\wren_a[3]~q ),
	.global_clock_enable(\global_clock_enable~0_combout ),
	.a_ram_data_in_bus_58(\ccc|a_ram_data_in_bus[58]~q ),
	.wraddress_a_bus_21(\ccc|wraddress_a_bus[21]~q ),
	.wraddress_a_bus_22(\ccc|wraddress_a_bus[22]~q ),
	.wraddress_a_bus_23(\ccc|wraddress_a_bus[23]~q ),
	.wraddress_a_bus_24(\ccc|wraddress_a_bus[24]~q ),
	.wraddress_a_bus_11(\ccc|wraddress_a_bus[11]~q ),
	.wraddress_a_bus_26(\ccc|wraddress_a_bus[26]~q ),
	.wraddress_a_bus_13(\ccc|wraddress_a_bus[13]~q ),
	.rdaddress_a_bus_21(\ccc|rdaddress_a_bus[21]~q ),
	.rdaddress_a_bus_22(\ccc|rdaddress_a_bus[22]~q ),
	.rdaddress_a_bus_23(\ccc|rdaddress_a_bus[23]~q ),
	.rdaddress_a_bus_24(\ccc|rdaddress_a_bus[24]~q ),
	.rdaddress_a_bus_11(\ccc|rdaddress_a_bus[11]~q ),
	.rdaddress_a_bus_26(\ccc|rdaddress_a_bus[26]~q ),
	.rdaddress_a_bus_13(\ccc|rdaddress_a_bus[13]~q ),
	.a_ram_data_in_bus_42(\ccc|a_ram_data_in_bus[42]~q ),
	.wraddress_a_bus_0(\ccc|wraddress_a_bus[0]~q ),
	.wraddress_a_bus_15(\ccc|wraddress_a_bus[15]~q ),
	.wraddress_a_bus_16(\ccc|wraddress_a_bus[16]~q ),
	.wraddress_a_bus_17(\ccc|wraddress_a_bus[17]~q ),
	.wraddress_a_bus_18(\ccc|wraddress_a_bus[18]~q ),
	.wraddress_a_bus_19(\ccc|wraddress_a_bus[19]~q ),
	.rdaddress_a_bus_0(\ccc|rdaddress_a_bus[0]~q ),
	.rdaddress_a_bus_15(\ccc|rdaddress_a_bus[15]~q ),
	.rdaddress_a_bus_16(\ccc|rdaddress_a_bus[16]~q ),
	.rdaddress_a_bus_17(\ccc|rdaddress_a_bus[17]~q ),
	.rdaddress_a_bus_18(\ccc|rdaddress_a_bus[18]~q ),
	.rdaddress_a_bus_19(\ccc|rdaddress_a_bus[19]~q ),
	.a_ram_data_in_bus_26(\ccc|a_ram_data_in_bus[26]~q ),
	.wraddress_a_bus_8(\ccc|wraddress_a_bus[8]~q ),
	.wraddress_a_bus_10(\ccc|wraddress_a_bus[10]~q ),
	.wraddress_a_bus_12(\ccc|wraddress_a_bus[12]~q ),
	.rdaddress_a_bus_8(\ccc|rdaddress_a_bus[8]~q ),
	.rdaddress_a_bus_10(\ccc|rdaddress_a_bus[10]~q ),
	.rdaddress_a_bus_12(\ccc|rdaddress_a_bus[12]~q ),
	.a_ram_data_in_bus_10(\ccc|a_ram_data_in_bus[10]~q ),
	.wraddress_a_bus_1(\ccc|wraddress_a_bus[1]~q ),
	.wraddress_a_bus_3(\ccc|wraddress_a_bus[3]~q ),
	.wraddress_a_bus_5(\ccc|wraddress_a_bus[5]~q ),
	.rdaddress_a_bus_1(\ccc|rdaddress_a_bus[1]~q ),
	.rdaddress_a_bus_3(\ccc|rdaddress_a_bus[3]~q ),
	.rdaddress_a_bus_5(\ccc|rdaddress_a_bus[5]~q ),
	.a_ram_data_in_bus_62(\ccc|a_ram_data_in_bus[62]~q ),
	.a_ram_data_in_bus_46(\ccc|a_ram_data_in_bus[46]~q ),
	.a_ram_data_in_bus_30(\ccc|a_ram_data_in_bus[30]~q ),
	.a_ram_data_in_bus_14(\ccc|a_ram_data_in_bus[14]~q ),
	.a_ram_data_in_bus_60(\ccc|a_ram_data_in_bus[60]~q ),
	.a_ram_data_in_bus_44(\ccc|a_ram_data_in_bus[44]~q ),
	.a_ram_data_in_bus_28(\ccc|a_ram_data_in_bus[28]~q ),
	.a_ram_data_in_bus_12(\ccc|a_ram_data_in_bus[12]~q ),
	.a_ram_data_in_bus_59(\ccc|a_ram_data_in_bus[59]~q ),
	.a_ram_data_in_bus_43(\ccc|a_ram_data_in_bus[43]~q ),
	.a_ram_data_in_bus_27(\ccc|a_ram_data_in_bus[27]~q ),
	.a_ram_data_in_bus_11(\ccc|a_ram_data_in_bus[11]~q ),
	.a_ram_data_in_bus_61(\ccc|a_ram_data_in_bus[61]~q ),
	.a_ram_data_in_bus_45(\ccc|a_ram_data_in_bus[45]~q ),
	.a_ram_data_in_bus_29(\ccc|a_ram_data_in_bus[29]~q ),
	.a_ram_data_in_bus_13(\ccc|a_ram_data_in_bus[13]~q ),
	.a_ram_data_in_bus_57(\ccc|a_ram_data_in_bus[57]~q ),
	.a_ram_data_in_bus_41(\ccc|a_ram_data_in_bus[41]~q ),
	.a_ram_data_in_bus_25(\ccc|a_ram_data_in_bus[25]~q ),
	.a_ram_data_in_bus_9(\ccc|a_ram_data_in_bus[9]~q ),
	.a_ram_data_in_bus_56(\ccc|a_ram_data_in_bus[56]~q ),
	.a_ram_data_in_bus_40(\ccc|a_ram_data_in_bus[40]~q ),
	.a_ram_data_in_bus_24(\ccc|a_ram_data_in_bus[24]~q ),
	.a_ram_data_in_bus_8(\ccc|a_ram_data_in_bus[8]~q ),
	.a_ram_data_in_bus_63(\ccc|a_ram_data_in_bus[63]~q ),
	.a_ram_data_in_bus_47(\ccc|a_ram_data_in_bus[47]~q ),
	.a_ram_data_in_bus_31(\ccc|a_ram_data_in_bus[31]~q ),
	.a_ram_data_in_bus_15(\ccc|a_ram_data_in_bus[15]~q ),
	.a_ram_data_in_bus_55(\ccc|a_ram_data_in_bus[55]~q ),
	.a_ram_data_in_bus_39(\ccc|a_ram_data_in_bus[39]~q ),
	.a_ram_data_in_bus_23(\ccc|a_ram_data_in_bus[23]~q ),
	.a_ram_data_in_bus_7(\ccc|a_ram_data_in_bus[7]~q ),
	.a_ram_data_in_bus_51(\ccc|a_ram_data_in_bus[51]~q ),
	.a_ram_data_in_bus_35(\ccc|a_ram_data_in_bus[35]~q ),
	.a_ram_data_in_bus_19(\ccc|a_ram_data_in_bus[19]~q ),
	.a_ram_data_in_bus_3(\ccc|a_ram_data_in_bus[3]~q ),
	.a_ram_data_in_bus_53(\ccc|a_ram_data_in_bus[53]~q ),
	.a_ram_data_in_bus_37(\ccc|a_ram_data_in_bus[37]~q ),
	.a_ram_data_in_bus_21(\ccc|a_ram_data_in_bus[21]~q ),
	.a_ram_data_in_bus_5(\ccc|a_ram_data_in_bus[5]~q ),
	.a_ram_data_in_bus_52(\ccc|a_ram_data_in_bus[52]~q ),
	.a_ram_data_in_bus_36(\ccc|a_ram_data_in_bus[36]~q ),
	.a_ram_data_in_bus_20(\ccc|a_ram_data_in_bus[20]~q ),
	.a_ram_data_in_bus_4(\ccc|a_ram_data_in_bus[4]~q ),
	.a_ram_data_in_bus_54(\ccc|a_ram_data_in_bus[54]~q ),
	.a_ram_data_in_bus_38(\ccc|a_ram_data_in_bus[38]~q ),
	.a_ram_data_in_bus_22(\ccc|a_ram_data_in_bus[22]~q ),
	.a_ram_data_in_bus_6(\ccc|a_ram_data_in_bus[6]~q ),
	.a_ram_data_in_bus_50(\ccc|a_ram_data_in_bus[50]~q ),
	.a_ram_data_in_bus_34(\ccc|a_ram_data_in_bus[34]~q ),
	.a_ram_data_in_bus_18(\ccc|a_ram_data_in_bus[18]~q ),
	.a_ram_data_in_bus_2(\ccc|a_ram_data_in_bus[2]~q ),
	.a_ram_data_in_bus_49(\ccc|a_ram_data_in_bus[49]~q ),
	.a_ram_data_in_bus_33(\ccc|a_ram_data_in_bus[33]~q ),
	.a_ram_data_in_bus_17(\ccc|a_ram_data_in_bus[17]~q ),
	.a_ram_data_in_bus_1(\ccc|a_ram_data_in_bus[1]~q ),
	.a_ram_data_in_bus_48(\ccc|a_ram_data_in_bus[48]~q ),
	.a_ram_data_in_bus_32(\ccc|a_ram_data_in_bus[32]~q ),
	.a_ram_data_in_bus_16(\ccc|a_ram_data_in_bus[16]~q ),
	.a_ram_data_in_bus_0(\ccc|a_ram_data_in_bus[0]~q ),
	.clk(clk));

fft_asj_fft_cnt_ctrl_fft_120 ccc(
	.ram_in_reg_1_6(\ram_cxb_wr_data|ram_in_reg[6][1]~q ),
	.ram_in_reg_1_5(\ram_cxb_wr_data|ram_in_reg[5][1]~q ),
	.ram_in_reg_1_4(\ram_cxb_wr_data|ram_in_reg[4][1]~q ),
	.ram_in_reg_1_7(\ram_cxb_wr_data|ram_in_reg[7][1]~q ),
	.ram_in_reg_0_6(\ram_cxb_wr_data|ram_in_reg[6][0]~q ),
	.ram_in_reg_0_5(\ram_cxb_wr_data|ram_in_reg[5][0]~q ),
	.ram_in_reg_0_4(\ram_cxb_wr_data|ram_in_reg[4][0]~q ),
	.ram_in_reg_0_7(\ram_cxb_wr_data|ram_in_reg[7][0]~q ),
	.ram_in_reg_7_6(\ram_cxb_wr_data|ram_in_reg[6][7]~q ),
	.ram_in_reg_7_5(\ram_cxb_wr_data|ram_in_reg[5][7]~q ),
	.ram_in_reg_7_4(\ram_cxb_wr_data|ram_in_reg[4][7]~q ),
	.ram_in_reg_7_7(\ram_cxb_wr_data|ram_in_reg[7][7]~q ),
	.ram_in_reg_6_6(\ram_cxb_wr_data|ram_in_reg[6][6]~q ),
	.ram_in_reg_6_5(\ram_cxb_wr_data|ram_in_reg[5][6]~q ),
	.ram_in_reg_6_4(\ram_cxb_wr_data|ram_in_reg[4][6]~q ),
	.ram_in_reg_6_7(\ram_cxb_wr_data|ram_in_reg[7][6]~q ),
	.ram_in_reg_5_6(\ram_cxb_wr_data|ram_in_reg[6][5]~q ),
	.ram_in_reg_5_5(\ram_cxb_wr_data|ram_in_reg[5][5]~q ),
	.ram_in_reg_5_4(\ram_cxb_wr_data|ram_in_reg[4][5]~q ),
	.ram_in_reg_5_7(\ram_cxb_wr_data|ram_in_reg[7][5]~q ),
	.ram_in_reg_4_6(\ram_cxb_wr_data|ram_in_reg[6][4]~q ),
	.ram_in_reg_4_5(\ram_cxb_wr_data|ram_in_reg[5][4]~q ),
	.ram_in_reg_4_4(\ram_cxb_wr_data|ram_in_reg[4][4]~q ),
	.ram_in_reg_4_7(\ram_cxb_wr_data|ram_in_reg[7][4]~q ),
	.ram_in_reg_3_6(\ram_cxb_wr_data|ram_in_reg[6][3]~q ),
	.ram_in_reg_3_5(\ram_cxb_wr_data|ram_in_reg[5][3]~q ),
	.ram_in_reg_3_4(\ram_cxb_wr_data|ram_in_reg[4][3]~q ),
	.ram_in_reg_3_7(\ram_cxb_wr_data|ram_in_reg[7][3]~q ),
	.ram_in_reg_2_6(\ram_cxb_wr_data|ram_in_reg[6][2]~q ),
	.ram_in_reg_2_5(\ram_cxb_wr_data|ram_in_reg[5][2]~q ),
	.ram_in_reg_2_4(\ram_cxb_wr_data|ram_in_reg[4][2]~q ),
	.ram_in_reg_2_7(\ram_cxb_wr_data|ram_in_reg[7][2]~q ),
	.ram_in_reg_1_2(\ram_cxb_wr_data|ram_in_reg[2][1]~q ),
	.ram_in_reg_1_1(\ram_cxb_wr_data|ram_in_reg[1][1]~q ),
	.ram_in_reg_1_0(\ram_cxb_wr_data|ram_in_reg[0][1]~q ),
	.ram_in_reg_1_3(\ram_cxb_wr_data|ram_in_reg[3][1]~q ),
	.ram_in_reg_0_2(\ram_cxb_wr_data|ram_in_reg[2][0]~q ),
	.ram_in_reg_0_1(\ram_cxb_wr_data|ram_in_reg[1][0]~q ),
	.ram_in_reg_0_0(\ram_cxb_wr_data|ram_in_reg[0][0]~q ),
	.ram_in_reg_0_3(\ram_cxb_wr_data|ram_in_reg[3][0]~q ),
	.ram_in_reg_7_2(\ram_cxb_wr_data|ram_in_reg[2][7]~q ),
	.ram_in_reg_7_1(\ram_cxb_wr_data|ram_in_reg[1][7]~q ),
	.ram_in_reg_7_0(\ram_cxb_wr_data|ram_in_reg[0][7]~q ),
	.ram_in_reg_7_3(\ram_cxb_wr_data|ram_in_reg[3][7]~q ),
	.ram_in_reg_6_2(\ram_cxb_wr_data|ram_in_reg[2][6]~q ),
	.ram_in_reg_6_1(\ram_cxb_wr_data|ram_in_reg[1][6]~q ),
	.ram_in_reg_6_0(\ram_cxb_wr_data|ram_in_reg[0][6]~q ),
	.ram_in_reg_6_3(\ram_cxb_wr_data|ram_in_reg[3][6]~q ),
	.ram_in_reg_5_2(\ram_cxb_wr_data|ram_in_reg[2][5]~q ),
	.ram_in_reg_5_1(\ram_cxb_wr_data|ram_in_reg[1][5]~q ),
	.ram_in_reg_5_0(\ram_cxb_wr_data|ram_in_reg[0][5]~q ),
	.ram_in_reg_5_3(\ram_cxb_wr_data|ram_in_reg[3][5]~q ),
	.ram_in_reg_4_2(\ram_cxb_wr_data|ram_in_reg[2][4]~q ),
	.ram_in_reg_4_1(\ram_cxb_wr_data|ram_in_reg[1][4]~q ),
	.ram_in_reg_4_0(\ram_cxb_wr_data|ram_in_reg[0][4]~q ),
	.ram_in_reg_4_3(\ram_cxb_wr_data|ram_in_reg[3][4]~q ),
	.ram_in_reg_3_2(\ram_cxb_wr_data|ram_in_reg[2][3]~q ),
	.ram_in_reg_3_1(\ram_cxb_wr_data|ram_in_reg[1][3]~q ),
	.ram_in_reg_3_0(\ram_cxb_wr_data|ram_in_reg[0][3]~q ),
	.ram_in_reg_3_3(\ram_cxb_wr_data|ram_in_reg[3][3]~q ),
	.ram_in_reg_2_2(\ram_cxb_wr_data|ram_in_reg[2][2]~q ),
	.ram_in_reg_2_1(\ram_cxb_wr_data|ram_in_reg[1][2]~q ),
	.ram_in_reg_2_0(\ram_cxb_wr_data|ram_in_reg[0][2]~q ),
	.ram_in_reg_2_3(\ram_cxb_wr_data|ram_in_reg[3][2]~q ),
	.q_b_10(\dat_B|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[10] ),
	.q_b_101(\dat_A|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[10] ),
	.q_b_102(\dat_B|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[10] ),
	.q_b_103(\dat_A|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[10] ),
	.q_b_104(\dat_B|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[10] ),
	.q_b_105(\dat_A|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[10] ),
	.q_b_106(\dat_B|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[10] ),
	.q_b_107(\dat_A|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[10] ),
	.q_b_14(\dat_B|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[14] ),
	.q_b_141(\dat_A|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[14] ),
	.q_b_142(\dat_B|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[14] ),
	.q_b_143(\dat_A|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[14] ),
	.q_b_144(\dat_B|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[14] ),
	.q_b_145(\dat_A|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[14] ),
	.q_b_146(\dat_B|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[14] ),
	.q_b_147(\dat_A|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[14] ),
	.q_b_12(\dat_B|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[12] ),
	.q_b_121(\dat_A|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[12] ),
	.q_b_122(\dat_B|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[12] ),
	.q_b_123(\dat_A|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[12] ),
	.q_b_124(\dat_B|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[12] ),
	.q_b_125(\dat_A|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[12] ),
	.q_b_126(\dat_B|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[12] ),
	.q_b_127(\dat_A|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[12] ),
	.q_b_11(\dat_B|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[11] ),
	.q_b_111(\dat_A|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[11] ),
	.q_b_112(\dat_B|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[11] ),
	.q_b_113(\dat_A|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[11] ),
	.q_b_114(\dat_B|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[11] ),
	.q_b_115(\dat_A|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[11] ),
	.q_b_116(\dat_B|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[11] ),
	.q_b_117(\dat_A|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[11] ),
	.q_b_13(\dat_B|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[13] ),
	.q_b_131(\dat_A|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[13] ),
	.q_b_132(\dat_B|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[13] ),
	.q_b_133(\dat_A|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[13] ),
	.q_b_134(\dat_B|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[13] ),
	.q_b_135(\dat_A|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[13] ),
	.q_b_136(\dat_B|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[13] ),
	.q_b_137(\dat_A|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[13] ),
	.q_b_9(\dat_B|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[9] ),
	.q_b_91(\dat_A|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[9] ),
	.q_b_92(\dat_B|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[9] ),
	.q_b_93(\dat_A|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[9] ),
	.q_b_94(\dat_B|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[9] ),
	.q_b_95(\dat_A|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[9] ),
	.q_b_96(\dat_B|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[9] ),
	.q_b_97(\dat_A|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[9] ),
	.q_b_8(\dat_B|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[8] ),
	.q_b_81(\dat_A|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[8] ),
	.q_b_82(\dat_B|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[8] ),
	.q_b_83(\dat_A|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[8] ),
	.q_b_84(\dat_B|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[8] ),
	.q_b_85(\dat_A|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[8] ),
	.q_b_86(\dat_B|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[8] ),
	.q_b_87(\dat_A|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[8] ),
	.q_b_15(\dat_B|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[15] ),
	.q_b_151(\dat_A|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[15] ),
	.q_b_152(\dat_B|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[15] ),
	.q_b_153(\dat_A|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[15] ),
	.q_b_154(\dat_B|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[15] ),
	.q_b_155(\dat_A|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[15] ),
	.q_b_156(\dat_B|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[15] ),
	.q_b_157(\dat_A|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[15] ),
	.q_b_7(\dat_B|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[7] ),
	.q_b_71(\dat_A|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[7] ),
	.q_b_72(\dat_B|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[7] ),
	.q_b_73(\dat_A|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[7] ),
	.q_b_74(\dat_B|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[7] ),
	.q_b_75(\dat_A|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[7] ),
	.q_b_76(\dat_B|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[7] ),
	.q_b_77(\dat_A|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[7] ),
	.q_b_3(\dat_B|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[3] ),
	.q_b_31(\dat_A|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[3] ),
	.q_b_32(\dat_B|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[3] ),
	.q_b_33(\dat_A|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[3] ),
	.q_b_34(\dat_B|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[3] ),
	.q_b_35(\dat_A|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[3] ),
	.q_b_36(\dat_B|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[3] ),
	.q_b_37(\dat_A|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[3] ),
	.q_b_5(\dat_B|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[5] ),
	.q_b_51(\dat_A|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[5] ),
	.q_b_52(\dat_B|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[5] ),
	.q_b_53(\dat_A|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[5] ),
	.q_b_54(\dat_B|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[5] ),
	.q_b_55(\dat_A|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[5] ),
	.q_b_56(\dat_B|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[5] ),
	.q_b_57(\dat_A|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[5] ),
	.q_b_4(\dat_B|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[4] ),
	.q_b_41(\dat_A|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[4] ),
	.q_b_42(\dat_B|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[4] ),
	.q_b_43(\dat_A|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[4] ),
	.q_b_44(\dat_B|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[4] ),
	.q_b_45(\dat_A|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[4] ),
	.q_b_46(\dat_B|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[4] ),
	.q_b_47(\dat_A|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[4] ),
	.q_b_6(\dat_B|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[6] ),
	.q_b_61(\dat_A|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[6] ),
	.q_b_62(\dat_B|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[6] ),
	.q_b_63(\dat_A|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[6] ),
	.q_b_64(\dat_B|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[6] ),
	.q_b_65(\dat_A|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[6] ),
	.q_b_66(\dat_B|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[6] ),
	.q_b_67(\dat_A|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[6] ),
	.q_b_2(\dat_B|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[2] ),
	.q_b_21(\dat_A|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[2] ),
	.q_b_22(\dat_B|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[2] ),
	.q_b_23(\dat_A|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[2] ),
	.q_b_24(\dat_B|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[2] ),
	.q_b_25(\dat_A|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[2] ),
	.q_b_26(\dat_B|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[2] ),
	.q_b_27(\dat_A|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[2] ),
	.q_b_1(\dat_B|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[1] ),
	.q_b_16(\dat_A|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[1] ),
	.q_b_17(\dat_B|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[1] ),
	.q_b_18(\dat_A|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[1] ),
	.q_b_19(\dat_B|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[1] ),
	.q_b_110(\dat_A|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[1] ),
	.q_b_118(\dat_B|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[1] ),
	.q_b_119(\dat_A|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[1] ),
	.q_b_0(\dat_B|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[0] ),
	.q_b_01(\dat_A|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[0] ),
	.q_b_02(\dat_B|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[0] ),
	.q_b_03(\dat_A|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[0] ),
	.q_b_04(\dat_B|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[0] ),
	.q_b_05(\dat_A|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[0] ),
	.q_b_06(\dat_B|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[0] ),
	.q_b_07(\dat_A|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[0] ),
	.global_clock_enable(\global_clock_enable~0_combout ),
	.ram_in_reg_0_01(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[0][0]~q ),
	.ram_in_reg_1_21(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[2][1]~q ),
	.ram_in_reg_2_01(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[0][2]~q ),
	.ram_in_reg_3_21(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[2][3]~q ),
	.ram_in_reg_4_01(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[0][4]~q ),
	.ram_in_reg_5_21(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[2][5]~q ),
	.ram_in_reg_6_01(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[0][6]~q ),
	.ram_in_reg_0_11(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[1][0]~q ),
	.ram_in_reg_1_11(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[1][1]~q ),
	.ram_in_reg_2_11(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[1][2]~q ),
	.ram_in_reg_3_11(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[1][3]~q ),
	.ram_in_reg_4_11(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[1][4]~q ),
	.ram_in_reg_5_11(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[1][5]~q ),
	.ram_in_reg_1_01(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[0][1]~q ),
	.ram_in_reg_3_01(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[0][3]~q ),
	.ram_in_reg_5_01(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[0][5]~q ),
	.ram_in_reg_1_31(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[3][1]~q ),
	.ram_in_reg_3_31(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[3][3]~q ),
	.ram_in_reg_5_31(\gen_wrsw_2:ram_cxb_wr|ram_in_reg[3][5]~q ),
	.ram_data_out0_10(\ccc|ram_data_out0[10]~q ),
	.ram_data_out1_10(\ccc|ram_data_out1[10]~q ),
	.ram_data_out2_10(\ccc|ram_data_out2[10]~q ),
	.ram_data_out3_10(\ccc|ram_data_out3[10]~q ),
	.ram_data_out0_14(\ccc|ram_data_out0[14]~q ),
	.ram_data_out1_14(\ccc|ram_data_out1[14]~q ),
	.ram_data_out2_14(\ccc|ram_data_out2[14]~q ),
	.ram_data_out3_14(\ccc|ram_data_out3[14]~q ),
	.ram_data_out0_12(\ccc|ram_data_out0[12]~q ),
	.ram_data_out1_12(\ccc|ram_data_out1[12]~q ),
	.ram_data_out2_12(\ccc|ram_data_out2[12]~q ),
	.ram_data_out3_12(\ccc|ram_data_out3[12]~q ),
	.ram_data_out0_11(\ccc|ram_data_out0[11]~q ),
	.ram_data_out1_11(\ccc|ram_data_out1[11]~q ),
	.ram_data_out2_11(\ccc|ram_data_out2[11]~q ),
	.ram_data_out3_11(\ccc|ram_data_out3[11]~q ),
	.ram_data_out0_13(\ccc|ram_data_out0[13]~q ),
	.ram_data_out1_13(\ccc|ram_data_out1[13]~q ),
	.ram_data_out2_13(\ccc|ram_data_out2[13]~q ),
	.ram_data_out3_13(\ccc|ram_data_out3[13]~q ),
	.ram_data_out0_9(\ccc|ram_data_out0[9]~q ),
	.ram_data_out1_9(\ccc|ram_data_out1[9]~q ),
	.ram_data_out2_9(\ccc|ram_data_out2[9]~q ),
	.ram_data_out3_9(\ccc|ram_data_out3[9]~q ),
	.ram_data_out0_8(\ccc|ram_data_out0[8]~q ),
	.ram_data_out1_8(\ccc|ram_data_out1[8]~q ),
	.ram_data_out2_8(\ccc|ram_data_out2[8]~q ),
	.ram_data_out3_8(\ccc|ram_data_out3[8]~q ),
	.ram_data_out0_15(\ccc|ram_data_out0[15]~q ),
	.ram_data_out1_15(\ccc|ram_data_out1[15]~q ),
	.ram_data_out2_15(\ccc|ram_data_out2[15]~q ),
	.ram_data_out3_15(\ccc|ram_data_out3[15]~q ),
	.ram_data_out0_7(\ccc|ram_data_out0[7]~q ),
	.ram_data_out1_7(\ccc|ram_data_out1[7]~q ),
	.ram_data_out2_7(\ccc|ram_data_out2[7]~q ),
	.ram_data_out3_7(\ccc|ram_data_out3[7]~q ),
	.ram_data_out0_3(\ccc|ram_data_out0[3]~q ),
	.ram_data_out1_3(\ccc|ram_data_out1[3]~q ),
	.ram_data_out2_3(\ccc|ram_data_out2[3]~q ),
	.ram_data_out3_3(\ccc|ram_data_out3[3]~q ),
	.ram_data_out0_5(\ccc|ram_data_out0[5]~q ),
	.ram_data_out1_5(\ccc|ram_data_out1[5]~q ),
	.ram_data_out2_5(\ccc|ram_data_out2[5]~q ),
	.ram_data_out3_5(\ccc|ram_data_out3[5]~q ),
	.ram_data_out0_4(\ccc|ram_data_out0[4]~q ),
	.ram_data_out1_4(\ccc|ram_data_out1[4]~q ),
	.ram_data_out2_4(\ccc|ram_data_out2[4]~q ),
	.ram_data_out3_4(\ccc|ram_data_out3[4]~q ),
	.ram_data_out0_6(\ccc|ram_data_out0[6]~q ),
	.ram_data_out1_6(\ccc|ram_data_out1[6]~q ),
	.ram_data_out2_6(\ccc|ram_data_out2[6]~q ),
	.ram_data_out3_6(\ccc|ram_data_out3[6]~q ),
	.ram_data_out0_2(\ccc|ram_data_out0[2]~q ),
	.ram_data_out1_2(\ccc|ram_data_out1[2]~q ),
	.ram_data_out2_2(\ccc|ram_data_out2[2]~q ),
	.ram_data_out3_2(\ccc|ram_data_out3[2]~q ),
	.ram_data_out0_1(\ccc|ram_data_out0[1]~q ),
	.ram_data_out1_1(\ccc|ram_data_out1[1]~q ),
	.ram_data_out2_1(\ccc|ram_data_out2[1]~q ),
	.ram_data_out3_1(\ccc|ram_data_out3[1]~q ),
	.ram_data_out0_0(\ccc|ram_data_out0[0]~q ),
	.ram_data_out1_0(\ccc|ram_data_out1[0]~q ),
	.ram_data_out2_0(\ccc|ram_data_out2[0]~q ),
	.ram_data_out3_0(\ccc|ram_data_out3[0]~q ),
	.data_rdy_vec_10(\data_rdy_vec[10]~q ),
	.ram_a_not_b_vec_10(\ram_a_not_b_vec[10]~q ),
	.b_ram_data_in_bus_58(\ccc|b_ram_data_in_bus[58]~q ),
	.wraddress_b_bus_21(\ccc|wraddress_b_bus[21]~q ),
	.wraddress_b_bus_22(\ccc|wraddress_b_bus[22]~q ),
	.wraddress_b_bus_23(\ccc|wraddress_b_bus[23]~q ),
	.wraddress_b_bus_24(\ccc|wraddress_b_bus[24]~q ),
	.wraddress_b_bus_11(\ccc|wraddress_b_bus[11]~q ),
	.wraddress_b_bus_26(\ccc|wraddress_b_bus[26]~q ),
	.wraddress_b_bus_13(\ccc|wraddress_b_bus[13]~q ),
	.rdaddress_b_bus_21(\ccc|rdaddress_b_bus[21]~q ),
	.rdaddress_b_bus_22(\ccc|rdaddress_b_bus[22]~q ),
	.rdaddress_b_bus_23(\ccc|rdaddress_b_bus[23]~q ),
	.rdaddress_b_bus_24(\ccc|rdaddress_b_bus[24]~q ),
	.rdaddress_b_bus_11(\ccc|rdaddress_b_bus[11]~q ),
	.rdaddress_b_bus_26(\ccc|rdaddress_b_bus[26]~q ),
	.rdaddress_b_bus_13(\ccc|rdaddress_b_bus[13]~q ),
	.a_ram_data_in_bus_58(\ccc|a_ram_data_in_bus[58]~q ),
	.wraddress_a_bus_21(\ccc|wraddress_a_bus[21]~q ),
	.wraddress_a_bus_22(\ccc|wraddress_a_bus[22]~q ),
	.wraddress_a_bus_23(\ccc|wraddress_a_bus[23]~q ),
	.wraddress_a_bus_24(\ccc|wraddress_a_bus[24]~q ),
	.wraddress_a_bus_11(\ccc|wraddress_a_bus[11]~q ),
	.wraddress_a_bus_26(\ccc|wraddress_a_bus[26]~q ),
	.wraddress_a_bus_13(\ccc|wraddress_a_bus[13]~q ),
	.rdaddress_a_bus_21(\ccc|rdaddress_a_bus[21]~q ),
	.rdaddress_a_bus_22(\ccc|rdaddress_a_bus[22]~q ),
	.rdaddress_a_bus_23(\ccc|rdaddress_a_bus[23]~q ),
	.rdaddress_a_bus_24(\ccc|rdaddress_a_bus[24]~q ),
	.rdaddress_a_bus_11(\ccc|rdaddress_a_bus[11]~q ),
	.rdaddress_a_bus_26(\ccc|rdaddress_a_bus[26]~q ),
	.rdaddress_a_bus_13(\ccc|rdaddress_a_bus[13]~q ),
	.b_ram_data_in_bus_42(\ccc|b_ram_data_in_bus[42]~q ),
	.wraddress_b_bus_0(\ccc|wraddress_b_bus[0]~q ),
	.wraddress_b_bus_15(\ccc|wraddress_b_bus[15]~q ),
	.wraddress_b_bus_16(\ccc|wraddress_b_bus[16]~q ),
	.wraddress_b_bus_17(\ccc|wraddress_b_bus[17]~q ),
	.wraddress_b_bus_18(\ccc|wraddress_b_bus[18]~q ),
	.wraddress_b_bus_19(\ccc|wraddress_b_bus[19]~q ),
	.rdaddress_b_bus_0(\ccc|rdaddress_b_bus[0]~q ),
	.rdaddress_b_bus_15(\ccc|rdaddress_b_bus[15]~q ),
	.rdaddress_b_bus_16(\ccc|rdaddress_b_bus[16]~q ),
	.rdaddress_b_bus_17(\ccc|rdaddress_b_bus[17]~q ),
	.rdaddress_b_bus_18(\ccc|rdaddress_b_bus[18]~q ),
	.rdaddress_b_bus_19(\ccc|rdaddress_b_bus[19]~q ),
	.a_ram_data_in_bus_42(\ccc|a_ram_data_in_bus[42]~q ),
	.wraddress_a_bus_0(\ccc|wraddress_a_bus[0]~q ),
	.wraddress_a_bus_15(\ccc|wraddress_a_bus[15]~q ),
	.wraddress_a_bus_16(\ccc|wraddress_a_bus[16]~q ),
	.wraddress_a_bus_17(\ccc|wraddress_a_bus[17]~q ),
	.wraddress_a_bus_18(\ccc|wraddress_a_bus[18]~q ),
	.wraddress_a_bus_19(\ccc|wraddress_a_bus[19]~q ),
	.rdaddress_a_bus_0(\ccc|rdaddress_a_bus[0]~q ),
	.rdaddress_a_bus_15(\ccc|rdaddress_a_bus[15]~q ),
	.rdaddress_a_bus_16(\ccc|rdaddress_a_bus[16]~q ),
	.rdaddress_a_bus_17(\ccc|rdaddress_a_bus[17]~q ),
	.rdaddress_a_bus_18(\ccc|rdaddress_a_bus[18]~q ),
	.rdaddress_a_bus_19(\ccc|rdaddress_a_bus[19]~q ),
	.b_ram_data_in_bus_26(\ccc|b_ram_data_in_bus[26]~q ),
	.wraddress_b_bus_8(\ccc|wraddress_b_bus[8]~q ),
	.wraddress_b_bus_10(\ccc|wraddress_b_bus[10]~q ),
	.wraddress_b_bus_12(\ccc|wraddress_b_bus[12]~q ),
	.rdaddress_b_bus_8(\ccc|rdaddress_b_bus[8]~q ),
	.rdaddress_b_bus_10(\ccc|rdaddress_b_bus[10]~q ),
	.rdaddress_b_bus_12(\ccc|rdaddress_b_bus[12]~q ),
	.a_ram_data_in_bus_26(\ccc|a_ram_data_in_bus[26]~q ),
	.wraddress_a_bus_8(\ccc|wraddress_a_bus[8]~q ),
	.wraddress_a_bus_10(\ccc|wraddress_a_bus[10]~q ),
	.wraddress_a_bus_12(\ccc|wraddress_a_bus[12]~q ),
	.rdaddress_a_bus_8(\ccc|rdaddress_a_bus[8]~q ),
	.rdaddress_a_bus_10(\ccc|rdaddress_a_bus[10]~q ),
	.rdaddress_a_bus_12(\ccc|rdaddress_a_bus[12]~q ),
	.b_ram_data_in_bus_10(\ccc|b_ram_data_in_bus[10]~q ),
	.wraddress_b_bus_1(\ccc|wraddress_b_bus[1]~q ),
	.wraddress_b_bus_3(\ccc|wraddress_b_bus[3]~q ),
	.wraddress_b_bus_5(\ccc|wraddress_b_bus[5]~q ),
	.rdaddress_b_bus_1(\ccc|rdaddress_b_bus[1]~q ),
	.rdaddress_b_bus_3(\ccc|rdaddress_b_bus[3]~q ),
	.rdaddress_b_bus_5(\ccc|rdaddress_b_bus[5]~q ),
	.a_ram_data_in_bus_10(\ccc|a_ram_data_in_bus[10]~q ),
	.wraddress_a_bus_1(\ccc|wraddress_a_bus[1]~q ),
	.wraddress_a_bus_3(\ccc|wraddress_a_bus[3]~q ),
	.wraddress_a_bus_5(\ccc|wraddress_a_bus[5]~q ),
	.rdaddress_a_bus_1(\ccc|rdaddress_a_bus[1]~q ),
	.rdaddress_a_bus_3(\ccc|rdaddress_a_bus[3]~q ),
	.rdaddress_a_bus_5(\ccc|rdaddress_a_bus[5]~q ),
	.b_ram_data_in_bus_62(\ccc|b_ram_data_in_bus[62]~q ),
	.a_ram_data_in_bus_62(\ccc|a_ram_data_in_bus[62]~q ),
	.b_ram_data_in_bus_46(\ccc|b_ram_data_in_bus[46]~q ),
	.a_ram_data_in_bus_46(\ccc|a_ram_data_in_bus[46]~q ),
	.b_ram_data_in_bus_30(\ccc|b_ram_data_in_bus[30]~q ),
	.a_ram_data_in_bus_30(\ccc|a_ram_data_in_bus[30]~q ),
	.b_ram_data_in_bus_14(\ccc|b_ram_data_in_bus[14]~q ),
	.a_ram_data_in_bus_14(\ccc|a_ram_data_in_bus[14]~q ),
	.b_ram_data_in_bus_60(\ccc|b_ram_data_in_bus[60]~q ),
	.a_ram_data_in_bus_60(\ccc|a_ram_data_in_bus[60]~q ),
	.b_ram_data_in_bus_44(\ccc|b_ram_data_in_bus[44]~q ),
	.a_ram_data_in_bus_44(\ccc|a_ram_data_in_bus[44]~q ),
	.b_ram_data_in_bus_28(\ccc|b_ram_data_in_bus[28]~q ),
	.a_ram_data_in_bus_28(\ccc|a_ram_data_in_bus[28]~q ),
	.b_ram_data_in_bus_12(\ccc|b_ram_data_in_bus[12]~q ),
	.a_ram_data_in_bus_12(\ccc|a_ram_data_in_bus[12]~q ),
	.b_ram_data_in_bus_59(\ccc|b_ram_data_in_bus[59]~q ),
	.a_ram_data_in_bus_59(\ccc|a_ram_data_in_bus[59]~q ),
	.b_ram_data_in_bus_43(\ccc|b_ram_data_in_bus[43]~q ),
	.a_ram_data_in_bus_43(\ccc|a_ram_data_in_bus[43]~q ),
	.b_ram_data_in_bus_27(\ccc|b_ram_data_in_bus[27]~q ),
	.a_ram_data_in_bus_27(\ccc|a_ram_data_in_bus[27]~q ),
	.b_ram_data_in_bus_11(\ccc|b_ram_data_in_bus[11]~q ),
	.a_ram_data_in_bus_11(\ccc|a_ram_data_in_bus[11]~q ),
	.b_ram_data_in_bus_61(\ccc|b_ram_data_in_bus[61]~q ),
	.a_ram_data_in_bus_61(\ccc|a_ram_data_in_bus[61]~q ),
	.b_ram_data_in_bus_45(\ccc|b_ram_data_in_bus[45]~q ),
	.a_ram_data_in_bus_45(\ccc|a_ram_data_in_bus[45]~q ),
	.b_ram_data_in_bus_29(\ccc|b_ram_data_in_bus[29]~q ),
	.a_ram_data_in_bus_29(\ccc|a_ram_data_in_bus[29]~q ),
	.b_ram_data_in_bus_13(\ccc|b_ram_data_in_bus[13]~q ),
	.a_ram_data_in_bus_13(\ccc|a_ram_data_in_bus[13]~q ),
	.b_ram_data_in_bus_57(\ccc|b_ram_data_in_bus[57]~q ),
	.a_ram_data_in_bus_57(\ccc|a_ram_data_in_bus[57]~q ),
	.b_ram_data_in_bus_41(\ccc|b_ram_data_in_bus[41]~q ),
	.a_ram_data_in_bus_41(\ccc|a_ram_data_in_bus[41]~q ),
	.b_ram_data_in_bus_25(\ccc|b_ram_data_in_bus[25]~q ),
	.a_ram_data_in_bus_25(\ccc|a_ram_data_in_bus[25]~q ),
	.b_ram_data_in_bus_9(\ccc|b_ram_data_in_bus[9]~q ),
	.a_ram_data_in_bus_9(\ccc|a_ram_data_in_bus[9]~q ),
	.b_ram_data_in_bus_56(\ccc|b_ram_data_in_bus[56]~q ),
	.a_ram_data_in_bus_56(\ccc|a_ram_data_in_bus[56]~q ),
	.b_ram_data_in_bus_40(\ccc|b_ram_data_in_bus[40]~q ),
	.a_ram_data_in_bus_40(\ccc|a_ram_data_in_bus[40]~q ),
	.b_ram_data_in_bus_24(\ccc|b_ram_data_in_bus[24]~q ),
	.a_ram_data_in_bus_24(\ccc|a_ram_data_in_bus[24]~q ),
	.b_ram_data_in_bus_8(\ccc|b_ram_data_in_bus[8]~q ),
	.a_ram_data_in_bus_8(\ccc|a_ram_data_in_bus[8]~q ),
	.b_ram_data_in_bus_63(\ccc|b_ram_data_in_bus[63]~q ),
	.a_ram_data_in_bus_63(\ccc|a_ram_data_in_bus[63]~q ),
	.b_ram_data_in_bus_47(\ccc|b_ram_data_in_bus[47]~q ),
	.a_ram_data_in_bus_47(\ccc|a_ram_data_in_bus[47]~q ),
	.b_ram_data_in_bus_31(\ccc|b_ram_data_in_bus[31]~q ),
	.a_ram_data_in_bus_31(\ccc|a_ram_data_in_bus[31]~q ),
	.b_ram_data_in_bus_15(\ccc|b_ram_data_in_bus[15]~q ),
	.a_ram_data_in_bus_15(\ccc|a_ram_data_in_bus[15]~q ),
	.b_ram_data_in_bus_55(\ccc|b_ram_data_in_bus[55]~q ),
	.a_ram_data_in_bus_55(\ccc|a_ram_data_in_bus[55]~q ),
	.b_ram_data_in_bus_39(\ccc|b_ram_data_in_bus[39]~q ),
	.a_ram_data_in_bus_39(\ccc|a_ram_data_in_bus[39]~q ),
	.b_ram_data_in_bus_23(\ccc|b_ram_data_in_bus[23]~q ),
	.a_ram_data_in_bus_23(\ccc|a_ram_data_in_bus[23]~q ),
	.b_ram_data_in_bus_7(\ccc|b_ram_data_in_bus[7]~q ),
	.a_ram_data_in_bus_7(\ccc|a_ram_data_in_bus[7]~q ),
	.b_ram_data_in_bus_51(\ccc|b_ram_data_in_bus[51]~q ),
	.a_ram_data_in_bus_51(\ccc|a_ram_data_in_bus[51]~q ),
	.b_ram_data_in_bus_35(\ccc|b_ram_data_in_bus[35]~q ),
	.a_ram_data_in_bus_35(\ccc|a_ram_data_in_bus[35]~q ),
	.b_ram_data_in_bus_19(\ccc|b_ram_data_in_bus[19]~q ),
	.a_ram_data_in_bus_19(\ccc|a_ram_data_in_bus[19]~q ),
	.b_ram_data_in_bus_3(\ccc|b_ram_data_in_bus[3]~q ),
	.a_ram_data_in_bus_3(\ccc|a_ram_data_in_bus[3]~q ),
	.b_ram_data_in_bus_53(\ccc|b_ram_data_in_bus[53]~q ),
	.a_ram_data_in_bus_53(\ccc|a_ram_data_in_bus[53]~q ),
	.b_ram_data_in_bus_37(\ccc|b_ram_data_in_bus[37]~q ),
	.a_ram_data_in_bus_37(\ccc|a_ram_data_in_bus[37]~q ),
	.b_ram_data_in_bus_21(\ccc|b_ram_data_in_bus[21]~q ),
	.a_ram_data_in_bus_21(\ccc|a_ram_data_in_bus[21]~q ),
	.b_ram_data_in_bus_5(\ccc|b_ram_data_in_bus[5]~q ),
	.a_ram_data_in_bus_5(\ccc|a_ram_data_in_bus[5]~q ),
	.b_ram_data_in_bus_52(\ccc|b_ram_data_in_bus[52]~q ),
	.a_ram_data_in_bus_52(\ccc|a_ram_data_in_bus[52]~q ),
	.b_ram_data_in_bus_36(\ccc|b_ram_data_in_bus[36]~q ),
	.a_ram_data_in_bus_36(\ccc|a_ram_data_in_bus[36]~q ),
	.b_ram_data_in_bus_20(\ccc|b_ram_data_in_bus[20]~q ),
	.a_ram_data_in_bus_20(\ccc|a_ram_data_in_bus[20]~q ),
	.b_ram_data_in_bus_4(\ccc|b_ram_data_in_bus[4]~q ),
	.a_ram_data_in_bus_4(\ccc|a_ram_data_in_bus[4]~q ),
	.b_ram_data_in_bus_54(\ccc|b_ram_data_in_bus[54]~q ),
	.a_ram_data_in_bus_54(\ccc|a_ram_data_in_bus[54]~q ),
	.b_ram_data_in_bus_38(\ccc|b_ram_data_in_bus[38]~q ),
	.a_ram_data_in_bus_38(\ccc|a_ram_data_in_bus[38]~q ),
	.b_ram_data_in_bus_22(\ccc|b_ram_data_in_bus[22]~q ),
	.a_ram_data_in_bus_22(\ccc|a_ram_data_in_bus[22]~q ),
	.b_ram_data_in_bus_6(\ccc|b_ram_data_in_bus[6]~q ),
	.a_ram_data_in_bus_6(\ccc|a_ram_data_in_bus[6]~q ),
	.b_ram_data_in_bus_50(\ccc|b_ram_data_in_bus[50]~q ),
	.a_ram_data_in_bus_50(\ccc|a_ram_data_in_bus[50]~q ),
	.b_ram_data_in_bus_34(\ccc|b_ram_data_in_bus[34]~q ),
	.a_ram_data_in_bus_34(\ccc|a_ram_data_in_bus[34]~q ),
	.b_ram_data_in_bus_18(\ccc|b_ram_data_in_bus[18]~q ),
	.a_ram_data_in_bus_18(\ccc|a_ram_data_in_bus[18]~q ),
	.b_ram_data_in_bus_2(\ccc|b_ram_data_in_bus[2]~q ),
	.a_ram_data_in_bus_2(\ccc|a_ram_data_in_bus[2]~q ),
	.b_ram_data_in_bus_49(\ccc|b_ram_data_in_bus[49]~q ),
	.a_ram_data_in_bus_49(\ccc|a_ram_data_in_bus[49]~q ),
	.b_ram_data_in_bus_33(\ccc|b_ram_data_in_bus[33]~q ),
	.a_ram_data_in_bus_33(\ccc|a_ram_data_in_bus[33]~q ),
	.b_ram_data_in_bus_17(\ccc|b_ram_data_in_bus[17]~q ),
	.a_ram_data_in_bus_17(\ccc|a_ram_data_in_bus[17]~q ),
	.b_ram_data_in_bus_1(\ccc|b_ram_data_in_bus[1]~q ),
	.a_ram_data_in_bus_1(\ccc|a_ram_data_in_bus[1]~q ),
	.b_ram_data_in_bus_48(\ccc|b_ram_data_in_bus[48]~q ),
	.a_ram_data_in_bus_48(\ccc|a_ram_data_in_bus[48]~q ),
	.b_ram_data_in_bus_32(\ccc|b_ram_data_in_bus[32]~q ),
	.a_ram_data_in_bus_32(\ccc|a_ram_data_in_bus[32]~q ),
	.b_ram_data_in_bus_16(\ccc|b_ram_data_in_bus[16]~q ),
	.a_ram_data_in_bus_16(\ccc|a_ram_data_in_bus[16]~q ),
	.b_ram_data_in_bus_0(\ccc|b_ram_data_in_bus[0]~q ),
	.a_ram_data_in_bus_0(\ccc|a_ram_data_in_bus[0]~q ),
	.ram_a_not_b_vec_1(\ram_a_not_b_vec[1]~q ),
	.data_in_r_2(\writer|data_in_r[2]~q ),
	.wr_address_i_int_0(\writer|wr_address_i_int[0]~q ),
	.wr_address_i_int_1(\writer|wr_address_i_int[1]~q ),
	.wr_address_i_int_2(\writer|wr_address_i_int[2]~q ),
	.wr_address_i_int_3(\writer|wr_address_i_int[3]~q ),
	.wr_address_i_int_4(\writer|wr_address_i_int[4]~q ),
	.wr_address_i_int_5(\writer|wr_address_i_int[5]~q ),
	.wr_address_i_int_6(\writer|wr_address_i_int[6]~q ),
	.ram_a_not_b_vec_7(\ram_a_not_b_vec[7]~q ),
	.ram_in_reg_0_02(\ram_cxb_rd|ram_in_reg[0][0]~q ),
	.ram_in_reg_1_02(\ram_cxb_rd|ram_in_reg[0][1]~q ),
	.ram_in_reg_2_02(\ram_cxb_rd|ram_in_reg[0][2]~q ),
	.ram_in_reg_3_02(\ram_cxb_rd|ram_in_reg[0][3]~q ),
	.ram_in_reg_4_02(\ram_cxb_rd|ram_in_reg[0][4]~q ),
	.ram_in_reg_5_02(\ram_cxb_rd|ram_in_reg[0][5]~q ),
	.tdl_arr_6_1(\gen_wrsw_2:k_delay|tdl_arr[1][6]~q ),
	.ram_in_reg_0_12(\ram_cxb_rd|ram_in_reg[1][0]~q ),
	.ram_in_reg_1_12(\ram_cxb_rd|ram_in_reg[1][1]~q ),
	.ram_in_reg_2_12(\ram_cxb_rd|ram_in_reg[1][2]~q ),
	.ram_in_reg_3_12(\ram_cxb_rd|ram_in_reg[1][3]~q ),
	.ram_in_reg_4_12(\ram_cxb_rd|ram_in_reg[1][4]~q ),
	.ram_in_reg_5_12(\ram_cxb_rd|ram_in_reg[1][5]~q ),
	.ram_in_reg_1_22(\ram_cxb_rd|ram_in_reg[2][1]~q ),
	.ram_in_reg_3_22(\ram_cxb_rd|ram_in_reg[2][3]~q ),
	.ram_in_reg_5_22(\ram_cxb_rd|ram_in_reg[2][5]~q ),
	.ram_in_reg_1_32(\ram_cxb_rd|ram_in_reg[3][1]~q ),
	.ram_in_reg_3_32(\ram_cxb_rd|ram_in_reg[3][3]~q ),
	.ram_in_reg_5_32(\ram_cxb_rd|ram_in_reg[3][5]~q ),
	.data_in_r_6(\writer|data_in_r[6]~q ),
	.data_in_r_4(\writer|data_in_r[4]~q ),
	.data_in_r_3(\writer|data_in_r[3]~q ),
	.data_in_r_5(\writer|data_in_r[5]~q ),
	.data_in_r_1(\writer|data_in_r[1]~q ),
	.data_in_r_0(\writer|data_in_r[0]~q ),
	.data_in_r_7(\writer|data_in_r[7]~q ),
	.data_in_i_7(\writer|data_in_i[7]~q ),
	.data_in_i_3(\writer|data_in_i[3]~q ),
	.data_in_i_5(\writer|data_in_i[5]~q ),
	.data_in_i_4(\writer|data_in_i[4]~q ),
	.data_in_i_6(\writer|data_in_i[6]~q ),
	.data_in_i_2(\writer|data_in_i[2]~q ),
	.data_in_i_1(\writer|data_in_i[1]~q ),
	.data_in_i_0(\writer|data_in_i[0]~q ),
	.clk(clk));

fft_asj_fft_in_write_sgl_fft_120 writer(
	.data_rdy_int1(\writer|data_rdy_int~q ),
	.wren_0(\writer|wren[0]~q ),
	.wren_1(\writer|wren[1]~q ),
	.wren_2(\writer|wren[2]~q ),
	.wren_3(\writer|wren[3]~q ),
	.core_real_in_2(\core_real_in[2]~q ),
	.core_real_in_6(\core_real_in[6]~q ),
	.core_real_in_4(\core_real_in[4]~q ),
	.core_real_in_3(\core_real_in[3]~q ),
	.core_real_in_5(\core_real_in[5]~q ),
	.core_real_in_1(\core_real_in[1]~q ),
	.core_real_in_0(\core_real_in[0]~q ),
	.core_real_in_7(\core_real_in[7]~q ),
	.core_imag_in_7(\core_imag_in[7]~q ),
	.core_imag_in_3(\core_imag_in[3]~q ),
	.core_imag_in_5(\core_imag_in[5]~q ),
	.core_imag_in_4(\core_imag_in[4]~q ),
	.core_imag_in_6(\core_imag_in[6]~q ),
	.core_imag_in_2(\core_imag_in[2]~q ),
	.core_imag_in_1(\core_imag_in[1]~q ),
	.core_imag_in_0(\core_imag_in[0]~q ),
	.anb1(\writer|anb~q ),
	.send_sop_s(\auk_dsp_atlantic_sink_1|send_sop_s~q ),
	.global_clock_enable(\global_clock_enable~0_combout ),
	.next_block1(\writer|next_block~q ),
	.data_in_r_2(\writer|data_in_r[2]~q ),
	.wr_address_i_int_0(\writer|wr_address_i_int[0]~q ),
	.wr_address_i_int_1(\writer|wr_address_i_int[1]~q ),
	.wr_address_i_int_2(\writer|wr_address_i_int[2]~q ),
	.wr_address_i_int_3(\writer|wr_address_i_int[3]~q ),
	.wr_address_i_int_4(\writer|wr_address_i_int[4]~q ),
	.wr_address_i_int_5(\writer|wr_address_i_int[5]~q ),
	.wr_address_i_int_6(\writer|wr_address_i_int[6]~q ),
	.data_in_r_6(\writer|data_in_r[6]~q ),
	.data_in_r_4(\writer|data_in_r[4]~q ),
	.data_in_r_3(\writer|data_in_r[3]~q ),
	.data_in_r_5(\writer|data_in_r[5]~q ),
	.data_in_r_1(\writer|data_in_r[1]~q ),
	.data_in_r_0(\writer|data_in_r[0]~q ),
	.data_in_r_7(\writer|data_in_r[7]~q ),
	.data_in_i_7(\writer|data_in_i[7]~q ),
	.data_in_i_3(\writer|data_in_i[3]~q ),
	.data_in_i_5(\writer|data_in_i[5]~q ),
	.data_in_i_4(\writer|data_in_i[4]~q ),
	.data_in_i_6(\writer|data_in_i[6]~q ),
	.data_in_i_2(\writer|data_in_i[2]~q ),
	.data_in_i_1(\writer|data_in_i[1]~q ),
	.data_in_i_0(\writer|data_in_i[0]~q ),
	.clk(clk),
	.reset_n(reset_n));

fft_asj_fft_wrengen_fft_120 sel_we(
	.global_clock_enable(\global_clock_enable~0_combout ),
	.wc_i1(\sel_we|wc_i~q ),
	.wd_i1(\sel_we|wd_i~q ),
	.ram_a_not_b_vec_26(\ram_a_not_b_vec[26]~q ),
	.p_cd_en_2(\p_cd_en[2]~q ),
	.p_cd_en_0(\p_cd_en[0]~q ),
	.p_cd_en_1(\p_cd_en[1]~q ),
	.clk(clk),
	.reset_n(reset_n));

fft_asj_fft_tdl_bit_rst_fft_120_6 delay_ctrl_np(
	.global_clock_enable(\global_clock_enable~0_combout ),
	.next_pass_i(\gen_gt256_mk:ctrl|next_pass_i~q ),
	.tdl_arr_5(\delay_ctrl_np|tdl_arr[5]~q ),
	.next_pass_vec_2(\gen_dft_2:bfpdft|next_pass_vec[2]~q ),
	.tdl_arr_9(\delay_ctrl_np|tdl_arr[9]~q ),
	.clk(clk),
	.reset_n(reset_n));

fft_asj_fft_m_k_counter_fft_120 \gen_gt256_mk:ctrl (
	.blk_done_int1(\gen_gt256_mk:ctrl|blk_done_int~q ),
	.source_valid_ctrl_sop(\source_valid_ctrl_sop~1_combout ),
	.stall_reg(\auk_dsp_interface_controller_1|stall_reg~q ),
	.source_stall_int_d(\auk_dsp_atlantic_source_1|source_stall_int_d~q ),
	.global_clock_enable(\global_clock_enable~0_combout ),
	.p_2(\gen_gt256_mk:ctrl|p[2]~q ),
	.p_0(\gen_gt256_mk:ctrl|p[0]~q ),
	.p_1(\gen_gt256_mk:ctrl|p[1]~q ),
	.tdl_arr_4(\gen_dft_2:bfpdft|gen_cont:delay_next_blk|tdl_arr[4]~q ),
	.data_rdy_vec_4(\data_rdy_vec[4]~q ),
	.next_pass_i1(\gen_gt256_mk:ctrl|next_pass_i~q ),
	.Equal0(\gen_gt256_mk:ctrl|Equal0~0_combout ),
	.tdl_arr_3(\gen_dft_2:bfpdft|gen_cont:delay_next_blk|tdl_arr[3]~q ),
	.k_count_0(\gen_gt256_mk:ctrl|k_count[0]~q ),
	.k_count_2(\gen_gt256_mk:ctrl|k_count[2]~q ),
	.k_count_4(\gen_gt256_mk:ctrl|k_count[4]~q ),
	.k_count_1(\gen_gt256_mk:ctrl|k_count[1]~q ),
	.k_count_3(\gen_gt256_mk:ctrl|k_count[3]~q ),
	.k_count_5(\gen_gt256_mk:ctrl|k_count[5]~q ),
	.k_count_6(\gen_gt256_mk:ctrl|k_count[6]~q ),
	.clk(clk),
	.reset_n(reset_n));

fft_auk_dspip_avalon_streaming_controller_fft_120 auk_dsp_interface_controller_1(
	.at_source_valid_s(at_source_valid_s),
	.source_packet_error_0(\auk_dsp_interface_controller_1|source_packet_error[0]~q ),
	.source_packet_error_1(\auk_dsp_interface_controller_1|source_packet_error[1]~q ),
	.valid_ctrl_int(\auk_dsp_atlantic_source_1|valid_ctrl_int~q ),
	.master_sink_ena(\master_sink_ena~q ),
	.source_stall_reg1(\auk_dsp_interface_controller_1|source_stall_reg~q ),
	.sink_stall_reg1(\auk_dsp_interface_controller_1|sink_stall_reg~q ),
	.sink_ready_ctrl(\auk_dsp_interface_controller_1|sink_ready_ctrl~0_combout ),
	.sink_stall(\auk_dsp_atlantic_sink_1|sink_stall~combout ),
	.packet_error_s_0(\auk_dsp_atlantic_sink_1|packet_error_s[0]~q ),
	.packet_error_s_1(\auk_dsp_atlantic_sink_1|packet_error_s[1]~q ),
	.Mux3(\auk_dsp_atlantic_source_1|Mux3~0_combout ),
	.stall_reg1(\auk_dsp_interface_controller_1|stall_reg~q ),
	.Mux0(\auk_dsp_atlantic_source_1|Mux0~0_combout ),
	.Mux01(\auk_dsp_atlantic_source_1|Mux0~2_combout ),
	.clk(clk),
	.reset_n(reset_n),
	.source_ready(source_ready));

fft_auk_dspip_avalon_streaming_source_fft_120 auk_dsp_atlantic_source_1(
	.data_count({\data_count_sig[8]~q ,\data_count_sig[7]~q ,\data_count_sig[6]~q ,\data_count_sig[5]~q ,\data_count_sig[4]~q ,\data_count_sig[3]~q ,\data_count_sig[2]~q ,\data_count_sig[1]~q ,\data_count_sig[0]~q }),
	.at_source_error_0(at_source_error_0),
	.at_source_error_1(at_source_error_1),
	.at_source_sop_s1(at_source_sop_s),
	.at_source_eop_s1(at_source_eop_s),
	.at_source_valid_s1(at_source_valid_s),
	.at_source_data_0(at_source_data_0),
	.at_source_data_1(at_source_data_1),
	.at_source_data_2(at_source_data_2),
	.at_source_data_3(at_source_data_3),
	.at_source_data_4(at_source_data_4),
	.at_source_data_5(at_source_data_5),
	.at_source_data_14(at_source_data_14),
	.at_source_data_15(at_source_data_15),
	.at_source_data_16(at_source_data_16),
	.at_source_data_17(at_source_data_17),
	.at_source_data_18(at_source_data_18),
	.at_source_data_19(at_source_data_19),
	.at_source_data_20(at_source_data_20),
	.at_source_data_21(at_source_data_21),
	.at_source_data_6(at_source_data_6),
	.at_source_data_7(at_source_data_7),
	.at_source_data_8(at_source_data_8),
	.at_source_data_9(at_source_data_9),
	.at_source_data_10(at_source_data_10),
	.at_source_data_11(at_source_data_11),
	.at_source_data_12(at_source_data_12),
	.at_source_data_13(at_source_data_13),
	.source_packet_error_0(\auk_dsp_interface_controller_1|source_packet_error[0]~q ),
	.source_packet_error_1(\auk_dsp_interface_controller_1|source_packet_error[1]~q ),
	.valid_ctrl_int2(\auk_dsp_atlantic_source_1|valid_ctrl_int~q ),
	.source_stall_reg(\auk_dsp_interface_controller_1|source_stall_reg~q ),
	.master_source_ena(\master_source_ena~q ),
	.source_valid_ctrl_sop(\source_valid_ctrl_sop~0_combout ),
	.Mux3(\auk_dsp_atlantic_source_1|Mux3~0_combout ),
	.source_valid_ctrl_sop1(\source_valid_ctrl_sop~1_combout ),
	.stall_reg(\auk_dsp_interface_controller_1|stall_reg~q ),
	.source_stall_int_d1(\auk_dsp_atlantic_source_1|source_stall_int_d~q ),
	.data({\fft_real_out[7]~q ,\fft_real_out[6]~q ,\fft_real_out[5]~q ,\fft_real_out[4]~q ,\fft_real_out[3]~q ,\fft_real_out[2]~q ,\fft_real_out[1]~q ,\fft_real_out[0]~q ,\fft_imag_out[7]~q ,\fft_imag_out[6]~q ,\fft_imag_out[5]~q ,\fft_imag_out[4]~q ,\fft_imag_out[3]~q ,
\fft_imag_out[2]~q ,\fft_imag_out[1]~q ,\fft_imag_out[0]~q ,\exponent_out[5]~q ,\exponent_out[4]~q ,\exponent_out[3]~q ,\exponent_out[2]~q ,\exponent_out[1]~q ,\exponent_out[0]~q }),
	.Mux0(\auk_dsp_atlantic_source_1|Mux0~0_combout ),
	.Mux01(\auk_dsp_atlantic_source_1|Mux0~2_combout ),
	.clk(clk),
	.reset_n(reset_n),
	.source_ready(source_ready));

fft_auk_dspip_avalon_streaming_sink_fft_120 auk_dsp_atlantic_sink_1(
	.q_b_2(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.q_b_10(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[10] ),
	.q_b_6(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.q_b_14(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[14] ),
	.q_b_4(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.q_b_12(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[12] ),
	.q_b_3(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.q_b_11(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[11] ),
	.q_b_5(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.q_b_13(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[13] ),
	.q_b_1(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.q_b_9(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[9] ),
	.q_b_0(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.q_b_8(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[8] ),
	.q_b_7(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.q_b_15(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[15] ),
	.at_sink_ready_s1(at_sink_ready_s),
	.sink_ready_ctrl(\auk_dsp_interface_controller_1|sink_ready_ctrl~0_combout ),
	.sink_stall1(\auk_dsp_atlantic_sink_1|sink_stall~combout ),
	.packet_error_s_0(\auk_dsp_atlantic_sink_1|packet_error_s[0]~q ),
	.packet_error_s_1(\auk_dsp_atlantic_sink_1|packet_error_s[1]~q ),
	.send_sop_s1(\auk_dsp_atlantic_sink_1|send_sop_s~q ),
	.send_eop_s1(\auk_dsp_atlantic_sink_1|send_eop_s~q ),
	.clk(clk),
	.reset_n(reset_n),
	.sink_error_0(sink_error_0),
	.sink_error_1(sink_error_1),
	.sink_valid(sink_valid),
	.sink_sop(sink_sop),
	.sink_eop(sink_eop),
	.at_sink_data({sink_real[7],sink_real[6],sink_real[5],sink_real[4],sink_real[3],sink_real[2],sink_real[1],sink_real[0],sink_imag[7],sink_imag[6],sink_imag[5],sink_imag[4],sink_imag[3],sink_imag[2],sink_imag[1],sink_imag[0]}));

dffeas \data_count_sig[3] (
	.clk(clk),
	.d(\data_count_sig[3]~15_combout ),
	.asdata(GND_port),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\data_count_sig[0]~18_combout ),
	.ena(\data_count_sig[0]~20_combout ),
	.q(\data_count_sig[3]~q ),
	.prn(vcc));
defparam \data_count_sig[3] .is_wysiwyg = "true";
defparam \data_count_sig[3] .power_up = "low";

dffeas \data_count_sig[2] (
	.clk(clk),
	.d(\data_count_sig[2]~13_combout ),
	.asdata(GND_port),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\data_count_sig[0]~18_combout ),
	.ena(\data_count_sig[0]~20_combout ),
	.q(\data_count_sig[2]~q ),
	.prn(vcc));
defparam \data_count_sig[2] .is_wysiwyg = "true";
defparam \data_count_sig[2] .power_up = "low";

dffeas \data_count_sig[1] (
	.clk(clk),
	.d(\data_count_sig[1]~11_combout ),
	.asdata(GND_port),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\data_count_sig[0]~18_combout ),
	.ena(\data_count_sig[0]~20_combout ),
	.q(\data_count_sig[1]~q ),
	.prn(vcc));
defparam \data_count_sig[1] .is_wysiwyg = "true";
defparam \data_count_sig[1] .power_up = "low";

dffeas \data_count_sig[0] (
	.clk(clk),
	.d(\data_count_sig[0]~9_combout ),
	.asdata(\master_source_sop~q ),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\data_count_sig[0]~18_combout ),
	.ena(\data_count_sig[0]~20_combout ),
	.q(\data_count_sig[0]~q ),
	.prn(vcc));
defparam \data_count_sig[0] .is_wysiwyg = "true";
defparam \data_count_sig[0] .power_up = "low";

dffeas \data_count_sig[6] (
	.clk(clk),
	.d(\data_count_sig[6]~25_combout ),
	.asdata(GND_port),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\data_count_sig[0]~18_combout ),
	.ena(\data_count_sig[0]~20_combout ),
	.q(\data_count_sig[6]~q ),
	.prn(vcc));
defparam \data_count_sig[6] .is_wysiwyg = "true";
defparam \data_count_sig[6] .power_up = "low";

dffeas \data_count_sig[7] (
	.clk(clk),
	.d(\data_count_sig[7]~27_combout ),
	.asdata(GND_port),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\data_count_sig[0]~18_combout ),
	.ena(\data_count_sig[0]~20_combout ),
	.q(\data_count_sig[7]~q ),
	.prn(vcc));
defparam \data_count_sig[7] .is_wysiwyg = "true";
defparam \data_count_sig[7] .power_up = "low";

dffeas \data_count_sig[4] (
	.clk(clk),
	.d(\data_count_sig[4]~21_combout ),
	.asdata(GND_port),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\data_count_sig[0]~18_combout ),
	.ena(\data_count_sig[0]~20_combout ),
	.q(\data_count_sig[4]~q ),
	.prn(vcc));
defparam \data_count_sig[4] .is_wysiwyg = "true";
defparam \data_count_sig[4] .power_up = "low";

dffeas \data_count_sig[5] (
	.clk(clk),
	.d(\data_count_sig[5]~23_combout ),
	.asdata(GND_port),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\data_count_sig[0]~18_combout ),
	.ena(\data_count_sig[0]~20_combout ),
	.q(\data_count_sig[5]~q ),
	.prn(vcc));
defparam \data_count_sig[5] .is_wysiwyg = "true";
defparam \data_count_sig[5] .power_up = "low";

dffeas \data_count_sig[8] (
	.clk(clk),
	.d(\data_count_sig[8]~29_combout ),
	.asdata(GND_port),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\data_count_sig[0]~18_combout ),
	.ena(\data_count_sig[0]~20_combout ),
	.q(\data_count_sig[8]~q ),
	.prn(vcc));
defparam \data_count_sig[8] .is_wysiwyg = "true";
defparam \data_count_sig[8] .power_up = "low";

cycloneiii_lcell_comb \data_count_sig[0]~9 (
	.dataa(\data_count_sig[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\data_count_sig[0]~9_combout ),
	.cout(\data_count_sig[0]~10 ));
defparam \data_count_sig[0]~9 .lut_mask = 16'h55AA;
defparam \data_count_sig[0]~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \data_count_sig[1]~11 (
	.dataa(\data_count_sig[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\data_count_sig[0]~10 ),
	.combout(\data_count_sig[1]~11_combout ),
	.cout(\data_count_sig[1]~12 ));
defparam \data_count_sig[1]~11 .lut_mask = 16'h5A5F;
defparam \data_count_sig[1]~11 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \data_count_sig[2]~13 (
	.dataa(\data_count_sig[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\data_count_sig[1]~12 ),
	.combout(\data_count_sig[2]~13_combout ),
	.cout(\data_count_sig[2]~14 ));
defparam \data_count_sig[2]~13 .lut_mask = 16'h5AAF;
defparam \data_count_sig[2]~13 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \data_count_sig[3]~15 (
	.dataa(\data_count_sig[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\data_count_sig[2]~14 ),
	.combout(\data_count_sig[3]~15_combout ),
	.cout(\data_count_sig[3]~16 ));
defparam \data_count_sig[3]~15 .lut_mask = 16'h5A5F;
defparam \data_count_sig[3]~15 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \data_count_sig[4]~21 (
	.dataa(\data_count_sig[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\data_count_sig[3]~16 ),
	.combout(\data_count_sig[4]~21_combout ),
	.cout(\data_count_sig[4]~22 ));
defparam \data_count_sig[4]~21 .lut_mask = 16'h5AAF;
defparam \data_count_sig[4]~21 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \data_count_sig[5]~23 (
	.dataa(\data_count_sig[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\data_count_sig[4]~22 ),
	.combout(\data_count_sig[5]~23_combout ),
	.cout(\data_count_sig[5]~24 ));
defparam \data_count_sig[5]~23 .lut_mask = 16'h5A5F;
defparam \data_count_sig[5]~23 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \data_count_sig[6]~25 (
	.dataa(\data_count_sig[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\data_count_sig[5]~24 ),
	.combout(\data_count_sig[6]~25_combout ),
	.cout(\data_count_sig[6]~26 ));
defparam \data_count_sig[6]~25 .lut_mask = 16'h5AAF;
defparam \data_count_sig[6]~25 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \data_count_sig[7]~27 (
	.dataa(\data_count_sig[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\data_count_sig[6]~26 ),
	.combout(\data_count_sig[7]~27_combout ),
	.cout(\data_count_sig[7]~28 ));
defparam \data_count_sig[7]~27 .lut_mask = 16'h5A5F;
defparam \data_count_sig[7]~27 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \data_count_sig[8]~29 (
	.dataa(\data_count_sig[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\data_count_sig[7]~28 ),
	.combout(\data_count_sig[8]~29_combout ),
	.cout());
defparam \data_count_sig[8]~29 .lut_mask = 16'h5A5A;
defparam \data_count_sig[8]~29 .sum_lutc_input = "cin";

dffeas fft_dirn_stream(
	.clk(clk),
	.d(\fft_dirn_stream~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_dirn_stream~q ),
	.prn(vcc));
defparam fft_dirn_stream.is_wysiwyg = "true";
defparam fft_dirn_stream.power_up = "low";

dffeas \fft_s2_cur.WAIT_FOR_LPP_INPUT (
	.clk(clk),
	.d(\Selector20~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_s2_cur.WAIT_FOR_LPP_INPUT~q ),
	.prn(vcc));
defparam \fft_s2_cur.WAIT_FOR_LPP_INPUT .is_wysiwyg = "true";
defparam \fft_s2_cur.WAIT_FOR_LPP_INPUT .power_up = "low";

dffeas fft_dirn_held_o2(
	.clk(clk),
	.d(\fft_dirn_held_o2~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_dirn_held_o2~q ),
	.prn(vcc));
defparam fft_dirn_held_o2.is_wysiwyg = "true";
defparam fft_dirn_held_o2.power_up = "low";

dffeas \fft_s2_cur.LPP_C_OUTPUT (
	.clk(clk),
	.d(\Selector22~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_s2_cur.LPP_C_OUTPUT~q ),
	.prn(vcc));
defparam \fft_s2_cur.LPP_C_OUTPUT .is_wysiwyg = "true";
defparam \fft_s2_cur.LPP_C_OUTPUT .power_up = "low";

dffeas \lpp_count_offset[0] (
	.clk(clk),
	.d(\lpp_count_offset[0]~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\lpp_count_offset[0]~12_combout ),
	.q(\lpp_count_offset[0]~q ),
	.prn(vcc));
defparam \lpp_count_offset[0] .is_wysiwyg = "true";
defparam \lpp_count_offset[0] .power_up = "low";

dffeas \lpp_count_offset[1] (
	.clk(clk),
	.d(\lpp_count_offset[1]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\lpp_count_offset[0]~12_combout ),
	.q(\lpp_count_offset[1]~q ),
	.prn(vcc));
defparam \lpp_count_offset[1] .is_wysiwyg = "true";
defparam \lpp_count_offset[1] .power_up = "low";

dffeas \lpp_count_offset[2] (
	.clk(clk),
	.d(\lpp_count_offset[2]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\lpp_count_offset[0]~12_combout ),
	.q(\lpp_count_offset[2]~q ),
	.prn(vcc));
defparam \lpp_count_offset[2] .is_wysiwyg = "true";
defparam \lpp_count_offset[2] .power_up = "low";

dffeas \lpp_count_offset[3] (
	.clk(clk),
	.d(\lpp_count_offset[3]~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\lpp_count_offset[0]~12_combout ),
	.q(\lpp_count_offset[3]~q ),
	.prn(vcc));
defparam \lpp_count_offset[3] .is_wysiwyg = "true";
defparam \lpp_count_offset[3] .power_up = "low";

dffeas \lpp_count_offset[4] (
	.clk(clk),
	.d(\lpp_count_offset[4]~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\lpp_count_offset[0]~12_combout ),
	.q(\lpp_count_offset[4]~q ),
	.prn(vcc));
defparam \lpp_count_offset[4] .is_wysiwyg = "true";
defparam \lpp_count_offset[4] .power_up = "low";

dffeas \lpp_count_offset[5] (
	.clk(clk),
	.d(\lpp_count_offset[5]~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\lpp_count_offset[0]~12_combout ),
	.q(\lpp_count_offset[5]~q ),
	.prn(vcc));
defparam \lpp_count_offset[5] .is_wysiwyg = "true";
defparam \lpp_count_offset[5] .power_up = "low";

dffeas \lpp_count_offset[6] (
	.clk(clk),
	.d(\lpp_count_offset[6]~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\lpp_count_offset[0]~12_combout ),
	.q(\lpp_count_offset[6]~q ),
	.prn(vcc));
defparam \lpp_count_offset[6] .is_wysiwyg = "true";
defparam \lpp_count_offset[6] .power_up = "low";

dffeas \lpp_count_offset[7] (
	.clk(clk),
	.d(\lpp_count_offset[7]~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\lpp_count_offset[0]~12_combout ),
	.q(\lpp_count_offset[7]~q ),
	.prn(vcc));
defparam \lpp_count_offset[7] .is_wysiwyg = "true";
defparam \lpp_count_offset[7] .power_up = "low";

dffeas \lpp_count_offset[8] (
	.clk(clk),
	.d(\lpp_count_offset[8]~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\lpp_count_offset[0]~12_combout ),
	.q(\lpp_count_offset[8]~q ),
	.prn(vcc));
defparam \lpp_count_offset[8] .is_wysiwyg = "true";
defparam \lpp_count_offset[8] .power_up = "low";

dffeas fft_dirn_held_o(
	.clk(clk),
	.d(\fft_dirn_held_o~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_dirn_held_o~q ),
	.prn(vcc));
defparam fft_dirn_held_o.is_wysiwyg = "true";
defparam fft_dirn_held_o.power_up = "low";

dffeas \lpp_count[0] (
	.clk(clk),
	.d(\Selector14~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_count[0]~q ),
	.prn(vcc));
defparam \lpp_count[0] .is_wysiwyg = "true";
defparam \lpp_count[0] .power_up = "low";

cycloneiii_lcell_comb \lpp_count_offset[0]~9 (
	.dataa(\lpp_count[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\lpp_count_offset[0]~9_combout ),
	.cout(\lpp_count_offset[0]~10 ));
defparam \lpp_count_offset[0]~9 .lut_mask = 16'h55AA;
defparam \lpp_count_offset[0]~9 .sum_lutc_input = "datac";

dffeas \lpp_count[1] (
	.clk(clk),
	.d(\lpp_count~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_count[1]~q ),
	.prn(vcc));
defparam \lpp_count[1] .is_wysiwyg = "true";
defparam \lpp_count[1] .power_up = "low";

cycloneiii_lcell_comb \lpp_count_offset[1]~13 (
	.dataa(\lpp_count[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\lpp_count_offset[0]~10 ),
	.combout(\lpp_count_offset[1]~13_combout ),
	.cout(\lpp_count_offset[1]~14 ));
defparam \lpp_count_offset[1]~13 .lut_mask = 16'h5A5F;
defparam \lpp_count_offset[1]~13 .sum_lutc_input = "cin";

dffeas \lpp_count[2] (
	.clk(clk),
	.d(\Selector13~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_count[2]~q ),
	.prn(vcc));
defparam \lpp_count[2] .is_wysiwyg = "true";
defparam \lpp_count[2] .power_up = "low";

cycloneiii_lcell_comb \lpp_count_offset[2]~15 (
	.dataa(\lpp_count[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\lpp_count_offset[1]~14 ),
	.combout(\lpp_count_offset[2]~15_combout ),
	.cout(\lpp_count_offset[2]~16 ));
defparam \lpp_count_offset[2]~15 .lut_mask = 16'h5AAF;
defparam \lpp_count_offset[2]~15 .sum_lutc_input = "cin";

dffeas \lpp_count[3] (
	.clk(clk),
	.d(\Selector12~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_count[3]~q ),
	.prn(vcc));
defparam \lpp_count[3] .is_wysiwyg = "true";
defparam \lpp_count[3] .power_up = "low";

cycloneiii_lcell_comb \lpp_count_offset[3]~17 (
	.dataa(\lpp_count[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\lpp_count_offset[2]~16 ),
	.combout(\lpp_count_offset[3]~17_combout ),
	.cout(\lpp_count_offset[3]~18 ));
defparam \lpp_count_offset[3]~17 .lut_mask = 16'h5A5F;
defparam \lpp_count_offset[3]~17 .sum_lutc_input = "cin";

dffeas \lpp_count[4] (
	.clk(clk),
	.d(\Selector11~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_count[4]~q ),
	.prn(vcc));
defparam \lpp_count[4] .is_wysiwyg = "true";
defparam \lpp_count[4] .power_up = "low";

cycloneiii_lcell_comb \lpp_count_offset[4]~19 (
	.dataa(\lpp_count[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\lpp_count_offset[3]~18 ),
	.combout(\lpp_count_offset[4]~19_combout ),
	.cout(\lpp_count_offset[4]~20 ));
defparam \lpp_count_offset[4]~19 .lut_mask = 16'h5AAF;
defparam \lpp_count_offset[4]~19 .sum_lutc_input = "cin";

dffeas \lpp_count[5] (
	.clk(clk),
	.d(\Selector10~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_count[5]~q ),
	.prn(vcc));
defparam \lpp_count[5] .is_wysiwyg = "true";
defparam \lpp_count[5] .power_up = "low";

cycloneiii_lcell_comb \lpp_count_offset[5]~21 (
	.dataa(\lpp_count[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\lpp_count_offset[4]~20 ),
	.combout(\lpp_count_offset[5]~21_combout ),
	.cout(\lpp_count_offset[5]~22 ));
defparam \lpp_count_offset[5]~21 .lut_mask = 16'h5A5F;
defparam \lpp_count_offset[5]~21 .sum_lutc_input = "cin";

dffeas \lpp_count[6] (
	.clk(clk),
	.d(\Selector9~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_count[6]~q ),
	.prn(vcc));
defparam \lpp_count[6] .is_wysiwyg = "true";
defparam \lpp_count[6] .power_up = "low";

cycloneiii_lcell_comb \lpp_count_offset[6]~23 (
	.dataa(\lpp_count[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\lpp_count_offset[5]~22 ),
	.combout(\lpp_count_offset[6]~23_combout ),
	.cout(\lpp_count_offset[6]~24 ));
defparam \lpp_count_offset[6]~23 .lut_mask = 16'h5AAF;
defparam \lpp_count_offset[6]~23 .sum_lutc_input = "cin";

dffeas \lpp_count[7] (
	.clk(clk),
	.d(\Selector8~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_count[7]~q ),
	.prn(vcc));
defparam \lpp_count[7] .is_wysiwyg = "true";
defparam \lpp_count[7] .power_up = "low";

cycloneiii_lcell_comb \lpp_count_offset[7]~25 (
	.dataa(\lpp_count[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\lpp_count_offset[6]~24 ),
	.combout(\lpp_count_offset[7]~25_combout ),
	.cout(\lpp_count_offset[7]~26 ));
defparam \lpp_count_offset[7]~25 .lut_mask = 16'h5A5F;
defparam \lpp_count_offset[7]~25 .sum_lutc_input = "cin";

dffeas \lpp_count[8] (
	.clk(clk),
	.d(\Selector7~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_count[8]~q ),
	.prn(vcc));
defparam \lpp_count[8] .is_wysiwyg = "true";
defparam \lpp_count[8] .power_up = "low";

cycloneiii_lcell_comb \lpp_count_offset[8]~27 (
	.dataa(\lpp_count[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\lpp_count_offset[7]~26 ),
	.combout(\lpp_count_offset[8]~27_combout ),
	.cout());
defparam \lpp_count_offset[8]~27 .lut_mask = 16'h5A5A;
defparam \lpp_count_offset[8]~27 .sum_lutc_input = "cin";

dffeas \lpp_ram_data_out_sw[1][1] (
	.clk(clk),
	.d(\lpp_ram_data_out_sw[1][1]~2_combout ),
	.asdata(\Mux30~3_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\gen_radix_2_last_pass:delay_mid|tdl_arr[4]~q ),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out_sw[1][1]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out_sw[1][1] .is_wysiwyg = "true";
defparam \lpp_ram_data_out_sw[1][1] .power_up = "low";

dffeas \lpp_ram_data_out_sw[0][1] (
	.clk(clk),
	.d(\lpp_ram_data_out_sw[0][1]~3_combout ),
	.asdata(\Mux30~3_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\gen_radix_2_last_pass:delay_mid|tdl_arr[4]~q ),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out_sw[0][1]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out_sw[0][1] .is_wysiwyg = "true";
defparam \lpp_ram_data_out_sw[0][1] .power_up = "low";

dffeas \lpp_ram_data_out_sw[1][0] (
	.clk(clk),
	.d(\lpp_ram_data_out_sw[1][0]~30_combout ),
	.asdata(\Mux31~3_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\gen_radix_2_last_pass:delay_mid|tdl_arr[4]~q ),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out_sw[1][0]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out_sw[1][0] .is_wysiwyg = "true";
defparam \lpp_ram_data_out_sw[1][0] .power_up = "low";

dffeas \lpp_ram_data_out_sw[0][0] (
	.clk(clk),
	.d(\lpp_ram_data_out_sw[0][0]~31_combout ),
	.asdata(\Mux31~3_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\gen_radix_2_last_pass:delay_mid|tdl_arr[4]~q ),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out_sw[0][0]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out_sw[0][0] .is_wysiwyg = "true";
defparam \lpp_ram_data_out_sw[0][0] .power_up = "low";

dffeas \lpp_ram_data_out_sw[1][7] (
	.clk(clk),
	.d(\lpp_ram_data_out_sw[1][7]~26_combout ),
	.asdata(\Mux24~3_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\gen_radix_2_last_pass:delay_mid|tdl_arr[4]~q ),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out_sw[1][7]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out_sw[1][7] .is_wysiwyg = "true";
defparam \lpp_ram_data_out_sw[1][7] .power_up = "low";

dffeas \lpp_ram_data_out_sw[0][7] (
	.clk(clk),
	.d(\lpp_ram_data_out_sw[0][7]~27_combout ),
	.asdata(\Mux24~3_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\gen_radix_2_last_pass:delay_mid|tdl_arr[4]~q ),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out_sw[0][7]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out_sw[0][7] .is_wysiwyg = "true";
defparam \lpp_ram_data_out_sw[0][7] .power_up = "low";

dffeas \lpp_ram_data_out_sw[1][6] (
	.clk(clk),
	.d(\lpp_ram_data_out_sw[1][6]~22_combout ),
	.asdata(\Mux25~3_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\gen_radix_2_last_pass:delay_mid|tdl_arr[4]~q ),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out_sw[1][6]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out_sw[1][6] .is_wysiwyg = "true";
defparam \lpp_ram_data_out_sw[1][6] .power_up = "low";

dffeas \lpp_ram_data_out_sw[0][6] (
	.clk(clk),
	.d(\lpp_ram_data_out_sw[0][6]~23_combout ),
	.asdata(\Mux25~3_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\gen_radix_2_last_pass:delay_mid|tdl_arr[4]~q ),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out_sw[0][6]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out_sw[0][6] .is_wysiwyg = "true";
defparam \lpp_ram_data_out_sw[0][6] .power_up = "low";

dffeas \lpp_ram_data_out_sw[1][5] (
	.clk(clk),
	.d(\lpp_ram_data_out_sw[1][5]~18_combout ),
	.asdata(\Mux26~3_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\gen_radix_2_last_pass:delay_mid|tdl_arr[4]~q ),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out_sw[1][5]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out_sw[1][5] .is_wysiwyg = "true";
defparam \lpp_ram_data_out_sw[1][5] .power_up = "low";

dffeas \lpp_ram_data_out_sw[0][5] (
	.clk(clk),
	.d(\lpp_ram_data_out_sw[0][5]~19_combout ),
	.asdata(\Mux26~3_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\gen_radix_2_last_pass:delay_mid|tdl_arr[4]~q ),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out_sw[0][5]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out_sw[0][5] .is_wysiwyg = "true";
defparam \lpp_ram_data_out_sw[0][5] .power_up = "low";

dffeas \lpp_ram_data_out_sw[1][4] (
	.clk(clk),
	.d(\lpp_ram_data_out_sw[1][4]~14_combout ),
	.asdata(\Mux27~3_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\gen_radix_2_last_pass:delay_mid|tdl_arr[4]~q ),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out_sw[1][4]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out_sw[1][4] .is_wysiwyg = "true";
defparam \lpp_ram_data_out_sw[1][4] .power_up = "low";

dffeas \lpp_ram_data_out_sw[0][4] (
	.clk(clk),
	.d(\lpp_ram_data_out_sw[0][4]~15_combout ),
	.asdata(\Mux27~3_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\gen_radix_2_last_pass:delay_mid|tdl_arr[4]~q ),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out_sw[0][4]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out_sw[0][4] .is_wysiwyg = "true";
defparam \lpp_ram_data_out_sw[0][4] .power_up = "low";

dffeas \lpp_ram_data_out_sw[1][3] (
	.clk(clk),
	.d(\lpp_ram_data_out_sw[1][3]~10_combout ),
	.asdata(\Mux28~3_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\gen_radix_2_last_pass:delay_mid|tdl_arr[4]~q ),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out_sw[1][3]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out_sw[1][3] .is_wysiwyg = "true";
defparam \lpp_ram_data_out_sw[1][3] .power_up = "low";

dffeas \lpp_ram_data_out_sw[0][3] (
	.clk(clk),
	.d(\lpp_ram_data_out_sw[0][3]~11_combout ),
	.asdata(\Mux28~3_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\gen_radix_2_last_pass:delay_mid|tdl_arr[4]~q ),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out_sw[0][3]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out_sw[0][3] .is_wysiwyg = "true";
defparam \lpp_ram_data_out_sw[0][3] .power_up = "low";

dffeas \lpp_ram_data_out_sw[1][2] (
	.clk(clk),
	.d(\lpp_ram_data_out_sw[1][2]~6_combout ),
	.asdata(\Mux29~3_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\gen_radix_2_last_pass:delay_mid|tdl_arr[4]~q ),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out_sw[1][2]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out_sw[1][2] .is_wysiwyg = "true";
defparam \lpp_ram_data_out_sw[1][2] .power_up = "low";

dffeas \lpp_ram_data_out_sw[0][2] (
	.clk(clk),
	.d(\lpp_ram_data_out_sw[0][2]~7_combout ),
	.asdata(\Mux29~3_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\gen_radix_2_last_pass:delay_mid|tdl_arr[4]~q ),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out_sw[0][2]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out_sw[0][2] .is_wysiwyg = "true";
defparam \lpp_ram_data_out_sw[0][2] .power_up = "low";

dffeas \lpp_ram_data_out_sw[1][9] (
	.clk(clk),
	.d(\lpp_ram_data_out_sw[1][9]~0_combout ),
	.asdata(\Mux22~3_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\gen_radix_2_last_pass:delay_mid|tdl_arr[4]~q ),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out_sw[1][9]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out_sw[1][9] .is_wysiwyg = "true";
defparam \lpp_ram_data_out_sw[1][9] .power_up = "low";

dffeas \lpp_ram_data_out_sw[0][9] (
	.clk(clk),
	.d(\lpp_ram_data_out_sw[0][9]~1_combout ),
	.asdata(\Mux22~3_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\gen_radix_2_last_pass:delay_mid|tdl_arr[4]~q ),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out_sw[0][9]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out_sw[0][9] .is_wysiwyg = "true";
defparam \lpp_ram_data_out_sw[0][9] .power_up = "low";

dffeas \lpp_ram_data_out_sw[1][8] (
	.clk(clk),
	.d(\lpp_ram_data_out_sw[1][8]~28_combout ),
	.asdata(\Mux23~3_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\gen_radix_2_last_pass:delay_mid|tdl_arr[4]~q ),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out_sw[1][8]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out_sw[1][8] .is_wysiwyg = "true";
defparam \lpp_ram_data_out_sw[1][8] .power_up = "low";

dffeas \lpp_ram_data_out_sw[0][8] (
	.clk(clk),
	.d(\lpp_ram_data_out_sw[0][8]~29_combout ),
	.asdata(\Mux23~3_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\gen_radix_2_last_pass:delay_mid|tdl_arr[4]~q ),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out_sw[0][8]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out_sw[0][8] .is_wysiwyg = "true";
defparam \lpp_ram_data_out_sw[0][8] .power_up = "low";

dffeas \lpp_ram_data_out_sw[1][15] (
	.clk(clk),
	.d(\lpp_ram_data_out_sw[1][15]~24_combout ),
	.asdata(\Mux16~3_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\gen_radix_2_last_pass:delay_mid|tdl_arr[4]~q ),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out_sw[1][15]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out_sw[1][15] .is_wysiwyg = "true";
defparam \lpp_ram_data_out_sw[1][15] .power_up = "low";

dffeas \lpp_ram_data_out_sw[0][15] (
	.clk(clk),
	.d(\lpp_ram_data_out_sw[0][15]~25_combout ),
	.asdata(\Mux16~3_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\gen_radix_2_last_pass:delay_mid|tdl_arr[4]~q ),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out_sw[0][15]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out_sw[0][15] .is_wysiwyg = "true";
defparam \lpp_ram_data_out_sw[0][15] .power_up = "low";

dffeas \lpp_ram_data_out_sw[1][14] (
	.clk(clk),
	.d(\lpp_ram_data_out_sw[1][14]~20_combout ),
	.asdata(\Mux17~3_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\gen_radix_2_last_pass:delay_mid|tdl_arr[4]~q ),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out_sw[1][14]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out_sw[1][14] .is_wysiwyg = "true";
defparam \lpp_ram_data_out_sw[1][14] .power_up = "low";

dffeas \lpp_ram_data_out_sw[0][14] (
	.clk(clk),
	.d(\lpp_ram_data_out_sw[0][14]~21_combout ),
	.asdata(\Mux17~3_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\gen_radix_2_last_pass:delay_mid|tdl_arr[4]~q ),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out_sw[0][14]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out_sw[0][14] .is_wysiwyg = "true";
defparam \lpp_ram_data_out_sw[0][14] .power_up = "low";

dffeas \lpp_ram_data_out_sw[1][13] (
	.clk(clk),
	.d(\lpp_ram_data_out_sw[1][13]~16_combout ),
	.asdata(\Mux18~3_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\gen_radix_2_last_pass:delay_mid|tdl_arr[4]~q ),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out_sw[1][13]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out_sw[1][13] .is_wysiwyg = "true";
defparam \lpp_ram_data_out_sw[1][13] .power_up = "low";

dffeas \lpp_ram_data_out_sw[0][13] (
	.clk(clk),
	.d(\lpp_ram_data_out_sw[0][13]~17_combout ),
	.asdata(\Mux18~3_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\gen_radix_2_last_pass:delay_mid|tdl_arr[4]~q ),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out_sw[0][13]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out_sw[0][13] .is_wysiwyg = "true";
defparam \lpp_ram_data_out_sw[0][13] .power_up = "low";

dffeas \lpp_ram_data_out_sw[1][12] (
	.clk(clk),
	.d(\lpp_ram_data_out_sw[1][12]~12_combout ),
	.asdata(\Mux19~3_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\gen_radix_2_last_pass:delay_mid|tdl_arr[4]~q ),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out_sw[1][12]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out_sw[1][12] .is_wysiwyg = "true";
defparam \lpp_ram_data_out_sw[1][12] .power_up = "low";

dffeas \lpp_ram_data_out_sw[0][12] (
	.clk(clk),
	.d(\lpp_ram_data_out_sw[0][12]~13_combout ),
	.asdata(\Mux19~3_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\gen_radix_2_last_pass:delay_mid|tdl_arr[4]~q ),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out_sw[0][12]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out_sw[0][12] .is_wysiwyg = "true";
defparam \lpp_ram_data_out_sw[0][12] .power_up = "low";

dffeas \lpp_ram_data_out_sw[1][11] (
	.clk(clk),
	.d(\lpp_ram_data_out_sw[1][11]~8_combout ),
	.asdata(\Mux20~3_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\gen_radix_2_last_pass:delay_mid|tdl_arr[4]~q ),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out_sw[1][11]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out_sw[1][11] .is_wysiwyg = "true";
defparam \lpp_ram_data_out_sw[1][11] .power_up = "low";

dffeas \lpp_ram_data_out_sw[0][11] (
	.clk(clk),
	.d(\lpp_ram_data_out_sw[0][11]~9_combout ),
	.asdata(\Mux20~3_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\gen_radix_2_last_pass:delay_mid|tdl_arr[4]~q ),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out_sw[0][11]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out_sw[0][11] .is_wysiwyg = "true";
defparam \lpp_ram_data_out_sw[0][11] .power_up = "low";

dffeas \lpp_ram_data_out_sw[1][10] (
	.clk(clk),
	.d(\lpp_ram_data_out_sw[1][10]~4_combout ),
	.asdata(\Mux21~3_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\gen_radix_2_last_pass:delay_mid|tdl_arr[4]~q ),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out_sw[1][10]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out_sw[1][10] .is_wysiwyg = "true";
defparam \lpp_ram_data_out_sw[1][10] .power_up = "low";

dffeas \lpp_ram_data_out_sw[0][10] (
	.clk(clk),
	.d(\lpp_ram_data_out_sw[0][10]~5_combout ),
	.asdata(\Mux21~3_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\gen_radix_2_last_pass:delay_mid|tdl_arr[4]~q ),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out_sw[0][10]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out_sw[0][10] .is_wysiwyg = "true";
defparam \lpp_ram_data_out_sw[0][10] .power_up = "low";

cycloneiii_lcell_comb \Add2~0 (
	.dataa(\lpp_count[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add2~0_combout ),
	.cout(\Add2~1 ));
defparam \Add2~0 .lut_mask = 16'h55AA;
defparam \Add2~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add2~2 (
	.dataa(\lpp_count[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~1 ),
	.combout(\Add2~2_combout ),
	.cout(\Add2~3 ));
defparam \Add2~2 .lut_mask = 16'h5A5F;
defparam \Add2~2 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add2~4 (
	.dataa(\lpp_count[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~3 ),
	.combout(\Add2~4_combout ),
	.cout(\Add2~5 ));
defparam \Add2~4 .lut_mask = 16'h5AAF;
defparam \Add2~4 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add2~6 (
	.dataa(\lpp_count[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~5 ),
	.combout(\Add2~6_combout ),
	.cout(\Add2~7 ));
defparam \Add2~6 .lut_mask = 16'h5A5F;
defparam \Add2~6 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add2~8 (
	.dataa(\lpp_count[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~7 ),
	.combout(\Add2~8_combout ),
	.cout(\Add2~9 ));
defparam \Add2~8 .lut_mask = 16'h5AAF;
defparam \Add2~8 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add2~10 (
	.dataa(\lpp_count[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~9 ),
	.combout(\Add2~10_combout ),
	.cout(\Add2~11 ));
defparam \Add2~10 .lut_mask = 16'h5A5F;
defparam \Add2~10 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add2~12 (
	.dataa(\lpp_count[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~11 ),
	.combout(\Add2~12_combout ),
	.cout(\Add2~13 ));
defparam \Add2~12 .lut_mask = 16'h5AAF;
defparam \Add2~12 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add2~14 (
	.dataa(\lpp_count[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~13 ),
	.combout(\Add2~14_combout ),
	.cout(\Add2~15 ));
defparam \Add2~14 .lut_mask = 16'h5A5F;
defparam \Add2~14 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add2~16 (
	.dataa(\lpp_count[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add2~15 ),
	.combout(\Add2~16_combout ),
	.cout());
defparam \Add2~16 .lut_mask = 16'h5A5A;
defparam \Add2~16 .sum_lutc_input = "cin";

dffeas \lpp_ram_data_out[2][1] (
	.clk(clk),
	.d(\lpp_ram_data_out~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[2][1]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[2][1] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[2][1] .power_up = "low";

dffeas \lpp_ram_data_out[1][1] (
	.clk(clk),
	.d(\lpp_ram_data_out~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[1][1]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[1][1] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[1][1] .power_up = "low";

dffeas \lpp_ram_data_out[0][1] (
	.clk(clk),
	.d(\lpp_ram_data_out~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[0][1]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[0][1] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[0][1] .power_up = "low";

dffeas \lpp_ram_data_out[3][1] (
	.clk(clk),
	.d(\lpp_ram_data_out~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[3][1]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[3][1] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[3][1] .power_up = "low";

cycloneiii_lcell_comb \lpp_ram_data_out_sw[1][1]~2 (
	.dataa(\Mux30~0_combout ),
	.datab(\Mux30~1_combout ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out_sw[1][1]~2_combout ),
	.cout());
defparam \lpp_ram_data_out_sw[1][1]~2 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out_sw[1][1]~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out_sw[0][1]~3 (
	.dataa(\Mux30~1_combout ),
	.datab(\Mux30~0_combout ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out_sw[0][1]~3_combout ),
	.cout());
defparam \lpp_ram_data_out_sw[0][1]~3 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out_sw[0][1]~3 .sum_lutc_input = "datac";

dffeas \lpp_ram_data_out[2][0] (
	.clk(clk),
	.d(\lpp_ram_data_out~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[2][0]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[2][0] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[2][0] .power_up = "low";

dffeas \lpp_ram_data_out[1][0] (
	.clk(clk),
	.d(\lpp_ram_data_out~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[1][0]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[1][0] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[1][0] .power_up = "low";

dffeas \lpp_ram_data_out[0][0] (
	.clk(clk),
	.d(\lpp_ram_data_out~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[0][0]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[0][0] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[0][0] .power_up = "low";

dffeas \lpp_ram_data_out[3][0] (
	.clk(clk),
	.d(\lpp_ram_data_out~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[3][0]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[3][0] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[3][0] .power_up = "low";

cycloneiii_lcell_comb \lpp_ram_data_out_sw[1][0]~30 (
	.dataa(\Mux31~0_combout ),
	.datab(\Mux31~1_combout ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out_sw[1][0]~30_combout ),
	.cout());
defparam \lpp_ram_data_out_sw[1][0]~30 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out_sw[1][0]~30 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out_sw[0][0]~31 (
	.dataa(\Mux31~1_combout ),
	.datab(\Mux31~0_combout ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out_sw[0][0]~31_combout ),
	.cout());
defparam \lpp_ram_data_out_sw[0][0]~31 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out_sw[0][0]~31 .sum_lutc_input = "datac";

dffeas \lpp_ram_data_out[2][7] (
	.clk(clk),
	.d(\lpp_ram_data_out~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[2][7]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[2][7] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[2][7] .power_up = "low";

dffeas \lpp_ram_data_out[1][7] (
	.clk(clk),
	.d(\lpp_ram_data_out~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[1][7]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[1][7] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[1][7] .power_up = "low";

dffeas \lpp_ram_data_out[0][7] (
	.clk(clk),
	.d(\lpp_ram_data_out~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[0][7]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[0][7] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[0][7] .power_up = "low";

dffeas \lpp_ram_data_out[3][7] (
	.clk(clk),
	.d(\lpp_ram_data_out~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[3][7]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[3][7] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[3][7] .power_up = "low";

cycloneiii_lcell_comb \lpp_ram_data_out_sw[1][7]~26 (
	.dataa(\Mux24~0_combout ),
	.datab(\Mux24~1_combout ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out_sw[1][7]~26_combout ),
	.cout());
defparam \lpp_ram_data_out_sw[1][7]~26 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out_sw[1][7]~26 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out_sw[0][7]~27 (
	.dataa(\Mux24~1_combout ),
	.datab(\Mux24~0_combout ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out_sw[0][7]~27_combout ),
	.cout());
defparam \lpp_ram_data_out_sw[0][7]~27 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out_sw[0][7]~27 .sum_lutc_input = "datac";

dffeas \lpp_ram_data_out[2][6] (
	.clk(clk),
	.d(\lpp_ram_data_out~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[2][6]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[2][6] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[2][6] .power_up = "low";

dffeas \lpp_ram_data_out[1][6] (
	.clk(clk),
	.d(\lpp_ram_data_out~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[1][6]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[1][6] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[1][6] .power_up = "low";

dffeas \lpp_ram_data_out[0][6] (
	.clk(clk),
	.d(\lpp_ram_data_out~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[0][6]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[0][6] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[0][6] .power_up = "low";

dffeas \lpp_ram_data_out[3][6] (
	.clk(clk),
	.d(\lpp_ram_data_out~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[3][6]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[3][6] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[3][6] .power_up = "low";

cycloneiii_lcell_comb \lpp_ram_data_out_sw[1][6]~22 (
	.dataa(\Mux25~0_combout ),
	.datab(\Mux25~1_combout ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out_sw[1][6]~22_combout ),
	.cout());
defparam \lpp_ram_data_out_sw[1][6]~22 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out_sw[1][6]~22 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out_sw[0][6]~23 (
	.dataa(\Mux25~1_combout ),
	.datab(\Mux25~0_combout ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out_sw[0][6]~23_combout ),
	.cout());
defparam \lpp_ram_data_out_sw[0][6]~23 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out_sw[0][6]~23 .sum_lutc_input = "datac";

dffeas \lpp_ram_data_out[2][5] (
	.clk(clk),
	.d(\lpp_ram_data_out~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[2][5]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[2][5] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[2][5] .power_up = "low";

dffeas \lpp_ram_data_out[1][5] (
	.clk(clk),
	.d(\lpp_ram_data_out~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[1][5]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[1][5] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[1][5] .power_up = "low";

dffeas \lpp_ram_data_out[0][5] (
	.clk(clk),
	.d(\lpp_ram_data_out~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[0][5]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[0][5] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[0][5] .power_up = "low";

dffeas \lpp_ram_data_out[3][5] (
	.clk(clk),
	.d(\lpp_ram_data_out~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[3][5]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[3][5] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[3][5] .power_up = "low";

cycloneiii_lcell_comb \lpp_ram_data_out_sw[1][5]~18 (
	.dataa(\Mux26~0_combout ),
	.datab(\Mux26~1_combout ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out_sw[1][5]~18_combout ),
	.cout());
defparam \lpp_ram_data_out_sw[1][5]~18 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out_sw[1][5]~18 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out_sw[0][5]~19 (
	.dataa(\Mux26~1_combout ),
	.datab(\Mux26~0_combout ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out_sw[0][5]~19_combout ),
	.cout());
defparam \lpp_ram_data_out_sw[0][5]~19 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out_sw[0][5]~19 .sum_lutc_input = "datac";

dffeas \lpp_ram_data_out[2][4] (
	.clk(clk),
	.d(\lpp_ram_data_out~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[2][4]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[2][4] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[2][4] .power_up = "low";

dffeas \lpp_ram_data_out[1][4] (
	.clk(clk),
	.d(\lpp_ram_data_out~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[1][4]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[1][4] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[1][4] .power_up = "low";

dffeas \lpp_ram_data_out[0][4] (
	.clk(clk),
	.d(\lpp_ram_data_out~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[0][4]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[0][4] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[0][4] .power_up = "low";

dffeas \lpp_ram_data_out[3][4] (
	.clk(clk),
	.d(\lpp_ram_data_out~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[3][4]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[3][4] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[3][4] .power_up = "low";

cycloneiii_lcell_comb \lpp_ram_data_out_sw[1][4]~14 (
	.dataa(\Mux27~0_combout ),
	.datab(\Mux27~1_combout ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out_sw[1][4]~14_combout ),
	.cout());
defparam \lpp_ram_data_out_sw[1][4]~14 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out_sw[1][4]~14 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out_sw[0][4]~15 (
	.dataa(\Mux27~1_combout ),
	.datab(\Mux27~0_combout ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out_sw[0][4]~15_combout ),
	.cout());
defparam \lpp_ram_data_out_sw[0][4]~15 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out_sw[0][4]~15 .sum_lutc_input = "datac";

dffeas \lpp_ram_data_out[2][3] (
	.clk(clk),
	.d(\lpp_ram_data_out~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[2][3]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[2][3] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[2][3] .power_up = "low";

dffeas \lpp_ram_data_out[1][3] (
	.clk(clk),
	.d(\lpp_ram_data_out~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[1][3]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[1][3] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[1][3] .power_up = "low";

dffeas \lpp_ram_data_out[0][3] (
	.clk(clk),
	.d(\lpp_ram_data_out~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[0][3]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[0][3] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[0][3] .power_up = "low";

dffeas \lpp_ram_data_out[3][3] (
	.clk(clk),
	.d(\lpp_ram_data_out~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[3][3]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[3][3] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[3][3] .power_up = "low";

cycloneiii_lcell_comb \lpp_ram_data_out_sw[1][3]~10 (
	.dataa(\Mux28~0_combout ),
	.datab(\Mux28~1_combout ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out_sw[1][3]~10_combout ),
	.cout());
defparam \lpp_ram_data_out_sw[1][3]~10 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out_sw[1][3]~10 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out_sw[0][3]~11 (
	.dataa(\Mux28~1_combout ),
	.datab(\Mux28~0_combout ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out_sw[0][3]~11_combout ),
	.cout());
defparam \lpp_ram_data_out_sw[0][3]~11 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out_sw[0][3]~11 .sum_lutc_input = "datac";

dffeas \lpp_ram_data_out[2][2] (
	.clk(clk),
	.d(\lpp_ram_data_out~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[2][2]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[2][2] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[2][2] .power_up = "low";

dffeas \lpp_ram_data_out[1][2] (
	.clk(clk),
	.d(\lpp_ram_data_out~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[1][2]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[1][2] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[1][2] .power_up = "low";

dffeas \lpp_ram_data_out[0][2] (
	.clk(clk),
	.d(\lpp_ram_data_out~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[0][2]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[0][2] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[0][2] .power_up = "low";

dffeas \lpp_ram_data_out[3][2] (
	.clk(clk),
	.d(\lpp_ram_data_out~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[3][2]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[3][2] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[3][2] .power_up = "low";

cycloneiii_lcell_comb \lpp_ram_data_out_sw[1][2]~6 (
	.dataa(\Mux29~0_combout ),
	.datab(\Mux29~1_combout ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out_sw[1][2]~6_combout ),
	.cout());
defparam \lpp_ram_data_out_sw[1][2]~6 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out_sw[1][2]~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out_sw[0][2]~7 (
	.dataa(\Mux29~1_combout ),
	.datab(\Mux29~0_combout ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out_sw[0][2]~7_combout ),
	.cout());
defparam \lpp_ram_data_out_sw[0][2]~7 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out_sw[0][2]~7 .sum_lutc_input = "datac";

dffeas \lpp_ram_data_out[2][9] (
	.clk(clk),
	.d(\lpp_ram_data_out~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[2][9]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[2][9] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[2][9] .power_up = "low";

dffeas \lpp_ram_data_out[1][9] (
	.clk(clk),
	.d(\lpp_ram_data_out~33_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[1][9]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[1][9] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[1][9] .power_up = "low";

dffeas \lpp_ram_data_out[0][9] (
	.clk(clk),
	.d(\lpp_ram_data_out~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[0][9]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[0][9] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[0][9] .power_up = "low";

dffeas \lpp_ram_data_out[3][9] (
	.clk(clk),
	.d(\lpp_ram_data_out~35_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[3][9]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[3][9] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[3][9] .power_up = "low";

cycloneiii_lcell_comb \lpp_ram_data_out_sw[1][9]~0 (
	.dataa(\Mux22~0_combout ),
	.datab(\Mux22~1_combout ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out_sw[1][9]~0_combout ),
	.cout());
defparam \lpp_ram_data_out_sw[1][9]~0 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out_sw[1][9]~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out_sw[0][9]~1 (
	.dataa(\Mux22~1_combout ),
	.datab(\Mux22~0_combout ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out_sw[0][9]~1_combout ),
	.cout());
defparam \lpp_ram_data_out_sw[0][9]~1 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out_sw[0][9]~1 .sum_lutc_input = "datac";

dffeas \lpp_ram_data_out[2][8] (
	.clk(clk),
	.d(\lpp_ram_data_out~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[2][8]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[2][8] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[2][8] .power_up = "low";

dffeas \lpp_ram_data_out[1][8] (
	.clk(clk),
	.d(\lpp_ram_data_out~37_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[1][8]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[1][8] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[1][8] .power_up = "low";

dffeas \lpp_ram_data_out[0][8] (
	.clk(clk),
	.d(\lpp_ram_data_out~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[0][8]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[0][8] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[0][8] .power_up = "low";

dffeas \lpp_ram_data_out[3][8] (
	.clk(clk),
	.d(\lpp_ram_data_out~39_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[3][8]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[3][8] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[3][8] .power_up = "low";

cycloneiii_lcell_comb \lpp_ram_data_out_sw[1][8]~28 (
	.dataa(\Mux23~0_combout ),
	.datab(\Mux23~1_combout ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out_sw[1][8]~28_combout ),
	.cout());
defparam \lpp_ram_data_out_sw[1][8]~28 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out_sw[1][8]~28 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out_sw[0][8]~29 (
	.dataa(\Mux23~1_combout ),
	.datab(\Mux23~0_combout ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out_sw[0][8]~29_combout ),
	.cout());
defparam \lpp_ram_data_out_sw[0][8]~29 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out_sw[0][8]~29 .sum_lutc_input = "datac";

dffeas \lpp_ram_data_out[2][15] (
	.clk(clk),
	.d(\lpp_ram_data_out~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[2][15]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[2][15] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[2][15] .power_up = "low";

dffeas \lpp_ram_data_out[1][15] (
	.clk(clk),
	.d(\lpp_ram_data_out~41_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[1][15]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[1][15] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[1][15] .power_up = "low";

dffeas \lpp_ram_data_out[0][15] (
	.clk(clk),
	.d(\lpp_ram_data_out~42_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[0][15]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[0][15] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[0][15] .power_up = "low";

dffeas \lpp_ram_data_out[3][15] (
	.clk(clk),
	.d(\lpp_ram_data_out~43_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[3][15]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[3][15] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[3][15] .power_up = "low";

cycloneiii_lcell_comb \lpp_ram_data_out_sw[1][15]~24 (
	.dataa(\Mux16~0_combout ),
	.datab(\Mux16~1_combout ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out_sw[1][15]~24_combout ),
	.cout());
defparam \lpp_ram_data_out_sw[1][15]~24 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out_sw[1][15]~24 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out_sw[0][15]~25 (
	.dataa(\Mux16~1_combout ),
	.datab(\Mux16~0_combout ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out_sw[0][15]~25_combout ),
	.cout());
defparam \lpp_ram_data_out_sw[0][15]~25 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out_sw[0][15]~25 .sum_lutc_input = "datac";

dffeas \lpp_ram_data_out[2][14] (
	.clk(clk),
	.d(\lpp_ram_data_out~44_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[2][14]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[2][14] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[2][14] .power_up = "low";

dffeas \lpp_ram_data_out[1][14] (
	.clk(clk),
	.d(\lpp_ram_data_out~45_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[1][14]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[1][14] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[1][14] .power_up = "low";

dffeas \lpp_ram_data_out[0][14] (
	.clk(clk),
	.d(\lpp_ram_data_out~46_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[0][14]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[0][14] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[0][14] .power_up = "low";

dffeas \lpp_ram_data_out[3][14] (
	.clk(clk),
	.d(\lpp_ram_data_out~47_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[3][14]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[3][14] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[3][14] .power_up = "low";

cycloneiii_lcell_comb \lpp_ram_data_out_sw[1][14]~20 (
	.dataa(\Mux17~0_combout ),
	.datab(\Mux17~1_combout ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out_sw[1][14]~20_combout ),
	.cout());
defparam \lpp_ram_data_out_sw[1][14]~20 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out_sw[1][14]~20 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out_sw[0][14]~21 (
	.dataa(\Mux17~1_combout ),
	.datab(\Mux17~0_combout ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out_sw[0][14]~21_combout ),
	.cout());
defparam \lpp_ram_data_out_sw[0][14]~21 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out_sw[0][14]~21 .sum_lutc_input = "datac";

dffeas \lpp_ram_data_out[2][13] (
	.clk(clk),
	.d(\lpp_ram_data_out~48_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[2][13]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[2][13] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[2][13] .power_up = "low";

dffeas \lpp_ram_data_out[1][13] (
	.clk(clk),
	.d(\lpp_ram_data_out~49_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[1][13]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[1][13] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[1][13] .power_up = "low";

dffeas \lpp_ram_data_out[0][13] (
	.clk(clk),
	.d(\lpp_ram_data_out~50_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[0][13]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[0][13] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[0][13] .power_up = "low";

dffeas \lpp_ram_data_out[3][13] (
	.clk(clk),
	.d(\lpp_ram_data_out~51_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[3][13]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[3][13] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[3][13] .power_up = "low";

cycloneiii_lcell_comb \lpp_ram_data_out_sw[1][13]~16 (
	.dataa(\Mux18~0_combout ),
	.datab(\Mux18~1_combout ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out_sw[1][13]~16_combout ),
	.cout());
defparam \lpp_ram_data_out_sw[1][13]~16 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out_sw[1][13]~16 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out_sw[0][13]~17 (
	.dataa(\Mux18~1_combout ),
	.datab(\Mux18~0_combout ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out_sw[0][13]~17_combout ),
	.cout());
defparam \lpp_ram_data_out_sw[0][13]~17 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out_sw[0][13]~17 .sum_lutc_input = "datac";

dffeas \lpp_ram_data_out[2][12] (
	.clk(clk),
	.d(\lpp_ram_data_out~52_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[2][12]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[2][12] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[2][12] .power_up = "low";

dffeas \lpp_ram_data_out[1][12] (
	.clk(clk),
	.d(\lpp_ram_data_out~53_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[1][12]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[1][12] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[1][12] .power_up = "low";

dffeas \lpp_ram_data_out[0][12] (
	.clk(clk),
	.d(\lpp_ram_data_out~54_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[0][12]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[0][12] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[0][12] .power_up = "low";

dffeas \lpp_ram_data_out[3][12] (
	.clk(clk),
	.d(\lpp_ram_data_out~55_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[3][12]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[3][12] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[3][12] .power_up = "low";

cycloneiii_lcell_comb \lpp_ram_data_out_sw[1][12]~12 (
	.dataa(\Mux19~0_combout ),
	.datab(\Mux19~1_combout ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out_sw[1][12]~12_combout ),
	.cout());
defparam \lpp_ram_data_out_sw[1][12]~12 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out_sw[1][12]~12 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out_sw[0][12]~13 (
	.dataa(\Mux19~1_combout ),
	.datab(\Mux19~0_combout ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out_sw[0][12]~13_combout ),
	.cout());
defparam \lpp_ram_data_out_sw[0][12]~13 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out_sw[0][12]~13 .sum_lutc_input = "datac";

dffeas \lpp_ram_data_out[2][11] (
	.clk(clk),
	.d(\lpp_ram_data_out~56_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[2][11]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[2][11] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[2][11] .power_up = "low";

dffeas \lpp_ram_data_out[1][11] (
	.clk(clk),
	.d(\lpp_ram_data_out~57_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[1][11]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[1][11] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[1][11] .power_up = "low";

dffeas \lpp_ram_data_out[0][11] (
	.clk(clk),
	.d(\lpp_ram_data_out~58_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[0][11]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[0][11] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[0][11] .power_up = "low";

dffeas \lpp_ram_data_out[3][11] (
	.clk(clk),
	.d(\lpp_ram_data_out~59_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[3][11]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[3][11] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[3][11] .power_up = "low";

cycloneiii_lcell_comb \lpp_ram_data_out_sw[1][11]~8 (
	.dataa(\Mux20~0_combout ),
	.datab(\Mux20~1_combout ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out_sw[1][11]~8_combout ),
	.cout());
defparam \lpp_ram_data_out_sw[1][11]~8 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out_sw[1][11]~8 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out_sw[0][11]~9 (
	.dataa(\Mux20~1_combout ),
	.datab(\Mux20~0_combout ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out_sw[0][11]~9_combout ),
	.cout());
defparam \lpp_ram_data_out_sw[0][11]~9 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out_sw[0][11]~9 .sum_lutc_input = "datac";

dffeas \lpp_ram_data_out[2][10] (
	.clk(clk),
	.d(\lpp_ram_data_out~60_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[2][10]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[2][10] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[2][10] .power_up = "low";

dffeas \lpp_ram_data_out[1][10] (
	.clk(clk),
	.d(\lpp_ram_data_out~61_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[1][10]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[1][10] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[1][10] .power_up = "low";

dffeas \lpp_ram_data_out[0][10] (
	.clk(clk),
	.d(\lpp_ram_data_out~62_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[0][10]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[0][10] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[0][10] .power_up = "low";

dffeas \lpp_ram_data_out[3][10] (
	.clk(clk),
	.d(\lpp_ram_data_out~63_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[3][10]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[3][10] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[3][10] .power_up = "low";

cycloneiii_lcell_comb \lpp_ram_data_out_sw[1][10]~4 (
	.dataa(\Mux21~0_combout ),
	.datab(\Mux21~1_combout ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out_sw[1][10]~4_combout ),
	.cout());
defparam \lpp_ram_data_out_sw[1][10]~4 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out_sw[1][10]~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out_sw[0][10]~5 (
	.dataa(\Mux21~1_combout ),
	.datab(\Mux21~0_combout ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out_sw[0][10]~5_combout ),
	.cout());
defparam \lpp_ram_data_out_sw[0][10]~5 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out_sw[0][10]~5 .sum_lutc_input = "datac";

dffeas fft_dirn(
	.clk(clk),
	.d(\fft_dirn~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_dirn~q ),
	.prn(vcc));
defparam fft_dirn.is_wysiwyg = "true";
defparam fft_dirn.power_up = "low";

dffeas lpp_sel(
	.clk(clk),
	.d(\lpp_sel~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\lpp_sel~q ),
	.prn(vcc));
defparam lpp_sel.is_wysiwyg = "true";
defparam lpp_sel.power_up = "low";

dffeas \wren_b[0] (
	.clk(clk),
	.d(\wren_b~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\wren_b[0]~q ),
	.prn(vcc));
defparam \wren_b[0] .is_wysiwyg = "true";
defparam \wren_b[0] .power_up = "low";

dffeas \wren_a[0] (
	.clk(clk),
	.d(\wren_a~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\global_clock_enable~0_combout ),
	.q(\wren_a[0]~q ),
	.prn(vcc));
defparam \wren_a[0] .is_wysiwyg = "true";
defparam \wren_a[0] .power_up = "low";

dffeas \wren_b[1] (
	.clk(clk),
	.d(\wren_b~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\wren_b[1]~q ),
	.prn(vcc));
defparam \wren_b[1] .is_wysiwyg = "true";
defparam \wren_b[1] .power_up = "low";

dffeas \wren_a[1] (
	.clk(clk),
	.d(\wren_a~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\global_clock_enable~0_combout ),
	.q(\wren_a[1]~q ),
	.prn(vcc));
defparam \wren_a[1] .is_wysiwyg = "true";
defparam \wren_a[1] .power_up = "low";

dffeas \wren_b[2] (
	.clk(clk),
	.d(\wren_b~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\wren_b[2]~q ),
	.prn(vcc));
defparam \wren_b[2] .is_wysiwyg = "true";
defparam \wren_b[2] .power_up = "low";

dffeas \wren_a[2] (
	.clk(clk),
	.d(\wren_a~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\global_clock_enable~0_combout ),
	.q(\wren_a[2]~q ),
	.prn(vcc));
defparam \wren_a[2] .is_wysiwyg = "true";
defparam \wren_a[2] .power_up = "low";

dffeas \wren_b[3] (
	.clk(clk),
	.d(\wren_b~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\wren_b[3]~q ),
	.prn(vcc));
defparam \wren_b[3] .is_wysiwyg = "true";
defparam \wren_b[3] .power_up = "low";

dffeas \wren_a[3] (
	.clk(clk),
	.d(\wren_a~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\global_clock_enable~0_combout ),
	.q(\wren_a[3]~q ),
	.prn(vcc));
defparam \wren_a[3] .is_wysiwyg = "true";
defparam \wren_a[3] .power_up = "low";

dffeas \core_real_in[2] (
	.clk(clk),
	.d(\core_real_in~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\core_real_in[2]~q ),
	.prn(vcc));
defparam \core_real_in[2] .is_wysiwyg = "true";
defparam \core_real_in[2] .power_up = "low";

dffeas \core_real_in[6] (
	.clk(clk),
	.d(\core_real_in~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\core_real_in[6]~q ),
	.prn(vcc));
defparam \core_real_in[6] .is_wysiwyg = "true";
defparam \core_real_in[6] .power_up = "low";

dffeas \core_real_in[4] (
	.clk(clk),
	.d(\core_real_in~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\core_real_in[4]~q ),
	.prn(vcc));
defparam \core_real_in[4] .is_wysiwyg = "true";
defparam \core_real_in[4] .power_up = "low";

dffeas \core_real_in[3] (
	.clk(clk),
	.d(\core_real_in~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\core_real_in[3]~q ),
	.prn(vcc));
defparam \core_real_in[3] .is_wysiwyg = "true";
defparam \core_real_in[3] .power_up = "low";

dffeas \core_real_in[5] (
	.clk(clk),
	.d(\core_real_in~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\core_real_in[5]~q ),
	.prn(vcc));
defparam \core_real_in[5] .is_wysiwyg = "true";
defparam \core_real_in[5] .power_up = "low";

dffeas \core_real_in[1] (
	.clk(clk),
	.d(\core_real_in~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\core_real_in[1]~q ),
	.prn(vcc));
defparam \core_real_in[1] .is_wysiwyg = "true";
defparam \core_real_in[1] .power_up = "low";

dffeas \core_real_in[0] (
	.clk(clk),
	.d(\core_real_in~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\core_real_in[0]~q ),
	.prn(vcc));
defparam \core_real_in[0] .is_wysiwyg = "true";
defparam \core_real_in[0] .power_up = "low";

dffeas \core_real_in[7] (
	.clk(clk),
	.d(\core_real_in~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\core_real_in[7]~q ),
	.prn(vcc));
defparam \core_real_in[7] .is_wysiwyg = "true";
defparam \core_real_in[7] .power_up = "low";

dffeas \core_imag_in[7] (
	.clk(clk),
	.d(\core_imag_in~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\core_imag_in[7]~q ),
	.prn(vcc));
defparam \core_imag_in[7] .is_wysiwyg = "true";
defparam \core_imag_in[7] .power_up = "low";

dffeas \core_imag_in[3] (
	.clk(clk),
	.d(\core_imag_in~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\core_imag_in[3]~q ),
	.prn(vcc));
defparam \core_imag_in[3] .is_wysiwyg = "true";
defparam \core_imag_in[3] .power_up = "low";

dffeas \core_imag_in[5] (
	.clk(clk),
	.d(\core_imag_in~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\core_imag_in[5]~q ),
	.prn(vcc));
defparam \core_imag_in[5] .is_wysiwyg = "true";
defparam \core_imag_in[5] .power_up = "low";

dffeas \core_imag_in[4] (
	.clk(clk),
	.d(\core_imag_in~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\core_imag_in[4]~q ),
	.prn(vcc));
defparam \core_imag_in[4] .is_wysiwyg = "true";
defparam \core_imag_in[4] .power_up = "low";

dffeas \core_imag_in[6] (
	.clk(clk),
	.d(\core_imag_in~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\core_imag_in[6]~q ),
	.prn(vcc));
defparam \core_imag_in[6] .is_wysiwyg = "true";
defparam \core_imag_in[6] .power_up = "low";

dffeas \core_imag_in[2] (
	.clk(clk),
	.d(\core_imag_in~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\core_imag_in[2]~q ),
	.prn(vcc));
defparam \core_imag_in[2] .is_wysiwyg = "true";
defparam \core_imag_in[2] .power_up = "low";

dffeas \core_imag_in[1] (
	.clk(clk),
	.d(\core_imag_in~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\core_imag_in[1]~q ),
	.prn(vcc));
defparam \core_imag_in[1] .is_wysiwyg = "true";
defparam \core_imag_in[1] .power_up = "low";

dffeas \core_imag_in[0] (
	.clk(clk),
	.d(\core_imag_in~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\core_imag_in[0]~q ),
	.prn(vcc));
defparam \core_imag_in[0] .is_wysiwyg = "true";
defparam \core_imag_in[0] .power_up = "low";

dffeas master_sink_ena(
	.clk(clk),
	.d(reset_n),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\master_sink_ena~q ),
	.prn(vcc));
defparam master_sink_ena.is_wysiwyg = "true";
defparam master_sink_ena.power_up = "low";

dffeas master_source_ena(
	.clk(clk),
	.d(\master_source_ena~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\master_source_ena~q ),
	.prn(vcc));
defparam master_source_ena.is_wysiwyg = "true";
defparam master_source_ena.power_up = "low";

dffeas sink_ready_ctrl_d(
	.clk(clk),
	.d(\auk_dsp_interface_controller_1|sink_ready_ctrl~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sink_ready_ctrl_d~q ),
	.prn(vcc));
defparam sink_ready_ctrl_d.is_wysiwyg = "true";
defparam sink_ready_ctrl_d.power_up = "low";

dffeas sop(
	.clk(clk),
	.d(\sop~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sop~q ),
	.prn(vcc));
defparam sop.is_wysiwyg = "true";
defparam sop.power_up = "low";

cycloneiii_lcell_comb \source_valid_ctrl_sop~0 (
	.dataa(\auk_dsp_interface_controller_1|sink_stall_reg~q ),
	.datab(\sink_ready_ctrl_d~q ),
	.datac(\auk_dsp_atlantic_sink_1|send_sop_s~q ),
	.datad(\sop~q ),
	.cin(gnd),
	.combout(\source_valid_ctrl_sop~0_combout ),
	.cout());
defparam \source_valid_ctrl_sop~0 .lut_mask = 16'hBFFF;
defparam \source_valid_ctrl_sop~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \source_valid_ctrl_sop~1 (
	.dataa(gnd),
	.datab(\sink_ready_ctrl_d~q ),
	.datac(\auk_dsp_atlantic_sink_1|send_sop_s~q ),
	.datad(\sop~q ),
	.cin(gnd),
	.combout(\source_valid_ctrl_sop~1_combout ),
	.cout());
defparam \source_valid_ctrl_sop~1 .lut_mask = 16'h3FFF;
defparam \source_valid_ctrl_sop~1 .sum_lutc_input = "datac";

dffeas \exponent_out[0] (
	.clk(clk),
	.d(\exponent_out~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\exponent_out[0]~q ),
	.prn(vcc));
defparam \exponent_out[0] .is_wysiwyg = "true";
defparam \exponent_out[0] .power_up = "low";

dffeas \exponent_out[1] (
	.clk(clk),
	.d(\exponent_out~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\exponent_out[1]~q ),
	.prn(vcc));
defparam \exponent_out[1] .is_wysiwyg = "true";
defparam \exponent_out[1] .power_up = "low";

dffeas \exponent_out[2] (
	.clk(clk),
	.d(\exponent_out~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\exponent_out[2]~q ),
	.prn(vcc));
defparam \exponent_out[2] .is_wysiwyg = "true";
defparam \exponent_out[2] .power_up = "low";

dffeas \exponent_out[3] (
	.clk(clk),
	.d(\exponent_out~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\exponent_out[3]~q ),
	.prn(vcc));
defparam \exponent_out[3] .is_wysiwyg = "true";
defparam \exponent_out[3] .power_up = "low";

dffeas \exponent_out[4] (
	.clk(clk),
	.d(\exponent_out~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\exponent_out[4]~q ),
	.prn(vcc));
defparam \exponent_out[4] .is_wysiwyg = "true";
defparam \exponent_out[4] .power_up = "low";

dffeas \exponent_out[5] (
	.clk(clk),
	.d(\exponent_out~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\exponent_out[5]~q ),
	.prn(vcc));
defparam \exponent_out[5] .is_wysiwyg = "true";
defparam \exponent_out[5] .power_up = "low";

dffeas \fft_real_out[0] (
	.clk(clk),
	.d(\fft_real_out~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_real_out[0]~q ),
	.prn(vcc));
defparam \fft_real_out[0] .is_wysiwyg = "true";
defparam \fft_real_out[0] .power_up = "low";

dffeas \fft_real_out[1] (
	.clk(clk),
	.d(\fft_real_out~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_real_out[1]~q ),
	.prn(vcc));
defparam \fft_real_out[1] .is_wysiwyg = "true";
defparam \fft_real_out[1] .power_up = "low";

dffeas \fft_real_out[2] (
	.clk(clk),
	.d(\fft_real_out~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_real_out[2]~q ),
	.prn(vcc));
defparam \fft_real_out[2] .is_wysiwyg = "true";
defparam \fft_real_out[2] .power_up = "low";

dffeas \fft_real_out[3] (
	.clk(clk),
	.d(\fft_real_out~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_real_out[3]~q ),
	.prn(vcc));
defparam \fft_real_out[3] .is_wysiwyg = "true";
defparam \fft_real_out[3] .power_up = "low";

dffeas \fft_real_out[4] (
	.clk(clk),
	.d(\fft_real_out~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_real_out[4]~q ),
	.prn(vcc));
defparam \fft_real_out[4] .is_wysiwyg = "true";
defparam \fft_real_out[4] .power_up = "low";

dffeas \fft_real_out[5] (
	.clk(clk),
	.d(\fft_real_out~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_real_out[5]~q ),
	.prn(vcc));
defparam \fft_real_out[5] .is_wysiwyg = "true";
defparam \fft_real_out[5] .power_up = "low";

dffeas \fft_real_out[6] (
	.clk(clk),
	.d(\fft_real_out~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_real_out[6]~q ),
	.prn(vcc));
defparam \fft_real_out[6] .is_wysiwyg = "true";
defparam \fft_real_out[6] .power_up = "low";

dffeas \fft_real_out[7] (
	.clk(clk),
	.d(\fft_real_out~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_real_out[7]~q ),
	.prn(vcc));
defparam \fft_real_out[7] .is_wysiwyg = "true";
defparam \fft_real_out[7] .power_up = "low";

dffeas \fft_imag_out[0] (
	.clk(clk),
	.d(\fft_imag_out~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_imag_out[0]~q ),
	.prn(vcc));
defparam \fft_imag_out[0] .is_wysiwyg = "true";
defparam \fft_imag_out[0] .power_up = "low";

dffeas \fft_imag_out[1] (
	.clk(clk),
	.d(\fft_imag_out~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_imag_out[1]~q ),
	.prn(vcc));
defparam \fft_imag_out[1] .is_wysiwyg = "true";
defparam \fft_imag_out[1] .power_up = "low";

dffeas \fft_imag_out[2] (
	.clk(clk),
	.d(\fft_imag_out~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_imag_out[2]~q ),
	.prn(vcc));
defparam \fft_imag_out[2] .is_wysiwyg = "true";
defparam \fft_imag_out[2] .power_up = "low";

dffeas \fft_imag_out[3] (
	.clk(clk),
	.d(\fft_imag_out~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_imag_out[3]~q ),
	.prn(vcc));
defparam \fft_imag_out[3] .is_wysiwyg = "true";
defparam \fft_imag_out[3] .power_up = "low";

dffeas \fft_imag_out[4] (
	.clk(clk),
	.d(\fft_imag_out~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_imag_out[4]~q ),
	.prn(vcc));
defparam \fft_imag_out[4] .is_wysiwyg = "true";
defparam \fft_imag_out[4] .power_up = "low";

dffeas \fft_imag_out[5] (
	.clk(clk),
	.d(\fft_imag_out~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_imag_out[5]~q ),
	.prn(vcc));
defparam \fft_imag_out[5] .is_wysiwyg = "true";
defparam \fft_imag_out[5] .power_up = "low";

dffeas \fft_imag_out[6] (
	.clk(clk),
	.d(\fft_imag_out~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_imag_out[6]~q ),
	.prn(vcc));
defparam \fft_imag_out[6] .is_wysiwyg = "true";
defparam \fft_imag_out[6] .power_up = "low";

dffeas \fft_imag_out[7] (
	.clk(clk),
	.d(\fft_imag_out~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_imag_out[7]~q ),
	.prn(vcc));
defparam \fft_imag_out[7] .is_wysiwyg = "true";
defparam \fft_imag_out[7] .power_up = "low";

cycloneiii_lcell_comb \global_clock_enable~0 (
	.dataa(\auk_dsp_atlantic_source_1|source_stall_int_d~q ),
	.datab(\source_valid_ctrl_sop~1_combout ),
	.datac(gnd),
	.datad(\auk_dsp_interface_controller_1|stall_reg~q ),
	.cin(gnd),
	.combout(\global_clock_enable~0_combout ),
	.cout());
defparam \global_clock_enable~0 .lut_mask = 16'hDD11;
defparam \global_clock_enable~0 .sum_lutc_input = "datac";

dffeas oe(
	.clk(clk),
	.d(\val_out~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\oe~q ),
	.prn(vcc));
defparam oe.is_wysiwyg = "true";
defparam oe.power_up = "low";

cycloneiii_lcell_comb \master_source_ena~0 (
	.dataa(reset_n),
	.datab(\oe~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\master_source_ena~0_combout ),
	.cout());
defparam \master_source_ena~0 .lut_mask = 16'hEEEE;
defparam \master_source_ena~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sop~0 (
	.dataa(\auk_dsp_atlantic_sink_1|send_eop_s~q ),
	.datab(\sink_ready_ctrl_d~q ),
	.datac(\auk_dsp_atlantic_sink_1|send_sop_s~q ),
	.datad(\sop~q ),
	.cin(gnd),
	.combout(\sop~0_combout ),
	.cout());
defparam \sop~0 .lut_mask = 16'hF7D5;
defparam \sop~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Equal0~0 (
	.dataa(\data_count_sig[0]~q ),
	.datab(\data_count_sig[1]~q ),
	.datac(\data_count_sig[2]~q ),
	.datad(\data_count_sig[3]~q ),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
defparam \Equal0~0 .lut_mask = 16'h7FFF;
defparam \Equal0~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Equal0~1 (
	.dataa(\data_count_sig[4]~q ),
	.datab(\data_count_sig[5]~q ),
	.datac(\data_count_sig[6]~q ),
	.datad(\data_count_sig[7]~q ),
	.cin(gnd),
	.combout(\Equal0~1_combout ),
	.cout());
defparam \Equal0~1 .lut_mask = 16'h7FFF;
defparam \Equal0~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \LessThan0~0 (
	.dataa(\data_count_sig[0]~q ),
	.datab(\data_count_sig[1]~q ),
	.datac(\data_count_sig[2]~q ),
	.datad(\data_count_sig[3]~q ),
	.cin(gnd),
	.combout(\LessThan0~0_combout ),
	.cout());
defparam \LessThan0~0 .lut_mask = 16'h7FFF;
defparam \LessThan0~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \LessThan0~1 (
	.dataa(\data_count_sig[4]~q ),
	.datab(\data_count_sig[5]~q ),
	.datac(\data_count_sig[6]~q ),
	.datad(\data_count_sig[7]~q ),
	.cin(gnd),
	.combout(\LessThan0~1_combout ),
	.cout());
defparam \LessThan0~1 .lut_mask = 16'h7FFF;
defparam \LessThan0~1 .sum_lutc_input = "datac";

dffeas master_source_sop(
	.clk(clk),
	.d(\master_source_sop~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\master_source_sop~q ),
	.prn(vcc));
defparam master_source_sop.is_wysiwyg = "true";
defparam master_source_sop.power_up = "low";

cycloneiii_lcell_comb \data_count_sig[0]~17 (
	.dataa(\LessThan0~0_combout ),
	.datab(\LessThan0~1_combout ),
	.datac(\data_count_sig[8]~q ),
	.datad(\master_source_sop~q ),
	.cin(gnd),
	.combout(\data_count_sig[0]~17_combout ),
	.cout());
defparam \data_count_sig[0]~17 .lut_mask = 16'hEFFF;
defparam \data_count_sig[0]~17 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \data_count_sig[0]~18 (
	.dataa(\Equal0~0_combout ),
	.datab(\Equal0~1_combout ),
	.datac(\data_count_sig[8]~q ),
	.datad(\data_count_sig[0]~17_combout ),
	.cin(gnd),
	.combout(\data_count_sig[0]~18_combout ),
	.cout());
defparam \data_count_sig[0]~18 .lut_mask = 16'hEFFF;
defparam \data_count_sig[0]~18 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \data_count_sig[0]~19 (
	.dataa(\data_count_sig[8]~q ),
	.datab(\master_source_sop~q ),
	.datac(\Equal0~0_combout ),
	.datad(\Equal0~1_combout ),
	.cin(gnd),
	.combout(\data_count_sig[0]~19_combout ),
	.cout());
defparam \data_count_sig[0]~19 .lut_mask = 16'hFFF7;
defparam \data_count_sig[0]~19 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \data_count_sig[0]~20 (
	.dataa(\auk_dsp_atlantic_source_1|source_stall_int_d~q ),
	.datab(\source_valid_ctrl_sop~1_combout ),
	.datac(\auk_dsp_interface_controller_1|stall_reg~q ),
	.datad(\data_count_sig[0]~19_combout ),
	.cin(gnd),
	.combout(\data_count_sig[0]~20_combout ),
	.cout());
defparam \data_count_sig[0]~20 .lut_mask = 16'hD1FF;
defparam \data_count_sig[0]~20 .sum_lutc_input = "datac";

dffeas \blk_exp_accum[0] (
	.clk(clk),
	.d(\Selector5~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\blk_exp_accum[0]~q ),
	.prn(vcc));
defparam \blk_exp_accum[0] .is_wysiwyg = "true";
defparam \blk_exp_accum[0] .power_up = "low";

cycloneiii_lcell_comb \exponent_out~0 (
	.dataa(reset_n),
	.datab(\oe~q ),
	.datac(\blk_exp_accum[0]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\exponent_out~0_combout ),
	.cout());
defparam \exponent_out~0 .lut_mask = 16'hFEFE;
defparam \exponent_out~0 .sum_lutc_input = "datac";

dffeas \blk_exp_accum[1] (
	.clk(clk),
	.d(\Selector4~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\blk_exp_accum[1]~q ),
	.prn(vcc));
defparam \blk_exp_accum[1] .is_wysiwyg = "true";
defparam \blk_exp_accum[1] .power_up = "low";

cycloneiii_lcell_comb \exponent_out~1 (
	.dataa(reset_n),
	.datab(\oe~q ),
	.datac(\blk_exp_accum[1]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\exponent_out~1_combout ),
	.cout());
defparam \exponent_out~1 .lut_mask = 16'hFEFE;
defparam \exponent_out~1 .sum_lutc_input = "datac";

dffeas \blk_exp_accum[2] (
	.clk(clk),
	.d(\Selector3~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\blk_exp_accum[2]~q ),
	.prn(vcc));
defparam \blk_exp_accum[2] .is_wysiwyg = "true";
defparam \blk_exp_accum[2] .power_up = "low";

cycloneiii_lcell_comb \exponent_out~2 (
	.dataa(reset_n),
	.datab(\oe~q ),
	.datac(\blk_exp_accum[2]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\exponent_out~2_combout ),
	.cout());
defparam \exponent_out~2 .lut_mask = 16'hFEFE;
defparam \exponent_out~2 .sum_lutc_input = "datac";

dffeas \blk_exp_accum[3] (
	.clk(clk),
	.d(\Selector2~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\blk_exp_accum[3]~q ),
	.prn(vcc));
defparam \blk_exp_accum[3] .is_wysiwyg = "true";
defparam \blk_exp_accum[3] .power_up = "low";

cycloneiii_lcell_comb \exponent_out~3 (
	.dataa(reset_n),
	.datab(\oe~q ),
	.datac(\blk_exp_accum[3]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\exponent_out~3_combout ),
	.cout());
defparam \exponent_out~3 .lut_mask = 16'hFEFE;
defparam \exponent_out~3 .sum_lutc_input = "datac";

dffeas \blk_exp_accum[4] (
	.clk(clk),
	.d(\Selector1~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\blk_exp_accum[4]~q ),
	.prn(vcc));
defparam \blk_exp_accum[4] .is_wysiwyg = "true";
defparam \blk_exp_accum[4] .power_up = "low";

cycloneiii_lcell_comb \exponent_out~4 (
	.dataa(reset_n),
	.datab(\oe~q ),
	.datac(\blk_exp_accum[4]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\exponent_out~4_combout ),
	.cout());
defparam \exponent_out~4 .lut_mask = 16'hFEFE;
defparam \exponent_out~4 .sum_lutc_input = "datac";

dffeas \blk_exp_accum[5] (
	.clk(clk),
	.d(\Selector0~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\blk_exp_accum[5]~q ),
	.prn(vcc));
defparam \blk_exp_accum[5] .is_wysiwyg = "true";
defparam \blk_exp_accum[5] .power_up = "low";

cycloneiii_lcell_comb \exponent_out~5 (
	.dataa(reset_n),
	.datab(\oe~q ),
	.datac(\blk_exp_accum[5]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\exponent_out~5_combout ),
	.cout());
defparam \exponent_out~5 .lut_mask = 16'hFEFE;
defparam \exponent_out~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \fft_real_out~0 (
	.dataa(\master_source_ena~0_combout ),
	.datab(\gen_radix_2_last_pass:lpp_r2|data_imag_o[0]~q ),
	.datac(\gen_radix_2_last_pass:lpp_r2|data_real_o[0]~q ),
	.datad(\fft_dirn_stream~q ),
	.cin(gnd),
	.combout(\fft_real_out~0_combout ),
	.cout());
defparam \fft_real_out~0 .lut_mask = 16'hFAFC;
defparam \fft_real_out~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \fft_real_out~1 (
	.dataa(\master_source_ena~0_combout ),
	.datab(\gen_radix_2_last_pass:lpp_r2|data_imag_o[1]~q ),
	.datac(\gen_radix_2_last_pass:lpp_r2|data_real_o[1]~q ),
	.datad(\fft_dirn_stream~q ),
	.cin(gnd),
	.combout(\fft_real_out~1_combout ),
	.cout());
defparam \fft_real_out~1 .lut_mask = 16'hFAFC;
defparam \fft_real_out~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \fft_real_out~2 (
	.dataa(\master_source_ena~0_combout ),
	.datab(\gen_radix_2_last_pass:lpp_r2|data_imag_o[2]~q ),
	.datac(\gen_radix_2_last_pass:lpp_r2|data_real_o[2]~q ),
	.datad(\fft_dirn_stream~q ),
	.cin(gnd),
	.combout(\fft_real_out~2_combout ),
	.cout());
defparam \fft_real_out~2 .lut_mask = 16'hFAFC;
defparam \fft_real_out~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \fft_real_out~3 (
	.dataa(\master_source_ena~0_combout ),
	.datab(\gen_radix_2_last_pass:lpp_r2|data_imag_o[3]~q ),
	.datac(\gen_radix_2_last_pass:lpp_r2|data_real_o[3]~q ),
	.datad(\fft_dirn_stream~q ),
	.cin(gnd),
	.combout(\fft_real_out~3_combout ),
	.cout());
defparam \fft_real_out~3 .lut_mask = 16'hFAFC;
defparam \fft_real_out~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \fft_real_out~4 (
	.dataa(\master_source_ena~0_combout ),
	.datab(\gen_radix_2_last_pass:lpp_r2|data_imag_o[4]~q ),
	.datac(\gen_radix_2_last_pass:lpp_r2|data_real_o[4]~q ),
	.datad(\fft_dirn_stream~q ),
	.cin(gnd),
	.combout(\fft_real_out~4_combout ),
	.cout());
defparam \fft_real_out~4 .lut_mask = 16'hFAFC;
defparam \fft_real_out~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \fft_real_out~5 (
	.dataa(\master_source_ena~0_combout ),
	.datab(\gen_radix_2_last_pass:lpp_r2|data_imag_o[5]~q ),
	.datac(\gen_radix_2_last_pass:lpp_r2|data_real_o[5]~q ),
	.datad(\fft_dirn_stream~q ),
	.cin(gnd),
	.combout(\fft_real_out~5_combout ),
	.cout());
defparam \fft_real_out~5 .lut_mask = 16'hFAFC;
defparam \fft_real_out~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \fft_real_out~6 (
	.dataa(\master_source_ena~0_combout ),
	.datab(\gen_radix_2_last_pass:lpp_r2|data_imag_o[6]~q ),
	.datac(\gen_radix_2_last_pass:lpp_r2|data_real_o[6]~q ),
	.datad(\fft_dirn_stream~q ),
	.cin(gnd),
	.combout(\fft_real_out~6_combout ),
	.cout());
defparam \fft_real_out~6 .lut_mask = 16'hFAFC;
defparam \fft_real_out~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \fft_real_out~7 (
	.dataa(\master_source_ena~0_combout ),
	.datab(\gen_radix_2_last_pass:lpp_r2|data_imag_o[7]~q ),
	.datac(\gen_radix_2_last_pass:lpp_r2|data_real_o[7]~q ),
	.datad(\fft_dirn_stream~q ),
	.cin(gnd),
	.combout(\fft_real_out~7_combout ),
	.cout());
defparam \fft_real_out~7 .lut_mask = 16'hFAFC;
defparam \fft_real_out~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \fft_imag_out~0 (
	.dataa(\master_source_ena~0_combout ),
	.datab(\gen_radix_2_last_pass:lpp_r2|data_real_o[0]~q ),
	.datac(\gen_radix_2_last_pass:lpp_r2|data_imag_o[0]~q ),
	.datad(\fft_dirn_stream~q ),
	.cin(gnd),
	.combout(\fft_imag_out~0_combout ),
	.cout());
defparam \fft_imag_out~0 .lut_mask = 16'hFAFC;
defparam \fft_imag_out~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \fft_imag_out~1 (
	.dataa(\master_source_ena~0_combout ),
	.datab(\gen_radix_2_last_pass:lpp_r2|data_real_o[1]~q ),
	.datac(\gen_radix_2_last_pass:lpp_r2|data_imag_o[1]~q ),
	.datad(\fft_dirn_stream~q ),
	.cin(gnd),
	.combout(\fft_imag_out~1_combout ),
	.cout());
defparam \fft_imag_out~1 .lut_mask = 16'hFAFC;
defparam \fft_imag_out~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \fft_imag_out~2 (
	.dataa(\master_source_ena~0_combout ),
	.datab(\gen_radix_2_last_pass:lpp_r2|data_real_o[2]~q ),
	.datac(\gen_radix_2_last_pass:lpp_r2|data_imag_o[2]~q ),
	.datad(\fft_dirn_stream~q ),
	.cin(gnd),
	.combout(\fft_imag_out~2_combout ),
	.cout());
defparam \fft_imag_out~2 .lut_mask = 16'hFAFC;
defparam \fft_imag_out~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \fft_imag_out~3 (
	.dataa(\master_source_ena~0_combout ),
	.datab(\gen_radix_2_last_pass:lpp_r2|data_real_o[3]~q ),
	.datac(\gen_radix_2_last_pass:lpp_r2|data_imag_o[3]~q ),
	.datad(\fft_dirn_stream~q ),
	.cin(gnd),
	.combout(\fft_imag_out~3_combout ),
	.cout());
defparam \fft_imag_out~3 .lut_mask = 16'hFAFC;
defparam \fft_imag_out~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \fft_imag_out~4 (
	.dataa(\master_source_ena~0_combout ),
	.datab(\gen_radix_2_last_pass:lpp_r2|data_real_o[4]~q ),
	.datac(\gen_radix_2_last_pass:lpp_r2|data_imag_o[4]~q ),
	.datad(\fft_dirn_stream~q ),
	.cin(gnd),
	.combout(\fft_imag_out~4_combout ),
	.cout());
defparam \fft_imag_out~4 .lut_mask = 16'hFAFC;
defparam \fft_imag_out~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \fft_imag_out~5 (
	.dataa(\master_source_ena~0_combout ),
	.datab(\gen_radix_2_last_pass:lpp_r2|data_real_o[5]~q ),
	.datac(\gen_radix_2_last_pass:lpp_r2|data_imag_o[5]~q ),
	.datad(\fft_dirn_stream~q ),
	.cin(gnd),
	.combout(\fft_imag_out~5_combout ),
	.cout());
defparam \fft_imag_out~5 .lut_mask = 16'hFAFC;
defparam \fft_imag_out~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \fft_imag_out~6 (
	.dataa(\master_source_ena~0_combout ),
	.datab(\gen_radix_2_last_pass:lpp_r2|data_real_o[6]~q ),
	.datac(\gen_radix_2_last_pass:lpp_r2|data_imag_o[6]~q ),
	.datad(\fft_dirn_stream~q ),
	.cin(gnd),
	.combout(\fft_imag_out~6_combout ),
	.cout());
defparam \fft_imag_out~6 .lut_mask = 16'hFAFC;
defparam \fft_imag_out~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \fft_imag_out~7 (
	.dataa(\master_source_ena~0_combout ),
	.datab(\gen_radix_2_last_pass:lpp_r2|data_real_o[7]~q ),
	.datac(\gen_radix_2_last_pass:lpp_r2|data_imag_o[7]~q ),
	.datad(\fft_dirn_stream~q ),
	.cin(gnd),
	.combout(\fft_imag_out~7_combout ),
	.cout());
defparam \fft_imag_out~7 .lut_mask = 16'hFAFC;
defparam \fft_imag_out~7 .sum_lutc_input = "datac";

dffeas \fft_s2_cur.IDLE (
	.clk(clk),
	.d(reset_n),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\fft_s2_cur.IDLE~0_combout ),
	.q(\fft_s2_cur.IDLE~q ),
	.prn(vcc));
defparam \fft_s2_cur.IDLE .is_wysiwyg = "true";
defparam \fft_s2_cur.IDLE .power_up = "low";

cycloneiii_lcell_comb \val_out~1 (
	.dataa(\fft_s2_cur.WAIT_FOR_LPP_INPUT~q ),
	.datab(gnd),
	.datac(reset_n),
	.datad(\fft_s2_cur.IDLE~q ),
	.cin(gnd),
	.combout(\val_out~1_combout ),
	.cout());
defparam \val_out~1 .lut_mask = 16'hFFF5;
defparam \val_out~1 .sum_lutc_input = "datac";

dffeas sop_out(
	.clk(clk),
	.d(\sop_out~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\sop_out~q ),
	.prn(vcc));
defparam sop_out.is_wysiwyg = "true";
defparam sop_out.power_up = "low";

cycloneiii_lcell_comb \master_source_sop~0 (
	.dataa(reset_n),
	.datab(\oe~q ),
	.datac(\sop_out~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\master_source_sop~0_combout ),
	.cout());
defparam \master_source_sop~0 .lut_mask = 16'hFEFE;
defparam \master_source_sop~0 .sum_lutc_input = "datac";

dffeas \fft_s2_cur.FIRST_LPP_C (
	.clk(clk),
	.d(\fft_s2_cur~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_s2_cur.FIRST_LPP_C~q ),
	.prn(vcc));
defparam \fft_s2_cur.FIRST_LPP_C .is_wysiwyg = "true";
defparam \fft_s2_cur.FIRST_LPP_C .power_up = "low";

cycloneiii_lcell_comb \Selector5~0 (
	.dataa(\gen_dft_2:bfpc|blk_exp[0]~q ),
	.datab(\blk_exp_accum[0]~q ),
	.datac(\fft_s2_cur.IDLE~q ),
	.datad(\fft_s2_cur.FIRST_LPP_C~q ),
	.cin(gnd),
	.combout(\Selector5~0_combout ),
	.cout());
defparam \Selector5~0 .lut_mask = 16'hFAFC;
defparam \Selector5~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector4~0 (
	.dataa(\gen_dft_2:bfpc|blk_exp[1]~q ),
	.datab(\blk_exp_accum[1]~q ),
	.datac(\fft_s2_cur.IDLE~q ),
	.datad(\fft_s2_cur.FIRST_LPP_C~q ),
	.cin(gnd),
	.combout(\Selector4~0_combout ),
	.cout());
defparam \Selector4~0 .lut_mask = 16'hFAFC;
defparam \Selector4~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector3~0 (
	.dataa(\gen_dft_2:bfpc|blk_exp[2]~q ),
	.datab(\blk_exp_accum[2]~q ),
	.datac(\fft_s2_cur.IDLE~q ),
	.datad(\fft_s2_cur.FIRST_LPP_C~q ),
	.cin(gnd),
	.combout(\Selector3~0_combout ),
	.cout());
defparam \Selector3~0 .lut_mask = 16'hFAFC;
defparam \Selector3~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector2~0 (
	.dataa(\gen_dft_2:bfpc|blk_exp[3]~q ),
	.datab(\blk_exp_accum[3]~q ),
	.datac(\fft_s2_cur.IDLE~q ),
	.datad(\fft_s2_cur.FIRST_LPP_C~q ),
	.cin(gnd),
	.combout(\Selector2~0_combout ),
	.cout());
defparam \Selector2~0 .lut_mask = 16'hFAFC;
defparam \Selector2~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector1~0 (
	.dataa(\gen_dft_2:bfpc|blk_exp[4]~q ),
	.datab(\blk_exp_accum[4]~q ),
	.datac(\fft_s2_cur.IDLE~q ),
	.datad(\fft_s2_cur.FIRST_LPP_C~q ),
	.cin(gnd),
	.combout(\Selector1~0_combout ),
	.cout());
defparam \Selector1~0 .lut_mask = 16'hFAFC;
defparam \Selector1~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector0~0 (
	.dataa(\gen_dft_2:bfpc|blk_exp[5]~q ),
	.datab(\blk_exp_accum[5]~q ),
	.datac(\fft_s2_cur.IDLE~q ),
	.datad(\fft_s2_cur.FIRST_LPP_C~q ),
	.cin(gnd),
	.combout(\Selector0~0_combout ),
	.cout());
defparam \Selector0~0 .lut_mask = 16'hFAFC;
defparam \Selector0~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \fft_dirn_stream~0 (
	.dataa(\fft_dirn_held_o2~q ),
	.datab(\fft_dirn_stream~q ),
	.datac(gnd),
	.datad(\fft_s2_cur.FIRST_LPP_C~q ),
	.cin(gnd),
	.combout(\fft_dirn_stream~0_combout ),
	.cout());
defparam \fft_dirn_stream~0 .lut_mask = 16'hAACC;
defparam \fft_dirn_stream~0 .sum_lutc_input = "datac";

dffeas \fft_s2_cur.LAST_LPP_C (
	.clk(clk),
	.d(\fft_s2_cur.IDLE~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\fft_s2_cur.IDLE~0_combout ),
	.q(\fft_s2_cur.LAST_LPP_C~q ),
	.prn(vcc));
defparam \fft_s2_cur.LAST_LPP_C .is_wysiwyg = "true";
defparam \fft_s2_cur.LAST_LPP_C .power_up = "low";

cycloneiii_lcell_comb \Selector20~0 (
	.dataa(\fft_s2_cur.WAIT_FOR_LPP_INPUT~q ),
	.datab(\fft_s2_cur.LAST_LPP_C~q ),
	.datac(\delay_lpp_en|tdl_arr[3]~q ),
	.datad(\fft_s2_cur.IDLE~q ),
	.cin(gnd),
	.combout(\Selector20~0_combout ),
	.cout());
defparam \Selector20~0 .lut_mask = 16'hEFFF;
defparam \Selector20~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Equal4~0 (
	.dataa(\lpp_count_offset[0]~q ),
	.datab(\lpp_count_offset[1]~q ),
	.datac(\lpp_count_offset[2]~q ),
	.datad(\lpp_count_offset[3]~q ),
	.cin(gnd),
	.combout(\Equal4~0_combout ),
	.cout());
defparam \Equal4~0 .lut_mask = 16'h7FFF;
defparam \Equal4~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Equal4~1 (
	.dataa(\lpp_count_offset[4]~q ),
	.datab(\lpp_count_offset[5]~q ),
	.datac(\lpp_count_offset[6]~q ),
	.datad(\lpp_count_offset[7]~q ),
	.cin(gnd),
	.combout(\Equal4~1_combout ),
	.cout());
defparam \Equal4~1 .lut_mask = 16'h7FFF;
defparam \Equal4~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Equal4~2 (
	.dataa(\Equal4~0_combout ),
	.datab(\Equal4~1_combout ),
	.datac(gnd),
	.datad(\lpp_count_offset[8]~q ),
	.cin(gnd),
	.combout(\Equal4~2_combout ),
	.cout());
defparam \Equal4~2 .lut_mask = 16'hEEFF;
defparam \Equal4~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \fft_s2_cur.IDLE~0 (
	.dataa(\global_clock_enable~0_combout ),
	.datab(reset_n),
	.datac(\fft_s2_cur.LPP_C_OUTPUT~q ),
	.datad(\Equal4~2_combout ),
	.cin(gnd),
	.combout(\fft_s2_cur.IDLE~0_combout ),
	.cout());
defparam \fft_s2_cur.IDLE~0 .lut_mask = 16'hBFFF;
defparam \fft_s2_cur.IDLE~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sop_out~0 (
	.dataa(reset_n),
	.datab(\fft_s2_cur.FIRST_LPP_C~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sop_out~0_combout ),
	.cout());
defparam \sop_out~0 .lut_mask = 16'hEEEE;
defparam \sop_out~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \fft_s2_cur~9 (
	.dataa(reset_n),
	.datab(\delay_lpp_en|tdl_arr[3]~q ),
	.datac(\fft_s2_cur.WAIT_FOR_LPP_INPUT~q ),
	.datad(\fft_s2_cur.LAST_LPP_C~q ),
	.cin(gnd),
	.combout(\fft_s2_cur~9_combout ),
	.cout());
defparam \fft_s2_cur~9 .lut_mask = 16'hFFFE;
defparam \fft_s2_cur~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \fft_dirn_held_o2~0 (
	.dataa(\fft_dirn_held_o~q ),
	.datab(\fft_dirn_held_o2~q ),
	.datac(gnd),
	.datad(\gen_gt256_mk:ctrl|blk_done_int~q ),
	.cin(gnd),
	.combout(\fft_dirn_held_o2~0_combout ),
	.cout());
defparam \fft_dirn_held_o2~0 .lut_mask = 16'hAACC;
defparam \fft_dirn_held_o2~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \fft_s2_cur.IDLE~1 (
	.dataa(reset_n),
	.datab(\fft_s2_cur.LPP_C_OUTPUT~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fft_s2_cur.IDLE~1_combout ),
	.cout());
defparam \fft_s2_cur.IDLE~1 .lut_mask = 16'hEEEE;
defparam \fft_s2_cur.IDLE~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector22~0 (
	.dataa(\fft_s2_cur.FIRST_LPP_C~q ),
	.datab(\fft_s2_cur.LPP_C_OUTPUT~q ),
	.datac(\Equal4~2_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector22~0_combout ),
	.cout());
defparam \Selector22~0 .lut_mask = 16'hFEFE;
defparam \Selector22~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_count_offset[0]~11 (
	.dataa(reset_n),
	.datab(\fft_s2_cur.WAIT_FOR_LPP_INPUT~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\lpp_count_offset[0]~11_combout ),
	.cout());
defparam \lpp_count_offset[0]~11 .lut_mask = 16'hEEEE;
defparam \lpp_count_offset[0]~11 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_count_offset[0]~12 (
	.dataa(\auk_dsp_atlantic_source_1|source_stall_int_d~q ),
	.datab(\source_valid_ctrl_sop~1_combout ),
	.datac(\auk_dsp_interface_controller_1|stall_reg~q ),
	.datad(\lpp_count_offset[0]~11_combout ),
	.cin(gnd),
	.combout(\lpp_count_offset[0]~12_combout ),
	.cout());
defparam \lpp_count_offset[0]~12 .lut_mask = 16'hD1FF;
defparam \lpp_count_offset[0]~12 .sum_lutc_input = "datac";

dffeas fft_dirn_held(
	.clk(clk),
	.d(\fft_dirn_held~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_dirn_held~q ),
	.prn(vcc));
defparam fft_dirn_held.is_wysiwyg = "true";
defparam fft_dirn_held.power_up = "low";

cycloneiii_lcell_comb \fft_dirn_held_o~0 (
	.dataa(\fft_dirn_held~q ),
	.datab(\fft_dirn_held_o~q ),
	.datac(gnd),
	.datad(\writer|next_block~q ),
	.cin(gnd),
	.combout(\fft_dirn_held_o~0_combout ),
	.cout());
defparam \fft_dirn_held_o~0 .lut_mask = 16'hAACC;
defparam \fft_dirn_held_o~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector14~0 (
	.dataa(\fft_s2_cur.WAIT_FOR_LPP_INPUT~q ),
	.datab(\fft_s2_cur.IDLE~q ),
	.datac(\Add2~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector14~0_combout ),
	.cout());
defparam \Selector14~0 .lut_mask = 16'hFEFE;
defparam \Selector14~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_count~0 (
	.dataa(\fft_s2_cur.IDLE~q ),
	.datab(\Add2~2_combout ),
	.datac(gnd),
	.datad(\fft_s2_cur.WAIT_FOR_LPP_INPUT~q ),
	.cin(gnd),
	.combout(\lpp_count~0_combout ),
	.cout());
defparam \lpp_count~0 .lut_mask = 16'hEEFF;
defparam \lpp_count~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector13~0 (
	.dataa(\fft_s2_cur.WAIT_FOR_LPP_INPUT~q ),
	.datab(\fft_s2_cur.IDLE~q ),
	.datac(\Add2~4_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector13~0_combout ),
	.cout());
defparam \Selector13~0 .lut_mask = 16'hFEFE;
defparam \Selector13~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector12~0 (
	.dataa(\fft_s2_cur.WAIT_FOR_LPP_INPUT~q ),
	.datab(\fft_s2_cur.IDLE~q ),
	.datac(\Add2~6_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector12~0_combout ),
	.cout());
defparam \Selector12~0 .lut_mask = 16'hFEFE;
defparam \Selector12~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector11~0 (
	.dataa(\fft_s2_cur.WAIT_FOR_LPP_INPUT~q ),
	.datab(\fft_s2_cur.IDLE~q ),
	.datac(\Add2~8_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector11~0_combout ),
	.cout());
defparam \Selector11~0 .lut_mask = 16'hFEFE;
defparam \Selector11~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector10~0 (
	.dataa(\fft_s2_cur.WAIT_FOR_LPP_INPUT~q ),
	.datab(\fft_s2_cur.IDLE~q ),
	.datac(\Add2~10_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector10~0_combout ),
	.cout());
defparam \Selector10~0 .lut_mask = 16'hFEFE;
defparam \Selector10~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector9~0 (
	.dataa(\fft_s2_cur.WAIT_FOR_LPP_INPUT~q ),
	.datab(\fft_s2_cur.IDLE~q ),
	.datac(\Add2~12_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector9~0_combout ),
	.cout());
defparam \Selector9~0 .lut_mask = 16'hFEFE;
defparam \Selector9~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector8~0 (
	.dataa(\fft_s2_cur.WAIT_FOR_LPP_INPUT~q ),
	.datab(\fft_s2_cur.IDLE~q ),
	.datac(\Add2~14_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector8~0_combout ),
	.cout());
defparam \Selector8~0 .lut_mask = 16'hFEFE;
defparam \Selector8~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector7~0 (
	.dataa(\fft_s2_cur.WAIT_FOR_LPP_INPUT~q ),
	.datab(\fft_s2_cur.IDLE~q ),
	.datac(\Add2~16_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector7~0_combout ),
	.cout());
defparam \Selector7~0 .lut_mask = 16'hFEFE;
defparam \Selector7~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux30~0 (
	.dataa(\lpp_ram_data_out[2][1]~q ),
	.datab(\lpp_ram_data_out[1][1]~q ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.cin(gnd),
	.combout(\Mux30~0_combout ),
	.cout());
defparam \Mux30~0 .lut_mask = 16'hAACC;
defparam \Mux30~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux30~1 (
	.dataa(\lpp_ram_data_out[0][1]~q ),
	.datab(\lpp_ram_data_out[3][1]~q ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.cin(gnd),
	.combout(\Mux30~1_combout ),
	.cout());
defparam \Mux30~1 .lut_mask = 16'hAACC;
defparam \Mux30~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux30~2 (
	.dataa(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.datab(\lpp_ram_data_out[2][1]~q ),
	.datac(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.datad(\lpp_ram_data_out[0][1]~q ),
	.cin(gnd),
	.combout(\Mux30~2_combout ),
	.cout());
defparam \Mux30~2 .lut_mask = 16'hFFDE;
defparam \Mux30~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux30~3 (
	.dataa(\lpp_ram_data_out[1][1]~q ),
	.datab(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.datac(\Mux30~2_combout ),
	.datad(\lpp_ram_data_out[3][1]~q ),
	.cin(gnd),
	.combout(\Mux30~3_combout ),
	.cout());
defparam \Mux30~3 .lut_mask = 16'hFFBE;
defparam \Mux30~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux31~0 (
	.dataa(\lpp_ram_data_out[2][0]~q ),
	.datab(\lpp_ram_data_out[1][0]~q ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.cin(gnd),
	.combout(\Mux31~0_combout ),
	.cout());
defparam \Mux31~0 .lut_mask = 16'hAACC;
defparam \Mux31~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux31~1 (
	.dataa(\lpp_ram_data_out[0][0]~q ),
	.datab(\lpp_ram_data_out[3][0]~q ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.cin(gnd),
	.combout(\Mux31~1_combout ),
	.cout());
defparam \Mux31~1 .lut_mask = 16'hAACC;
defparam \Mux31~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux31~2 (
	.dataa(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.datab(\lpp_ram_data_out[1][0]~q ),
	.datac(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.datad(\lpp_ram_data_out[0][0]~q ),
	.cin(gnd),
	.combout(\Mux31~2_combout ),
	.cout());
defparam \Mux31~2 .lut_mask = 16'hFFDE;
defparam \Mux31~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux31~3 (
	.dataa(\lpp_ram_data_out[2][0]~q ),
	.datab(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.datac(\Mux31~2_combout ),
	.datad(\lpp_ram_data_out[3][0]~q ),
	.cin(gnd),
	.combout(\Mux31~3_combout ),
	.cout());
defparam \Mux31~3 .lut_mask = 16'hFFBE;
defparam \Mux31~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux24~0 (
	.dataa(\lpp_ram_data_out[2][7]~q ),
	.datab(\lpp_ram_data_out[1][7]~q ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.cin(gnd),
	.combout(\Mux24~0_combout ),
	.cout());
defparam \Mux24~0 .lut_mask = 16'hAACC;
defparam \Mux24~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux24~1 (
	.dataa(\lpp_ram_data_out[0][7]~q ),
	.datab(\lpp_ram_data_out[3][7]~q ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.cin(gnd),
	.combout(\Mux24~1_combout ),
	.cout());
defparam \Mux24~1 .lut_mask = 16'hAACC;
defparam \Mux24~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux24~2 (
	.dataa(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.datab(\lpp_ram_data_out[2][7]~q ),
	.datac(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.datad(\lpp_ram_data_out[0][7]~q ),
	.cin(gnd),
	.combout(\Mux24~2_combout ),
	.cout());
defparam \Mux24~2 .lut_mask = 16'hFFDE;
defparam \Mux24~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux24~3 (
	.dataa(\lpp_ram_data_out[1][7]~q ),
	.datab(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.datac(\Mux24~2_combout ),
	.datad(\lpp_ram_data_out[3][7]~q ),
	.cin(gnd),
	.combout(\Mux24~3_combout ),
	.cout());
defparam \Mux24~3 .lut_mask = 16'hFFBE;
defparam \Mux24~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux25~0 (
	.dataa(\lpp_ram_data_out[2][6]~q ),
	.datab(\lpp_ram_data_out[1][6]~q ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.cin(gnd),
	.combout(\Mux25~0_combout ),
	.cout());
defparam \Mux25~0 .lut_mask = 16'hAACC;
defparam \Mux25~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux25~1 (
	.dataa(\lpp_ram_data_out[0][6]~q ),
	.datab(\lpp_ram_data_out[3][6]~q ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.cin(gnd),
	.combout(\Mux25~1_combout ),
	.cout());
defparam \Mux25~1 .lut_mask = 16'hAACC;
defparam \Mux25~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux25~2 (
	.dataa(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.datab(\lpp_ram_data_out[1][6]~q ),
	.datac(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.datad(\lpp_ram_data_out[0][6]~q ),
	.cin(gnd),
	.combout(\Mux25~2_combout ),
	.cout());
defparam \Mux25~2 .lut_mask = 16'hFFDE;
defparam \Mux25~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux25~3 (
	.dataa(\lpp_ram_data_out[2][6]~q ),
	.datab(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.datac(\Mux25~2_combout ),
	.datad(\lpp_ram_data_out[3][6]~q ),
	.cin(gnd),
	.combout(\Mux25~3_combout ),
	.cout());
defparam \Mux25~3 .lut_mask = 16'hFFBE;
defparam \Mux25~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux26~0 (
	.dataa(\lpp_ram_data_out[2][5]~q ),
	.datab(\lpp_ram_data_out[1][5]~q ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.cin(gnd),
	.combout(\Mux26~0_combout ),
	.cout());
defparam \Mux26~0 .lut_mask = 16'hAACC;
defparam \Mux26~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux26~1 (
	.dataa(\lpp_ram_data_out[0][5]~q ),
	.datab(\lpp_ram_data_out[3][5]~q ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.cin(gnd),
	.combout(\Mux26~1_combout ),
	.cout());
defparam \Mux26~1 .lut_mask = 16'hAACC;
defparam \Mux26~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux26~2 (
	.dataa(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.datab(\lpp_ram_data_out[2][5]~q ),
	.datac(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.datad(\lpp_ram_data_out[0][5]~q ),
	.cin(gnd),
	.combout(\Mux26~2_combout ),
	.cout());
defparam \Mux26~2 .lut_mask = 16'hFFDE;
defparam \Mux26~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux26~3 (
	.dataa(\lpp_ram_data_out[1][5]~q ),
	.datab(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.datac(\Mux26~2_combout ),
	.datad(\lpp_ram_data_out[3][5]~q ),
	.cin(gnd),
	.combout(\Mux26~3_combout ),
	.cout());
defparam \Mux26~3 .lut_mask = 16'hFFBE;
defparam \Mux26~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux27~0 (
	.dataa(\lpp_ram_data_out[2][4]~q ),
	.datab(\lpp_ram_data_out[1][4]~q ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.cin(gnd),
	.combout(\Mux27~0_combout ),
	.cout());
defparam \Mux27~0 .lut_mask = 16'hAACC;
defparam \Mux27~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux27~1 (
	.dataa(\lpp_ram_data_out[0][4]~q ),
	.datab(\lpp_ram_data_out[3][4]~q ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.cin(gnd),
	.combout(\Mux27~1_combout ),
	.cout());
defparam \Mux27~1 .lut_mask = 16'hAACC;
defparam \Mux27~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux27~2 (
	.dataa(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.datab(\lpp_ram_data_out[1][4]~q ),
	.datac(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.datad(\lpp_ram_data_out[0][4]~q ),
	.cin(gnd),
	.combout(\Mux27~2_combout ),
	.cout());
defparam \Mux27~2 .lut_mask = 16'hFFDE;
defparam \Mux27~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux27~3 (
	.dataa(\lpp_ram_data_out[2][4]~q ),
	.datab(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.datac(\Mux27~2_combout ),
	.datad(\lpp_ram_data_out[3][4]~q ),
	.cin(gnd),
	.combout(\Mux27~3_combout ),
	.cout());
defparam \Mux27~3 .lut_mask = 16'hFFBE;
defparam \Mux27~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux28~0 (
	.dataa(\lpp_ram_data_out[2][3]~q ),
	.datab(\lpp_ram_data_out[1][3]~q ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.cin(gnd),
	.combout(\Mux28~0_combout ),
	.cout());
defparam \Mux28~0 .lut_mask = 16'hAACC;
defparam \Mux28~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux28~1 (
	.dataa(\lpp_ram_data_out[0][3]~q ),
	.datab(\lpp_ram_data_out[3][3]~q ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.cin(gnd),
	.combout(\Mux28~1_combout ),
	.cout());
defparam \Mux28~1 .lut_mask = 16'hAACC;
defparam \Mux28~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux28~2 (
	.dataa(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.datab(\lpp_ram_data_out[2][3]~q ),
	.datac(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.datad(\lpp_ram_data_out[0][3]~q ),
	.cin(gnd),
	.combout(\Mux28~2_combout ),
	.cout());
defparam \Mux28~2 .lut_mask = 16'hFFDE;
defparam \Mux28~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux28~3 (
	.dataa(\lpp_ram_data_out[1][3]~q ),
	.datab(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.datac(\Mux28~2_combout ),
	.datad(\lpp_ram_data_out[3][3]~q ),
	.cin(gnd),
	.combout(\Mux28~3_combout ),
	.cout());
defparam \Mux28~3 .lut_mask = 16'hFFBE;
defparam \Mux28~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux29~0 (
	.dataa(\lpp_ram_data_out[2][2]~q ),
	.datab(\lpp_ram_data_out[1][2]~q ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.cin(gnd),
	.combout(\Mux29~0_combout ),
	.cout());
defparam \Mux29~0 .lut_mask = 16'hAACC;
defparam \Mux29~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux29~1 (
	.dataa(\lpp_ram_data_out[0][2]~q ),
	.datab(\lpp_ram_data_out[3][2]~q ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.cin(gnd),
	.combout(\Mux29~1_combout ),
	.cout());
defparam \Mux29~1 .lut_mask = 16'hAACC;
defparam \Mux29~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux29~2 (
	.dataa(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.datab(\lpp_ram_data_out[1][2]~q ),
	.datac(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.datad(\lpp_ram_data_out[0][2]~q ),
	.cin(gnd),
	.combout(\Mux29~2_combout ),
	.cout());
defparam \Mux29~2 .lut_mask = 16'hFFDE;
defparam \Mux29~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux29~3 (
	.dataa(\lpp_ram_data_out[2][2]~q ),
	.datab(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.datac(\Mux29~2_combout ),
	.datad(\lpp_ram_data_out[3][2]~q ),
	.cin(gnd),
	.combout(\Mux29~3_combout ),
	.cout());
defparam \Mux29~3 .lut_mask = 16'hFFBE;
defparam \Mux29~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux22~0 (
	.dataa(\lpp_ram_data_out[2][9]~q ),
	.datab(\lpp_ram_data_out[1][9]~q ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.cin(gnd),
	.combout(\Mux22~0_combout ),
	.cout());
defparam \Mux22~0 .lut_mask = 16'hAACC;
defparam \Mux22~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux22~1 (
	.dataa(\lpp_ram_data_out[0][9]~q ),
	.datab(\lpp_ram_data_out[3][9]~q ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.cin(gnd),
	.combout(\Mux22~1_combout ),
	.cout());
defparam \Mux22~1 .lut_mask = 16'hAACC;
defparam \Mux22~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux22~2 (
	.dataa(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.datab(\lpp_ram_data_out[2][9]~q ),
	.datac(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.datad(\lpp_ram_data_out[0][9]~q ),
	.cin(gnd),
	.combout(\Mux22~2_combout ),
	.cout());
defparam \Mux22~2 .lut_mask = 16'hFFDE;
defparam \Mux22~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux22~3 (
	.dataa(\lpp_ram_data_out[1][9]~q ),
	.datab(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.datac(\Mux22~2_combout ),
	.datad(\lpp_ram_data_out[3][9]~q ),
	.cin(gnd),
	.combout(\Mux22~3_combout ),
	.cout());
defparam \Mux22~3 .lut_mask = 16'hFFBE;
defparam \Mux22~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux23~0 (
	.dataa(\lpp_ram_data_out[2][8]~q ),
	.datab(\lpp_ram_data_out[1][8]~q ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.cin(gnd),
	.combout(\Mux23~0_combout ),
	.cout());
defparam \Mux23~0 .lut_mask = 16'hAACC;
defparam \Mux23~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux23~1 (
	.dataa(\lpp_ram_data_out[0][8]~q ),
	.datab(\lpp_ram_data_out[3][8]~q ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.cin(gnd),
	.combout(\Mux23~1_combout ),
	.cout());
defparam \Mux23~1 .lut_mask = 16'hAACC;
defparam \Mux23~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux23~2 (
	.dataa(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.datab(\lpp_ram_data_out[1][8]~q ),
	.datac(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.datad(\lpp_ram_data_out[0][8]~q ),
	.cin(gnd),
	.combout(\Mux23~2_combout ),
	.cout());
defparam \Mux23~2 .lut_mask = 16'hFFDE;
defparam \Mux23~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux23~3 (
	.dataa(\lpp_ram_data_out[2][8]~q ),
	.datab(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.datac(\Mux23~2_combout ),
	.datad(\lpp_ram_data_out[3][8]~q ),
	.cin(gnd),
	.combout(\Mux23~3_combout ),
	.cout());
defparam \Mux23~3 .lut_mask = 16'hFFBE;
defparam \Mux23~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux16~0 (
	.dataa(\lpp_ram_data_out[2][15]~q ),
	.datab(\lpp_ram_data_out[1][15]~q ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.cin(gnd),
	.combout(\Mux16~0_combout ),
	.cout());
defparam \Mux16~0 .lut_mask = 16'hAACC;
defparam \Mux16~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux16~1 (
	.dataa(\lpp_ram_data_out[0][15]~q ),
	.datab(\lpp_ram_data_out[3][15]~q ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.cin(gnd),
	.combout(\Mux16~1_combout ),
	.cout());
defparam \Mux16~1 .lut_mask = 16'hAACC;
defparam \Mux16~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux16~2 (
	.dataa(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.datab(\lpp_ram_data_out[2][15]~q ),
	.datac(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.datad(\lpp_ram_data_out[0][15]~q ),
	.cin(gnd),
	.combout(\Mux16~2_combout ),
	.cout());
defparam \Mux16~2 .lut_mask = 16'hFFDE;
defparam \Mux16~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux16~3 (
	.dataa(\lpp_ram_data_out[1][15]~q ),
	.datab(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.datac(\Mux16~2_combout ),
	.datad(\lpp_ram_data_out[3][15]~q ),
	.cin(gnd),
	.combout(\Mux16~3_combout ),
	.cout());
defparam \Mux16~3 .lut_mask = 16'hFFBE;
defparam \Mux16~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux17~0 (
	.dataa(\lpp_ram_data_out[2][14]~q ),
	.datab(\lpp_ram_data_out[1][14]~q ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.cin(gnd),
	.combout(\Mux17~0_combout ),
	.cout());
defparam \Mux17~0 .lut_mask = 16'hAACC;
defparam \Mux17~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux17~1 (
	.dataa(\lpp_ram_data_out[0][14]~q ),
	.datab(\lpp_ram_data_out[3][14]~q ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.cin(gnd),
	.combout(\Mux17~1_combout ),
	.cout());
defparam \Mux17~1 .lut_mask = 16'hAACC;
defparam \Mux17~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux17~2 (
	.dataa(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.datab(\lpp_ram_data_out[1][14]~q ),
	.datac(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.datad(\lpp_ram_data_out[0][14]~q ),
	.cin(gnd),
	.combout(\Mux17~2_combout ),
	.cout());
defparam \Mux17~2 .lut_mask = 16'hFFDE;
defparam \Mux17~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux17~3 (
	.dataa(\lpp_ram_data_out[2][14]~q ),
	.datab(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.datac(\Mux17~2_combout ),
	.datad(\lpp_ram_data_out[3][14]~q ),
	.cin(gnd),
	.combout(\Mux17~3_combout ),
	.cout());
defparam \Mux17~3 .lut_mask = 16'hFFBE;
defparam \Mux17~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux18~0 (
	.dataa(\lpp_ram_data_out[2][13]~q ),
	.datab(\lpp_ram_data_out[1][13]~q ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.cin(gnd),
	.combout(\Mux18~0_combout ),
	.cout());
defparam \Mux18~0 .lut_mask = 16'hAACC;
defparam \Mux18~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux18~1 (
	.dataa(\lpp_ram_data_out[0][13]~q ),
	.datab(\lpp_ram_data_out[3][13]~q ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.cin(gnd),
	.combout(\Mux18~1_combout ),
	.cout());
defparam \Mux18~1 .lut_mask = 16'hAACC;
defparam \Mux18~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux18~2 (
	.dataa(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.datab(\lpp_ram_data_out[2][13]~q ),
	.datac(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.datad(\lpp_ram_data_out[0][13]~q ),
	.cin(gnd),
	.combout(\Mux18~2_combout ),
	.cout());
defparam \Mux18~2 .lut_mask = 16'hFFDE;
defparam \Mux18~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux18~3 (
	.dataa(\lpp_ram_data_out[1][13]~q ),
	.datab(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.datac(\Mux18~2_combout ),
	.datad(\lpp_ram_data_out[3][13]~q ),
	.cin(gnd),
	.combout(\Mux18~3_combout ),
	.cout());
defparam \Mux18~3 .lut_mask = 16'hFFBE;
defparam \Mux18~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux19~0 (
	.dataa(\lpp_ram_data_out[2][12]~q ),
	.datab(\lpp_ram_data_out[1][12]~q ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.cin(gnd),
	.combout(\Mux19~0_combout ),
	.cout());
defparam \Mux19~0 .lut_mask = 16'hAACC;
defparam \Mux19~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux19~1 (
	.dataa(\lpp_ram_data_out[0][12]~q ),
	.datab(\lpp_ram_data_out[3][12]~q ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.cin(gnd),
	.combout(\Mux19~1_combout ),
	.cout());
defparam \Mux19~1 .lut_mask = 16'hAACC;
defparam \Mux19~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux19~2 (
	.dataa(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.datab(\lpp_ram_data_out[1][12]~q ),
	.datac(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.datad(\lpp_ram_data_out[0][12]~q ),
	.cin(gnd),
	.combout(\Mux19~2_combout ),
	.cout());
defparam \Mux19~2 .lut_mask = 16'hFFDE;
defparam \Mux19~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux19~3 (
	.dataa(\lpp_ram_data_out[2][12]~q ),
	.datab(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.datac(\Mux19~2_combout ),
	.datad(\lpp_ram_data_out[3][12]~q ),
	.cin(gnd),
	.combout(\Mux19~3_combout ),
	.cout());
defparam \Mux19~3 .lut_mask = 16'hFFBE;
defparam \Mux19~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux20~0 (
	.dataa(\lpp_ram_data_out[2][11]~q ),
	.datab(\lpp_ram_data_out[1][11]~q ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.cin(gnd),
	.combout(\Mux20~0_combout ),
	.cout());
defparam \Mux20~0 .lut_mask = 16'hAACC;
defparam \Mux20~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux20~1 (
	.dataa(\lpp_ram_data_out[0][11]~q ),
	.datab(\lpp_ram_data_out[3][11]~q ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.cin(gnd),
	.combout(\Mux20~1_combout ),
	.cout());
defparam \Mux20~1 .lut_mask = 16'hAACC;
defparam \Mux20~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux20~2 (
	.dataa(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.datab(\lpp_ram_data_out[2][11]~q ),
	.datac(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.datad(\lpp_ram_data_out[0][11]~q ),
	.cin(gnd),
	.combout(\Mux20~2_combout ),
	.cout());
defparam \Mux20~2 .lut_mask = 16'hFFDE;
defparam \Mux20~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux20~3 (
	.dataa(\lpp_ram_data_out[1][11]~q ),
	.datab(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.datac(\Mux20~2_combout ),
	.datad(\lpp_ram_data_out[3][11]~q ),
	.cin(gnd),
	.combout(\Mux20~3_combout ),
	.cout());
defparam \Mux20~3 .lut_mask = 16'hFFBE;
defparam \Mux20~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux21~0 (
	.dataa(\lpp_ram_data_out[2][10]~q ),
	.datab(\lpp_ram_data_out[1][10]~q ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.cin(gnd),
	.combout(\Mux21~0_combout ),
	.cout());
defparam \Mux21~0 .lut_mask = 16'hAACC;
defparam \Mux21~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux21~1 (
	.dataa(\lpp_ram_data_out[0][10]~q ),
	.datab(\lpp_ram_data_out[3][10]~q ),
	.datac(gnd),
	.datad(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.cin(gnd),
	.combout(\Mux21~1_combout ),
	.cout());
defparam \Mux21~1 .lut_mask = 16'hAACC;
defparam \Mux21~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux21~2 (
	.dataa(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.datab(\lpp_ram_data_out[1][10]~q ),
	.datac(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.datad(\lpp_ram_data_out[0][10]~q ),
	.cin(gnd),
	.combout(\Mux21~2_combout ),
	.cout());
defparam \Mux21~2 .lut_mask = 16'hFFDE;
defparam \Mux21~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux21~3 (
	.dataa(\lpp_ram_data_out[2][10]~q ),
	.datab(\gen_radix_2_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.datac(\Mux21~2_combout ),
	.datad(\lpp_ram_data_out[3][10]~q ),
	.cin(gnd),
	.combout(\Mux21~3_combout ),
	.cout());
defparam \Mux21~3 .lut_mask = 16'hFFBE;
defparam \Mux21~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \fft_dirn_held~0 (
	.dataa(reset_n),
	.datab(\fft_dirn~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fft_dirn_held~0_combout ),
	.cout());
defparam \fft_dirn_held~0 .lut_mask = 16'hEEEE;
defparam \fft_dirn_held~0 .sum_lutc_input = "datac";

dffeas \data_rdy_vec[4] (
	.clk(clk),
	.d(\data_rdy_vec~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_rdy_vec[4]~q ),
	.prn(vcc));
defparam \data_rdy_vec[4] .is_wysiwyg = "true";
defparam \data_rdy_vec[4] .power_up = "low";

cycloneiii_lcell_comb \lpp_ram_data_out~0 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[1] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[1] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~0_combout ),
	.cout());
defparam \lpp_ram_data_out~0 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~1 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[1] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[1] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~1_combout ),
	.cout());
defparam \lpp_ram_data_out~1 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~2 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[1] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[1] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~2_combout ),
	.cout());
defparam \lpp_ram_data_out~2 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~3 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[1] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[1] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~3_combout ),
	.cout());
defparam \lpp_ram_data_out~3 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~4 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[0] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[0] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~4_combout ),
	.cout());
defparam \lpp_ram_data_out~4 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~5 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[0] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[0] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~5_combout ),
	.cout());
defparam \lpp_ram_data_out~5 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~6 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[0] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[0] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~6_combout ),
	.cout());
defparam \lpp_ram_data_out~6 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~7 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[0] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[0] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~7_combout ),
	.cout());
defparam \lpp_ram_data_out~7 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~8 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[7] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[7] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~8_combout ),
	.cout());
defparam \lpp_ram_data_out~8 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~8 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~9 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[7] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[7] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~9_combout ),
	.cout());
defparam \lpp_ram_data_out~9 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~10 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[7] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[7] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~10_combout ),
	.cout());
defparam \lpp_ram_data_out~10 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~10 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~11 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[7] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[7] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~11_combout ),
	.cout());
defparam \lpp_ram_data_out~11 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~11 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~12 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[6] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[6] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~12_combout ),
	.cout());
defparam \lpp_ram_data_out~12 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~12 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~13 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[6] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[6] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~13_combout ),
	.cout());
defparam \lpp_ram_data_out~13 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~13 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~14 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[6] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[6] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~14_combout ),
	.cout());
defparam \lpp_ram_data_out~14 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~14 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~15 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[6] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[6] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~15_combout ),
	.cout());
defparam \lpp_ram_data_out~15 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~15 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~16 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[5] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[5] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~16_combout ),
	.cout());
defparam \lpp_ram_data_out~16 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~16 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~17 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[5] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[5] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~17_combout ),
	.cout());
defparam \lpp_ram_data_out~17 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~17 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~18 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[5] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[5] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~18_combout ),
	.cout());
defparam \lpp_ram_data_out~18 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~18 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~19 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[5] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[5] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~19_combout ),
	.cout());
defparam \lpp_ram_data_out~19 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~19 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~20 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[4] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[4] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~20_combout ),
	.cout());
defparam \lpp_ram_data_out~20 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~20 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~21 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[4] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[4] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~21_combout ),
	.cout());
defparam \lpp_ram_data_out~21 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~21 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~22 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[4] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[4] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~22_combout ),
	.cout());
defparam \lpp_ram_data_out~22 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~22 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~23 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[4] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[4] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~23_combout ),
	.cout());
defparam \lpp_ram_data_out~23 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~23 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~24 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[3] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[3] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~24_combout ),
	.cout());
defparam \lpp_ram_data_out~24 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~24 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~25 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[3] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[3] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~25_combout ),
	.cout());
defparam \lpp_ram_data_out~25 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~25 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~26 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[3] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[3] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~26_combout ),
	.cout());
defparam \lpp_ram_data_out~26 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~26 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~27 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[3] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[3] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~27_combout ),
	.cout());
defparam \lpp_ram_data_out~27 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~27 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~28 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[2] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[2] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~28_combout ),
	.cout());
defparam \lpp_ram_data_out~28 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~28 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~29 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[2] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[2] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~29_combout ),
	.cout());
defparam \lpp_ram_data_out~29 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~29 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~30 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[2] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[2] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~30_combout ),
	.cout());
defparam \lpp_ram_data_out~30 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~30 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~31 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[2] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[2] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~31_combout ),
	.cout());
defparam \lpp_ram_data_out~31 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~31 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~32 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[9] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[9] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~32_combout ),
	.cout());
defparam \lpp_ram_data_out~32 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~32 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~33 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[9] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[9] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~33_combout ),
	.cout());
defparam \lpp_ram_data_out~33 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~33 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~34 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[9] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[9] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~34_combout ),
	.cout());
defparam \lpp_ram_data_out~34 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~34 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~35 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[9] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[9] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~35_combout ),
	.cout());
defparam \lpp_ram_data_out~35 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~35 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~36 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[8] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[8] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~36_combout ),
	.cout());
defparam \lpp_ram_data_out~36 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~36 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~37 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[8] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[8] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~37_combout ),
	.cout());
defparam \lpp_ram_data_out~37 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~37 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~38 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[8] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[8] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~38_combout ),
	.cout());
defparam \lpp_ram_data_out~38 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~38 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~39 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[8] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[8] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~39_combout ),
	.cout());
defparam \lpp_ram_data_out~39 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~39 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~40 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[15] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[15] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~40_combout ),
	.cout());
defparam \lpp_ram_data_out~40 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~40 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~41 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[15] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[15] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~41_combout ),
	.cout());
defparam \lpp_ram_data_out~41 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~41 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~42 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[15] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[15] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~42_combout ),
	.cout());
defparam \lpp_ram_data_out~42 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~42 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~43 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[15] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[15] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~43_combout ),
	.cout());
defparam \lpp_ram_data_out~43 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~43 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~44 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[14] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[14] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~44_combout ),
	.cout());
defparam \lpp_ram_data_out~44 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~44 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~45 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[14] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[14] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~45_combout ),
	.cout());
defparam \lpp_ram_data_out~45 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~45 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~46 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[14] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[14] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~46_combout ),
	.cout());
defparam \lpp_ram_data_out~46 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~46 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~47 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[14] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[14] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~47_combout ),
	.cout());
defparam \lpp_ram_data_out~47 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~47 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~48 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[13] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[13] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~48_combout ),
	.cout());
defparam \lpp_ram_data_out~48 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~48 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~49 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[13] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[13] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~49_combout ),
	.cout());
defparam \lpp_ram_data_out~49 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~49 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~50 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[13] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[13] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~50_combout ),
	.cout());
defparam \lpp_ram_data_out~50 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~50 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~51 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[13] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[13] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~51_combout ),
	.cout());
defparam \lpp_ram_data_out~51 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~51 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~52 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[12] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[12] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~52_combout ),
	.cout());
defparam \lpp_ram_data_out~52 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~52 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~53 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[12] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[12] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~53_combout ),
	.cout());
defparam \lpp_ram_data_out~53 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~53 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~54 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[12] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[12] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~54_combout ),
	.cout());
defparam \lpp_ram_data_out~54 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~54 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~55 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[12] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[12] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~55_combout ),
	.cout());
defparam \lpp_ram_data_out~55 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~55 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~56 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[11] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[11] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~56_combout ),
	.cout());
defparam \lpp_ram_data_out~56 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~56 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~57 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[11] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[11] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~57_combout ),
	.cout());
defparam \lpp_ram_data_out~57 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~57 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~58 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[11] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[11] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~58_combout ),
	.cout());
defparam \lpp_ram_data_out~58 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~58 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~59 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[11] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[11] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~59_combout ),
	.cout());
defparam \lpp_ram_data_out~59 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~59 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~60 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[10] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[10] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~60_combout ),
	.cout());
defparam \lpp_ram_data_out~60 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~60 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~61 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[10] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[10] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~61_combout ),
	.cout());
defparam \lpp_ram_data_out~61 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~61 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~62 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[10] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[10] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~62_combout ),
	.cout());
defparam \lpp_ram_data_out~62 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~62 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lpp_ram_data_out~63 (
	.dataa(\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[10] ),
	.datab(\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[10] ),
	.datac(gnd),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~63_combout ),
	.cout());
defparam \lpp_ram_data_out~63 .lut_mask = 16'hAACC;
defparam \lpp_ram_data_out~63 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \fft_dirn~0 (
	.dataa(inverse),
	.datab(\fft_dirn~q ),
	.datac(gnd),
	.datad(\auk_dsp_atlantic_sink_1|send_sop_s~q ),
	.cin(gnd),
	.combout(\fft_dirn~0_combout ),
	.cout());
defparam \fft_dirn~0 .lut_mask = 16'hAACC;
defparam \fft_dirn~0 .sum_lutc_input = "datac";

dffeas \data_rdy_vec[3] (
	.clk(clk),
	.d(\data_rdy_vec~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_rdy_vec[3]~q ),
	.prn(vcc));
defparam \data_rdy_vec[3] .is_wysiwyg = "true";
defparam \data_rdy_vec[3] .power_up = "low";

cycloneiii_lcell_comb \data_rdy_vec~0 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~0_combout ),
	.cout());
defparam \data_rdy_vec~0 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~0 .sum_lutc_input = "datac";

dffeas \wc_vec[6] (
	.clk(clk),
	.d(\wc_vec~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\wc_vec[6]~q ),
	.prn(vcc));
defparam \wc_vec[6] .is_wysiwyg = "true";
defparam \wc_vec[6] .power_up = "low";

dffeas \rdaddress_c_bus[0] (
	.clk(clk),
	.d(\rdaddress_c_bus~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\rdaddress_c_bus[0]~q ),
	.prn(vcc));
defparam \rdaddress_c_bus[0] .is_wysiwyg = "true";
defparam \rdaddress_c_bus[0] .power_up = "low";

dffeas \rdaddress_c_bus[15] (
	.clk(clk),
	.d(\rdaddress_c_bus~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\rdaddress_c_bus[15]~q ),
	.prn(vcc));
defparam \rdaddress_c_bus[15] .is_wysiwyg = "true";
defparam \rdaddress_c_bus[15] .power_up = "low";

dffeas \rdaddress_c_bus[16] (
	.clk(clk),
	.d(\rdaddress_c_bus~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\rdaddress_c_bus[16]~q ),
	.prn(vcc));
defparam \rdaddress_c_bus[16] .is_wysiwyg = "true";
defparam \rdaddress_c_bus[16] .power_up = "low";

dffeas \rdaddress_c_bus[10] (
	.clk(clk),
	.d(\rdaddress_c_bus~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\rdaddress_c_bus[10]~q ),
	.prn(vcc));
defparam \rdaddress_c_bus[10] .is_wysiwyg = "true";
defparam \rdaddress_c_bus[10] .power_up = "low";

dffeas \rdaddress_c_bus[11] (
	.clk(clk),
	.d(\rdaddress_c_bus~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\rdaddress_c_bus[11]~q ),
	.prn(vcc));
defparam \rdaddress_c_bus[11] .is_wysiwyg = "true";
defparam \rdaddress_c_bus[11] .power_up = "low";

dffeas \rdaddress_c_bus[12] (
	.clk(clk),
	.d(\rdaddress_c_bus~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\rdaddress_c_bus[12]~q ),
	.prn(vcc));
defparam \rdaddress_c_bus[12] .is_wysiwyg = "true";
defparam \rdaddress_c_bus[12] .power_up = "low";

dffeas \rdaddress_c_bus[13] (
	.clk(clk),
	.d(\rdaddress_c_bus~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\rdaddress_c_bus[13]~q ),
	.prn(vcc));
defparam \rdaddress_c_bus[13] .is_wysiwyg = "true";
defparam \rdaddress_c_bus[13] .power_up = "low";

dffeas \wd_vec[6] (
	.clk(clk),
	.d(\wd_vec~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\wd_vec[6]~q ),
	.prn(vcc));
defparam \wd_vec[6] .is_wysiwyg = "true";
defparam \wd_vec[6] .power_up = "low";

cycloneiii_lcell_comb \lpp_sel~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\gen_radix_2_last_pass:gen_lpp_addr|delay_en|tdl_arr[4]~q ),
	.datad(\lpp_sel~q ),
	.cin(gnd),
	.combout(\lpp_sel~0_combout ),
	.cout());
defparam \lpp_sel~0 .lut_mask = 16'h0FF0;
defparam \lpp_sel~0 .sum_lutc_input = "datac";

dffeas \rdaddress_c_bus[20] (
	.clk(clk),
	.d(\rdaddress_c_bus~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\rdaddress_c_bus[20]~q ),
	.prn(vcc));
defparam \rdaddress_c_bus[20] .is_wysiwyg = "true";
defparam \rdaddress_c_bus[20] .power_up = "low";

dffeas \data_rdy_vec[2] (
	.clk(clk),
	.d(\data_rdy_vec~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_rdy_vec[2]~q ),
	.prn(vcc));
defparam \data_rdy_vec[2] .is_wysiwyg = "true";
defparam \data_rdy_vec[2] .power_up = "low";

cycloneiii_lcell_comb \data_rdy_vec~1 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~1_combout ),
	.cout());
defparam \data_rdy_vec~1 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~1 .sum_lutc_input = "datac";

dffeas \wc_vec[5] (
	.clk(clk),
	.d(\wc_vec~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\wc_vec[5]~q ),
	.prn(vcc));
defparam \wc_vec[5] .is_wysiwyg = "true";
defparam \wc_vec[5] .power_up = "low";

cycloneiii_lcell_comb \wc_vec~0 (
	.dataa(reset_n),
	.datab(\wc_vec[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wc_vec~0_combout ),
	.cout());
defparam \wc_vec~0 .lut_mask = 16'hEEEE;
defparam \wc_vec~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rdaddress_c_bus~0 (
	.dataa(reset_n),
	.datab(\gen_radix_2_last_pass:ram_cxb_rd_lpp|ram_in_reg[0][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\rdaddress_c_bus~0_combout ),
	.cout());
defparam \rdaddress_c_bus~0 .lut_mask = 16'hEEEE;
defparam \rdaddress_c_bus~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rdaddress_c_bus~1 (
	.dataa(reset_n),
	.datab(\gen_radix_2_last_pass:ram_cxb_rd_lpp|ram_in_reg[0][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\rdaddress_c_bus~1_combout ),
	.cout());
defparam \rdaddress_c_bus~1 .lut_mask = 16'hEEEE;
defparam \rdaddress_c_bus~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rdaddress_c_bus~2 (
	.dataa(reset_n),
	.datab(\gen_radix_2_last_pass:ram_cxb_rd_lpp|ram_in_reg[0][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\rdaddress_c_bus~2_combout ),
	.cout());
defparam \rdaddress_c_bus~2 .lut_mask = 16'hEEEE;
defparam \rdaddress_c_bus~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rdaddress_c_bus~3 (
	.dataa(reset_n),
	.datab(\gen_radix_2_last_pass:ram_cxb_rd_lpp|ram_in_reg[0][3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\rdaddress_c_bus~3_combout ),
	.cout());
defparam \rdaddress_c_bus~3 .lut_mask = 16'hEEEE;
defparam \rdaddress_c_bus~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rdaddress_c_bus~4 (
	.dataa(reset_n),
	.datab(\gen_radix_2_last_pass:ram_cxb_rd_lpp|ram_in_reg[0][4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\rdaddress_c_bus~4_combout ),
	.cout());
defparam \rdaddress_c_bus~4 .lut_mask = 16'hEEEE;
defparam \rdaddress_c_bus~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rdaddress_c_bus~5 (
	.dataa(reset_n),
	.datab(\gen_radix_2_last_pass:ram_cxb_rd_lpp|ram_in_reg[0][5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\rdaddress_c_bus~5_combout ),
	.cout());
defparam \rdaddress_c_bus~5 .lut_mask = 16'hEEEE;
defparam \rdaddress_c_bus~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rdaddress_c_bus~6 (
	.dataa(\gen_radix_2_last_pass:ram_cxb_rd_lpp|ram_in_reg[1][6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\rdaddress_c_bus~6_combout ),
	.cout());
defparam \rdaddress_c_bus~6 .lut_mask = 16'hFF55;
defparam \rdaddress_c_bus~6 .sum_lutc_input = "datac";

dffeas \wd_vec[5] (
	.clk(clk),
	.d(\wd_vec~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\wd_vec[5]~q ),
	.prn(vcc));
defparam \wd_vec[5] .is_wysiwyg = "true";
defparam \wd_vec[5] .power_up = "low";

cycloneiii_lcell_comb \wd_vec~0 (
	.dataa(reset_n),
	.datab(\wd_vec[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wd_vec~0_combout ),
	.cout());
defparam \wd_vec~0 .lut_mask = 16'hEEEE;
defparam \wd_vec~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rdaddress_c_bus~7 (
	.dataa(reset_n),
	.datab(\gen_radix_2_last_pass:ram_cxb_rd_lpp|ram_in_reg[1][6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\rdaddress_c_bus~7_combout ),
	.cout());
defparam \rdaddress_c_bus~7 .lut_mask = 16'hEEEE;
defparam \rdaddress_c_bus~7 .sum_lutc_input = "datac";

dffeas \data_rdy_vec[1] (
	.clk(clk),
	.d(\data_rdy_vec~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_rdy_vec[1]~q ),
	.prn(vcc));
defparam \data_rdy_vec[1] .is_wysiwyg = "true";
defparam \data_rdy_vec[1] .power_up = "low";

cycloneiii_lcell_comb \data_rdy_vec~2 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~2_combout ),
	.cout());
defparam \data_rdy_vec~2 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~2 .sum_lutc_input = "datac";

dffeas \wc_vec[4] (
	.clk(clk),
	.d(\wc_vec~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\wc_vec[4]~q ),
	.prn(vcc));
defparam \wc_vec[4] .is_wysiwyg = "true";
defparam \wc_vec[4] .power_up = "low";

cycloneiii_lcell_comb \wc_vec~1 (
	.dataa(reset_n),
	.datab(\wc_vec[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wc_vec~1_combout ),
	.cout());
defparam \wc_vec~1 .lut_mask = 16'hEEEE;
defparam \wc_vec~1 .sum_lutc_input = "datac";

dffeas \wd_vec[4] (
	.clk(clk),
	.d(\wd_vec~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\wd_vec[4]~q ),
	.prn(vcc));
defparam \wd_vec[4] .is_wysiwyg = "true";
defparam \wd_vec[4] .power_up = "low";

cycloneiii_lcell_comb \wd_vec~1 (
	.dataa(reset_n),
	.datab(\wd_vec[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wd_vec~1_combout ),
	.cout());
defparam \wd_vec~1 .lut_mask = 16'hEEEE;
defparam \wd_vec~1 .sum_lutc_input = "datac";

dffeas \data_rdy_vec[0] (
	.clk(clk),
	.d(\data_rdy_vec~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_rdy_vec[0]~q ),
	.prn(vcc));
defparam \data_rdy_vec[0] .is_wysiwyg = "true";
defparam \data_rdy_vec[0] .power_up = "low";

cycloneiii_lcell_comb \data_rdy_vec~3 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~3_combout ),
	.cout());
defparam \data_rdy_vec~3 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~3 .sum_lutc_input = "datac";

dffeas \wc_vec[3] (
	.clk(clk),
	.d(\wc_vec~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\wc_vec[3]~q ),
	.prn(vcc));
defparam \wc_vec[3] .is_wysiwyg = "true";
defparam \wc_vec[3] .power_up = "low";

cycloneiii_lcell_comb \wc_vec~2 (
	.dataa(reset_n),
	.datab(\wc_vec[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wc_vec~2_combout ),
	.cout());
defparam \wc_vec~2 .lut_mask = 16'hEEEE;
defparam \wc_vec~2 .sum_lutc_input = "datac";

dffeas \wd_vec[3] (
	.clk(clk),
	.d(\wd_vec~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\wd_vec[3]~q ),
	.prn(vcc));
defparam \wd_vec[3] .is_wysiwyg = "true";
defparam \wd_vec[3] .power_up = "low";

cycloneiii_lcell_comb \wd_vec~2 (
	.dataa(reset_n),
	.datab(\wd_vec[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wd_vec~2_combout ),
	.cout());
defparam \wd_vec~2 .lut_mask = 16'hEEEE;
defparam \wd_vec~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \data_rdy_vec~4 (
	.dataa(reset_n),
	.datab(\writer|data_rdy_int~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~4_combout ),
	.cout());
defparam \data_rdy_vec~4 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~4 .sum_lutc_input = "datac";

dffeas \wc_vec[2] (
	.clk(clk),
	.d(\wc_vec~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\wc_vec[2]~q ),
	.prn(vcc));
defparam \wc_vec[2] .is_wysiwyg = "true";
defparam \wc_vec[2] .power_up = "low";

cycloneiii_lcell_comb \wc_vec~3 (
	.dataa(reset_n),
	.datab(\wc_vec[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wc_vec~3_combout ),
	.cout());
defparam \wc_vec~3 .lut_mask = 16'hEEEE;
defparam \wc_vec~3 .sum_lutc_input = "datac";

dffeas \wd_vec[2] (
	.clk(clk),
	.d(\wd_vec~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\wd_vec[2]~q ),
	.prn(vcc));
defparam \wd_vec[2] .is_wysiwyg = "true";
defparam \wd_vec[2] .power_up = "low";

cycloneiii_lcell_comb \wd_vec~3 (
	.dataa(reset_n),
	.datab(\wd_vec[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wd_vec~3_combout ),
	.cout());
defparam \wd_vec~3 .lut_mask = 16'hEEEE;
defparam \wd_vec~3 .sum_lutc_input = "datac";

dffeas \wc_vec[1] (
	.clk(clk),
	.d(\wc_vec~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\wc_vec[1]~q ),
	.prn(vcc));
defparam \wc_vec[1] .is_wysiwyg = "true";
defparam \wc_vec[1] .power_up = "low";

cycloneiii_lcell_comb \wc_vec~4 (
	.dataa(reset_n),
	.datab(\wc_vec[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wc_vec~4_combout ),
	.cout());
defparam \wc_vec~4 .lut_mask = 16'hEEEE;
defparam \wc_vec~4 .sum_lutc_input = "datac";

dffeas \p_tdl[18][0] (
	.clk(clk),
	.d(\p_tdl[17][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[18][0]~q ),
	.prn(vcc));
defparam \p_tdl[18][0] .is_wysiwyg = "true";
defparam \p_tdl[18][0] .power_up = "low";

dffeas \p_tdl[18][2] (
	.clk(clk),
	.d(\p_tdl[17][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[18][2]~q ),
	.prn(vcc));
defparam \p_tdl[18][2] .is_wysiwyg = "true";
defparam \p_tdl[18][2] .power_up = "low";

dffeas \p_tdl[18][1] (
	.clk(clk),
	.d(\p_tdl[17][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[18][1]~q ),
	.prn(vcc));
defparam \p_tdl[18][1] .is_wysiwyg = "true";
defparam \p_tdl[18][1] .power_up = "low";

dffeas \wd_vec[1] (
	.clk(clk),
	.d(\wd_vec~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\wd_vec[1]~q ),
	.prn(vcc));
defparam \wd_vec[1] .is_wysiwyg = "true";
defparam \wd_vec[1] .power_up = "low";

cycloneiii_lcell_comb \wd_vec~4 (
	.dataa(reset_n),
	.datab(\wd_vec[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wd_vec~4_combout ),
	.cout());
defparam \wd_vec~4 .lut_mask = 16'hEEEE;
defparam \wd_vec~4 .sum_lutc_input = "datac";

dffeas \wc_vec[0] (
	.clk(clk),
	.d(\wc_vec~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\wc_vec[0]~q ),
	.prn(vcc));
defparam \wc_vec[0] .is_wysiwyg = "true";
defparam \wc_vec[0] .power_up = "low";

cycloneiii_lcell_comb \wc_vec~5 (
	.dataa(reset_n),
	.datab(\wc_vec[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wc_vec~5_combout ),
	.cout());
defparam \wc_vec~5 .lut_mask = 16'hEEEE;
defparam \wc_vec~5 .sum_lutc_input = "datac";

dffeas \p_tdl[17][0] (
	.clk(clk),
	.d(\p_tdl[16][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[17][0]~q ),
	.prn(vcc));
defparam \p_tdl[17][0] .is_wysiwyg = "true";
defparam \p_tdl[17][0] .power_up = "low";

dffeas \p_tdl[17][2] (
	.clk(clk),
	.d(\p_tdl[16][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[17][2]~q ),
	.prn(vcc));
defparam \p_tdl[17][2] .is_wysiwyg = "true";
defparam \p_tdl[17][2] .power_up = "low";

dffeas \p_tdl[17][1] (
	.clk(clk),
	.d(\p_tdl[16][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[17][1]~q ),
	.prn(vcc));
defparam \p_tdl[17][1] .is_wysiwyg = "true";
defparam \p_tdl[17][1] .power_up = "low";

dffeas \wd_vec[0] (
	.clk(clk),
	.d(\wd_vec~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\wd_vec[0]~q ),
	.prn(vcc));
defparam \wd_vec[0] .is_wysiwyg = "true";
defparam \wd_vec[0] .power_up = "low";

cycloneiii_lcell_comb \wd_vec~5 (
	.dataa(reset_n),
	.datab(\wd_vec[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wd_vec~5_combout ),
	.cout());
defparam \wd_vec~5 .lut_mask = 16'hEEEE;
defparam \wd_vec~5 .sum_lutc_input = "datac";

dffeas \twiddle_data[0][0][0] (
	.clk(clk),
	.d(\twiddle_data~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data[0][0][0]~q ),
	.prn(vcc));
defparam \twiddle_data[0][0][0] .is_wysiwyg = "true";
defparam \twiddle_data[0][0][0] .power_up = "low";

dffeas \twiddle_data[0][0][1] (
	.clk(clk),
	.d(\twiddle_data~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data[0][0][1]~q ),
	.prn(vcc));
defparam \twiddle_data[0][0][1] .is_wysiwyg = "true";
defparam \twiddle_data[0][0][1] .power_up = "low";

dffeas \twiddle_data[0][0][2] (
	.clk(clk),
	.d(\twiddle_data~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data[0][0][2]~q ),
	.prn(vcc));
defparam \twiddle_data[0][0][2] .is_wysiwyg = "true";
defparam \twiddle_data[0][0][2] .power_up = "low";

dffeas \twiddle_data[0][0][3] (
	.clk(clk),
	.d(\twiddle_data~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data[0][0][3]~q ),
	.prn(vcc));
defparam \twiddle_data[0][0][3] .is_wysiwyg = "true";
defparam \twiddle_data[0][0][3] .power_up = "low";

dffeas \twiddle_data[0][0][4] (
	.clk(clk),
	.d(\twiddle_data~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data[0][0][4]~q ),
	.prn(vcc));
defparam \twiddle_data[0][0][4] .is_wysiwyg = "true";
defparam \twiddle_data[0][0][4] .power_up = "low";

dffeas \twiddle_data[0][0][5] (
	.clk(clk),
	.d(\twiddle_data~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data[0][0][5]~q ),
	.prn(vcc));
defparam \twiddle_data[0][0][5] .is_wysiwyg = "true";
defparam \twiddle_data[0][0][5] .power_up = "low";

dffeas \twiddle_data[0][0][6] (
	.clk(clk),
	.d(\twiddle_data~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data[0][0][6]~q ),
	.prn(vcc));
defparam \twiddle_data[0][0][6] .is_wysiwyg = "true";
defparam \twiddle_data[0][0][6] .power_up = "low";

dffeas \twiddle_data[0][0][7] (
	.clk(clk),
	.d(\twiddle_data~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data[0][0][7]~q ),
	.prn(vcc));
defparam \twiddle_data[0][0][7] .is_wysiwyg = "true";
defparam \twiddle_data[0][0][7] .power_up = "low";

dffeas \twiddle_data[0][1][0] (
	.clk(clk),
	.d(\twiddle_data~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data[0][1][0]~q ),
	.prn(vcc));
defparam \twiddle_data[0][1][0] .is_wysiwyg = "true";
defparam \twiddle_data[0][1][0] .power_up = "low";

dffeas \twiddle_data[0][1][1] (
	.clk(clk),
	.d(\twiddle_data~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data[0][1][1]~q ),
	.prn(vcc));
defparam \twiddle_data[0][1][1] .is_wysiwyg = "true";
defparam \twiddle_data[0][1][1] .power_up = "low";

dffeas \twiddle_data[0][1][2] (
	.clk(clk),
	.d(\twiddle_data~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data[0][1][2]~q ),
	.prn(vcc));
defparam \twiddle_data[0][1][2] .is_wysiwyg = "true";
defparam \twiddle_data[0][1][2] .power_up = "low";

dffeas \twiddle_data[0][1][3] (
	.clk(clk),
	.d(\twiddle_data~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data[0][1][3]~q ),
	.prn(vcc));
defparam \twiddle_data[0][1][3] .is_wysiwyg = "true";
defparam \twiddle_data[0][1][3] .power_up = "low";

dffeas \twiddle_data[0][1][4] (
	.clk(clk),
	.d(\twiddle_data~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data[0][1][4]~q ),
	.prn(vcc));
defparam \twiddle_data[0][1][4] .is_wysiwyg = "true";
defparam \twiddle_data[0][1][4] .power_up = "low";

dffeas \twiddle_data[0][1][5] (
	.clk(clk),
	.d(\twiddle_data~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data[0][1][5]~q ),
	.prn(vcc));
defparam \twiddle_data[0][1][5] .is_wysiwyg = "true";
defparam \twiddle_data[0][1][5] .power_up = "low";

dffeas \twiddle_data[0][1][6] (
	.clk(clk),
	.d(\twiddle_data~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data[0][1][6]~q ),
	.prn(vcc));
defparam \twiddle_data[0][1][6] .is_wysiwyg = "true";
defparam \twiddle_data[0][1][6] .power_up = "low";

dffeas \twiddle_data[0][1][7] (
	.clk(clk),
	.d(\twiddle_data~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data[0][1][7]~q ),
	.prn(vcc));
defparam \twiddle_data[0][1][7] .is_wysiwyg = "true";
defparam \twiddle_data[0][1][7] .power_up = "low";

dffeas \twiddle_data[1][0][0] (
	.clk(clk),
	.d(\twiddle_data~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data[1][0][0]~q ),
	.prn(vcc));
defparam \twiddle_data[1][0][0] .is_wysiwyg = "true";
defparam \twiddle_data[1][0][0] .power_up = "low";

dffeas \twiddle_data[1][0][1] (
	.clk(clk),
	.d(\twiddle_data~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data[1][0][1]~q ),
	.prn(vcc));
defparam \twiddle_data[1][0][1] .is_wysiwyg = "true";
defparam \twiddle_data[1][0][1] .power_up = "low";

dffeas \twiddle_data[1][0][2] (
	.clk(clk),
	.d(\twiddle_data~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data[1][0][2]~q ),
	.prn(vcc));
defparam \twiddle_data[1][0][2] .is_wysiwyg = "true";
defparam \twiddle_data[1][0][2] .power_up = "low";

dffeas \twiddle_data[1][0][3] (
	.clk(clk),
	.d(\twiddle_data~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data[1][0][3]~q ),
	.prn(vcc));
defparam \twiddle_data[1][0][3] .is_wysiwyg = "true";
defparam \twiddle_data[1][0][3] .power_up = "low";

dffeas \twiddle_data[1][0][4] (
	.clk(clk),
	.d(\twiddle_data~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data[1][0][4]~q ),
	.prn(vcc));
defparam \twiddle_data[1][0][4] .is_wysiwyg = "true";
defparam \twiddle_data[1][0][4] .power_up = "low";

dffeas \twiddle_data[1][0][5] (
	.clk(clk),
	.d(\twiddle_data~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data[1][0][5]~q ),
	.prn(vcc));
defparam \twiddle_data[1][0][5] .is_wysiwyg = "true";
defparam \twiddle_data[1][0][5] .power_up = "low";

dffeas \twiddle_data[1][0][6] (
	.clk(clk),
	.d(\twiddle_data~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data[1][0][6]~q ),
	.prn(vcc));
defparam \twiddle_data[1][0][6] .is_wysiwyg = "true";
defparam \twiddle_data[1][0][6] .power_up = "low";

dffeas \twiddle_data[1][0][7] (
	.clk(clk),
	.d(\twiddle_data~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data[1][0][7]~q ),
	.prn(vcc));
defparam \twiddle_data[1][0][7] .is_wysiwyg = "true";
defparam \twiddle_data[1][0][7] .power_up = "low";

dffeas \twiddle_data[1][1][0] (
	.clk(clk),
	.d(\twiddle_data~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data[1][1][0]~q ),
	.prn(vcc));
defparam \twiddle_data[1][1][0] .is_wysiwyg = "true";
defparam \twiddle_data[1][1][0] .power_up = "low";

dffeas \twiddle_data[1][1][1] (
	.clk(clk),
	.d(\twiddle_data~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data[1][1][1]~q ),
	.prn(vcc));
defparam \twiddle_data[1][1][1] .is_wysiwyg = "true";
defparam \twiddle_data[1][1][1] .power_up = "low";

dffeas \twiddle_data[1][1][2] (
	.clk(clk),
	.d(\twiddle_data~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data[1][1][2]~q ),
	.prn(vcc));
defparam \twiddle_data[1][1][2] .is_wysiwyg = "true";
defparam \twiddle_data[1][1][2] .power_up = "low";

dffeas \twiddle_data[1][1][3] (
	.clk(clk),
	.d(\twiddle_data~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data[1][1][3]~q ),
	.prn(vcc));
defparam \twiddle_data[1][1][3] .is_wysiwyg = "true";
defparam \twiddle_data[1][1][3] .power_up = "low";

dffeas \twiddle_data[1][1][4] (
	.clk(clk),
	.d(\twiddle_data~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data[1][1][4]~q ),
	.prn(vcc));
defparam \twiddle_data[1][1][4] .is_wysiwyg = "true";
defparam \twiddle_data[1][1][4] .power_up = "low";

dffeas \twiddle_data[1][1][5] (
	.clk(clk),
	.d(\twiddle_data~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data[1][1][5]~q ),
	.prn(vcc));
defparam \twiddle_data[1][1][5] .is_wysiwyg = "true";
defparam \twiddle_data[1][1][5] .power_up = "low";

dffeas \twiddle_data[1][1][6] (
	.clk(clk),
	.d(\twiddle_data~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data[1][1][6]~q ),
	.prn(vcc));
defparam \twiddle_data[1][1][6] .is_wysiwyg = "true";
defparam \twiddle_data[1][1][6] .power_up = "low";

dffeas \twiddle_data[1][1][7] (
	.clk(clk),
	.d(\twiddle_data~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data[1][1][7]~q ),
	.prn(vcc));
defparam \twiddle_data[1][1][7] .is_wysiwyg = "true";
defparam \twiddle_data[1][1][7] .power_up = "low";

dffeas \twiddle_data[2][0][0] (
	.clk(clk),
	.d(\twiddle_data~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data[2][0][0]~q ),
	.prn(vcc));
defparam \twiddle_data[2][0][0] .is_wysiwyg = "true";
defparam \twiddle_data[2][0][0] .power_up = "low";

dffeas \twiddle_data[2][0][1] (
	.clk(clk),
	.d(\twiddle_data~33_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data[2][0][1]~q ),
	.prn(vcc));
defparam \twiddle_data[2][0][1] .is_wysiwyg = "true";
defparam \twiddle_data[2][0][1] .power_up = "low";

dffeas \twiddle_data[2][0][2] (
	.clk(clk),
	.d(\twiddle_data~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data[2][0][2]~q ),
	.prn(vcc));
defparam \twiddle_data[2][0][2] .is_wysiwyg = "true";
defparam \twiddle_data[2][0][2] .power_up = "low";

dffeas \twiddle_data[2][0][3] (
	.clk(clk),
	.d(\twiddle_data~35_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data[2][0][3]~q ),
	.prn(vcc));
defparam \twiddle_data[2][0][3] .is_wysiwyg = "true";
defparam \twiddle_data[2][0][3] .power_up = "low";

dffeas \twiddle_data[2][0][4] (
	.clk(clk),
	.d(\twiddle_data~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data[2][0][4]~q ),
	.prn(vcc));
defparam \twiddle_data[2][0][4] .is_wysiwyg = "true";
defparam \twiddle_data[2][0][4] .power_up = "low";

dffeas \twiddle_data[2][0][5] (
	.clk(clk),
	.d(\twiddle_data~37_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data[2][0][5]~q ),
	.prn(vcc));
defparam \twiddle_data[2][0][5] .is_wysiwyg = "true";
defparam \twiddle_data[2][0][5] .power_up = "low";

dffeas \twiddle_data[2][0][6] (
	.clk(clk),
	.d(\twiddle_data~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data[2][0][6]~q ),
	.prn(vcc));
defparam \twiddle_data[2][0][6] .is_wysiwyg = "true";
defparam \twiddle_data[2][0][6] .power_up = "low";

dffeas \twiddle_data[2][0][7] (
	.clk(clk),
	.d(\twiddle_data~39_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data[2][0][7]~q ),
	.prn(vcc));
defparam \twiddle_data[2][0][7] .is_wysiwyg = "true";
defparam \twiddle_data[2][0][7] .power_up = "low";

dffeas \twiddle_data[2][1][0] (
	.clk(clk),
	.d(\twiddle_data~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data[2][1][0]~q ),
	.prn(vcc));
defparam \twiddle_data[2][1][0] .is_wysiwyg = "true";
defparam \twiddle_data[2][1][0] .power_up = "low";

dffeas \twiddle_data[2][1][1] (
	.clk(clk),
	.d(\twiddle_data~41_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data[2][1][1]~q ),
	.prn(vcc));
defparam \twiddle_data[2][1][1] .is_wysiwyg = "true";
defparam \twiddle_data[2][1][1] .power_up = "low";

dffeas \twiddle_data[2][1][2] (
	.clk(clk),
	.d(\twiddle_data~42_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data[2][1][2]~q ),
	.prn(vcc));
defparam \twiddle_data[2][1][2] .is_wysiwyg = "true";
defparam \twiddle_data[2][1][2] .power_up = "low";

dffeas \twiddle_data[2][1][3] (
	.clk(clk),
	.d(\twiddle_data~43_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data[2][1][3]~q ),
	.prn(vcc));
defparam \twiddle_data[2][1][3] .is_wysiwyg = "true";
defparam \twiddle_data[2][1][3] .power_up = "low";

dffeas \twiddle_data[2][1][4] (
	.clk(clk),
	.d(\twiddle_data~44_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data[2][1][4]~q ),
	.prn(vcc));
defparam \twiddle_data[2][1][4] .is_wysiwyg = "true";
defparam \twiddle_data[2][1][4] .power_up = "low";

dffeas \twiddle_data[2][1][5] (
	.clk(clk),
	.d(\twiddle_data~45_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data[2][1][5]~q ),
	.prn(vcc));
defparam \twiddle_data[2][1][5] .is_wysiwyg = "true";
defparam \twiddle_data[2][1][5] .power_up = "low";

dffeas \twiddle_data[2][1][6] (
	.clk(clk),
	.d(\twiddle_data~46_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data[2][1][6]~q ),
	.prn(vcc));
defparam \twiddle_data[2][1][6] .is_wysiwyg = "true";
defparam \twiddle_data[2][1][6] .power_up = "low";

dffeas \twiddle_data[2][1][7] (
	.clk(clk),
	.d(\twiddle_data~47_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data[2][1][7]~q ),
	.prn(vcc));
defparam \twiddle_data[2][1][7] .is_wysiwyg = "true";
defparam \twiddle_data[2][1][7] .power_up = "low";

cycloneiii_lcell_comb \wc_vec~6 (
	.dataa(reset_n),
	.datab(\sel_we|wc_i~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wc_vec~6_combout ),
	.cout());
defparam \wc_vec~6 .lut_mask = 16'hEEEE;
defparam \wc_vec~6 .sum_lutc_input = "datac";

dffeas \p_tdl[16][0] (
	.clk(clk),
	.d(\p_cd_en[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[16][0]~q ),
	.prn(vcc));
defparam \p_tdl[16][0] .is_wysiwyg = "true";
defparam \p_tdl[16][0] .power_up = "low";

dffeas \p_tdl[16][2] (
	.clk(clk),
	.d(\p_cd_en[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[16][2]~q ),
	.prn(vcc));
defparam \p_tdl[16][2] .is_wysiwyg = "true";
defparam \p_tdl[16][2] .power_up = "low";

dffeas \p_tdl[16][1] (
	.clk(clk),
	.d(\p_cd_en[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[16][1]~q ),
	.prn(vcc));
defparam \p_tdl[16][1] .is_wysiwyg = "true";
defparam \p_tdl[16][1] .power_up = "low";

cycloneiii_lcell_comb \wd_vec~6 (
	.dataa(reset_n),
	.datab(\sel_we|wd_i~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wd_vec~6_combout ),
	.cout());
defparam \wd_vec~6 .lut_mask = 16'hEEEE;
defparam \wd_vec~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \twiddle_data~0 (
	.dataa(\twrom|gen_M4K:cos_1n|gen_auto:altsyncram_component|auto_generated|q_a[0] ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data~0_combout ),
	.cout());
defparam \twiddle_data~0 .lut_mask = 16'hAAFF;
defparam \twiddle_data~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \twiddle_data~1 (
	.dataa(\twrom|gen_M4K:cos_1n|gen_auto:altsyncram_component|auto_generated|q_a[1] ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data~1_combout ),
	.cout());
defparam \twiddle_data~1 .lut_mask = 16'hAAFF;
defparam \twiddle_data~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \twiddle_data~2 (
	.dataa(\twrom|gen_M4K:cos_1n|gen_auto:altsyncram_component|auto_generated|q_a[2] ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data~2_combout ),
	.cout());
defparam \twiddle_data~2 .lut_mask = 16'hAAFF;
defparam \twiddle_data~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \twiddle_data~3 (
	.dataa(\twrom|gen_M4K:cos_1n|gen_auto:altsyncram_component|auto_generated|q_a[3] ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data~3_combout ),
	.cout());
defparam \twiddle_data~3 .lut_mask = 16'hAAFF;
defparam \twiddle_data~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \twiddle_data~4 (
	.dataa(\twrom|gen_M4K:cos_1n|gen_auto:altsyncram_component|auto_generated|q_a[4] ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data~4_combout ),
	.cout());
defparam \twiddle_data~4 .lut_mask = 16'hAAFF;
defparam \twiddle_data~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \twiddle_data~5 (
	.dataa(\twrom|gen_M4K:cos_1n|gen_auto:altsyncram_component|auto_generated|q_a[5] ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data~5_combout ),
	.cout());
defparam \twiddle_data~5 .lut_mask = 16'hAAFF;
defparam \twiddle_data~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \twiddle_data~6 (
	.dataa(\twrom|gen_M4K:cos_1n|gen_auto:altsyncram_component|auto_generated|q_a[6] ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data~6_combout ),
	.cout());
defparam \twiddle_data~6 .lut_mask = 16'hAAFF;
defparam \twiddle_data~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \twiddle_data~7 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:cos_1n|gen_auto:altsyncram_component|auto_generated|q_a[7] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~7_combout ),
	.cout());
defparam \twiddle_data~7 .lut_mask = 16'hEEEE;
defparam \twiddle_data~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \twiddle_data~8 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:sin_1n|gen_auto:altsyncram_component|auto_generated|q_a[0] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~8_combout ),
	.cout());
defparam \twiddle_data~8 .lut_mask = 16'hEEEE;
defparam \twiddle_data~8 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \twiddle_data~9 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:sin_1n|gen_auto:altsyncram_component|auto_generated|q_a[1] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~9_combout ),
	.cout());
defparam \twiddle_data~9 .lut_mask = 16'hEEEE;
defparam \twiddle_data~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \twiddle_data~10 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:sin_1n|gen_auto:altsyncram_component|auto_generated|q_a[2] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~10_combout ),
	.cout());
defparam \twiddle_data~10 .lut_mask = 16'hEEEE;
defparam \twiddle_data~10 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \twiddle_data~11 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:sin_1n|gen_auto:altsyncram_component|auto_generated|q_a[3] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~11_combout ),
	.cout());
defparam \twiddle_data~11 .lut_mask = 16'hEEEE;
defparam \twiddle_data~11 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \twiddle_data~12 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:sin_1n|gen_auto:altsyncram_component|auto_generated|q_a[4] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~12_combout ),
	.cout());
defparam \twiddle_data~12 .lut_mask = 16'hEEEE;
defparam \twiddle_data~12 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \twiddle_data~13 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:sin_1n|gen_auto:altsyncram_component|auto_generated|q_a[5] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~13_combout ),
	.cout());
defparam \twiddle_data~13 .lut_mask = 16'hEEEE;
defparam \twiddle_data~13 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \twiddle_data~14 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:sin_1n|gen_auto:altsyncram_component|auto_generated|q_a[6] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~14_combout ),
	.cout());
defparam \twiddle_data~14 .lut_mask = 16'hEEEE;
defparam \twiddle_data~14 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \twiddle_data~15 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:sin_1n|gen_auto:altsyncram_component|auto_generated|q_a[7] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~15_combout ),
	.cout());
defparam \twiddle_data~15 .lut_mask = 16'hEEEE;
defparam \twiddle_data~15 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \twiddle_data~16 (
	.dataa(\twrom|gen_M4K:cos_2n|gen_auto:altsyncram_component|auto_generated|q_a[0] ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data~16_combout ),
	.cout());
defparam \twiddle_data~16 .lut_mask = 16'hAAFF;
defparam \twiddle_data~16 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \twiddle_data~17 (
	.dataa(\twrom|gen_M4K:cos_2n|gen_auto:altsyncram_component|auto_generated|q_a[1] ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data~17_combout ),
	.cout());
defparam \twiddle_data~17 .lut_mask = 16'hAAFF;
defparam \twiddle_data~17 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \twiddle_data~18 (
	.dataa(\twrom|gen_M4K:cos_2n|gen_auto:altsyncram_component|auto_generated|q_a[2] ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data~18_combout ),
	.cout());
defparam \twiddle_data~18 .lut_mask = 16'hAAFF;
defparam \twiddle_data~18 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \twiddle_data~19 (
	.dataa(\twrom|gen_M4K:cos_2n|gen_auto:altsyncram_component|auto_generated|q_a[3] ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data~19_combout ),
	.cout());
defparam \twiddle_data~19 .lut_mask = 16'hAAFF;
defparam \twiddle_data~19 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \twiddle_data~20 (
	.dataa(\twrom|gen_M4K:cos_2n|gen_auto:altsyncram_component|auto_generated|q_a[4] ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data~20_combout ),
	.cout());
defparam \twiddle_data~20 .lut_mask = 16'hAAFF;
defparam \twiddle_data~20 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \twiddle_data~21 (
	.dataa(\twrom|gen_M4K:cos_2n|gen_auto:altsyncram_component|auto_generated|q_a[5] ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data~21_combout ),
	.cout());
defparam \twiddle_data~21 .lut_mask = 16'hAAFF;
defparam \twiddle_data~21 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \twiddle_data~22 (
	.dataa(\twrom|gen_M4K:cos_2n|gen_auto:altsyncram_component|auto_generated|q_a[6] ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data~22_combout ),
	.cout());
defparam \twiddle_data~22 .lut_mask = 16'hAAFF;
defparam \twiddle_data~22 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \twiddle_data~23 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:cos_2n|gen_auto:altsyncram_component|auto_generated|q_a[7] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~23_combout ),
	.cout());
defparam \twiddle_data~23 .lut_mask = 16'hEEEE;
defparam \twiddle_data~23 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \twiddle_data~24 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:sin_2n|gen_auto:altsyncram_component|auto_generated|q_a[0] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~24_combout ),
	.cout());
defparam \twiddle_data~24 .lut_mask = 16'hEEEE;
defparam \twiddle_data~24 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \twiddle_data~25 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:sin_2n|gen_auto:altsyncram_component|auto_generated|q_a[1] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~25_combout ),
	.cout());
defparam \twiddle_data~25 .lut_mask = 16'hEEEE;
defparam \twiddle_data~25 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \twiddle_data~26 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:sin_2n|gen_auto:altsyncram_component|auto_generated|q_a[2] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~26_combout ),
	.cout());
defparam \twiddle_data~26 .lut_mask = 16'hEEEE;
defparam \twiddle_data~26 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \twiddle_data~27 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:sin_2n|gen_auto:altsyncram_component|auto_generated|q_a[3] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~27_combout ),
	.cout());
defparam \twiddle_data~27 .lut_mask = 16'hEEEE;
defparam \twiddle_data~27 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \twiddle_data~28 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:sin_2n|gen_auto:altsyncram_component|auto_generated|q_a[4] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~28_combout ),
	.cout());
defparam \twiddle_data~28 .lut_mask = 16'hEEEE;
defparam \twiddle_data~28 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \twiddle_data~29 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:sin_2n|gen_auto:altsyncram_component|auto_generated|q_a[5] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~29_combout ),
	.cout());
defparam \twiddle_data~29 .lut_mask = 16'hEEEE;
defparam \twiddle_data~29 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \twiddle_data~30 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:sin_2n|gen_auto:altsyncram_component|auto_generated|q_a[6] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~30_combout ),
	.cout());
defparam \twiddle_data~30 .lut_mask = 16'hEEEE;
defparam \twiddle_data~30 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \twiddle_data~31 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:sin_2n|gen_auto:altsyncram_component|auto_generated|q_a[7] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~31_combout ),
	.cout());
defparam \twiddle_data~31 .lut_mask = 16'hEEEE;
defparam \twiddle_data~31 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \twiddle_data~32 (
	.dataa(\twrom|gen_M4K:cos_3n|gen_auto:altsyncram_component|auto_generated|q_a[0] ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data~32_combout ),
	.cout());
defparam \twiddle_data~32 .lut_mask = 16'hAAFF;
defparam \twiddle_data~32 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \twiddle_data~33 (
	.dataa(\twrom|gen_M4K:cos_3n|gen_auto:altsyncram_component|auto_generated|q_a[1] ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data~33_combout ),
	.cout());
defparam \twiddle_data~33 .lut_mask = 16'hAAFF;
defparam \twiddle_data~33 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \twiddle_data~34 (
	.dataa(\twrom|gen_M4K:cos_3n|gen_auto:altsyncram_component|auto_generated|q_a[2] ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data~34_combout ),
	.cout());
defparam \twiddle_data~34 .lut_mask = 16'hAAFF;
defparam \twiddle_data~34 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \twiddle_data~35 (
	.dataa(\twrom|gen_M4K:cos_3n|gen_auto:altsyncram_component|auto_generated|q_a[3] ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data~35_combout ),
	.cout());
defparam \twiddle_data~35 .lut_mask = 16'hAAFF;
defparam \twiddle_data~35 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \twiddle_data~36 (
	.dataa(\twrom|gen_M4K:cos_3n|gen_auto:altsyncram_component|auto_generated|q_a[4] ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data~36_combout ),
	.cout());
defparam \twiddle_data~36 .lut_mask = 16'hAAFF;
defparam \twiddle_data~36 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \twiddle_data~37 (
	.dataa(\twrom|gen_M4K:cos_3n|gen_auto:altsyncram_component|auto_generated|q_a[5] ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data~37_combout ),
	.cout());
defparam \twiddle_data~37 .lut_mask = 16'hAAFF;
defparam \twiddle_data~37 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \twiddle_data~38 (
	.dataa(\twrom|gen_M4K:cos_3n|gen_auto:altsyncram_component|auto_generated|q_a[6] ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data~38_combout ),
	.cout());
defparam \twiddle_data~38 .lut_mask = 16'hAAFF;
defparam \twiddle_data~38 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \twiddle_data~39 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:cos_3n|gen_auto:altsyncram_component|auto_generated|q_a[7] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~39_combout ),
	.cout());
defparam \twiddle_data~39 .lut_mask = 16'hEEEE;
defparam \twiddle_data~39 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \twiddle_data~40 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:sin_3n|gen_auto:altsyncram_component|auto_generated|q_a[0] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~40_combout ),
	.cout());
defparam \twiddle_data~40 .lut_mask = 16'hEEEE;
defparam \twiddle_data~40 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \twiddle_data~41 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:sin_3n|gen_auto:altsyncram_component|auto_generated|q_a[1] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~41_combout ),
	.cout());
defparam \twiddle_data~41 .lut_mask = 16'hEEEE;
defparam \twiddle_data~41 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \twiddle_data~42 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:sin_3n|gen_auto:altsyncram_component|auto_generated|q_a[2] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~42_combout ),
	.cout());
defparam \twiddle_data~42 .lut_mask = 16'hEEEE;
defparam \twiddle_data~42 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \twiddle_data~43 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:sin_3n|gen_auto:altsyncram_component|auto_generated|q_a[3] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~43_combout ),
	.cout());
defparam \twiddle_data~43 .lut_mask = 16'hEEEE;
defparam \twiddle_data~43 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \twiddle_data~44 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:sin_3n|gen_auto:altsyncram_component|auto_generated|q_a[4] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~44_combout ),
	.cout());
defparam \twiddle_data~44 .lut_mask = 16'hEEEE;
defparam \twiddle_data~44 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \twiddle_data~45 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:sin_3n|gen_auto:altsyncram_component|auto_generated|q_a[5] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~45_combout ),
	.cout());
defparam \twiddle_data~45 .lut_mask = 16'hEEEE;
defparam \twiddle_data~45 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \twiddle_data~46 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:sin_3n|gen_auto:altsyncram_component|auto_generated|q_a[6] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~46_combout ),
	.cout());
defparam \twiddle_data~46 .lut_mask = 16'hEEEE;
defparam \twiddle_data~46 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \twiddle_data~47 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:sin_3n|gen_auto:altsyncram_component|auto_generated|q_a[7] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~47_combout ),
	.cout());
defparam \twiddle_data~47 .lut_mask = 16'hEEEE;
defparam \twiddle_data~47 .sum_lutc_input = "datac";

dffeas en_slb(
	.clk(clk),
	.d(\en_slb~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\en_slb~q ),
	.prn(vcc));
defparam en_slb.is_wysiwyg = "true";
defparam en_slb.power_up = "low";

dffeas \ram_a_not_b_vec[26] (
	.clk(clk),
	.d(\ram_a_not_b_vec~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\ram_a_not_b_vec[26]~q ),
	.prn(vcc));
defparam \ram_a_not_b_vec[26] .is_wysiwyg = "true";
defparam \ram_a_not_b_vec[26] .power_up = "low";

dffeas \p_cd_en[2] (
	.clk(clk),
	.d(\p_tdl[14][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_cd_en[2]~q ),
	.prn(vcc));
defparam \p_cd_en[2] .is_wysiwyg = "true";
defparam \p_cd_en[2] .power_up = "low";

dffeas \p_cd_en[0] (
	.clk(clk),
	.d(\p_tdl[14][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_cd_en[0]~q ),
	.prn(vcc));
defparam \p_cd_en[0] .is_wysiwyg = "true";
defparam \p_cd_en[0] .power_up = "low";

dffeas \p_cd_en[1] (
	.clk(clk),
	.d(\p_tdl[14][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_cd_en[1]~q ),
	.prn(vcc));
defparam \p_cd_en[1] .is_wysiwyg = "true";
defparam \p_cd_en[1] .power_up = "low";

cycloneiii_lcell_comb \en_slb~0 (
	.dataa(\delay_ctrl_np|tdl_arr[9]~q ),
	.datab(\gen_gt256_mk:ctrl|p[1]~q ),
	.datac(\gen_gt256_mk:ctrl|p[2]~q ),
	.datad(\gen_gt256_mk:ctrl|p[0]~q ),
	.cin(gnd),
	.combout(\en_slb~0_combout ),
	.cout());
defparam \en_slb~0 .lut_mask = 16'hFEFF;
defparam \en_slb~0 .sum_lutc_input = "datac";

dffeas \ram_a_not_b_vec[25] (
	.clk(clk),
	.d(\ram_a_not_b_vec~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\ram_a_not_b_vec[25]~q ),
	.prn(vcc));
defparam \ram_a_not_b_vec[25] .is_wysiwyg = "true";
defparam \ram_a_not_b_vec[25] .power_up = "low";

cycloneiii_lcell_comb \ram_a_not_b_vec~0 (
	.dataa(\ram_a_not_b_vec[25]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\ram_a_not_b_vec~0_combout ),
	.cout());
defparam \ram_a_not_b_vec~0 .lut_mask = 16'hAAFF;
defparam \ram_a_not_b_vec~0 .sum_lutc_input = "datac";

dffeas \p_tdl[14][2] (
	.clk(clk),
	.d(\p_tdl[13][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[14][2]~q ),
	.prn(vcc));
defparam \p_tdl[14][2] .is_wysiwyg = "true";
defparam \p_tdl[14][2] .power_up = "low";

dffeas \p_tdl[14][0] (
	.clk(clk),
	.d(\p_tdl[13][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[14][0]~q ),
	.prn(vcc));
defparam \p_tdl[14][0] .is_wysiwyg = "true";
defparam \p_tdl[14][0] .power_up = "low";

dffeas \p_tdl[14][1] (
	.clk(clk),
	.d(\p_tdl[13][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[14][1]~q ),
	.prn(vcc));
defparam \p_tdl[14][1] .is_wysiwyg = "true";
defparam \p_tdl[14][1] .power_up = "low";

dffeas \ram_a_not_b_vec[24] (
	.clk(clk),
	.d(\ram_a_not_b_vec~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\ram_a_not_b_vec[24]~q ),
	.prn(vcc));
defparam \ram_a_not_b_vec[24] .is_wysiwyg = "true";
defparam \ram_a_not_b_vec[24] .power_up = "low";

cycloneiii_lcell_comb \ram_a_not_b_vec~1 (
	.dataa(\ram_a_not_b_vec[24]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\ram_a_not_b_vec~1_combout ),
	.cout());
defparam \ram_a_not_b_vec~1 .lut_mask = 16'hAAFF;
defparam \ram_a_not_b_vec~1 .sum_lutc_input = "datac";

dffeas \p_tdl[13][2] (
	.clk(clk),
	.d(\p_tdl[12][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[13][2]~q ),
	.prn(vcc));
defparam \p_tdl[13][2] .is_wysiwyg = "true";
defparam \p_tdl[13][2] .power_up = "low";

dffeas \p_tdl[13][0] (
	.clk(clk),
	.d(\p_tdl[12][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[13][0]~q ),
	.prn(vcc));
defparam \p_tdl[13][0] .is_wysiwyg = "true";
defparam \p_tdl[13][0] .power_up = "low";

dffeas \p_tdl[13][1] (
	.clk(clk),
	.d(\p_tdl[12][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[13][1]~q ),
	.prn(vcc));
defparam \p_tdl[13][1] .is_wysiwyg = "true";
defparam \p_tdl[13][1] .power_up = "low";

dffeas \ram_a_not_b_vec[23] (
	.clk(clk),
	.d(\ram_a_not_b_vec~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\ram_a_not_b_vec[23]~q ),
	.prn(vcc));
defparam \ram_a_not_b_vec[23] .is_wysiwyg = "true";
defparam \ram_a_not_b_vec[23] .power_up = "low";

cycloneiii_lcell_comb \ram_a_not_b_vec~2 (
	.dataa(\ram_a_not_b_vec[23]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\ram_a_not_b_vec~2_combout ),
	.cout());
defparam \ram_a_not_b_vec~2 .lut_mask = 16'hAAFF;
defparam \ram_a_not_b_vec~2 .sum_lutc_input = "datac";

dffeas \p_tdl[12][2] (
	.clk(clk),
	.d(\p_tdl[11][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[12][2]~q ),
	.prn(vcc));
defparam \p_tdl[12][2] .is_wysiwyg = "true";
defparam \p_tdl[12][2] .power_up = "low";

dffeas \p_tdl[12][0] (
	.clk(clk),
	.d(\p_tdl[11][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[12][0]~q ),
	.prn(vcc));
defparam \p_tdl[12][0] .is_wysiwyg = "true";
defparam \p_tdl[12][0] .power_up = "low";

dffeas \p_tdl[12][1] (
	.clk(clk),
	.d(\p_tdl[11][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[12][1]~q ),
	.prn(vcc));
defparam \p_tdl[12][1] .is_wysiwyg = "true";
defparam \p_tdl[12][1] .power_up = "low";

dffeas \sw_r_tdl[4][0] (
	.clk(clk),
	.d(\sw_r_tdl[3][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\sw_r_tdl[4][0]~q ),
	.prn(vcc));
defparam \sw_r_tdl[4][0] .is_wysiwyg = "true";
defparam \sw_r_tdl[4][0] .power_up = "low";

dffeas \sw_r_tdl[4][1] (
	.clk(clk),
	.d(\sw_r_tdl[3][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\sw_r_tdl[4][1]~q ),
	.prn(vcc));
defparam \sw_r_tdl[4][1] .is_wysiwyg = "true";
defparam \sw_r_tdl[4][1] .power_up = "low";

dffeas \ram_a_not_b_vec[22] (
	.clk(clk),
	.d(\ram_a_not_b_vec~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\ram_a_not_b_vec[22]~q ),
	.prn(vcc));
defparam \ram_a_not_b_vec[22] .is_wysiwyg = "true";
defparam \ram_a_not_b_vec[22] .power_up = "low";

cycloneiii_lcell_comb \ram_a_not_b_vec~3 (
	.dataa(\ram_a_not_b_vec[22]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\ram_a_not_b_vec~3_combout ),
	.cout());
defparam \ram_a_not_b_vec~3 .lut_mask = 16'hAAFF;
defparam \ram_a_not_b_vec~3 .sum_lutc_input = "datac";

dffeas \p_tdl[11][2] (
	.clk(clk),
	.d(\p_tdl[10][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[11][2]~q ),
	.prn(vcc));
defparam \p_tdl[11][2] .is_wysiwyg = "true";
defparam \p_tdl[11][2] .power_up = "low";

dffeas \p_tdl[11][0] (
	.clk(clk),
	.d(\p_tdl[10][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[11][0]~q ),
	.prn(vcc));
defparam \p_tdl[11][0] .is_wysiwyg = "true";
defparam \p_tdl[11][0] .power_up = "low";

dffeas \p_tdl[11][1] (
	.clk(clk),
	.d(\p_tdl[10][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[11][1]~q ),
	.prn(vcc));
defparam \p_tdl[11][1] .is_wysiwyg = "true";
defparam \p_tdl[11][1] .power_up = "low";

dffeas \data_rdy_vec[10] (
	.clk(clk),
	.d(\data_rdy_vec~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_rdy_vec[10]~q ),
	.prn(vcc));
defparam \data_rdy_vec[10] .is_wysiwyg = "true";
defparam \data_rdy_vec[10] .power_up = "low";

dffeas \ram_a_not_b_vec[10] (
	.clk(clk),
	.d(\ram_a_not_b_vec~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\ram_a_not_b_vec[10]~q ),
	.prn(vcc));
defparam \ram_a_not_b_vec[10] .is_wysiwyg = "true";
defparam \ram_a_not_b_vec[10] .power_up = "low";

dffeas \sw_r_tdl[3][0] (
	.clk(clk),
	.d(\sw_r_tdl[2][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\sw_r_tdl[3][0]~q ),
	.prn(vcc));
defparam \sw_r_tdl[3][0] .is_wysiwyg = "true";
defparam \sw_r_tdl[3][0] .power_up = "low";

dffeas \sw_r_tdl[3][1] (
	.clk(clk),
	.d(\sw_r_tdl[2][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\sw_r_tdl[3][1]~q ),
	.prn(vcc));
defparam \sw_r_tdl[3][1] .is_wysiwyg = "true";
defparam \sw_r_tdl[3][1] .power_up = "low";

dffeas \ram_a_not_b_vec[21] (
	.clk(clk),
	.d(\ram_a_not_b_vec~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\ram_a_not_b_vec[21]~q ),
	.prn(vcc));
defparam \ram_a_not_b_vec[21] .is_wysiwyg = "true";
defparam \ram_a_not_b_vec[21] .power_up = "low";

cycloneiii_lcell_comb \ram_a_not_b_vec~4 (
	.dataa(\ram_a_not_b_vec[21]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\ram_a_not_b_vec~4_combout ),
	.cout());
defparam \ram_a_not_b_vec~4 .lut_mask = 16'hAAFF;
defparam \ram_a_not_b_vec~4 .sum_lutc_input = "datac";

dffeas \p_tdl[10][2] (
	.clk(clk),
	.d(\p_tdl[9][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[10][2]~q ),
	.prn(vcc));
defparam \p_tdl[10][2] .is_wysiwyg = "true";
defparam \p_tdl[10][2] .power_up = "low";

dffeas \p_tdl[10][0] (
	.clk(clk),
	.d(\p_tdl[9][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[10][0]~q ),
	.prn(vcc));
defparam \p_tdl[10][0] .is_wysiwyg = "true";
defparam \p_tdl[10][0] .power_up = "low";

dffeas \p_tdl[10][1] (
	.clk(clk),
	.d(\p_tdl[9][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[10][1]~q ),
	.prn(vcc));
defparam \p_tdl[10][1] .is_wysiwyg = "true";
defparam \p_tdl[10][1] .power_up = "low";

dffeas \data_rdy_vec[9] (
	.clk(clk),
	.d(\data_rdy_vec~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_rdy_vec[9]~q ),
	.prn(vcc));
defparam \data_rdy_vec[9] .is_wysiwyg = "true";
defparam \data_rdy_vec[9] .power_up = "low";

cycloneiii_lcell_comb \data_rdy_vec~5 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~5_combout ),
	.cout());
defparam \data_rdy_vec~5 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~5 .sum_lutc_input = "datac";

dffeas \ram_a_not_b_vec[9] (
	.clk(clk),
	.d(\ram_a_not_b_vec~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\ram_a_not_b_vec[9]~q ),
	.prn(vcc));
defparam \ram_a_not_b_vec[9] .is_wysiwyg = "true";
defparam \ram_a_not_b_vec[9] .power_up = "low";

cycloneiii_lcell_comb \ram_a_not_b_vec~5 (
	.dataa(\ram_a_not_b_vec[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\ram_a_not_b_vec~5_combout ),
	.cout());
defparam \ram_a_not_b_vec~5 .lut_mask = 16'hAAFF;
defparam \ram_a_not_b_vec~5 .sum_lutc_input = "datac";

dffeas \sw_r_tdl[2][0] (
	.clk(clk),
	.d(\sw_r_tdl[1][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\sw_r_tdl[2][0]~q ),
	.prn(vcc));
defparam \sw_r_tdl[2][0] .is_wysiwyg = "true";
defparam \sw_r_tdl[2][0] .power_up = "low";

dffeas \sw_r_tdl[2][1] (
	.clk(clk),
	.d(\sw_r_tdl[1][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\sw_r_tdl[2][1]~q ),
	.prn(vcc));
defparam \sw_r_tdl[2][1] .is_wysiwyg = "true";
defparam \sw_r_tdl[2][1] .power_up = "low";

dffeas \ram_a_not_b_vec[20] (
	.clk(clk),
	.d(\ram_a_not_b_vec~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\ram_a_not_b_vec[20]~q ),
	.prn(vcc));
defparam \ram_a_not_b_vec[20] .is_wysiwyg = "true";
defparam \ram_a_not_b_vec[20] .power_up = "low";

cycloneiii_lcell_comb \ram_a_not_b_vec~6 (
	.dataa(\ram_a_not_b_vec[20]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\ram_a_not_b_vec~6_combout ),
	.cout());
defparam \ram_a_not_b_vec~6 .lut_mask = 16'hAAFF;
defparam \ram_a_not_b_vec~6 .sum_lutc_input = "datac";

dffeas \p_tdl[9][2] (
	.clk(clk),
	.d(\p_tdl[8][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[9][2]~q ),
	.prn(vcc));
defparam \p_tdl[9][2] .is_wysiwyg = "true";
defparam \p_tdl[9][2] .power_up = "low";

dffeas \p_tdl[9][0] (
	.clk(clk),
	.d(\p_tdl[8][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[9][0]~q ),
	.prn(vcc));
defparam \p_tdl[9][0] .is_wysiwyg = "true";
defparam \p_tdl[9][0] .power_up = "low";

dffeas \p_tdl[9][1] (
	.clk(clk),
	.d(\p_tdl[8][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[9][1]~q ),
	.prn(vcc));
defparam \p_tdl[9][1] .is_wysiwyg = "true";
defparam \p_tdl[9][1] .power_up = "low";

dffeas \ram_a_not_b_vec[29] (
	.clk(clk),
	.d(\ram_a_not_b_vec~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\ram_a_not_b_vec[29]~q ),
	.prn(vcc));
defparam \ram_a_not_b_vec[29] .is_wysiwyg = "true";
defparam \ram_a_not_b_vec[29] .power_up = "low";

dffeas \ram_a_not_b_vec[1] (
	.clk(clk),
	.d(\ram_a_not_b_vec~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\ram_a_not_b_vec[1]~q ),
	.prn(vcc));
defparam \ram_a_not_b_vec[1] .is_wysiwyg = "true";
defparam \ram_a_not_b_vec[1] .power_up = "low";

cycloneiii_lcell_comb \wren_b~0 (
	.dataa(\ram_a_not_b_vec[29]~q ),
	.datab(\writer|wren[0]~q ),
	.datac(gnd),
	.datad(\ram_a_not_b_vec[1]~q ),
	.cin(gnd),
	.combout(\wren_b~0_combout ),
	.cout());
defparam \wren_b~0 .lut_mask = 16'hAACC;
defparam \wren_b~0 .sum_lutc_input = "datac";

dffeas \ram_a_not_b_vec[7] (
	.clk(clk),
	.d(\ram_a_not_b_vec~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\ram_a_not_b_vec[7]~q ),
	.prn(vcc));
defparam \ram_a_not_b_vec[7] .is_wysiwyg = "true";
defparam \ram_a_not_b_vec[7] .power_up = "low";

cycloneiii_lcell_comb \wren_a~0 (
	.dataa(\writer|wren[0]~q ),
	.datab(\ram_a_not_b_vec[1]~q ),
	.datac(gnd),
	.datad(\ram_a_not_b_vec[29]~q ),
	.cin(gnd),
	.combout(\wren_a~0_combout ),
	.cout());
defparam \wren_a~0 .lut_mask = 16'h88BB;
defparam \wren_a~0 .sum_lutc_input = "datac";

dffeas \data_rdy_vec[8] (
	.clk(clk),
	.d(\data_rdy_vec~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_rdy_vec[8]~q ),
	.prn(vcc));
defparam \data_rdy_vec[8] .is_wysiwyg = "true";
defparam \data_rdy_vec[8] .power_up = "low";

cycloneiii_lcell_comb \data_rdy_vec~6 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~6_combout ),
	.cout());
defparam \data_rdy_vec~6 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~6 .sum_lutc_input = "datac";

dffeas \ram_a_not_b_vec[8] (
	.clk(clk),
	.d(\ram_a_not_b_vec~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\ram_a_not_b_vec[8]~q ),
	.prn(vcc));
defparam \ram_a_not_b_vec[8] .is_wysiwyg = "true";
defparam \ram_a_not_b_vec[8] .power_up = "low";

cycloneiii_lcell_comb \ram_a_not_b_vec~7 (
	.dataa(\ram_a_not_b_vec[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\ram_a_not_b_vec~7_combout ),
	.cout());
defparam \ram_a_not_b_vec~7 .lut_mask = 16'hAAFF;
defparam \ram_a_not_b_vec~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wren_b~1 (
	.dataa(\ram_a_not_b_vec[29]~q ),
	.datab(\writer|wren[1]~q ),
	.datac(gnd),
	.datad(\ram_a_not_b_vec[1]~q ),
	.cin(gnd),
	.combout(\wren_b~1_combout ),
	.cout());
defparam \wren_b~1 .lut_mask = 16'hAACC;
defparam \wren_b~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wren_a~1 (
	.dataa(\writer|wren[1]~q ),
	.datab(\ram_a_not_b_vec[1]~q ),
	.datac(gnd),
	.datad(\ram_a_not_b_vec[29]~q ),
	.cin(gnd),
	.combout(\wren_a~1_combout ),
	.cout());
defparam \wren_a~1 .lut_mask = 16'h88BB;
defparam \wren_a~1 .sum_lutc_input = "datac";

dffeas \sw_r_tdl[1][0] (
	.clk(clk),
	.d(\sw_r_tdl[0][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\sw_r_tdl[1][0]~q ),
	.prn(vcc));
defparam \sw_r_tdl[1][0] .is_wysiwyg = "true";
defparam \sw_r_tdl[1][0] .power_up = "low";

cycloneiii_lcell_comb \wren_b~2 (
	.dataa(\ram_a_not_b_vec[29]~q ),
	.datab(\writer|wren[2]~q ),
	.datac(gnd),
	.datad(\ram_a_not_b_vec[1]~q ),
	.cin(gnd),
	.combout(\wren_b~2_combout ),
	.cout());
defparam \wren_b~2 .lut_mask = 16'hAACC;
defparam \wren_b~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wren_a~2 (
	.dataa(\writer|wren[2]~q ),
	.datab(\ram_a_not_b_vec[1]~q ),
	.datac(gnd),
	.datad(\ram_a_not_b_vec[29]~q ),
	.cin(gnd),
	.combout(\wren_a~2_combout ),
	.cout());
defparam \wren_a~2 .lut_mask = 16'h88BB;
defparam \wren_a~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wren_b~3 (
	.dataa(\ram_a_not_b_vec[29]~q ),
	.datab(\writer|wren[3]~q ),
	.datac(gnd),
	.datad(\ram_a_not_b_vec[1]~q ),
	.cin(gnd),
	.combout(\wren_b~3_combout ),
	.cout());
defparam \wren_b~3 .lut_mask = 16'hAACC;
defparam \wren_b~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wren_a~3 (
	.dataa(\writer|wren[3]~q ),
	.datab(\ram_a_not_b_vec[1]~q ),
	.datac(gnd),
	.datad(\ram_a_not_b_vec[29]~q ),
	.cin(gnd),
	.combout(\wren_a~3_combout ),
	.cout());
defparam \wren_a~3 .lut_mask = 16'h88BB;
defparam \wren_a~3 .sum_lutc_input = "datac";

dffeas \sw_r_tdl[1][1] (
	.clk(clk),
	.d(\sw_r_tdl[0][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\sw_r_tdl[1][1]~q ),
	.prn(vcc));
defparam \sw_r_tdl[1][1] .is_wysiwyg = "true";
defparam \sw_r_tdl[1][1] .power_up = "low";

dffeas \ram_a_not_b_vec[19] (
	.clk(clk),
	.d(\ram_a_not_b_vec~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\ram_a_not_b_vec[19]~q ),
	.prn(vcc));
defparam \ram_a_not_b_vec[19] .is_wysiwyg = "true";
defparam \ram_a_not_b_vec[19] .power_up = "low";

cycloneiii_lcell_comb \ram_a_not_b_vec~8 (
	.dataa(\ram_a_not_b_vec[19]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\ram_a_not_b_vec~8_combout ),
	.cout());
defparam \ram_a_not_b_vec~8 .lut_mask = 16'hAAFF;
defparam \ram_a_not_b_vec~8 .sum_lutc_input = "datac";

dffeas \p_tdl[8][2] (
	.clk(clk),
	.d(\p_tdl[7][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[8][2]~q ),
	.prn(vcc));
defparam \p_tdl[8][2] .is_wysiwyg = "true";
defparam \p_tdl[8][2] .power_up = "low";

dffeas \p_tdl[8][0] (
	.clk(clk),
	.d(\p_tdl[7][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[8][0]~q ),
	.prn(vcc));
defparam \p_tdl[8][0] .is_wysiwyg = "true";
defparam \p_tdl[8][0] .power_up = "low";

dffeas \p_tdl[8][1] (
	.clk(clk),
	.d(\p_tdl[7][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[8][1]~q ),
	.prn(vcc));
defparam \p_tdl[8][1] .is_wysiwyg = "true";
defparam \p_tdl[8][1] .power_up = "low";

dffeas \ram_a_not_b_vec[28] (
	.clk(clk),
	.d(\ram_a_not_b_vec~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\ram_a_not_b_vec[28]~q ),
	.prn(vcc));
defparam \ram_a_not_b_vec[28] .is_wysiwyg = "true";
defparam \ram_a_not_b_vec[28] .power_up = "low";

cycloneiii_lcell_comb \ram_a_not_b_vec~9 (
	.dataa(\ram_a_not_b_vec[28]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\ram_a_not_b_vec~9_combout ),
	.cout());
defparam \ram_a_not_b_vec~9 .lut_mask = 16'hAAFF;
defparam \ram_a_not_b_vec~9 .sum_lutc_input = "datac";

dffeas \ram_a_not_b_vec[0] (
	.clk(clk),
	.d(\ram_a_not_b_vec~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\ram_a_not_b_vec[0]~q ),
	.prn(vcc));
defparam \ram_a_not_b_vec[0] .is_wysiwyg = "true";
defparam \ram_a_not_b_vec[0] .power_up = "low";

cycloneiii_lcell_comb \ram_a_not_b_vec~10 (
	.dataa(\ram_a_not_b_vec[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\ram_a_not_b_vec~10_combout ),
	.cout());
defparam \ram_a_not_b_vec~10 .lut_mask = 16'hAAFF;
defparam \ram_a_not_b_vec~10 .sum_lutc_input = "datac";

dffeas \ram_a_not_b_vec[6] (
	.clk(clk),
	.d(\ram_a_not_b_vec~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\ram_a_not_b_vec[6]~q ),
	.prn(vcc));
defparam \ram_a_not_b_vec[6] .is_wysiwyg = "true";
defparam \ram_a_not_b_vec[6] .power_up = "low";

cycloneiii_lcell_comb \ram_a_not_b_vec~11 (
	.dataa(\ram_a_not_b_vec[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\ram_a_not_b_vec~11_combout ),
	.cout());
defparam \ram_a_not_b_vec~11 .lut_mask = 16'hAAFF;
defparam \ram_a_not_b_vec~11 .sum_lutc_input = "datac";

dffeas \data_rdy_vec[7] (
	.clk(clk),
	.d(\data_rdy_vec~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_rdy_vec[7]~q ),
	.prn(vcc));
defparam \data_rdy_vec[7] .is_wysiwyg = "true";
defparam \data_rdy_vec[7] .power_up = "low";

cycloneiii_lcell_comb \data_rdy_vec~7 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~7_combout ),
	.cout());
defparam \data_rdy_vec~7 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_a_not_b_vec~12 (
	.dataa(\ram_a_not_b_vec[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\ram_a_not_b_vec~12_combout ),
	.cout());
defparam \ram_a_not_b_vec~12 .lut_mask = 16'hAAFF;
defparam \ram_a_not_b_vec~12 .sum_lutc_input = "datac";

dffeas \sw_r_tdl[0][0] (
	.clk(clk),
	.d(\rd_adgen|sw[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\sw_r_tdl[0][0]~q ),
	.prn(vcc));
defparam \sw_r_tdl[0][0] .is_wysiwyg = "true";
defparam \sw_r_tdl[0][0] .power_up = "low";

dffeas \sw_r_tdl[0][1] (
	.clk(clk),
	.d(\rd_adgen|sw[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\sw_r_tdl[0][1]~q ),
	.prn(vcc));
defparam \sw_r_tdl[0][1] .is_wysiwyg = "true";
defparam \sw_r_tdl[0][1] .power_up = "low";

dffeas \ram_a_not_b_vec[18] (
	.clk(clk),
	.d(\ram_a_not_b_vec~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\ram_a_not_b_vec[18]~q ),
	.prn(vcc));
defparam \ram_a_not_b_vec[18] .is_wysiwyg = "true";
defparam \ram_a_not_b_vec[18] .power_up = "low";

cycloneiii_lcell_comb \ram_a_not_b_vec~13 (
	.dataa(\ram_a_not_b_vec[18]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\ram_a_not_b_vec~13_combout ),
	.cout());
defparam \ram_a_not_b_vec~13 .lut_mask = 16'hAAFF;
defparam \ram_a_not_b_vec~13 .sum_lutc_input = "datac";

dffeas \p_tdl[7][2] (
	.clk(clk),
	.d(\p_tdl[6][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[7][2]~q ),
	.prn(vcc));
defparam \p_tdl[7][2] .is_wysiwyg = "true";
defparam \p_tdl[7][2] .power_up = "low";

dffeas \p_tdl[7][0] (
	.clk(clk),
	.d(\p_tdl[6][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[7][0]~q ),
	.prn(vcc));
defparam \p_tdl[7][0] .is_wysiwyg = "true";
defparam \p_tdl[7][0] .power_up = "low";

dffeas \p_tdl[7][1] (
	.clk(clk),
	.d(\p_tdl[6][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[7][1]~q ),
	.prn(vcc));
defparam \p_tdl[7][1] .is_wysiwyg = "true";
defparam \p_tdl[7][1] .power_up = "low";

dffeas \ram_a_not_b_vec[27] (
	.clk(clk),
	.d(\ram_a_not_b_vec~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\ram_a_not_b_vec[27]~q ),
	.prn(vcc));
defparam \ram_a_not_b_vec[27] .is_wysiwyg = "true";
defparam \ram_a_not_b_vec[27] .power_up = "low";

cycloneiii_lcell_comb \ram_a_not_b_vec~14 (
	.dataa(\ram_a_not_b_vec[27]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\ram_a_not_b_vec~14_combout ),
	.cout());
defparam \ram_a_not_b_vec~14 .lut_mask = 16'hAAFF;
defparam \ram_a_not_b_vec~14 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_a_not_b_vec~15 (
	.dataa(\writer|anb~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\ram_a_not_b_vec~15_combout ),
	.cout());
defparam \ram_a_not_b_vec~15 .lut_mask = 16'hAAFF;
defparam \ram_a_not_b_vec~15 .sum_lutc_input = "datac";

dffeas \data_imag_in_reg[2] (
	.clk(clk),
	.d(\data_imag_in_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_imag_in_reg[2]~q ),
	.prn(vcc));
defparam \data_imag_in_reg[2] .is_wysiwyg = "true";
defparam \data_imag_in_reg[2] .power_up = "low";

dffeas \data_real_in_reg[2] (
	.clk(clk),
	.d(\data_real_in_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_real_in_reg[2]~q ),
	.prn(vcc));
defparam \data_real_in_reg[2] .is_wysiwyg = "true";
defparam \data_real_in_reg[2] .power_up = "low";

cycloneiii_lcell_comb \core_real_in~0 (
	.dataa(\data_imag_in_reg[2]~q ),
	.datab(\data_real_in_reg[2]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_real_in~0_combout ),
	.cout());
defparam \core_real_in~0 .lut_mask = 16'hAACC;
defparam \core_real_in~0 .sum_lutc_input = "datac";

dffeas \ram_a_not_b_vec[5] (
	.clk(clk),
	.d(\ram_a_not_b_vec~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\ram_a_not_b_vec[5]~q ),
	.prn(vcc));
defparam \ram_a_not_b_vec[5] .is_wysiwyg = "true";
defparam \ram_a_not_b_vec[5] .power_up = "low";

cycloneiii_lcell_comb \ram_a_not_b_vec~16 (
	.dataa(\ram_a_not_b_vec[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\ram_a_not_b_vec~16_combout ),
	.cout());
defparam \ram_a_not_b_vec~16 .lut_mask = 16'hAAFF;
defparam \ram_a_not_b_vec~16 .sum_lutc_input = "datac";

dffeas \data_rdy_vec[6] (
	.clk(clk),
	.d(\data_rdy_vec~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_rdy_vec[6]~q ),
	.prn(vcc));
defparam \data_rdy_vec[6] .is_wysiwyg = "true";
defparam \data_rdy_vec[6] .power_up = "low";

cycloneiii_lcell_comb \data_rdy_vec~8 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~8_combout ),
	.cout());
defparam \data_rdy_vec~8 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~8 .sum_lutc_input = "datac";

dffeas \data_imag_in_reg[6] (
	.clk(clk),
	.d(\data_imag_in_reg~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_imag_in_reg[6]~q ),
	.prn(vcc));
defparam \data_imag_in_reg[6] .is_wysiwyg = "true";
defparam \data_imag_in_reg[6] .power_up = "low";

dffeas \data_real_in_reg[6] (
	.clk(clk),
	.d(\data_real_in_reg~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_real_in_reg[6]~q ),
	.prn(vcc));
defparam \data_real_in_reg[6] .is_wysiwyg = "true";
defparam \data_real_in_reg[6] .power_up = "low";

cycloneiii_lcell_comb \core_real_in~1 (
	.dataa(\data_imag_in_reg[6]~q ),
	.datab(\data_real_in_reg[6]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_real_in~1_combout ),
	.cout());
defparam \core_real_in~1 .lut_mask = 16'hAACC;
defparam \core_real_in~1 .sum_lutc_input = "datac";

dffeas \data_imag_in_reg[4] (
	.clk(clk),
	.d(\data_imag_in_reg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_imag_in_reg[4]~q ),
	.prn(vcc));
defparam \data_imag_in_reg[4] .is_wysiwyg = "true";
defparam \data_imag_in_reg[4] .power_up = "low";

dffeas \data_real_in_reg[4] (
	.clk(clk),
	.d(\data_real_in_reg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_real_in_reg[4]~q ),
	.prn(vcc));
defparam \data_real_in_reg[4] .is_wysiwyg = "true";
defparam \data_real_in_reg[4] .power_up = "low";

cycloneiii_lcell_comb \core_real_in~2 (
	.dataa(\data_imag_in_reg[4]~q ),
	.datab(\data_real_in_reg[4]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_real_in~2_combout ),
	.cout());
defparam \core_real_in~2 .lut_mask = 16'hAACC;
defparam \core_real_in~2 .sum_lutc_input = "datac";

dffeas \data_imag_in_reg[3] (
	.clk(clk),
	.d(\data_imag_in_reg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_imag_in_reg[3]~q ),
	.prn(vcc));
defparam \data_imag_in_reg[3] .is_wysiwyg = "true";
defparam \data_imag_in_reg[3] .power_up = "low";

dffeas \data_real_in_reg[3] (
	.clk(clk),
	.d(\data_real_in_reg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_real_in_reg[3]~q ),
	.prn(vcc));
defparam \data_real_in_reg[3] .is_wysiwyg = "true";
defparam \data_real_in_reg[3] .power_up = "low";

cycloneiii_lcell_comb \core_real_in~3 (
	.dataa(\data_imag_in_reg[3]~q ),
	.datab(\data_real_in_reg[3]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_real_in~3_combout ),
	.cout());
defparam \core_real_in~3 .lut_mask = 16'hAACC;
defparam \core_real_in~3 .sum_lutc_input = "datac";

dffeas \data_imag_in_reg[5] (
	.clk(clk),
	.d(\data_imag_in_reg~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_imag_in_reg[5]~q ),
	.prn(vcc));
defparam \data_imag_in_reg[5] .is_wysiwyg = "true";
defparam \data_imag_in_reg[5] .power_up = "low";

dffeas \data_real_in_reg[5] (
	.clk(clk),
	.d(\data_real_in_reg~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_real_in_reg[5]~q ),
	.prn(vcc));
defparam \data_real_in_reg[5] .is_wysiwyg = "true";
defparam \data_real_in_reg[5] .power_up = "low";

cycloneiii_lcell_comb \core_real_in~4 (
	.dataa(\data_imag_in_reg[5]~q ),
	.datab(\data_real_in_reg[5]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_real_in~4_combout ),
	.cout());
defparam \core_real_in~4 .lut_mask = 16'hAACC;
defparam \core_real_in~4 .sum_lutc_input = "datac";

dffeas \data_imag_in_reg[1] (
	.clk(clk),
	.d(\data_imag_in_reg~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_imag_in_reg[1]~q ),
	.prn(vcc));
defparam \data_imag_in_reg[1] .is_wysiwyg = "true";
defparam \data_imag_in_reg[1] .power_up = "low";

dffeas \data_real_in_reg[1] (
	.clk(clk),
	.d(\data_real_in_reg~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_real_in_reg[1]~q ),
	.prn(vcc));
defparam \data_real_in_reg[1] .is_wysiwyg = "true";
defparam \data_real_in_reg[1] .power_up = "low";

cycloneiii_lcell_comb \core_real_in~5 (
	.dataa(\data_imag_in_reg[1]~q ),
	.datab(\data_real_in_reg[1]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_real_in~5_combout ),
	.cout());
defparam \core_real_in~5 .lut_mask = 16'hAACC;
defparam \core_real_in~5 .sum_lutc_input = "datac";

dffeas \data_imag_in_reg[0] (
	.clk(clk),
	.d(\data_imag_in_reg~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_imag_in_reg[0]~q ),
	.prn(vcc));
defparam \data_imag_in_reg[0] .is_wysiwyg = "true";
defparam \data_imag_in_reg[0] .power_up = "low";

dffeas \data_real_in_reg[0] (
	.clk(clk),
	.d(\data_real_in_reg~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_real_in_reg[0]~q ),
	.prn(vcc));
defparam \data_real_in_reg[0] .is_wysiwyg = "true";
defparam \data_real_in_reg[0] .power_up = "low";

cycloneiii_lcell_comb \core_real_in~6 (
	.dataa(\data_imag_in_reg[0]~q ),
	.datab(\data_real_in_reg[0]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_real_in~6_combout ),
	.cout());
defparam \core_real_in~6 .lut_mask = 16'hAACC;
defparam \core_real_in~6 .sum_lutc_input = "datac";

dffeas \data_imag_in_reg[7] (
	.clk(clk),
	.d(\data_imag_in_reg~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_imag_in_reg[7]~q ),
	.prn(vcc));
defparam \data_imag_in_reg[7] .is_wysiwyg = "true";
defparam \data_imag_in_reg[7] .power_up = "low";

dffeas \data_real_in_reg[7] (
	.clk(clk),
	.d(\data_real_in_reg~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_real_in_reg[7]~q ),
	.prn(vcc));
defparam \data_real_in_reg[7] .is_wysiwyg = "true";
defparam \data_real_in_reg[7] .power_up = "low";

cycloneiii_lcell_comb \core_real_in~7 (
	.dataa(\data_imag_in_reg[7]~q ),
	.datab(\data_real_in_reg[7]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_real_in~7_combout ),
	.cout());
defparam \core_real_in~7 .lut_mask = 16'hAACC;
defparam \core_real_in~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \core_imag_in~0 (
	.dataa(\data_real_in_reg[7]~q ),
	.datab(\data_imag_in_reg[7]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_imag_in~0_combout ),
	.cout());
defparam \core_imag_in~0 .lut_mask = 16'hAACC;
defparam \core_imag_in~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \core_imag_in~1 (
	.dataa(\data_real_in_reg[3]~q ),
	.datab(\data_imag_in_reg[3]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_imag_in~1_combout ),
	.cout());
defparam \core_imag_in~1 .lut_mask = 16'hAACC;
defparam \core_imag_in~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \core_imag_in~2 (
	.dataa(\data_real_in_reg[5]~q ),
	.datab(\data_imag_in_reg[5]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_imag_in~2_combout ),
	.cout());
defparam \core_imag_in~2 .lut_mask = 16'hAACC;
defparam \core_imag_in~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \core_imag_in~3 (
	.dataa(\data_real_in_reg[4]~q ),
	.datab(\data_imag_in_reg[4]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_imag_in~3_combout ),
	.cout());
defparam \core_imag_in~3 .lut_mask = 16'hAACC;
defparam \core_imag_in~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \core_imag_in~4 (
	.dataa(\data_real_in_reg[6]~q ),
	.datab(\data_imag_in_reg[6]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_imag_in~4_combout ),
	.cout());
defparam \core_imag_in~4 .lut_mask = 16'hAACC;
defparam \core_imag_in~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \core_imag_in~5 (
	.dataa(\data_real_in_reg[2]~q ),
	.datab(\data_imag_in_reg[2]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_imag_in~5_combout ),
	.cout());
defparam \core_imag_in~5 .lut_mask = 16'hAACC;
defparam \core_imag_in~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \core_imag_in~6 (
	.dataa(\data_real_in_reg[1]~q ),
	.datab(\data_imag_in_reg[1]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_imag_in~6_combout ),
	.cout());
defparam \core_imag_in~6 .lut_mask = 16'hAACC;
defparam \core_imag_in~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \core_imag_in~7 (
	.dataa(\data_real_in_reg[0]~q ),
	.datab(\data_imag_in_reg[0]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_imag_in~7_combout ),
	.cout());
defparam \core_imag_in~7 .lut_mask = 16'hAACC;
defparam \core_imag_in~7 .sum_lutc_input = "datac";

dffeas \ram_a_not_b_vec[17] (
	.clk(clk),
	.d(\ram_a_not_b_vec~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\ram_a_not_b_vec[17]~q ),
	.prn(vcc));
defparam \ram_a_not_b_vec[17] .is_wysiwyg = "true";
defparam \ram_a_not_b_vec[17] .power_up = "low";

cycloneiii_lcell_comb \ram_a_not_b_vec~17 (
	.dataa(\ram_a_not_b_vec[17]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\ram_a_not_b_vec~17_combout ),
	.cout());
defparam \ram_a_not_b_vec~17 .lut_mask = 16'hAAFF;
defparam \ram_a_not_b_vec~17 .sum_lutc_input = "datac";

dffeas \p_tdl[6][2] (
	.clk(clk),
	.d(\p_tdl[5][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[6][2]~q ),
	.prn(vcc));
defparam \p_tdl[6][2] .is_wysiwyg = "true";
defparam \p_tdl[6][2] .power_up = "low";

dffeas \p_tdl[6][0] (
	.clk(clk),
	.d(\p_tdl[5][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[6][0]~q ),
	.prn(vcc));
defparam \p_tdl[6][0] .is_wysiwyg = "true";
defparam \p_tdl[6][0] .power_up = "low";

dffeas \p_tdl[6][1] (
	.clk(clk),
	.d(\p_tdl[5][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[6][1]~q ),
	.prn(vcc));
defparam \p_tdl[6][1] .is_wysiwyg = "true";
defparam \p_tdl[6][1] .power_up = "low";

cycloneiii_lcell_comb \ram_a_not_b_vec~18 (
	.dataa(\ram_a_not_b_vec[26]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\ram_a_not_b_vec~18_combout ),
	.cout());
defparam \ram_a_not_b_vec~18 .lut_mask = 16'hAAFF;
defparam \ram_a_not_b_vec~18 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \data_imag_in_reg~0 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_imag_in_reg~0_combout ),
	.cout());
defparam \data_imag_in_reg~0 .lut_mask = 16'hEEEE;
defparam \data_imag_in_reg~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \data_real_in_reg~0 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[10] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_real_in_reg~0_combout ),
	.cout());
defparam \data_real_in_reg~0 .lut_mask = 16'hEEEE;
defparam \data_real_in_reg~0 .sum_lutc_input = "datac";

dffeas \ram_a_not_b_vec[4] (
	.clk(clk),
	.d(\ram_a_not_b_vec~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\ram_a_not_b_vec[4]~q ),
	.prn(vcc));
defparam \ram_a_not_b_vec[4] .is_wysiwyg = "true";
defparam \ram_a_not_b_vec[4] .power_up = "low";

cycloneiii_lcell_comb \ram_a_not_b_vec~19 (
	.dataa(\ram_a_not_b_vec[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\ram_a_not_b_vec~19_combout ),
	.cout());
defparam \ram_a_not_b_vec~19 .lut_mask = 16'hAAFF;
defparam \ram_a_not_b_vec~19 .sum_lutc_input = "datac";

dffeas \data_rdy_vec[5] (
	.clk(clk),
	.d(\data_rdy_vec~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_rdy_vec[5]~q ),
	.prn(vcc));
defparam \data_rdy_vec[5] .is_wysiwyg = "true";
defparam \data_rdy_vec[5] .power_up = "low";

cycloneiii_lcell_comb \data_rdy_vec~9 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~9_combout ),
	.cout());
defparam \data_rdy_vec~9 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \data_imag_in_reg~1 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_imag_in_reg~1_combout ),
	.cout());
defparam \data_imag_in_reg~1 .lut_mask = 16'hEEEE;
defparam \data_imag_in_reg~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \data_real_in_reg~1 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[14] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_real_in_reg~1_combout ),
	.cout());
defparam \data_real_in_reg~1 .lut_mask = 16'hEEEE;
defparam \data_real_in_reg~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \data_imag_in_reg~2 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_imag_in_reg~2_combout ),
	.cout());
defparam \data_imag_in_reg~2 .lut_mask = 16'hEEEE;
defparam \data_imag_in_reg~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \data_real_in_reg~2 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[12] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_real_in_reg~2_combout ),
	.cout());
defparam \data_real_in_reg~2 .lut_mask = 16'hEEEE;
defparam \data_real_in_reg~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \data_imag_in_reg~3 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_imag_in_reg~3_combout ),
	.cout());
defparam \data_imag_in_reg~3 .lut_mask = 16'hEEEE;
defparam \data_imag_in_reg~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \data_real_in_reg~3 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[11] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_real_in_reg~3_combout ),
	.cout());
defparam \data_real_in_reg~3 .lut_mask = 16'hEEEE;
defparam \data_real_in_reg~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \data_imag_in_reg~4 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_imag_in_reg~4_combout ),
	.cout());
defparam \data_imag_in_reg~4 .lut_mask = 16'hEEEE;
defparam \data_imag_in_reg~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \data_real_in_reg~4 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[13] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_real_in_reg~4_combout ),
	.cout());
defparam \data_real_in_reg~4 .lut_mask = 16'hEEEE;
defparam \data_real_in_reg~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \data_imag_in_reg~5 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_imag_in_reg~5_combout ),
	.cout());
defparam \data_imag_in_reg~5 .lut_mask = 16'hEEEE;
defparam \data_imag_in_reg~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \data_real_in_reg~5 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[9] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_real_in_reg~5_combout ),
	.cout());
defparam \data_real_in_reg~5 .lut_mask = 16'hEEEE;
defparam \data_real_in_reg~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \data_imag_in_reg~6 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_imag_in_reg~6_combout ),
	.cout());
defparam \data_imag_in_reg~6 .lut_mask = 16'hEEEE;
defparam \data_imag_in_reg~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \data_real_in_reg~6 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[8] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_real_in_reg~6_combout ),
	.cout());
defparam \data_real_in_reg~6 .lut_mask = 16'hEEEE;
defparam \data_real_in_reg~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \data_imag_in_reg~7 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_imag_in_reg~7_combout ),
	.cout());
defparam \data_imag_in_reg~7 .lut_mask = 16'hEEEE;
defparam \data_imag_in_reg~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \data_real_in_reg~7 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[15] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_real_in_reg~7_combout ),
	.cout());
defparam \data_real_in_reg~7 .lut_mask = 16'hEEEE;
defparam \data_real_in_reg~7 .sum_lutc_input = "datac";

dffeas \ram_a_not_b_vec[16] (
	.clk(clk),
	.d(\ram_a_not_b_vec~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\ram_a_not_b_vec[16]~q ),
	.prn(vcc));
defparam \ram_a_not_b_vec[16] .is_wysiwyg = "true";
defparam \ram_a_not_b_vec[16] .power_up = "low";

cycloneiii_lcell_comb \ram_a_not_b_vec~20 (
	.dataa(\ram_a_not_b_vec[16]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\ram_a_not_b_vec~20_combout ),
	.cout());
defparam \ram_a_not_b_vec~20 .lut_mask = 16'hAAFF;
defparam \ram_a_not_b_vec~20 .sum_lutc_input = "datac";

dffeas \p_tdl[5][2] (
	.clk(clk),
	.d(\p_tdl[4][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[5][2]~q ),
	.prn(vcc));
defparam \p_tdl[5][2] .is_wysiwyg = "true";
defparam \p_tdl[5][2] .power_up = "low";

dffeas \p_tdl[5][0] (
	.clk(clk),
	.d(\p_tdl[4][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[5][0]~q ),
	.prn(vcc));
defparam \p_tdl[5][0] .is_wysiwyg = "true";
defparam \p_tdl[5][0] .power_up = "low";

dffeas \p_tdl[5][1] (
	.clk(clk),
	.d(\p_tdl[4][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[5][1]~q ),
	.prn(vcc));
defparam \p_tdl[5][1] .is_wysiwyg = "true";
defparam \p_tdl[5][1] .power_up = "low";

dffeas \ram_a_not_b_vec[3] (
	.clk(clk),
	.d(\ram_a_not_b_vec~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\ram_a_not_b_vec[3]~q ),
	.prn(vcc));
defparam \ram_a_not_b_vec[3] .is_wysiwyg = "true";
defparam \ram_a_not_b_vec[3] .power_up = "low";

cycloneiii_lcell_comb \ram_a_not_b_vec~21 (
	.dataa(\ram_a_not_b_vec[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\ram_a_not_b_vec~21_combout ),
	.cout());
defparam \ram_a_not_b_vec~21 .lut_mask = 16'hAAFF;
defparam \ram_a_not_b_vec~21 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \data_rdy_vec~10 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~10_combout ),
	.cout());
defparam \data_rdy_vec~10 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~10 .sum_lutc_input = "datac";

dffeas \ram_a_not_b_vec[15] (
	.clk(clk),
	.d(\ram_a_not_b_vec~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\ram_a_not_b_vec[15]~q ),
	.prn(vcc));
defparam \ram_a_not_b_vec[15] .is_wysiwyg = "true";
defparam \ram_a_not_b_vec[15] .power_up = "low";

cycloneiii_lcell_comb \ram_a_not_b_vec~22 (
	.dataa(\ram_a_not_b_vec[15]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\ram_a_not_b_vec~22_combout ),
	.cout());
defparam \ram_a_not_b_vec~22 .lut_mask = 16'hAAFF;
defparam \ram_a_not_b_vec~22 .sum_lutc_input = "datac";

dffeas \p_tdl[4][2] (
	.clk(clk),
	.d(\p_tdl[3][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[4][2]~q ),
	.prn(vcc));
defparam \p_tdl[4][2] .is_wysiwyg = "true";
defparam \p_tdl[4][2] .power_up = "low";

dffeas \p_tdl[4][0] (
	.clk(clk),
	.d(\p_tdl[3][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[4][0]~q ),
	.prn(vcc));
defparam \p_tdl[4][0] .is_wysiwyg = "true";
defparam \p_tdl[4][0] .power_up = "low";

dffeas \p_tdl[4][1] (
	.clk(clk),
	.d(\p_tdl[3][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[4][1]~q ),
	.prn(vcc));
defparam \p_tdl[4][1] .is_wysiwyg = "true";
defparam \p_tdl[4][1] .power_up = "low";

dffeas \ram_a_not_b_vec[2] (
	.clk(clk),
	.d(\ram_a_not_b_vec~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\ram_a_not_b_vec[2]~q ),
	.prn(vcc));
defparam \ram_a_not_b_vec[2] .is_wysiwyg = "true";
defparam \ram_a_not_b_vec[2] .power_up = "low";

cycloneiii_lcell_comb \ram_a_not_b_vec~23 (
	.dataa(\ram_a_not_b_vec[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\ram_a_not_b_vec~23_combout ),
	.cout());
defparam \ram_a_not_b_vec~23 .lut_mask = 16'hAAFF;
defparam \ram_a_not_b_vec~23 .sum_lutc_input = "datac";

dffeas \ram_a_not_b_vec[14] (
	.clk(clk),
	.d(\ram_a_not_b_vec~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\ram_a_not_b_vec[14]~q ),
	.prn(vcc));
defparam \ram_a_not_b_vec[14] .is_wysiwyg = "true";
defparam \ram_a_not_b_vec[14] .power_up = "low";

cycloneiii_lcell_comb \ram_a_not_b_vec~24 (
	.dataa(\ram_a_not_b_vec[14]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\ram_a_not_b_vec~24_combout ),
	.cout());
defparam \ram_a_not_b_vec~24 .lut_mask = 16'hAAFF;
defparam \ram_a_not_b_vec~24 .sum_lutc_input = "datac";

dffeas \p_tdl[3][2] (
	.clk(clk),
	.d(\p_tdl[2][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[3][2]~q ),
	.prn(vcc));
defparam \p_tdl[3][2] .is_wysiwyg = "true";
defparam \p_tdl[3][2] .power_up = "low";

dffeas \p_tdl[3][0] (
	.clk(clk),
	.d(\p_tdl[2][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[3][0]~q ),
	.prn(vcc));
defparam \p_tdl[3][0] .is_wysiwyg = "true";
defparam \p_tdl[3][0] .power_up = "low";

dffeas \p_tdl[3][1] (
	.clk(clk),
	.d(\p_tdl[2][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[3][1]~q ),
	.prn(vcc));
defparam \p_tdl[3][1] .is_wysiwyg = "true";
defparam \p_tdl[3][1] .power_up = "low";

cycloneiii_lcell_comb \ram_a_not_b_vec~25 (
	.dataa(\ram_a_not_b_vec[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\ram_a_not_b_vec~25_combout ),
	.cout());
defparam \ram_a_not_b_vec~25 .lut_mask = 16'hAAFF;
defparam \ram_a_not_b_vec~25 .sum_lutc_input = "datac";

dffeas \ram_a_not_b_vec[13] (
	.clk(clk),
	.d(\ram_a_not_b_vec~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\ram_a_not_b_vec[13]~q ),
	.prn(vcc));
defparam \ram_a_not_b_vec[13] .is_wysiwyg = "true";
defparam \ram_a_not_b_vec[13] .power_up = "low";

cycloneiii_lcell_comb \ram_a_not_b_vec~26 (
	.dataa(\ram_a_not_b_vec[13]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\ram_a_not_b_vec~26_combout ),
	.cout());
defparam \ram_a_not_b_vec~26 .lut_mask = 16'hAAFF;
defparam \ram_a_not_b_vec~26 .sum_lutc_input = "datac";

dffeas \p_tdl[2][2] (
	.clk(clk),
	.d(\p_tdl[1][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[2][2]~q ),
	.prn(vcc));
defparam \p_tdl[2][2] .is_wysiwyg = "true";
defparam \p_tdl[2][2] .power_up = "low";

dffeas \p_tdl[2][0] (
	.clk(clk),
	.d(\p_tdl[1][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[2][0]~q ),
	.prn(vcc));
defparam \p_tdl[2][0] .is_wysiwyg = "true";
defparam \p_tdl[2][0] .power_up = "low";

dffeas \p_tdl[2][1] (
	.clk(clk),
	.d(\p_tdl[1][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[2][1]~q ),
	.prn(vcc));
defparam \p_tdl[2][1] .is_wysiwyg = "true";
defparam \p_tdl[2][1] .power_up = "low";

dffeas \ram_a_not_b_vec[12] (
	.clk(clk),
	.d(\ram_a_not_b_vec~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\ram_a_not_b_vec[12]~q ),
	.prn(vcc));
defparam \ram_a_not_b_vec[12] .is_wysiwyg = "true";
defparam \ram_a_not_b_vec[12] .power_up = "low";

cycloneiii_lcell_comb \ram_a_not_b_vec~27 (
	.dataa(\ram_a_not_b_vec[12]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\ram_a_not_b_vec~27_combout ),
	.cout());
defparam \ram_a_not_b_vec~27 .lut_mask = 16'hAAFF;
defparam \ram_a_not_b_vec~27 .sum_lutc_input = "datac";

dffeas \p_tdl[1][2] (
	.clk(clk),
	.d(\p_tdl[0][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[1][2]~q ),
	.prn(vcc));
defparam \p_tdl[1][2] .is_wysiwyg = "true";
defparam \p_tdl[1][2] .power_up = "low";

dffeas \p_tdl[1][0] (
	.clk(clk),
	.d(\p_tdl[0][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[1][0]~q ),
	.prn(vcc));
defparam \p_tdl[1][0] .is_wysiwyg = "true";
defparam \p_tdl[1][0] .power_up = "low";

dffeas \p_tdl[1][1] (
	.clk(clk),
	.d(\p_tdl[0][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[1][1]~q ),
	.prn(vcc));
defparam \p_tdl[1][1] .is_wysiwyg = "true";
defparam \p_tdl[1][1] .power_up = "low";

dffeas \ram_a_not_b_vec[11] (
	.clk(clk),
	.d(\ram_a_not_b_vec~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\ram_a_not_b_vec[11]~q ),
	.prn(vcc));
defparam \ram_a_not_b_vec[11] .is_wysiwyg = "true";
defparam \ram_a_not_b_vec[11] .power_up = "low";

cycloneiii_lcell_comb \ram_a_not_b_vec~28 (
	.dataa(\ram_a_not_b_vec[11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\ram_a_not_b_vec~28_combout ),
	.cout());
defparam \ram_a_not_b_vec~28 .lut_mask = 16'hAAFF;
defparam \ram_a_not_b_vec~28 .sum_lutc_input = "datac";

dffeas \p_tdl[0][2] (
	.clk(clk),
	.d(\gen_gt256_mk:ctrl|p[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[0][2]~q ),
	.prn(vcc));
defparam \p_tdl[0][2] .is_wysiwyg = "true";
defparam \p_tdl[0][2] .power_up = "low";

dffeas \p_tdl[0][0] (
	.clk(clk),
	.d(\gen_gt256_mk:ctrl|p[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[0][0]~q ),
	.prn(vcc));
defparam \p_tdl[0][0] .is_wysiwyg = "true";
defparam \p_tdl[0][0] .power_up = "low";

dffeas \p_tdl[0][1] (
	.clk(clk),
	.d(\gen_gt256_mk:ctrl|p[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[0][1]~q ),
	.prn(vcc));
defparam \p_tdl[0][1] .is_wysiwyg = "true";
defparam \p_tdl[0][1] .power_up = "low";

cycloneiii_lcell_comb \ram_a_not_b_vec~29 (
	.dataa(\ram_a_not_b_vec[10]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\ram_a_not_b_vec~29_combout ),
	.cout());
defparam \ram_a_not_b_vec~29 .lut_mask = 16'hAAFF;
defparam \ram_a_not_b_vec~29 .sum_lutc_input = "datac";

endmodule

module fft_asj_fft_3dp_rom_fft_120 (
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_3,
	q_a_4,
	q_a_5,
	q_a_6,
	q_a_7,
	q_a_01,
	q_a_11,
	q_a_21,
	q_a_31,
	q_a_41,
	q_a_51,
	q_a_61,
	q_a_71,
	q_a_02,
	q_a_12,
	q_a_22,
	q_a_32,
	q_a_42,
	q_a_52,
	q_a_62,
	q_a_72,
	q_a_03,
	q_a_13,
	q_a_23,
	q_a_33,
	q_a_43,
	q_a_53,
	q_a_63,
	q_a_73,
	q_a_04,
	q_a_14,
	q_a_24,
	q_a_34,
	q_a_44,
	q_a_54,
	q_a_64,
	q_a_74,
	q_a_05,
	q_a_15,
	q_a_25,
	q_a_35,
	q_a_45,
	q_a_55,
	q_a_65,
	q_a_75,
	global_clock_enable,
	twad_tdl_0_6,
	twad_tdl_1_6,
	twad_tdl_2_6,
	twad_tdl_3_6,
	twad_tdl_4_6,
	twad_tdl_5_6,
	twad_tdl_6_6,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_a_0;
output 	q_a_1;
output 	q_a_2;
output 	q_a_3;
output 	q_a_4;
output 	q_a_5;
output 	q_a_6;
output 	q_a_7;
output 	q_a_01;
output 	q_a_11;
output 	q_a_21;
output 	q_a_31;
output 	q_a_41;
output 	q_a_51;
output 	q_a_61;
output 	q_a_71;
output 	q_a_02;
output 	q_a_12;
output 	q_a_22;
output 	q_a_32;
output 	q_a_42;
output 	q_a_52;
output 	q_a_62;
output 	q_a_72;
output 	q_a_03;
output 	q_a_13;
output 	q_a_23;
output 	q_a_33;
output 	q_a_43;
output 	q_a_53;
output 	q_a_63;
output 	q_a_73;
output 	q_a_04;
output 	q_a_14;
output 	q_a_24;
output 	q_a_34;
output 	q_a_44;
output 	q_a_54;
output 	q_a_64;
output 	q_a_74;
output 	q_a_05;
output 	q_a_15;
output 	q_a_25;
output 	q_a_35;
output 	q_a_45;
output 	q_a_55;
output 	q_a_65;
output 	q_a_75;
input 	global_clock_enable;
input 	twad_tdl_0_6;
input 	twad_tdl_1_6;
input 	twad_tdl_2_6;
input 	twad_tdl_3_6;
input 	twad_tdl_4_6;
input 	twad_tdl_5_6;
input 	twad_tdl_6_6;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_twid_rom_fft_120_2 \gen_M4K:cos_3n (
	.q_a_0(q_a_04),
	.q_a_1(q_a_14),
	.q_a_2(q_a_24),
	.q_a_3(q_a_34),
	.q_a_4(q_a_44),
	.q_a_5(q_a_54),
	.q_a_6(q_a_64),
	.q_a_7(q_a_74),
	.global_clock_enable(global_clock_enable),
	.twad_tdl_0_6(twad_tdl_0_6),
	.twad_tdl_1_6(twad_tdl_1_6),
	.twad_tdl_2_6(twad_tdl_2_6),
	.twad_tdl_3_6(twad_tdl_3_6),
	.twad_tdl_4_6(twad_tdl_4_6),
	.twad_tdl_5_6(twad_tdl_5_6),
	.twad_tdl_6_6(twad_tdl_6_6),
	.clk(clk));

fft_twid_rom_fft_120_1 \gen_M4K:cos_2n (
	.q_a_0(q_a_02),
	.q_a_1(q_a_12),
	.q_a_2(q_a_22),
	.q_a_3(q_a_32),
	.q_a_4(q_a_42),
	.q_a_5(q_a_52),
	.q_a_6(q_a_62),
	.q_a_7(q_a_72),
	.global_clock_enable(global_clock_enable),
	.twad_tdl_0_6(twad_tdl_0_6),
	.twad_tdl_1_6(twad_tdl_1_6),
	.twad_tdl_2_6(twad_tdl_2_6),
	.twad_tdl_3_6(twad_tdl_3_6),
	.twad_tdl_4_6(twad_tdl_4_6),
	.twad_tdl_5_6(twad_tdl_5_6),
	.twad_tdl_6_6(twad_tdl_6_6),
	.clk(clk));

fft_twid_rom_fft_120 \gen_M4K:cos_1n (
	.q_a_0(q_a_0),
	.q_a_1(q_a_1),
	.q_a_2(q_a_2),
	.q_a_3(q_a_3),
	.q_a_4(q_a_4),
	.q_a_5(q_a_5),
	.q_a_6(q_a_6),
	.q_a_7(q_a_7),
	.global_clock_enable(global_clock_enable),
	.twad_tdl_0_6(twad_tdl_0_6),
	.twad_tdl_1_6(twad_tdl_1_6),
	.twad_tdl_2_6(twad_tdl_2_6),
	.twad_tdl_3_6(twad_tdl_3_6),
	.twad_tdl_4_6(twad_tdl_4_6),
	.twad_tdl_5_6(twad_tdl_5_6),
	.twad_tdl_6_6(twad_tdl_6_6),
	.clk(clk));

fft_twid_rom_fft_120_5 \gen_M4K:sin_3n (
	.q_a_0(q_a_05),
	.q_a_1(q_a_15),
	.q_a_2(q_a_25),
	.q_a_3(q_a_35),
	.q_a_4(q_a_45),
	.q_a_5(q_a_55),
	.q_a_6(q_a_65),
	.q_a_7(q_a_75),
	.global_clock_enable(global_clock_enable),
	.twad_tdl_0_6(twad_tdl_0_6),
	.twad_tdl_1_6(twad_tdl_1_6),
	.twad_tdl_2_6(twad_tdl_2_6),
	.twad_tdl_3_6(twad_tdl_3_6),
	.twad_tdl_4_6(twad_tdl_4_6),
	.twad_tdl_5_6(twad_tdl_5_6),
	.twad_tdl_6_6(twad_tdl_6_6),
	.clk(clk));

fft_twid_rom_fft_120_4 \gen_M4K:sin_2n (
	.q_a_0(q_a_03),
	.q_a_1(q_a_13),
	.q_a_2(q_a_23),
	.q_a_3(q_a_33),
	.q_a_4(q_a_43),
	.q_a_5(q_a_53),
	.q_a_6(q_a_63),
	.q_a_7(q_a_73),
	.global_clock_enable(global_clock_enable),
	.twad_tdl_0_6(twad_tdl_0_6),
	.twad_tdl_1_6(twad_tdl_1_6),
	.twad_tdl_2_6(twad_tdl_2_6),
	.twad_tdl_3_6(twad_tdl_3_6),
	.twad_tdl_4_6(twad_tdl_4_6),
	.twad_tdl_5_6(twad_tdl_5_6),
	.twad_tdl_6_6(twad_tdl_6_6),
	.clk(clk));

fft_twid_rom_fft_120_3 \gen_M4K:sin_1n (
	.q_a_0(q_a_01),
	.q_a_1(q_a_11),
	.q_a_2(q_a_21),
	.q_a_3(q_a_31),
	.q_a_4(q_a_41),
	.q_a_5(q_a_51),
	.q_a_6(q_a_61),
	.q_a_7(q_a_71),
	.global_clock_enable(global_clock_enable),
	.twad_tdl_0_6(twad_tdl_0_6),
	.twad_tdl_1_6(twad_tdl_1_6),
	.twad_tdl_2_6(twad_tdl_2_6),
	.twad_tdl_3_6(twad_tdl_3_6),
	.twad_tdl_4_6(twad_tdl_4_6),
	.twad_tdl_5_6(twad_tdl_5_6),
	.twad_tdl_6_6(twad_tdl_6_6),
	.clk(clk));

endmodule

module fft_twid_rom_fft_120 (
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_3,
	q_a_4,
	q_a_5,
	q_a_6,
	q_a_7,
	global_clock_enable,
	twad_tdl_0_6,
	twad_tdl_1_6,
	twad_tdl_2_6,
	twad_tdl_3_6,
	twad_tdl_4_6,
	twad_tdl_5_6,
	twad_tdl_6_6,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_a_0;
output 	q_a_1;
output 	q_a_2;
output 	q_a_3;
output 	q_a_4;
output 	q_a_5;
output 	q_a_6;
output 	q_a_7;
input 	global_clock_enable;
input 	twad_tdl_0_6;
input 	twad_tdl_1_6;
input 	twad_tdl_2_6;
input 	twad_tdl_3_6;
input 	twad_tdl_4_6;
input 	twad_tdl_5_6;
input 	twad_tdl_6_6;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_altsyncram_1 \gen_auto:altsyncram_component (
	.q_a({q_a_unconnected_wire_15,q_a_unconnected_wire_14,q_a_unconnected_wire_13,q_a_unconnected_wire_12,q_a_unconnected_wire_11,q_a_unconnected_wire_10,q_a_unconnected_wire_9,q_a_unconnected_wire_8,q_a_7,q_a_6,q_a_5,q_a_4,q_a_3,q_a_2,q_a_1,q_a_0}),
	.clocken0(global_clock_enable),
	.address_a({twad_tdl_6_6,twad_tdl_5_6,twad_tdl_4_6,twad_tdl_3_6,twad_tdl_2_6,twad_tdl_1_6,twad_tdl_0_6}),
	.clock0(clk));

endmodule

module fft_altsyncram_1 (
	q_a,
	clocken0,
	address_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_a;
input 	clocken0;
input 	[6:0] address_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_altsyncram_b191 auto_generated(
	.q_a({q_a[7],q_a[6],q_a[5],q_a[4],q_a[3],q_a[2],q_a[1],q_a[0]}),
	.clocken0(clocken0),
	.address_a({address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.clock0(clock0));

endmodule

module fft_altsyncram_b191 (
	q_a,
	clocken0,
	address_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q_a;
input 	clocken0;
input 	[6:0] address_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTADATAOUT_bus;
wire [143:0] ram_block1a1_PORTADATAOUT_bus;
wire [143:0] ram_block1a2_PORTADATAOUT_bus;
wire [143:0] ram_block1a3_PORTADATAOUT_bus;
wire [143:0] ram_block1a4_PORTADATAOUT_bus;
wire [143:0] ram_block1a5_PORTADATAOUT_bus;
wire [143:0] ram_block1a6_PORTADATAOUT_bus;
wire [143:0] ram_block1a7_PORTADATAOUT_bus;

assign q_a[0] = ram_block1a0_PORTADATAOUT_bus[0];

assign q_a[1] = ram_block1a1_PORTADATAOUT_bus[0];

assign q_a[2] = ram_block1a2_PORTADATAOUT_bus[0];

assign q_a[3] = ram_block1a3_PORTADATAOUT_bus[0];

assign q_a[4] = ram_block1a4_PORTADATAOUT_bus[0];

assign q_a[5] = ram_block1a5_PORTADATAOUT_bus[0];

assign q_a[6] = ram_block1a6_PORTADATAOUT_bus[0];

assign q_a[7] = ram_block1a7_PORTADATAOUT_bus[0];

cycloneiii_ram_block ram_block1a0(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a0_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.init_file = "fft_1n512cos.hex";
defparam ram_block1a0.init_file_layout = "port_a";
defparam ram_block1a0.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_3dp_rom_fft_120:twrom|twid_rom_fft_120:\\gen_M4K:cos_1n|altsyncram:\\gen_auto:altsyncram_component|altsyncram_b191:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.operation_mode = "rom";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 7;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "clock0";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 127;
defparam ram_block1a0.port_a_logical_ram_depth = 128;
defparam ram_block1a0.port_a_logical_ram_width = 8;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.ram_block_type = "auto";
defparam ram_block1a0.mem_init0 = 128'h6633333364DB4B52AAAA56DB2631E0FF;

cycloneiii_ram_block ram_block1a1(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a1_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.init_file = "fft_1n512cos.hex";
defparam ram_block1a1.init_file_layout = "port_a";
defparam ram_block1a1.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_3dp_rom_fft_120:twrom|twid_rom_fft_120:\\gen_M4K:cos_1n|altsyncram:\\gen_auto:altsyncram_component|altsyncram_b191:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.operation_mode = "rom";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 7;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "clock0";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 127;
defparam ram_block1a1.port_a_logical_ram_depth = 128;
defparam ram_block1a1.port_a_logical_ram_width = 8;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.ram_block_type = "auto";
defparam ram_block1a1.mem_init0 = 128'hD2969696D24926C99999CE38E1F01FFF;

cycloneiii_ram_block ram_block1a2(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a2_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.init_file = "fft_1n512cos.hex";
defparam ram_block1a2.init_file_layout = "port_a";
defparam ram_block1a2.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_3dp_rom_fft_120:twrom|twid_rom_fft_120:\\gen_M4K:cos_1n|altsyncram:\\gen_auto:altsyncram_component|altsyncram_b191:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.operation_mode = "rom";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 7;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "clock0";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 127;
defparam ram_block1a2.port_a_logical_ram_depth = 128;
defparam ram_block1a2.port_a_logical_ram_width = 8;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.ram_block_type = "auto";
defparam ram_block1a2.mem_init0 = 128'h318E718E31C71E3878783E07E00FFFFF;

cycloneiii_ram_block ram_block1a3(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a3_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.init_file = "fft_1n512cos.hex";
defparam ram_block1a3.init_file_layout = "port_a";
defparam ram_block1a3.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_3dp_rom_fft_120:twrom|twid_rom_fft_120:\\gen_M4K:cos_1n|altsyncram:\\gen_auto:altsyncram_component|altsyncram_b191:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.operation_mode = "rom";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 7;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "clock0";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 127;
defparam ram_block1a3.port_a_logical_ram_depth = 128;
defparam ram_block1a3.port_a_logical_ram_width = 8;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.ram_block_type = "auto";
defparam ram_block1a3.mem_init0 = 128'h0F81F07E0FC0FE07F807FE001FFFFFFF;

cycloneiii_ram_block ram_block1a4(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a4_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.init_file = "fft_1n512cos.hex";
defparam ram_block1a4.init_file_layout = "port_a";
defparam ram_block1a4.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_3dp_rom_fft_120:twrom|twid_rom_fft_120:\\gen_M4K:cos_1n|altsyncram:\\gen_auto:altsyncram_component|altsyncram_b191:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.operation_mode = "rom";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 7;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "clock0";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 127;
defparam ram_block1a4.port_a_logical_ram_depth = 128;
defparam ram_block1a4.port_a_logical_ram_width = 8;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.ram_block_type = "auto";
defparam ram_block1a4.mem_init0 = 128'h007FF001FFC001FFF80001FFFFFFFFFF;

cycloneiii_ram_block ram_block1a5(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a5_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.init_file = "fft_1n512cos.hex";
defparam ram_block1a5.init_file_layout = "port_a";
defparam ram_block1a5.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_3dp_rom_fft_120:twrom|twid_rom_fft_120:\\gen_M4K:cos_1n|altsyncram:\\gen_auto:altsyncram_component|altsyncram_b191:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.operation_mode = "rom";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 7;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "clock0";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 127;
defparam ram_block1a5.port_a_logical_ram_depth = 128;
defparam ram_block1a5.port_a_logical_ram_width = 8;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.ram_block_type = "auto";
defparam ram_block1a5.mem_init0 = 128'h00000FFFFFC0000007FFFFFFFFFFFFFF;

cycloneiii_ram_block ram_block1a6(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a6_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.init_file = "fft_1n512cos.hex";
defparam ram_block1a6.init_file_layout = "port_a";
defparam ram_block1a6.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_3dp_rom_fft_120:twrom|twid_rom_fft_120:\\gen_M4K:cos_1n|altsyncram:\\gen_auto:altsyncram_component|altsyncram_b191:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.operation_mode = "rom";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 7;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "clock0";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 127;
defparam ram_block1a6.port_a_logical_ram_depth = 128;
defparam ram_block1a6.port_a_logical_ram_width = 8;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.ram_block_type = "auto";
defparam ram_block1a6.mem_init0 = 128'h00000000003FFFFFFFFFFFFFFFFFFFFF;

cycloneiii_ram_block ram_block1a7(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a7_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.init_file = "fft_1n512cos.hex";
defparam ram_block1a7.init_file_layout = "port_a";
defparam ram_block1a7.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_3dp_rom_fft_120:twrom|twid_rom_fft_120:\\gen_M4K:cos_1n|altsyncram:\\gen_auto:altsyncram_component|altsyncram_b191:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.operation_mode = "rom";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 7;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "clock0";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 127;
defparam ram_block1a7.port_a_logical_ram_depth = 128;
defparam ram_block1a7.port_a_logical_ram_width = 8;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.ram_block_type = "auto";
defparam ram_block1a7.mem_init0 = 128'h00000000000000000000000000000000;

endmodule

module fft_twid_rom_fft_120_1 (
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_3,
	q_a_4,
	q_a_5,
	q_a_6,
	q_a_7,
	global_clock_enable,
	twad_tdl_0_6,
	twad_tdl_1_6,
	twad_tdl_2_6,
	twad_tdl_3_6,
	twad_tdl_4_6,
	twad_tdl_5_6,
	twad_tdl_6_6,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_a_0;
output 	q_a_1;
output 	q_a_2;
output 	q_a_3;
output 	q_a_4;
output 	q_a_5;
output 	q_a_6;
output 	q_a_7;
input 	global_clock_enable;
input 	twad_tdl_0_6;
input 	twad_tdl_1_6;
input 	twad_tdl_2_6;
input 	twad_tdl_3_6;
input 	twad_tdl_4_6;
input 	twad_tdl_5_6;
input 	twad_tdl_6_6;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_altsyncram_2 \gen_auto:altsyncram_component (
	.q_a({q_a_unconnected_wire_15,q_a_unconnected_wire_14,q_a_unconnected_wire_13,q_a_unconnected_wire_12,q_a_unconnected_wire_11,q_a_unconnected_wire_10,q_a_unconnected_wire_9,q_a_unconnected_wire_8,q_a_7,q_a_6,q_a_5,q_a_4,q_a_3,q_a_2,q_a_1,q_a_0}),
	.clocken0(global_clock_enable),
	.address_a({twad_tdl_6_6,twad_tdl_5_6,twad_tdl_4_6,twad_tdl_3_6,twad_tdl_2_6,twad_tdl_1_6,twad_tdl_0_6}),
	.clock0(clk));

endmodule

module fft_altsyncram_2 (
	q_a,
	clocken0,
	address_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_a;
input 	clocken0;
input 	[6:0] address_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_altsyncram_c191 auto_generated(
	.q_a({q_a[7],q_a[6],q_a[5],q_a[4],q_a[3],q_a[2],q_a[1],q_a[0]}),
	.clocken0(clocken0),
	.address_a({address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.clock0(clock0));

endmodule

module fft_altsyncram_c191 (
	q_a,
	clocken0,
	address_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q_a;
input 	clocken0;
input 	[6:0] address_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTADATAOUT_bus;
wire [143:0] ram_block1a1_PORTADATAOUT_bus;
wire [143:0] ram_block1a2_PORTADATAOUT_bus;
wire [143:0] ram_block1a3_PORTADATAOUT_bus;
wire [143:0] ram_block1a4_PORTADATAOUT_bus;
wire [143:0] ram_block1a5_PORTADATAOUT_bus;
wire [143:0] ram_block1a6_PORTADATAOUT_bus;
wire [143:0] ram_block1a7_PORTADATAOUT_bus;

assign q_a[0] = ram_block1a0_PORTADATAOUT_bus[0];

assign q_a[1] = ram_block1a1_PORTADATAOUT_bus[0];

assign q_a[2] = ram_block1a2_PORTADATAOUT_bus[0];

assign q_a[3] = ram_block1a3_PORTADATAOUT_bus[0];

assign q_a[4] = ram_block1a4_PORTADATAOUT_bus[0];

assign q_a[5] = ram_block1a5_PORTADATAOUT_bus[0];

assign q_a[6] = ram_block1a6_PORTADATAOUT_bus[0];

assign q_a[7] = ram_block1a7_PORTADATAOUT_bus[0];

cycloneiii_ram_block ram_block1a0(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a0_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.init_file = "fft_2n512cos.hex";
defparam ram_block1a0.init_file_layout = "port_a";
defparam ram_block1a0.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_3dp_rom_fft_120:twrom|twid_rom_fft_120:\\gen_M4K:cos_2n|altsyncram:\\gen_auto:altsyncram_component|altsyncram_c191:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.operation_mode = "rom";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 7;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "clock0";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 127;
defparam ram_block1a0.port_a_logical_ram_depth = 128;
defparam ram_block1a0.port_a_logical_ram_width = 8;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.ram_block_type = "auto";
defparam ram_block1a0.mem_init0 = 128'hE3496E00736B554AA555AD9C00ED258F;

cycloneiii_ram_block ram_block1a1(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a1_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.init_file = "fft_2n512cos.hex";
defparam ram_block1a1.init_file_layout = "port_a";
defparam ram_block1a1.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_3dp_rom_fft_120:twrom|twid_rom_fft_120:\\gen_M4K:cos_2n|altsyncram:\\gen_auto:altsyncram_component|altsyncram_c191:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.operation_mode = "rom";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 7;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "clock0";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 127;
defparam ram_block1a1.port_a_logical_ram_depth = 128;
defparam ram_block1a1.port_a_logical_ram_width = 8;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.ram_block_type = "auto";
defparam ram_block1a1.mem_init0 = 128'h1F3B25555A4D998CC666C92955A49C7F;

cycloneiii_ram_block ram_block1a2(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a2_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.init_file = "fft_2n512cos.hex";
defparam ram_block1a2.init_file_layout = "port_a";
defparam ram_block1a2.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_3dp_rom_fft_120:twrom|twid_rom_fft_120:\\gen_M4K:cos_2n|altsyncram:\\gen_auto:altsyncram_component|altsyncram_c191:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.operation_mode = "rom";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 7;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "clock0";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 127;
defparam ram_block1a2.port_a_logical_ram_depth = 128;
defparam ram_block1a2.port_a_logical_ram_width = 8;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.ram_block_type = "auto";
defparam ram_block1a2.mem_init0 = 128'h00F8E33336DB4B5A52D25B64CC6383FF;

cycloneiii_ram_block ram_block1a3(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a3_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.init_file = "fft_2n512cos.hex";
defparam ram_block1a3.init_file_layout = "port_a";
defparam ram_block1a3.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_3dp_rom_fft_120:twrom|twid_rom_fft_120:\\gen_M4K:cos_2n|altsyncram:\\gen_auto:altsyncram_component|altsyncram_c191:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.operation_mode = "rom";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 7;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "clock0";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 127;
defparam ram_block1a3.port_a_logical_ram_depth = 128;
defparam ram_block1a3.port_a_logical_ram_width = 8;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.ram_block_type = "auto";
defparam ram_block1a3.mem_init0 = 128'h0007E0F0F1C738C631CE38E3C3E07FFF;

cycloneiii_ram_block ram_block1a4(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a4_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.init_file = "fft_2n512cos.hex";
defparam ram_block1a4.init_file_layout = "port_a";
defparam ram_block1a4.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_3dp_rom_fft_120:twrom|twid_rom_fft_120:\\gen_M4K:cos_2n|altsyncram:\\gen_auto:altsyncram_component|altsyncram_c191:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.operation_mode = "rom";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 7;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "clock0";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 127;
defparam ram_block1a4.port_a_logical_ram_depth = 128;
defparam ram_block1a4.port_a_logical_ram_width = 8;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.ram_block_type = "auto";
defparam ram_block1a4.mem_init0 = 128'h00001FF00FC0F83E0FC1F81FC01FFFFF;

cycloneiii_ram_block ram_block1a5(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a5_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.init_file = "fft_2n512cos.hex";
defparam ram_block1a5.init_file_layout = "port_a";
defparam ram_block1a5.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_3dp_rom_fft_120:twrom|twid_rom_fft_120:\\gen_M4K:cos_2n|altsyncram:\\gen_auto:altsyncram_component|altsyncram_c191:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.operation_mode = "rom";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 7;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "clock0";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 127;
defparam ram_block1a5.port_a_logical_ram_depth = 128;
defparam ram_block1a5.port_a_logical_ram_width = 8;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.ram_block_type = "auto";
defparam ram_block1a5.mem_init0 = 128'h0000000FFFC007FE003FF8003FFFFFFF;

cycloneiii_ram_block ram_block1a6(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a6_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.init_file = "fft_2n512cos.hex";
defparam ram_block1a6.init_file_layout = "port_a";
defparam ram_block1a6.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_3dp_rom_fft_120:twrom|twid_rom_fft_120:\\gen_M4K:cos_2n|altsyncram:\\gen_auto:altsyncram_component|altsyncram_c191:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.operation_mode = "rom";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 7;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "clock0";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 127;
defparam ram_block1a6.port_a_logical_ram_depth = 128;
defparam ram_block1a6.port_a_logical_ram_width = 8;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.ram_block_type = "auto";
defparam ram_block1a6.mem_init0 = 128'h00000000003FFFFE000007FFFFFFFFFF;

cycloneiii_ram_block ram_block1a7(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a7_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.init_file = "fft_2n512cos.hex";
defparam ram_block1a7.init_file_layout = "port_a";
defparam ram_block1a7.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_3dp_rom_fft_120:twrom|twid_rom_fft_120:\\gen_M4K:cos_2n|altsyncram:\\gen_auto:altsyncram_component|altsyncram_c191:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.operation_mode = "rom";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 7;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "clock0";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 127;
defparam ram_block1a7.port_a_logical_ram_depth = 128;
defparam ram_block1a7.port_a_logical_ram_width = 8;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.ram_block_type = "auto";
defparam ram_block1a7.mem_init0 = 128'hFFFFFFFFFFFFFFFE0000000000000000;

endmodule

module fft_twid_rom_fft_120_2 (
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_3,
	q_a_4,
	q_a_5,
	q_a_6,
	q_a_7,
	global_clock_enable,
	twad_tdl_0_6,
	twad_tdl_1_6,
	twad_tdl_2_6,
	twad_tdl_3_6,
	twad_tdl_4_6,
	twad_tdl_5_6,
	twad_tdl_6_6,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_a_0;
output 	q_a_1;
output 	q_a_2;
output 	q_a_3;
output 	q_a_4;
output 	q_a_5;
output 	q_a_6;
output 	q_a_7;
input 	global_clock_enable;
input 	twad_tdl_0_6;
input 	twad_tdl_1_6;
input 	twad_tdl_2_6;
input 	twad_tdl_3_6;
input 	twad_tdl_4_6;
input 	twad_tdl_5_6;
input 	twad_tdl_6_6;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_altsyncram_3 \gen_auto:altsyncram_component (
	.q_a({q_a_unconnected_wire_15,q_a_unconnected_wire_14,q_a_unconnected_wire_13,q_a_unconnected_wire_12,q_a_unconnected_wire_11,q_a_unconnected_wire_10,q_a_unconnected_wire_9,q_a_unconnected_wire_8,q_a_7,q_a_6,q_a_5,q_a_4,q_a_3,q_a_2,q_a_1,q_a_0}),
	.clocken0(global_clock_enable),
	.address_a({twad_tdl_6_6,twad_tdl_5_6,twad_tdl_4_6,twad_tdl_3_6,twad_tdl_2_6,twad_tdl_1_6,twad_tdl_0_6}),
	.clock0(clk));

endmodule

module fft_altsyncram_3 (
	q_a,
	clocken0,
	address_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_a;
input 	clocken0;
input 	[6:0] address_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_altsyncram_d191 auto_generated(
	.q_a({q_a[7],q_a[6],q_a[5],q_a[4],q_a[3],q_a[2],q_a[1],q_a[0]}),
	.clocken0(clocken0),
	.address_a({address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.clock0(clock0));

endmodule

module fft_altsyncram_d191 (
	q_a,
	clocken0,
	address_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q_a;
input 	clocken0;
input 	[6:0] address_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTADATAOUT_bus;
wire [143:0] ram_block1a1_PORTADATAOUT_bus;
wire [143:0] ram_block1a2_PORTADATAOUT_bus;
wire [143:0] ram_block1a3_PORTADATAOUT_bus;
wire [143:0] ram_block1a4_PORTADATAOUT_bus;
wire [143:0] ram_block1a5_PORTADATAOUT_bus;
wire [143:0] ram_block1a6_PORTADATAOUT_bus;
wire [143:0] ram_block1a7_PORTADATAOUT_bus;

assign q_a[0] = ram_block1a0_PORTADATAOUT_bus[0];

assign q_a[1] = ram_block1a1_PORTADATAOUT_bus[0];

assign q_a[2] = ram_block1a2_PORTADATAOUT_bus[0];

assign q_a[3] = ram_block1a3_PORTADATAOUT_bus[0];

assign q_a[4] = ram_block1a4_PORTADATAOUT_bus[0];

assign q_a[5] = ram_block1a5_PORTADATAOUT_bus[0];

assign q_a[6] = ram_block1a6_PORTADATAOUT_bus[0];

assign q_a[7] = ram_block1a7_PORTADATAOUT_bus[0];

cycloneiii_ram_block ram_block1a0(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a0_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.init_file = "fft_3n512cos.hex";
defparam ram_block1a0.init_file_layout = "port_a";
defparam ram_block1a0.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_3dp_rom_fft_120:twrom|twid_rom_fft_120:\\gen_M4K:cos_3n|altsyncram:\\gen_auto:altsyncram_component|altsyncram_d191:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.operation_mode = "rom";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 7;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "clock0";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 127;
defparam ram_block1a0.port_a_logical_ram_depth = 128;
defparam ram_block1a0.port_a_logical_ram_width = 8;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.ram_block_type = "auto";
defparam ram_block1a0.mem_init0 = 128'hD9871A9FD4FB206A60732499FF2A78A7;

cycloneiii_ram_block ram_block1a1(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a1_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.init_file = "fft_3n512cos.hex";
defparam ram_block1a1.init_file_layout = "port_a";
defparam ram_block1a1.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_3dp_rom_fft_120:twrom|twid_rom_fft_120:\\gen_M4K:cos_3n|altsyncram:\\gen_auto:altsyncram_component|altsyncram_d191:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.operation_mode = "rom";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 7;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "clock0";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 127;
defparam ram_block1a1.port_a_logical_ram_depth = 128;
defparam ram_block1a1.port_a_logical_ram_width = 8;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.ram_block_type = "auto";
defparam ram_block1a1.mem_init0 = 128'hE1F8F9B567076AB3800F1C780033559F;

cycloneiii_ram_block ram_block1a2(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a2_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.init_file = "fft_3n512cos.hex";
defparam ram_block1a2.init_file_layout = "port_a";
defparam ram_block1a2.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_3dp_rom_fft_120:twrom|twid_rom_fft_120:\\gen_M4K:cos_3n|altsyncram:\\gen_auto:altsyncram_component|altsyncram_d191:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.operation_mode = "rom";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 7;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "clock0";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 127;
defparam ram_block1a2.port_a_logical_ram_depth = 128;
defparam ram_block1a2.port_a_logical_ram_width = 8;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.ram_block_type = "auto";
defparam ram_block1a2.mem_init0 = 128'h54AAAD267800E6695555A952AA96CC7F;

cycloneiii_ram_block ram_block1a3(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a3_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.init_file = "fft_3n512cos.hex";
defparam ram_block1a3.init_file_layout = "port_a";
defparam ram_block1a3.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_3dp_rom_fft_120:twrom|twid_rom_fft_120:\\gen_M4K:cos_3n|altsyncram:\\gen_auto:altsyncram_component|altsyncram_d191:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.operation_mode = "rom";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 7;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "clock0";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 127;
defparam ram_block1a3.port_a_logical_ram_depth = 128;
defparam ram_block1a3.port_a_logical_ram_width = 8;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.ram_block_type = "auto";
defparam ram_block1a3.mem_init0 = 128'h993331C780001E18CCCC9B366671C3FF;

cycloneiii_ram_block ram_block1a4(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a4_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.init_file = "fft_3n512cos.hex";
defparam ram_block1a4.init_file_layout = "port_a";
defparam ram_block1a4.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_3dp_rom_fft_120:twrom|twid_rom_fft_120:\\gen_M4K:cos_3n|altsyncram:\\gen_auto:altsyncram_component|altsyncram_d191:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.operation_mode = "rom";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 7;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "clock0";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 127;
defparam ram_block1a4.port_a_logical_ram_depth = 128;
defparam ram_block1a4.port_a_logical_ram_width = 8;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.ram_block_type = "auto";
defparam ram_block1a4.mem_init0 = 128'hE1C3C1F8000001F83C3C78F1E1F03FFF;

cycloneiii_ram_block ram_block1a5(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a5_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.init_file = "fft_3n512cos.hex";
defparam ram_block1a5.init_file_layout = "port_a";
defparam ram_block1a5.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_3dp_rom_fft_120:twrom|twid_rom_fft_120:\\gen_M4K:cos_3n|altsyncram:\\gen_auto:altsyncram_component|altsyncram_d191:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.operation_mode = "rom";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 7;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "clock0";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 127;
defparam ram_block1a5.port_a_logical_ram_depth = 128;
defparam ram_block1a5.port_a_logical_ram_width = 8;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.ram_block_type = "auto";
defparam ram_block1a5.mem_init0 = 128'hFE03FE0000000007FC03F80FE00FFFFF;

cycloneiii_ram_block ram_block1a6(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a6_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.init_file = "fft_3n512cos.hex";
defparam ram_block1a6.init_file_layout = "port_a";
defparam ram_block1a6.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_3dp_rom_fft_120:twrom|twid_rom_fft_120:\\gen_M4K:cos_3n|altsyncram:\\gen_auto:altsyncram_component|altsyncram_d191:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.operation_mode = "rom";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 7;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "clock0";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 127;
defparam ram_block1a6.port_a_logical_ram_depth = 128;
defparam ram_block1a6.port_a_logical_ram_width = 8;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.ram_block_type = "auto";
defparam ram_block1a6.mem_init0 = 128'hFFFC00000000000003FFF8001FFFFFFF;

cycloneiii_ram_block ram_block1a7(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a7_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.init_file = "fft_3n512cos.hex";
defparam ram_block1a7.init_file_layout = "port_a";
defparam ram_block1a7.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_3dp_rom_fft_120:twrom|twid_rom_fft_120:\\gen_M4K:cos_3n|altsyncram:\\gen_auto:altsyncram_component|altsyncram_d191:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.operation_mode = "rom";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 7;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "clock0";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 127;
defparam ram_block1a7.port_a_logical_ram_depth = 128;
defparam ram_block1a7.port_a_logical_ram_width = 8;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.ram_block_type = "auto";
defparam ram_block1a7.mem_init0 = 128'hFFFFFFFFFFFFFFFFFFFFF80000000000;

endmodule

module fft_twid_rom_fft_120_3 (
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_3,
	q_a_4,
	q_a_5,
	q_a_6,
	q_a_7,
	global_clock_enable,
	twad_tdl_0_6,
	twad_tdl_1_6,
	twad_tdl_2_6,
	twad_tdl_3_6,
	twad_tdl_4_6,
	twad_tdl_5_6,
	twad_tdl_6_6,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_a_0;
output 	q_a_1;
output 	q_a_2;
output 	q_a_3;
output 	q_a_4;
output 	q_a_5;
output 	q_a_6;
output 	q_a_7;
input 	global_clock_enable;
input 	twad_tdl_0_6;
input 	twad_tdl_1_6;
input 	twad_tdl_2_6;
input 	twad_tdl_3_6;
input 	twad_tdl_4_6;
input 	twad_tdl_5_6;
input 	twad_tdl_6_6;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_altsyncram_4 \gen_auto:altsyncram_component (
	.q_a({q_a_unconnected_wire_15,q_a_unconnected_wire_14,q_a_unconnected_wire_13,q_a_unconnected_wire_12,q_a_unconnected_wire_11,q_a_unconnected_wire_10,q_a_unconnected_wire_9,q_a_unconnected_wire_8,q_a_7,q_a_6,q_a_5,q_a_4,q_a_3,q_a_2,q_a_1,q_a_0}),
	.clocken0(global_clock_enable),
	.address_a({twad_tdl_6_6,twad_tdl_5_6,twad_tdl_4_6,twad_tdl_3_6,twad_tdl_2_6,twad_tdl_1_6,twad_tdl_0_6}),
	.clock0(clk));

endmodule

module fft_altsyncram_4 (
	q_a,
	clocken0,
	address_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_a;
input 	clocken0;
input 	[6:0] address_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_altsyncram_g191 auto_generated(
	.q_a({q_a[7],q_a[6],q_a[5],q_a[4],q_a[3],q_a[2],q_a[1],q_a[0]}),
	.clocken0(clocken0),
	.address_a({address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.clock0(clock0));

endmodule

module fft_altsyncram_g191 (
	q_a,
	clocken0,
	address_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q_a;
input 	clocken0;
input 	[6:0] address_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTADATAOUT_bus;
wire [143:0] ram_block1a1_PORTADATAOUT_bus;
wire [143:0] ram_block1a2_PORTADATAOUT_bus;
wire [143:0] ram_block1a3_PORTADATAOUT_bus;
wire [143:0] ram_block1a4_PORTADATAOUT_bus;
wire [143:0] ram_block1a5_PORTADATAOUT_bus;
wire [143:0] ram_block1a6_PORTADATAOUT_bus;
wire [143:0] ram_block1a7_PORTADATAOUT_bus;

assign q_a[0] = ram_block1a0_PORTADATAOUT_bus[0];

assign q_a[1] = ram_block1a1_PORTADATAOUT_bus[0];

assign q_a[2] = ram_block1a2_PORTADATAOUT_bus[0];

assign q_a[3] = ram_block1a3_PORTADATAOUT_bus[0];

assign q_a[4] = ram_block1a4_PORTADATAOUT_bus[0];

assign q_a[5] = ram_block1a5_PORTADATAOUT_bus[0];

assign q_a[6] = ram_block1a6_PORTADATAOUT_bus[0];

assign q_a[7] = ram_block1a7_PORTADATAOUT_bus[0];

cycloneiii_ram_block ram_block1a0(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a0_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.init_file = "fft_1n512sin.hex";
defparam ram_block1a0.init_file_layout = "port_a";
defparam ram_block1a0.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_3dp_rom_fft_120:twrom|twid_rom_fft_120:\\gen_M4K:sin_1n|altsyncram:\\gen_auto:altsyncram_component|altsyncram_g191:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.operation_mode = "rom";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 7;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "clock0";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 127;
defparam ram_block1a0.port_a_logical_ram_depth = 128;
defparam ram_block1a0.port_a_logical_ram_width = 8;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.ram_block_type = "auto";
defparam ram_block1a0.mem_init0 = 128'hFE0F18C9B6D4AAAA95A5B64D999998CC;

cycloneiii_ram_block ram_block1a1(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a1_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.init_file = "fft_1n512sin.hex";
defparam ram_block1a1.init_file_layout = "port_a";
defparam ram_block1a1.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_3dp_rom_fft_120:twrom|twid_rom_fft_120:\\gen_M4K:sin_1n|altsyncram:\\gen_auto:altsyncram_component|altsyncram_g191:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.operation_mode = "rom";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 7;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "clock0";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 127;
defparam ram_block1a1.port_a_logical_ram_depth = 128;
defparam ram_block1a1.port_a_logical_ram_width = 8;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.ram_block_type = "auto";
defparam ram_block1a1.mem_init0 = 128'hFFF01F0E38E7333326C92496D2D2D296;

cycloneiii_ram_block ram_block1a2(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a2_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.init_file = "fft_1n512sin.hex";
defparam ram_block1a2.init_file_layout = "port_a";
defparam ram_block1a2.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_3dp_rom_fft_120:twrom|twid_rom_fft_120:\\gen_M4K:sin_1n|altsyncram:\\gen_auto:altsyncram_component|altsyncram_g191:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.operation_mode = "rom";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 7;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "clock0";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 127;
defparam ram_block1a2.port_a_logical_ram_depth = 128;
defparam ram_block1a2.port_a_logical_ram_width = 8;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.ram_block_type = "auto";
defparam ram_block1a2.mem_init0 = 128'hFFFFE00FC0F83C3C38F1C718E31CE318;

cycloneiii_ram_block ram_block1a3(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a3_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.init_file = "fft_1n512sin.hex";
defparam ram_block1a3.init_file_layout = "port_a";
defparam ram_block1a3.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_3dp_rom_fft_120:twrom|twid_rom_fft_120:\\gen_M4K:sin_1n|altsyncram:\\gen_auto:altsyncram_component|altsyncram_g191:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.operation_mode = "rom";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 7;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "clock0";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 127;
defparam ram_block1a3.port_a_logical_ram_depth = 128;
defparam ram_block1a3.port_a_logical_ram_width = 8;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.ram_block_type = "auto";
defparam ram_block1a3.mem_init0 = 128'hFFFFFFF000FFC03FC0FE07E0FC1F03E0;

cycloneiii_ram_block ram_block1a4(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a4_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.init_file = "fft_1n512sin.hex";
defparam ram_block1a4.init_file_layout = "port_a";
defparam ram_block1a4.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_3dp_rom_fft_120:twrom|twid_rom_fft_120:\\gen_M4K:sin_1n|altsyncram:\\gen_auto:altsyncram_component|altsyncram_g191:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.operation_mode = "rom";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 7;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "clock0";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 127;
defparam ram_block1a4.port_a_logical_ram_depth = 128;
defparam ram_block1a4.port_a_logical_ram_width = 8;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.ram_block_type = "auto";
defparam ram_block1a4.mem_init0 = 128'hFFFFFFFFFF00003FFF0007FF001FFC00;

cycloneiii_ram_block ram_block1a5(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a5_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.init_file = "fft_1n512sin.hex";
defparam ram_block1a5.init_file_layout = "port_a";
defparam ram_block1a5.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_3dp_rom_fft_120:twrom|twid_rom_fft_120:\\gen_M4K:sin_1n|altsyncram:\\gen_auto:altsyncram_component|altsyncram_g191:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.operation_mode = "rom";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 7;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "clock0";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 127;
defparam ram_block1a5.port_a_logical_ram_depth = 128;
defparam ram_block1a5.port_a_logical_ram_width = 8;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.ram_block_type = "auto";
defparam ram_block1a5.mem_init0 = 128'hFFFFFFFFFFFFFFC0000007FFFFE00000;

cycloneiii_ram_block ram_block1a6(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a6_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.init_file = "fft_1n512sin.hex";
defparam ram_block1a6.init_file_layout = "port_a";
defparam ram_block1a6.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_3dp_rom_fft_120:twrom|twid_rom_fft_120:\\gen_M4K:sin_1n|altsyncram:\\gen_auto:altsyncram_component|altsyncram_g191:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.operation_mode = "rom";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 7;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "clock0";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 127;
defparam ram_block1a6.port_a_logical_ram_depth = 128;
defparam ram_block1a6.port_a_logical_ram_width = 8;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.ram_block_type = "auto";
defparam ram_block1a6.mem_init0 = 128'hFFFFFFFFFFFFFFFFFFFFF80000000000;

cycloneiii_ram_block ram_block1a7(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a7_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.init_file = "fft_1n512sin.hex";
defparam ram_block1a7.init_file_layout = "port_a";
defparam ram_block1a7.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_3dp_rom_fft_120:twrom|twid_rom_fft_120:\\gen_M4K:sin_1n|altsyncram:\\gen_auto:altsyncram_component|altsyncram_g191:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.operation_mode = "rom";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 7;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "clock0";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 127;
defparam ram_block1a7.port_a_logical_ram_depth = 128;
defparam ram_block1a7.port_a_logical_ram_width = 8;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.ram_block_type = "auto";
defparam ram_block1a7.mem_init0 = 128'h00000000000000000000000000000000;

endmodule

module fft_twid_rom_fft_120_4 (
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_3,
	q_a_4,
	q_a_5,
	q_a_6,
	q_a_7,
	global_clock_enable,
	twad_tdl_0_6,
	twad_tdl_1_6,
	twad_tdl_2_6,
	twad_tdl_3_6,
	twad_tdl_4_6,
	twad_tdl_5_6,
	twad_tdl_6_6,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_a_0;
output 	q_a_1;
output 	q_a_2;
output 	q_a_3;
output 	q_a_4;
output 	q_a_5;
output 	q_a_6;
output 	q_a_7;
input 	global_clock_enable;
input 	twad_tdl_0_6;
input 	twad_tdl_1_6;
input 	twad_tdl_2_6;
input 	twad_tdl_3_6;
input 	twad_tdl_4_6;
input 	twad_tdl_5_6;
input 	twad_tdl_6_6;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_altsyncram_5 \gen_auto:altsyncram_component (
	.q_a({q_a_unconnected_wire_15,q_a_unconnected_wire_14,q_a_unconnected_wire_13,q_a_unconnected_wire_12,q_a_unconnected_wire_11,q_a_unconnected_wire_10,q_a_unconnected_wire_9,q_a_unconnected_wire_8,q_a_7,q_a_6,q_a_5,q_a_4,q_a_3,q_a_2,q_a_1,q_a_0}),
	.clocken0(global_clock_enable),
	.address_a({twad_tdl_6_6,twad_tdl_5_6,twad_tdl_4_6,twad_tdl_3_6,twad_tdl_2_6,twad_tdl_1_6,twad_tdl_0_6}),
	.clock0(clk));

endmodule

module fft_altsyncram_5 (
	q_a,
	clocken0,
	address_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_a;
input 	clocken0;
input 	[6:0] address_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_altsyncram_h191 auto_generated(
	.q_a({q_a[7],q_a[6],q_a[5],q_a[4],q_a[3],q_a[2],q_a[1],q_a[0]}),
	.clocken0(clocken0),
	.address_a({address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.clock0(clock0));

endmodule

module fft_altsyncram_h191 (
	q_a,
	clocken0,
	address_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q_a;
input 	clocken0;
input 	[6:0] address_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTADATAOUT_bus;
wire [143:0] ram_block1a1_PORTADATAOUT_bus;
wire [143:0] ram_block1a2_PORTADATAOUT_bus;
wire [143:0] ram_block1a3_PORTADATAOUT_bus;
wire [143:0] ram_block1a4_PORTADATAOUT_bus;
wire [143:0] ram_block1a5_PORTADATAOUT_bus;
wire [143:0] ram_block1a6_PORTADATAOUT_bus;
wire [143:0] ram_block1a7_PORTADATAOUT_bus;

assign q_a[0] = ram_block1a0_PORTADATAOUT_bus[0];

assign q_a[1] = ram_block1a1_PORTADATAOUT_bus[0];

assign q_a[2] = ram_block1a2_PORTADATAOUT_bus[0];

assign q_a[3] = ram_block1a3_PORTADATAOUT_bus[0];

assign q_a[4] = ram_block1a4_PORTADATAOUT_bus[0];

assign q_a[5] = ram_block1a5_PORTADATAOUT_bus[0];

assign q_a[6] = ram_block1a6_PORTADATAOUT_bus[0];

assign q_a[7] = ram_block1a7_PORTADATAOUT_bus[0];

cycloneiii_ram_block ram_block1a0(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a0_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.init_file = "fft_2n512sin.hex";
defparam ram_block1a0.init_file_layout = "port_a";
defparam ram_block1a0.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_3dp_rom_fft_120:twrom|twid_rom_fft_120:\\gen_M4K:sin_2n|altsyncram:\\gen_auto:altsyncram_component|altsyncram_h191:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.operation_mode = "rom";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 7;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "clock0";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 127;
defparam ram_block1a0.port_a_logical_ram_depth = 128;
defparam ram_block1a0.port_a_logical_ram_width = 8;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.ram_block_type = "auto";
defparam ram_block1a0.mem_init0 = 128'hA555AD9C00ED258FE3496E00736B554A;

cycloneiii_ram_block ram_block1a1(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a1_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.init_file = "fft_2n512sin.hex";
defparam ram_block1a1.init_file_layout = "port_a";
defparam ram_block1a1.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_3dp_rom_fft_120:twrom|twid_rom_fft_120:\\gen_M4K:sin_2n|altsyncram:\\gen_auto:altsyncram_component|altsyncram_h191:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.operation_mode = "rom";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 7;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "clock0";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 127;
defparam ram_block1a1.port_a_logical_ram_depth = 128;
defparam ram_block1a1.port_a_logical_ram_width = 8;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.ram_block_type = "auto";
defparam ram_block1a1.mem_init0 = 128'hC666C92955A49C7FFC724B552926CCC6;

cycloneiii_ram_block ram_block1a2(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a2_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.init_file = "fft_2n512sin.hex";
defparam ram_block1a2.init_file_layout = "port_a";
defparam ram_block1a2.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_3dp_rom_fft_120:twrom|twid_rom_fft_120:\\gen_M4K:sin_2n|altsyncram:\\gen_auto:altsyncram_component|altsyncram_h191:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.operation_mode = "rom";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 7;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "clock0";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 127;
defparam ram_block1a2.port_a_logical_ram_depth = 128;
defparam ram_block1a2.port_a_logical_ram_width = 8;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.ram_block_type = "auto";
defparam ram_block1a2.mem_init0 = 128'h52D25B64CC6383FFFF838C664DB49694;

cycloneiii_ram_block ram_block1a3(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a3_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.init_file = "fft_2n512sin.hex";
defparam ram_block1a3.init_file_layout = "port_a";
defparam ram_block1a3.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_3dp_rom_fft_120:twrom|twid_rom_fft_120:\\gen_M4K:sin_2n|altsyncram:\\gen_auto:altsyncram_component|altsyncram_h191:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.operation_mode = "rom";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 7;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "clock0";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 127;
defparam ram_block1a3.port_a_logical_ram_depth = 128;
defparam ram_block1a3.port_a_logical_ram_width = 8;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.ram_block_type = "auto";
defparam ram_block1a3.mem_init0 = 128'h31CE38E3C3E07FFFFFFC0F878E38E718;

cycloneiii_ram_block ram_block1a4(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a4_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.init_file = "fft_2n512sin.hex";
defparam ram_block1a4.init_file_layout = "port_a";
defparam ram_block1a4.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_3dp_rom_fft_120:twrom|twid_rom_fft_120:\\gen_M4K:sin_2n|altsyncram:\\gen_auto:altsyncram_component|altsyncram_h191:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.operation_mode = "rom";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 7;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "clock0";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 127;
defparam ram_block1a4.port_a_logical_ram_depth = 128;
defparam ram_block1a4.port_a_logical_ram_width = 8;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.ram_block_type = "auto";
defparam ram_block1a4.mem_init0 = 128'h0FC1F81FC01FFFFFFFFFF007F03F07E0;

cycloneiii_ram_block ram_block1a5(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a5_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.init_file = "fft_2n512sin.hex";
defparam ram_block1a5.init_file_layout = "port_a";
defparam ram_block1a5.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_3dp_rom_fft_120:twrom|twid_rom_fft_120:\\gen_M4K:sin_2n|altsyncram:\\gen_auto:altsyncram_component|altsyncram_h191:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.operation_mode = "rom";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 7;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "clock0";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 127;
defparam ram_block1a5.port_a_logical_ram_depth = 128;
defparam ram_block1a5.port_a_logical_ram_width = 8;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.ram_block_type = "auto";
defparam ram_block1a5.mem_init0 = 128'h003FF8003FFFFFFFFFFFFFF8003FF800;

cycloneiii_ram_block ram_block1a6(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a6_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.init_file = "fft_2n512sin.hex";
defparam ram_block1a6.init_file_layout = "port_a";
defparam ram_block1a6.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_3dp_rom_fft_120:twrom|twid_rom_fft_120:\\gen_M4K:sin_2n|altsyncram:\\gen_auto:altsyncram_component|altsyncram_h191:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.operation_mode = "rom";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 7;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "clock0";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 127;
defparam ram_block1a6.port_a_logical_ram_depth = 128;
defparam ram_block1a6.port_a_logical_ram_width = 8;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.ram_block_type = "auto";
defparam ram_block1a6.mem_init0 = 128'h000007FFFFFFFFFFFFFFFFFFFFC00000;

cycloneiii_ram_block ram_block1a7(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a7_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.init_file = "fft_2n512sin.hex";
defparam ram_block1a7.init_file_layout = "port_a";
defparam ram_block1a7.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_3dp_rom_fft_120:twrom|twid_rom_fft_120:\\gen_M4K:sin_2n|altsyncram:\\gen_auto:altsyncram_component|altsyncram_h191:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.operation_mode = "rom";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 7;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "clock0";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 127;
defparam ram_block1a7.port_a_logical_ram_depth = 128;
defparam ram_block1a7.port_a_logical_ram_width = 8;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.ram_block_type = "auto";
defparam ram_block1a7.mem_init0 = 128'h00000000000000000000000000000000;

endmodule

module fft_twid_rom_fft_120_5 (
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_3,
	q_a_4,
	q_a_5,
	q_a_6,
	q_a_7,
	global_clock_enable,
	twad_tdl_0_6,
	twad_tdl_1_6,
	twad_tdl_2_6,
	twad_tdl_3_6,
	twad_tdl_4_6,
	twad_tdl_5_6,
	twad_tdl_6_6,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_a_0;
output 	q_a_1;
output 	q_a_2;
output 	q_a_3;
output 	q_a_4;
output 	q_a_5;
output 	q_a_6;
output 	q_a_7;
input 	global_clock_enable;
input 	twad_tdl_0_6;
input 	twad_tdl_1_6;
input 	twad_tdl_2_6;
input 	twad_tdl_3_6;
input 	twad_tdl_4_6;
input 	twad_tdl_5_6;
input 	twad_tdl_6_6;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_altsyncram_6 \gen_auto:altsyncram_component (
	.q_a({q_a_unconnected_wire_15,q_a_unconnected_wire_14,q_a_unconnected_wire_13,q_a_unconnected_wire_12,q_a_unconnected_wire_11,q_a_unconnected_wire_10,q_a_unconnected_wire_9,q_a_unconnected_wire_8,q_a_7,q_a_6,q_a_5,q_a_4,q_a_3,q_a_2,q_a_1,q_a_0}),
	.clocken0(global_clock_enable),
	.address_a({twad_tdl_6_6,twad_tdl_5_6,twad_tdl_4_6,twad_tdl_3_6,twad_tdl_2_6,twad_tdl_1_6,twad_tdl_0_6}),
	.clock0(clk));

endmodule

module fft_altsyncram_6 (
	q_a,
	clocken0,
	address_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_a;
input 	clocken0;
input 	[6:0] address_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_altsyncram_i191 auto_generated(
	.q_a({q_a[7],q_a[6],q_a[5],q_a[4],q_a[3],q_a[2],q_a[1],q_a[0]}),
	.clocken0(clocken0),
	.address_a({address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.clock0(clock0));

endmodule

module fft_altsyncram_i191 (
	q_a,
	clocken0,
	address_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q_a;
input 	clocken0;
input 	[6:0] address_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTADATAOUT_bus;
wire [143:0] ram_block1a1_PORTADATAOUT_bus;
wire [143:0] ram_block1a2_PORTADATAOUT_bus;
wire [143:0] ram_block1a3_PORTADATAOUT_bus;
wire [143:0] ram_block1a4_PORTADATAOUT_bus;
wire [143:0] ram_block1a5_PORTADATAOUT_bus;
wire [143:0] ram_block1a6_PORTADATAOUT_bus;
wire [143:0] ram_block1a7_PORTADATAOUT_bus;

assign q_a[0] = ram_block1a0_PORTADATAOUT_bus[0];

assign q_a[1] = ram_block1a1_PORTADATAOUT_bus[0];

assign q_a[2] = ram_block1a2_PORTADATAOUT_bus[0];

assign q_a[3] = ram_block1a3_PORTADATAOUT_bus[0];

assign q_a[4] = ram_block1a4_PORTADATAOUT_bus[0];

assign q_a[5] = ram_block1a5_PORTADATAOUT_bus[0];

assign q_a[6] = ram_block1a6_PORTADATAOUT_bus[0];

assign q_a[7] = ram_block1a7_PORTADATAOUT_bus[0];

cycloneiii_ram_block ram_block1a0(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a0_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.init_file = "fft_3n512sin.hex";
defparam ram_block1a0.init_file_layout = "port_a";
defparam ram_block1a0.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_3dp_rom_fft_120:twrom|twid_rom_fft_120:\\gen_M4K:sin_3n|altsyncram:\\gen_auto:altsyncram_component|altsyncram_i191:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.operation_mode = "rom";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 7;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "clock0";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 127;
defparam ram_block1a0.port_a_logical_ram_depth = 128;
defparam ram_block1a0.port_a_logical_ram_width = 8;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.ram_block_type = "auto";
defparam ram_block1a0.mem_init0 = 128'hCA3CA9FF32499C0CAC09BE57F2B1C336;

cycloneiii_ram_block ram_block1a1(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a1_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.init_file = "fft_3n512sin.hex";
defparam ram_block1a1.init_file_layout = "port_a";
defparam ram_block1a1.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_3dp_rom_fft_120:twrom|twid_rom_fft_120:\\gen_M4K:sin_3n|altsyncram:\\gen_auto:altsyncram_component|altsyncram_i191:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.operation_mode = "rom";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 7;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "clock0";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 127;
defparam ram_block1a1.port_a_logical_ram_depth = 128;
defparam ram_block1a1.port_a_logical_ram_width = 8;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.ram_block_type = "auto";
defparam ram_block1a1.mem_init0 = 128'h396931FF0E387C0F36A47F9AA98FFC38;

cycloneiii_ram_block ram_block1a2(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a2_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.init_file = "fft_3n512sin.hex";
defparam ram_block1a2.init_file_layout = "port_a";
defparam ram_block1a2.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_3dp_rom_fft_120:twrom|twid_rom_fft_120:\\gen_M4K:sin_3n|altsyncram:\\gen_auto:altsyncram_component|altsyncram_i191:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.operation_mode = "rom";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 7;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "clock0";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 127;
defparam ram_block1a2.port_a_logical_ram_depth = 128;
defparam ram_block1a2.port_a_logical_ram_width = 8;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.ram_block_type = "auto";
defparam ram_block1a2.mem_init0 = 128'h071B6B55AB52A95A9263FFE332D5556A;

cycloneiii_ram_block ram_block1a3(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a3_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.init_file = "fft_3n512sin.hex";
defparam ram_block1a3.init_file_layout = "port_a";
defparam ram_block1a3.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_3dp_rom_fft_120:twrom|twid_rom_fft_120:\\gen_M4K:sin_3n|altsyncram:\\gen_auto:altsyncram_component|altsyncram_i191:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.operation_mode = "rom";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 7;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "clock0";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 127;
defparam ram_block1a3.port_a_logical_ram_depth = 128;
defparam ram_block1a3.port_a_logical_ram_width = 8;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.ram_block_type = "auto";
defparam ram_block1a3.mem_init0 = 128'h00F8E73366C99B398E1FFFFC3CE6664C;

cycloneiii_ram_block ram_block1a4(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a4_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.init_file = "fft_3n512sin.hex";
defparam ram_block1a4.init_file_layout = "port_a";
defparam ram_block1a4.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_3dp_rom_fft_120:twrom|twid_rom_fft_120:\\gen_M4K:sin_3n|altsyncram:\\gen_auto:altsyncram_component|altsyncram_i191:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.operation_mode = "rom";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 7;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "clock0";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 127;
defparam ram_block1a4.port_a_logical_ram_depth = 128;
defparam ram_block1a4.port_a_logical_ram_width = 8;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.ram_block_type = "auto";
defparam ram_block1a4.mem_init0 = 128'h0007E0F0E1C7870781FFFFFFC0F87870;

cycloneiii_ram_block ram_block1a5(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a5_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.init_file = "fft_3n512sin.hex";
defparam ram_block1a5.init_file_layout = "port_a";
defparam ram_block1a5.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_3dp_rom_fft_120:twrom|twid_rom_fft_120:\\gen_M4K:sin_3n|altsyncram:\\gen_auto:altsyncram_component|altsyncram_i191:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.operation_mode = "rom";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 7;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "clock0";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 127;
defparam ram_block1a5.port_a_logical_ram_depth = 128;
defparam ram_block1a5.port_a_logical_ram_width = 8;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.ram_block_type = "auto";
defparam ram_block1a5.mem_init0 = 128'h00001FF01FC07F007FFFFFFFFF007F80;

cycloneiii_ram_block ram_block1a6(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a6_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.init_file = "fft_3n512sin.hex";
defparam ram_block1a6.init_file_layout = "port_a";
defparam ram_block1a6.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_3dp_rom_fft_120:twrom|twid_rom_fft_120:\\gen_M4K:sin_3n|altsyncram:\\gen_auto:altsyncram_component|altsyncram_i191:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.operation_mode = "rom";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 7;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "clock0";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 127;
defparam ram_block1a6.port_a_logical_ram_depth = 128;
defparam ram_block1a6.port_a_logical_ram_width = 8;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.ram_block_type = "auto";
defparam ram_block1a6.mem_init0 = 128'h0000000FFFC000FFFFFFFFFFFFFF8000;

cycloneiii_ram_block ram_block1a7(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a7_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.init_file = "fft_3n512sin.hex";
defparam ram_block1a7.init_file_layout = "port_a";
defparam ram_block1a7.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_3dp_rom_fft_120:twrom|twid_rom_fft_120:\\gen_M4K:sin_3n|altsyncram:\\gen_auto:altsyncram_component|altsyncram_i191:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.operation_mode = "rom";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 7;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "clock0";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 127;
defparam ram_block1a7.port_a_logical_ram_depth = 128;
defparam ram_block1a7.port_a_logical_ram_width = 8;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.ram_block_type = "auto";
defparam ram_block1a7.mem_init0 = 128'hFFFFFFFFFFC000000000000000000000;

endmodule

module fft_asj_fft_4dp_ram_fft_120 (
	q_b_1,
	q_b_11,
	q_b_12,
	q_b_13,
	q_b_0,
	q_b_01,
	q_b_02,
	q_b_03,
	q_b_7,
	q_b_71,
	q_b_72,
	q_b_73,
	q_b_6,
	q_b_61,
	q_b_62,
	q_b_63,
	q_b_5,
	q_b_51,
	q_b_52,
	q_b_53,
	q_b_4,
	q_b_41,
	q_b_42,
	q_b_43,
	q_b_3,
	q_b_31,
	q_b_32,
	q_b_33,
	q_b_2,
	q_b_21,
	q_b_22,
	q_b_23,
	q_b_9,
	q_b_91,
	q_b_92,
	q_b_93,
	q_b_8,
	q_b_81,
	q_b_82,
	q_b_83,
	q_b_15,
	q_b_151,
	q_b_152,
	q_b_153,
	q_b_14,
	q_b_141,
	q_b_142,
	q_b_143,
	q_b_131,
	q_b_132,
	q_b_133,
	q_b_134,
	q_b_121,
	q_b_122,
	q_b_123,
	q_b_124,
	q_b_111,
	q_b_112,
	q_b_113,
	q_b_114,
	q_b_10,
	q_b_101,
	q_b_102,
	q_b_103,
	ram_in_reg_1_6,
	ram_in_reg_1_5,
	ram_in_reg_1_4,
	ram_in_reg_1_7,
	ram_in_reg_0_6,
	ram_in_reg_0_5,
	ram_in_reg_0_4,
	ram_in_reg_0_7,
	ram_in_reg_7_6,
	ram_in_reg_7_5,
	ram_in_reg_7_4,
	ram_in_reg_7_7,
	ram_in_reg_6_6,
	ram_in_reg_6_5,
	ram_in_reg_6_4,
	ram_in_reg_6_7,
	ram_in_reg_5_6,
	ram_in_reg_5_5,
	ram_in_reg_5_4,
	ram_in_reg_5_7,
	ram_in_reg_4_6,
	ram_in_reg_4_5,
	ram_in_reg_4_4,
	ram_in_reg_4_7,
	ram_in_reg_3_6,
	ram_in_reg_3_5,
	ram_in_reg_3_4,
	ram_in_reg_3_7,
	ram_in_reg_2_6,
	ram_in_reg_2_5,
	ram_in_reg_2_4,
	ram_in_reg_2_7,
	ram_in_reg_1_2,
	ram_in_reg_1_1,
	ram_in_reg_1_0,
	ram_in_reg_1_3,
	ram_in_reg_0_2,
	ram_in_reg_0_1,
	ram_in_reg_0_0,
	ram_in_reg_0_3,
	ram_in_reg_7_2,
	ram_in_reg_7_1,
	ram_in_reg_7_0,
	ram_in_reg_7_3,
	ram_in_reg_6_2,
	ram_in_reg_6_1,
	ram_in_reg_6_0,
	ram_in_reg_6_3,
	ram_in_reg_5_2,
	ram_in_reg_5_1,
	ram_in_reg_5_0,
	ram_in_reg_5_3,
	ram_in_reg_4_2,
	ram_in_reg_4_1,
	ram_in_reg_4_0,
	ram_in_reg_4_3,
	ram_in_reg_3_2,
	ram_in_reg_3_1,
	ram_in_reg_3_0,
	ram_in_reg_3_3,
	ram_in_reg_2_2,
	ram_in_reg_2_1,
	ram_in_reg_2_0,
	ram_in_reg_2_3,
	global_clock_enable,
	wc_vec_6,
	ram_in_reg_0_01,
	ram_in_reg_1_21,
	ram_in_reg_2_01,
	ram_in_reg_3_21,
	ram_in_reg_4_01,
	ram_in_reg_5_21,
	ram_in_reg_6_01,
	rdaddress_c_bus_0,
	rdaddress_c_bus_15,
	rdaddress_c_bus_16,
	rdaddress_c_bus_10,
	rdaddress_c_bus_11,
	rdaddress_c_bus_12,
	rdaddress_c_bus_13,
	ram_in_reg_0_11,
	ram_in_reg_1_11,
	ram_in_reg_2_11,
	ram_in_reg_3_11,
	ram_in_reg_4_11,
	ram_in_reg_5_11,
	rdaddress_c_bus_20,
	ram_in_reg_1_01,
	ram_in_reg_3_01,
	ram_in_reg_5_01,
	ram_in_reg_1_31,
	ram_in_reg_3_31,
	ram_in_reg_5_31,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_1;
output 	q_b_11;
output 	q_b_12;
output 	q_b_13;
output 	q_b_0;
output 	q_b_01;
output 	q_b_02;
output 	q_b_03;
output 	q_b_7;
output 	q_b_71;
output 	q_b_72;
output 	q_b_73;
output 	q_b_6;
output 	q_b_61;
output 	q_b_62;
output 	q_b_63;
output 	q_b_5;
output 	q_b_51;
output 	q_b_52;
output 	q_b_53;
output 	q_b_4;
output 	q_b_41;
output 	q_b_42;
output 	q_b_43;
output 	q_b_3;
output 	q_b_31;
output 	q_b_32;
output 	q_b_33;
output 	q_b_2;
output 	q_b_21;
output 	q_b_22;
output 	q_b_23;
output 	q_b_9;
output 	q_b_91;
output 	q_b_92;
output 	q_b_93;
output 	q_b_8;
output 	q_b_81;
output 	q_b_82;
output 	q_b_83;
output 	q_b_15;
output 	q_b_151;
output 	q_b_152;
output 	q_b_153;
output 	q_b_14;
output 	q_b_141;
output 	q_b_142;
output 	q_b_143;
output 	q_b_131;
output 	q_b_132;
output 	q_b_133;
output 	q_b_134;
output 	q_b_121;
output 	q_b_122;
output 	q_b_123;
output 	q_b_124;
output 	q_b_111;
output 	q_b_112;
output 	q_b_113;
output 	q_b_114;
output 	q_b_10;
output 	q_b_101;
output 	q_b_102;
output 	q_b_103;
input 	ram_in_reg_1_6;
input 	ram_in_reg_1_5;
input 	ram_in_reg_1_4;
input 	ram_in_reg_1_7;
input 	ram_in_reg_0_6;
input 	ram_in_reg_0_5;
input 	ram_in_reg_0_4;
input 	ram_in_reg_0_7;
input 	ram_in_reg_7_6;
input 	ram_in_reg_7_5;
input 	ram_in_reg_7_4;
input 	ram_in_reg_7_7;
input 	ram_in_reg_6_6;
input 	ram_in_reg_6_5;
input 	ram_in_reg_6_4;
input 	ram_in_reg_6_7;
input 	ram_in_reg_5_6;
input 	ram_in_reg_5_5;
input 	ram_in_reg_5_4;
input 	ram_in_reg_5_7;
input 	ram_in_reg_4_6;
input 	ram_in_reg_4_5;
input 	ram_in_reg_4_4;
input 	ram_in_reg_4_7;
input 	ram_in_reg_3_6;
input 	ram_in_reg_3_5;
input 	ram_in_reg_3_4;
input 	ram_in_reg_3_7;
input 	ram_in_reg_2_6;
input 	ram_in_reg_2_5;
input 	ram_in_reg_2_4;
input 	ram_in_reg_2_7;
input 	ram_in_reg_1_2;
input 	ram_in_reg_1_1;
input 	ram_in_reg_1_0;
input 	ram_in_reg_1_3;
input 	ram_in_reg_0_2;
input 	ram_in_reg_0_1;
input 	ram_in_reg_0_0;
input 	ram_in_reg_0_3;
input 	ram_in_reg_7_2;
input 	ram_in_reg_7_1;
input 	ram_in_reg_7_0;
input 	ram_in_reg_7_3;
input 	ram_in_reg_6_2;
input 	ram_in_reg_6_1;
input 	ram_in_reg_6_0;
input 	ram_in_reg_6_3;
input 	ram_in_reg_5_2;
input 	ram_in_reg_5_1;
input 	ram_in_reg_5_0;
input 	ram_in_reg_5_3;
input 	ram_in_reg_4_2;
input 	ram_in_reg_4_1;
input 	ram_in_reg_4_0;
input 	ram_in_reg_4_3;
input 	ram_in_reg_3_2;
input 	ram_in_reg_3_1;
input 	ram_in_reg_3_0;
input 	ram_in_reg_3_3;
input 	ram_in_reg_2_2;
input 	ram_in_reg_2_1;
input 	ram_in_reg_2_0;
input 	ram_in_reg_2_3;
input 	global_clock_enable;
input 	wc_vec_6;
input 	ram_in_reg_0_01;
input 	ram_in_reg_1_21;
input 	ram_in_reg_2_01;
input 	ram_in_reg_3_21;
input 	ram_in_reg_4_01;
input 	ram_in_reg_5_21;
input 	ram_in_reg_6_01;
input 	rdaddress_c_bus_0;
input 	rdaddress_c_bus_15;
input 	rdaddress_c_bus_16;
input 	rdaddress_c_bus_10;
input 	rdaddress_c_bus_11;
input 	rdaddress_c_bus_12;
input 	rdaddress_c_bus_13;
input 	ram_in_reg_0_11;
input 	ram_in_reg_1_11;
input 	ram_in_reg_2_11;
input 	ram_in_reg_3_11;
input 	ram_in_reg_4_11;
input 	ram_in_reg_5_11;
input 	rdaddress_c_bus_20;
input 	ram_in_reg_1_01;
input 	ram_in_reg_3_01;
input 	ram_in_reg_5_01;
input 	ram_in_reg_1_31;
input 	ram_in_reg_3_31;
input 	ram_in_reg_5_31;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_asj_fft_data_ram_fft_120_3 \gen_rams:3:dat_A (
	.q_b_1(q_b_13),
	.q_b_0(q_b_03),
	.q_b_7(q_b_73),
	.q_b_6(q_b_63),
	.q_b_5(q_b_53),
	.q_b_4(q_b_43),
	.q_b_3(q_b_33),
	.q_b_2(q_b_23),
	.q_b_9(q_b_93),
	.q_b_8(q_b_83),
	.q_b_15(q_b_153),
	.q_b_14(q_b_143),
	.q_b_13(q_b_134),
	.q_b_12(q_b_124),
	.q_b_11(q_b_114),
	.q_b_10(q_b_103),
	.ram_in_reg_1_7(ram_in_reg_1_7),
	.ram_in_reg_0_7(ram_in_reg_0_7),
	.ram_in_reg_7_7(ram_in_reg_7_7),
	.ram_in_reg_6_7(ram_in_reg_6_7),
	.ram_in_reg_5_7(ram_in_reg_5_7),
	.ram_in_reg_4_7(ram_in_reg_4_7),
	.ram_in_reg_3_7(ram_in_reg_3_7),
	.ram_in_reg_2_7(ram_in_reg_2_7),
	.ram_in_reg_1_3(ram_in_reg_1_3),
	.ram_in_reg_0_3(ram_in_reg_0_3),
	.ram_in_reg_7_3(ram_in_reg_7_3),
	.ram_in_reg_6_3(ram_in_reg_6_3),
	.ram_in_reg_5_3(ram_in_reg_5_3),
	.ram_in_reg_4_3(ram_in_reg_4_3),
	.ram_in_reg_3_3(ram_in_reg_3_3),
	.ram_in_reg_2_3(ram_in_reg_2_3),
	.global_clock_enable(global_clock_enable),
	.wc_vec_6(wc_vec_6),
	.ram_in_reg_6_0(ram_in_reg_6_01),
	.rdaddress_c_bus_0(rdaddress_c_bus_0),
	.rdaddress_c_bus_15(rdaddress_c_bus_15),
	.rdaddress_c_bus_16(rdaddress_c_bus_16),
	.rdaddress_c_bus_10(rdaddress_c_bus_10),
	.rdaddress_c_bus_11(rdaddress_c_bus_11),
	.rdaddress_c_bus_12(rdaddress_c_bus_12),
	.ram_in_reg_0_1(ram_in_reg_0_11),
	.ram_in_reg_2_1(ram_in_reg_2_11),
	.ram_in_reg_4_1(ram_in_reg_4_11),
	.rdaddress_c_bus_20(rdaddress_c_bus_20),
	.ram_in_reg_1_31(ram_in_reg_1_31),
	.ram_in_reg_3_31(ram_in_reg_3_31),
	.ram_in_reg_5_31(ram_in_reg_5_31),
	.clk(clk));

fft_asj_fft_data_ram_fft_120_2 \gen_rams:2:dat_A (
	.q_b_1(q_b_1),
	.q_b_0(q_b_0),
	.q_b_7(q_b_7),
	.q_b_6(q_b_6),
	.q_b_5(q_b_5),
	.q_b_4(q_b_4),
	.q_b_3(q_b_3),
	.q_b_2(q_b_2),
	.q_b_9(q_b_9),
	.q_b_8(q_b_8),
	.q_b_15(q_b_15),
	.q_b_14(q_b_14),
	.q_b_13(q_b_131),
	.q_b_12(q_b_121),
	.q_b_11(q_b_111),
	.q_b_10(q_b_10),
	.ram_in_reg_1_6(ram_in_reg_1_6),
	.ram_in_reg_0_6(ram_in_reg_0_6),
	.ram_in_reg_7_6(ram_in_reg_7_6),
	.ram_in_reg_6_6(ram_in_reg_6_6),
	.ram_in_reg_5_6(ram_in_reg_5_6),
	.ram_in_reg_4_6(ram_in_reg_4_6),
	.ram_in_reg_3_6(ram_in_reg_3_6),
	.ram_in_reg_2_6(ram_in_reg_2_6),
	.ram_in_reg_1_2(ram_in_reg_1_2),
	.ram_in_reg_0_2(ram_in_reg_0_2),
	.ram_in_reg_7_2(ram_in_reg_7_2),
	.ram_in_reg_6_2(ram_in_reg_6_2),
	.ram_in_reg_5_2(ram_in_reg_5_2),
	.ram_in_reg_4_2(ram_in_reg_4_2),
	.ram_in_reg_3_2(ram_in_reg_3_2),
	.ram_in_reg_2_2(ram_in_reg_2_2),
	.global_clock_enable(global_clock_enable),
	.wc_vec_6(wc_vec_6),
	.ram_in_reg_0_0(ram_in_reg_0_01),
	.ram_in_reg_1_21(ram_in_reg_1_21),
	.ram_in_reg_2_0(ram_in_reg_2_01),
	.ram_in_reg_3_21(ram_in_reg_3_21),
	.ram_in_reg_4_0(ram_in_reg_4_01),
	.ram_in_reg_5_21(ram_in_reg_5_21),
	.ram_in_reg_6_0(ram_in_reg_6_01),
	.rdaddress_c_bus_0(rdaddress_c_bus_0),
	.rdaddress_c_bus_15(rdaddress_c_bus_15),
	.rdaddress_c_bus_16(rdaddress_c_bus_16),
	.rdaddress_c_bus_10(rdaddress_c_bus_10),
	.rdaddress_c_bus_11(rdaddress_c_bus_11),
	.rdaddress_c_bus_12(rdaddress_c_bus_12),
	.rdaddress_c_bus_13(rdaddress_c_bus_13),
	.clk(clk));

fft_asj_fft_data_ram_fft_120_1 \gen_rams:1:dat_A (
	.q_b_1(q_b_11),
	.q_b_0(q_b_01),
	.q_b_7(q_b_71),
	.q_b_6(q_b_61),
	.q_b_5(q_b_51),
	.q_b_4(q_b_41),
	.q_b_3(q_b_31),
	.q_b_2(q_b_21),
	.q_b_9(q_b_91),
	.q_b_8(q_b_81),
	.q_b_15(q_b_151),
	.q_b_14(q_b_141),
	.q_b_13(q_b_132),
	.q_b_12(q_b_122),
	.q_b_11(q_b_112),
	.q_b_10(q_b_101),
	.ram_in_reg_1_5(ram_in_reg_1_5),
	.ram_in_reg_0_5(ram_in_reg_0_5),
	.ram_in_reg_7_5(ram_in_reg_7_5),
	.ram_in_reg_6_5(ram_in_reg_6_5),
	.ram_in_reg_5_5(ram_in_reg_5_5),
	.ram_in_reg_4_5(ram_in_reg_4_5),
	.ram_in_reg_3_5(ram_in_reg_3_5),
	.ram_in_reg_2_5(ram_in_reg_2_5),
	.ram_in_reg_1_1(ram_in_reg_1_1),
	.ram_in_reg_0_1(ram_in_reg_0_1),
	.ram_in_reg_7_1(ram_in_reg_7_1),
	.ram_in_reg_6_1(ram_in_reg_6_1),
	.ram_in_reg_5_1(ram_in_reg_5_1),
	.ram_in_reg_4_1(ram_in_reg_4_1),
	.ram_in_reg_3_1(ram_in_reg_3_1),
	.ram_in_reg_2_1(ram_in_reg_2_1),
	.global_clock_enable(global_clock_enable),
	.wc_vec_6(wc_vec_6),
	.ram_in_reg_6_0(ram_in_reg_6_01),
	.rdaddress_c_bus_0(rdaddress_c_bus_0),
	.rdaddress_c_bus_15(rdaddress_c_bus_15),
	.rdaddress_c_bus_16(rdaddress_c_bus_16),
	.rdaddress_c_bus_10(rdaddress_c_bus_10),
	.rdaddress_c_bus_11(rdaddress_c_bus_11),
	.rdaddress_c_bus_12(rdaddress_c_bus_12),
	.ram_in_reg_0_11(ram_in_reg_0_11),
	.ram_in_reg_1_11(ram_in_reg_1_11),
	.ram_in_reg_2_11(ram_in_reg_2_11),
	.ram_in_reg_3_11(ram_in_reg_3_11),
	.ram_in_reg_4_11(ram_in_reg_4_11),
	.ram_in_reg_5_11(ram_in_reg_5_11),
	.rdaddress_c_bus_20(rdaddress_c_bus_20),
	.clk(clk));

fft_asj_fft_data_ram_fft_120 \gen_rams:0:dat_A (
	.q_b_1(q_b_12),
	.q_b_0(q_b_02),
	.q_b_7(q_b_72),
	.q_b_6(q_b_62),
	.q_b_5(q_b_52),
	.q_b_4(q_b_42),
	.q_b_3(q_b_32),
	.q_b_2(q_b_22),
	.q_b_9(q_b_92),
	.q_b_8(q_b_82),
	.q_b_15(q_b_152),
	.q_b_14(q_b_142),
	.q_b_13(q_b_133),
	.q_b_12(q_b_123),
	.q_b_11(q_b_113),
	.q_b_10(q_b_102),
	.ram_in_reg_1_4(ram_in_reg_1_4),
	.ram_in_reg_0_4(ram_in_reg_0_4),
	.ram_in_reg_7_4(ram_in_reg_7_4),
	.ram_in_reg_6_4(ram_in_reg_6_4),
	.ram_in_reg_5_4(ram_in_reg_5_4),
	.ram_in_reg_4_4(ram_in_reg_4_4),
	.ram_in_reg_3_4(ram_in_reg_3_4),
	.ram_in_reg_2_4(ram_in_reg_2_4),
	.ram_in_reg_1_0(ram_in_reg_1_0),
	.ram_in_reg_0_0(ram_in_reg_0_0),
	.ram_in_reg_7_0(ram_in_reg_7_0),
	.ram_in_reg_6_0(ram_in_reg_6_0),
	.ram_in_reg_5_0(ram_in_reg_5_0),
	.ram_in_reg_4_0(ram_in_reg_4_0),
	.ram_in_reg_3_0(ram_in_reg_3_0),
	.ram_in_reg_2_0(ram_in_reg_2_0),
	.global_clock_enable(global_clock_enable),
	.wc_vec_6(wc_vec_6),
	.ram_in_reg_0_01(ram_in_reg_0_01),
	.ram_in_reg_2_01(ram_in_reg_2_01),
	.ram_in_reg_4_01(ram_in_reg_4_01),
	.ram_in_reg_6_01(ram_in_reg_6_01),
	.rdaddress_c_bus_0(rdaddress_c_bus_0),
	.rdaddress_c_bus_15(rdaddress_c_bus_15),
	.rdaddress_c_bus_16(rdaddress_c_bus_16),
	.rdaddress_c_bus_10(rdaddress_c_bus_10),
	.rdaddress_c_bus_11(rdaddress_c_bus_11),
	.rdaddress_c_bus_12(rdaddress_c_bus_12),
	.rdaddress_c_bus_13(rdaddress_c_bus_13),
	.ram_in_reg_1_01(ram_in_reg_1_01),
	.ram_in_reg_3_01(ram_in_reg_3_01),
	.ram_in_reg_5_01(ram_in_reg_5_01),
	.clk(clk));

endmodule

module fft_asj_fft_data_ram_fft_120 (
	q_b_1,
	q_b_0,
	q_b_7,
	q_b_6,
	q_b_5,
	q_b_4,
	q_b_3,
	q_b_2,
	q_b_9,
	q_b_8,
	q_b_15,
	q_b_14,
	q_b_13,
	q_b_12,
	q_b_11,
	q_b_10,
	ram_in_reg_1_4,
	ram_in_reg_0_4,
	ram_in_reg_7_4,
	ram_in_reg_6_4,
	ram_in_reg_5_4,
	ram_in_reg_4_4,
	ram_in_reg_3_4,
	ram_in_reg_2_4,
	ram_in_reg_1_0,
	ram_in_reg_0_0,
	ram_in_reg_7_0,
	ram_in_reg_6_0,
	ram_in_reg_5_0,
	ram_in_reg_4_0,
	ram_in_reg_3_0,
	ram_in_reg_2_0,
	global_clock_enable,
	wc_vec_6,
	ram_in_reg_0_01,
	ram_in_reg_2_01,
	ram_in_reg_4_01,
	ram_in_reg_6_01,
	rdaddress_c_bus_0,
	rdaddress_c_bus_15,
	rdaddress_c_bus_16,
	rdaddress_c_bus_10,
	rdaddress_c_bus_11,
	rdaddress_c_bus_12,
	rdaddress_c_bus_13,
	ram_in_reg_1_01,
	ram_in_reg_3_01,
	ram_in_reg_5_01,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_1;
output 	q_b_0;
output 	q_b_7;
output 	q_b_6;
output 	q_b_5;
output 	q_b_4;
output 	q_b_3;
output 	q_b_2;
output 	q_b_9;
output 	q_b_8;
output 	q_b_15;
output 	q_b_14;
output 	q_b_13;
output 	q_b_12;
output 	q_b_11;
output 	q_b_10;
input 	ram_in_reg_1_4;
input 	ram_in_reg_0_4;
input 	ram_in_reg_7_4;
input 	ram_in_reg_6_4;
input 	ram_in_reg_5_4;
input 	ram_in_reg_4_4;
input 	ram_in_reg_3_4;
input 	ram_in_reg_2_4;
input 	ram_in_reg_1_0;
input 	ram_in_reg_0_0;
input 	ram_in_reg_7_0;
input 	ram_in_reg_6_0;
input 	ram_in_reg_5_0;
input 	ram_in_reg_4_0;
input 	ram_in_reg_3_0;
input 	ram_in_reg_2_0;
input 	global_clock_enable;
input 	wc_vec_6;
input 	ram_in_reg_0_01;
input 	ram_in_reg_2_01;
input 	ram_in_reg_4_01;
input 	ram_in_reg_6_01;
input 	rdaddress_c_bus_0;
input 	rdaddress_c_bus_15;
input 	rdaddress_c_bus_16;
input 	rdaddress_c_bus_10;
input 	rdaddress_c_bus_11;
input 	rdaddress_c_bus_12;
input 	rdaddress_c_bus_13;
input 	ram_in_reg_1_01;
input 	ram_in_reg_3_01;
input 	ram_in_reg_5_01;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_altsyncram_7 \gen_M4K:altsyncram_component (
	.q_b({q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.data_a({ram_in_reg_7_0,ram_in_reg_6_0,ram_in_reg_5_0,ram_in_reg_4_0,ram_in_reg_3_0,ram_in_reg_2_0,ram_in_reg_1_0,ram_in_reg_0_0,ram_in_reg_7_4,ram_in_reg_6_4,ram_in_reg_5_4,ram_in_reg_4_4,ram_in_reg_3_4,ram_in_reg_2_4,ram_in_reg_1_4,ram_in_reg_0_4}),
	.clocken0(global_clock_enable),
	.wren_a(wc_vec_6),
	.address_a({ram_in_reg_6_01,ram_in_reg_5_01,ram_in_reg_4_01,ram_in_reg_3_01,ram_in_reg_2_01,ram_in_reg_1_01,ram_in_reg_0_01}),
	.address_b({rdaddress_c_bus_13,rdaddress_c_bus_12,rdaddress_c_bus_11,rdaddress_c_bus_10,rdaddress_c_bus_16,rdaddress_c_bus_15,rdaddress_c_bus_0}),
	.clock0(clk));

endmodule

module fft_altsyncram_7 (
	q_b,
	data_a,
	clocken0,
	wren_a,
	address_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	[15:0] data_a;
input 	clocken0;
input 	wren_a;
input 	[6:0] address_a;
input 	[6:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_altsyncram_lmu3 auto_generated(
	.q_b({q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.data_a({data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.clocken0(clocken0),
	.wren_a(wren_a),
	.address_a({address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.clock0(clock0));

endmodule

module fft_altsyncram_lmu3 (
	q_b,
	data_a,
	clocken0,
	wren_a,
	address_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	[15:0] data_a;
input 	clocken0;
input 	wren_a;
input 	[6:0] address_a;
input 	[6:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

cycloneiii_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "old";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 7;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 127;
defparam ram_block1a1.port_a_logical_ram_depth = 128;
defparam ram_block1a1.port_a_logical_ram_width = 16;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 7;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "clock0";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 127;
defparam ram_block1a1.port_b_logical_ram_depth = 128;
defparam ram_block1a1.port_b_logical_ram_width = 16;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "old";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 7;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 127;
defparam ram_block1a0.port_a_logical_ram_depth = 128;
defparam ram_block1a0.port_a_logical_ram_width = 16;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 7;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "clock0";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 127;
defparam ram_block1a0.port_b_logical_ram_depth = 128;
defparam ram_block1a0.port_b_logical_ram_width = 16;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "old";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 7;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 127;
defparam ram_block1a7.port_a_logical_ram_depth = 128;
defparam ram_block1a7.port_a_logical_ram_width = 16;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 7;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "clock0";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 127;
defparam ram_block1a7.port_b_logical_ram_depth = 128;
defparam ram_block1a7.port_b_logical_ram_width = 16;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "old";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 7;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 127;
defparam ram_block1a6.port_a_logical_ram_depth = 128;
defparam ram_block1a6.port_a_logical_ram_width = 16;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 7;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "clock0";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 127;
defparam ram_block1a6.port_b_logical_ram_depth = 128;
defparam ram_block1a6.port_b_logical_ram_width = 16;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "old";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 7;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 127;
defparam ram_block1a5.port_a_logical_ram_depth = 128;
defparam ram_block1a5.port_a_logical_ram_width = 16;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 7;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "clock0";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 127;
defparam ram_block1a5.port_b_logical_ram_depth = 128;
defparam ram_block1a5.port_b_logical_ram_width = 16;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "old";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 7;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 127;
defparam ram_block1a4.port_a_logical_ram_depth = 128;
defparam ram_block1a4.port_a_logical_ram_width = 16;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 7;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "clock0";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 127;
defparam ram_block1a4.port_b_logical_ram_depth = 128;
defparam ram_block1a4.port_b_logical_ram_width = 16;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "old";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 7;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 127;
defparam ram_block1a3.port_a_logical_ram_depth = 128;
defparam ram_block1a3.port_a_logical_ram_width = 16;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 7;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "clock0";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 127;
defparam ram_block1a3.port_b_logical_ram_depth = 128;
defparam ram_block1a3.port_b_logical_ram_width = 16;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "old";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 7;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 127;
defparam ram_block1a2.port_a_logical_ram_depth = 128;
defparam ram_block1a2.port_a_logical_ram_width = 16;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 7;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "clock0";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 127;
defparam ram_block1a2.port_b_logical_ram_depth = 128;
defparam ram_block1a2.port_b_logical_ram_width = 16;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.clk0_output_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "old";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 7;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 127;
defparam ram_block1a9.port_a_logical_ram_depth = 128;
defparam ram_block1a9.port_a_logical_ram_width = 16;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 7;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "clock0";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 127;
defparam ram_block1a9.port_b_logical_ram_depth = 128;
defparam ram_block1a9.port_b_logical_ram_width = 16;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.clk0_output_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "old";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 7;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 127;
defparam ram_block1a8.port_a_logical_ram_depth = 128;
defparam ram_block1a8.port_a_logical_ram_width = 16;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 7;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "clock0";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 127;
defparam ram_block1a8.port_b_logical_ram_depth = 128;
defparam ram_block1a8.port_b_logical_ram_width = 16;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.clk0_output_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "old";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 7;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 127;
defparam ram_block1a15.port_a_logical_ram_depth = 128;
defparam ram_block1a15.port_a_logical_ram_width = 16;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 7;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "clock0";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 127;
defparam ram_block1a15.port_b_logical_ram_depth = 128;
defparam ram_block1a15.port_b_logical_ram_width = 16;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.clk0_output_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "old";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 7;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 127;
defparam ram_block1a14.port_a_logical_ram_depth = 128;
defparam ram_block1a14.port_a_logical_ram_width = 16;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 7;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "clock0";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 127;
defparam ram_block1a14.port_b_logical_ram_depth = 128;
defparam ram_block1a14.port_b_logical_ram_width = 16;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.clk0_output_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "old";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 7;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 127;
defparam ram_block1a13.port_a_logical_ram_depth = 128;
defparam ram_block1a13.port_a_logical_ram_width = 16;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 7;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "clock0";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 127;
defparam ram_block1a13.port_b_logical_ram_depth = 128;
defparam ram_block1a13.port_b_logical_ram_width = 16;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.clk0_output_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "old";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 7;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 127;
defparam ram_block1a12.port_a_logical_ram_depth = 128;
defparam ram_block1a12.port_a_logical_ram_width = 16;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 7;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "clock0";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 127;
defparam ram_block1a12.port_b_logical_ram_depth = 128;
defparam ram_block1a12.port_b_logical_ram_width = 16;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.clk0_output_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "old";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 7;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 127;
defparam ram_block1a11.port_a_logical_ram_depth = 128;
defparam ram_block1a11.port_a_logical_ram_width = 16;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 7;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "clock0";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 127;
defparam ram_block1a11.port_b_logical_ram_depth = 128;
defparam ram_block1a11.port_b_logical_ram_width = 16;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.clk0_output_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "old";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 7;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 127;
defparam ram_block1a10.port_a_logical_ram_depth = 128;
defparam ram_block1a10.port_a_logical_ram_width = 16;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 7;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "clock0";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 127;
defparam ram_block1a10.port_b_logical_ram_depth = 128;
defparam ram_block1a10.port_b_logical_ram_width = 16;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";

endmodule

module fft_asj_fft_data_ram_fft_120_1 (
	q_b_1,
	q_b_0,
	q_b_7,
	q_b_6,
	q_b_5,
	q_b_4,
	q_b_3,
	q_b_2,
	q_b_9,
	q_b_8,
	q_b_15,
	q_b_14,
	q_b_13,
	q_b_12,
	q_b_11,
	q_b_10,
	ram_in_reg_1_5,
	ram_in_reg_0_5,
	ram_in_reg_7_5,
	ram_in_reg_6_5,
	ram_in_reg_5_5,
	ram_in_reg_4_5,
	ram_in_reg_3_5,
	ram_in_reg_2_5,
	ram_in_reg_1_1,
	ram_in_reg_0_1,
	ram_in_reg_7_1,
	ram_in_reg_6_1,
	ram_in_reg_5_1,
	ram_in_reg_4_1,
	ram_in_reg_3_1,
	ram_in_reg_2_1,
	global_clock_enable,
	wc_vec_6,
	ram_in_reg_6_0,
	rdaddress_c_bus_0,
	rdaddress_c_bus_15,
	rdaddress_c_bus_16,
	rdaddress_c_bus_10,
	rdaddress_c_bus_11,
	rdaddress_c_bus_12,
	ram_in_reg_0_11,
	ram_in_reg_1_11,
	ram_in_reg_2_11,
	ram_in_reg_3_11,
	ram_in_reg_4_11,
	ram_in_reg_5_11,
	rdaddress_c_bus_20,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_1;
output 	q_b_0;
output 	q_b_7;
output 	q_b_6;
output 	q_b_5;
output 	q_b_4;
output 	q_b_3;
output 	q_b_2;
output 	q_b_9;
output 	q_b_8;
output 	q_b_15;
output 	q_b_14;
output 	q_b_13;
output 	q_b_12;
output 	q_b_11;
output 	q_b_10;
input 	ram_in_reg_1_5;
input 	ram_in_reg_0_5;
input 	ram_in_reg_7_5;
input 	ram_in_reg_6_5;
input 	ram_in_reg_5_5;
input 	ram_in_reg_4_5;
input 	ram_in_reg_3_5;
input 	ram_in_reg_2_5;
input 	ram_in_reg_1_1;
input 	ram_in_reg_0_1;
input 	ram_in_reg_7_1;
input 	ram_in_reg_6_1;
input 	ram_in_reg_5_1;
input 	ram_in_reg_4_1;
input 	ram_in_reg_3_1;
input 	ram_in_reg_2_1;
input 	global_clock_enable;
input 	wc_vec_6;
input 	ram_in_reg_6_0;
input 	rdaddress_c_bus_0;
input 	rdaddress_c_bus_15;
input 	rdaddress_c_bus_16;
input 	rdaddress_c_bus_10;
input 	rdaddress_c_bus_11;
input 	rdaddress_c_bus_12;
input 	ram_in_reg_0_11;
input 	ram_in_reg_1_11;
input 	ram_in_reg_2_11;
input 	ram_in_reg_3_11;
input 	ram_in_reg_4_11;
input 	ram_in_reg_5_11;
input 	rdaddress_c_bus_20;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_altsyncram_8 \gen_M4K:altsyncram_component (
	.q_b({q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.data_a({ram_in_reg_7_1,ram_in_reg_6_1,ram_in_reg_5_1,ram_in_reg_4_1,ram_in_reg_3_1,ram_in_reg_2_1,ram_in_reg_1_1,ram_in_reg_0_1,ram_in_reg_7_5,ram_in_reg_6_5,ram_in_reg_5_5,ram_in_reg_4_5,ram_in_reg_3_5,ram_in_reg_2_5,ram_in_reg_1_5,ram_in_reg_0_5}),
	.clocken0(global_clock_enable),
	.wren_a(wc_vec_6),
	.address_a({ram_in_reg_6_0,ram_in_reg_5_11,ram_in_reg_4_11,ram_in_reg_3_11,ram_in_reg_2_11,ram_in_reg_1_11,ram_in_reg_0_11}),
	.address_b({rdaddress_c_bus_20,rdaddress_c_bus_12,rdaddress_c_bus_11,rdaddress_c_bus_10,rdaddress_c_bus_16,rdaddress_c_bus_15,rdaddress_c_bus_0}),
	.clock0(clk));

endmodule

module fft_altsyncram_8 (
	q_b,
	data_a,
	clocken0,
	wren_a,
	address_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	[15:0] data_a;
input 	clocken0;
input 	wren_a;
input 	[6:0] address_a;
input 	[6:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_altsyncram_lmu3_1 auto_generated(
	.q_b({q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.data_a({data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.clocken0(clocken0),
	.wren_a(wren_a),
	.address_a({address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.clock0(clock0));

endmodule

module fft_altsyncram_lmu3_1 (
	q_b,
	data_a,
	clocken0,
	wren_a,
	address_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	[15:0] data_a;
input 	clocken0;
input 	wren_a;
input 	[6:0] address_a;
input 	[6:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

cycloneiii_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "old";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 7;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 127;
defparam ram_block1a1.port_a_logical_ram_depth = 128;
defparam ram_block1a1.port_a_logical_ram_width = 16;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 7;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "clock0";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 127;
defparam ram_block1a1.port_b_logical_ram_depth = 128;
defparam ram_block1a1.port_b_logical_ram_width = 16;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "old";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 7;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 127;
defparam ram_block1a0.port_a_logical_ram_depth = 128;
defparam ram_block1a0.port_a_logical_ram_width = 16;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 7;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "clock0";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 127;
defparam ram_block1a0.port_b_logical_ram_depth = 128;
defparam ram_block1a0.port_b_logical_ram_width = 16;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "old";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 7;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 127;
defparam ram_block1a7.port_a_logical_ram_depth = 128;
defparam ram_block1a7.port_a_logical_ram_width = 16;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 7;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "clock0";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 127;
defparam ram_block1a7.port_b_logical_ram_depth = 128;
defparam ram_block1a7.port_b_logical_ram_width = 16;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "old";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 7;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 127;
defparam ram_block1a6.port_a_logical_ram_depth = 128;
defparam ram_block1a6.port_a_logical_ram_width = 16;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 7;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "clock0";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 127;
defparam ram_block1a6.port_b_logical_ram_depth = 128;
defparam ram_block1a6.port_b_logical_ram_width = 16;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "old";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 7;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 127;
defparam ram_block1a5.port_a_logical_ram_depth = 128;
defparam ram_block1a5.port_a_logical_ram_width = 16;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 7;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "clock0";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 127;
defparam ram_block1a5.port_b_logical_ram_depth = 128;
defparam ram_block1a5.port_b_logical_ram_width = 16;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "old";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 7;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 127;
defparam ram_block1a4.port_a_logical_ram_depth = 128;
defparam ram_block1a4.port_a_logical_ram_width = 16;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 7;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "clock0";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 127;
defparam ram_block1a4.port_b_logical_ram_depth = 128;
defparam ram_block1a4.port_b_logical_ram_width = 16;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "old";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 7;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 127;
defparam ram_block1a3.port_a_logical_ram_depth = 128;
defparam ram_block1a3.port_a_logical_ram_width = 16;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 7;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "clock0";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 127;
defparam ram_block1a3.port_b_logical_ram_depth = 128;
defparam ram_block1a3.port_b_logical_ram_width = 16;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "old";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 7;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 127;
defparam ram_block1a2.port_a_logical_ram_depth = 128;
defparam ram_block1a2.port_a_logical_ram_width = 16;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 7;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "clock0";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 127;
defparam ram_block1a2.port_b_logical_ram_depth = 128;
defparam ram_block1a2.port_b_logical_ram_width = 16;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.clk0_output_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "old";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 7;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 127;
defparam ram_block1a9.port_a_logical_ram_depth = 128;
defparam ram_block1a9.port_a_logical_ram_width = 16;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 7;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "clock0";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 127;
defparam ram_block1a9.port_b_logical_ram_depth = 128;
defparam ram_block1a9.port_b_logical_ram_width = 16;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.clk0_output_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "old";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 7;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 127;
defparam ram_block1a8.port_a_logical_ram_depth = 128;
defparam ram_block1a8.port_a_logical_ram_width = 16;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 7;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "clock0";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 127;
defparam ram_block1a8.port_b_logical_ram_depth = 128;
defparam ram_block1a8.port_b_logical_ram_width = 16;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.clk0_output_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "old";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 7;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 127;
defparam ram_block1a15.port_a_logical_ram_depth = 128;
defparam ram_block1a15.port_a_logical_ram_width = 16;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 7;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "clock0";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 127;
defparam ram_block1a15.port_b_logical_ram_depth = 128;
defparam ram_block1a15.port_b_logical_ram_width = 16;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.clk0_output_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "old";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 7;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 127;
defparam ram_block1a14.port_a_logical_ram_depth = 128;
defparam ram_block1a14.port_a_logical_ram_width = 16;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 7;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "clock0";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 127;
defparam ram_block1a14.port_b_logical_ram_depth = 128;
defparam ram_block1a14.port_b_logical_ram_width = 16;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.clk0_output_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "old";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 7;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 127;
defparam ram_block1a13.port_a_logical_ram_depth = 128;
defparam ram_block1a13.port_a_logical_ram_width = 16;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 7;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "clock0";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 127;
defparam ram_block1a13.port_b_logical_ram_depth = 128;
defparam ram_block1a13.port_b_logical_ram_width = 16;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.clk0_output_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "old";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 7;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 127;
defparam ram_block1a12.port_a_logical_ram_depth = 128;
defparam ram_block1a12.port_a_logical_ram_width = 16;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 7;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "clock0";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 127;
defparam ram_block1a12.port_b_logical_ram_depth = 128;
defparam ram_block1a12.port_b_logical_ram_width = 16;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.clk0_output_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "old";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 7;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 127;
defparam ram_block1a11.port_a_logical_ram_depth = 128;
defparam ram_block1a11.port_a_logical_ram_width = 16;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 7;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "clock0";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 127;
defparam ram_block1a11.port_b_logical_ram_depth = 128;
defparam ram_block1a11.port_b_logical_ram_width = 16;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.clk0_output_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "old";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 7;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 127;
defparam ram_block1a10.port_a_logical_ram_depth = 128;
defparam ram_block1a10.port_a_logical_ram_width = 16;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 7;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "clock0";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 127;
defparam ram_block1a10.port_b_logical_ram_depth = 128;
defparam ram_block1a10.port_b_logical_ram_width = 16;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";

endmodule

module fft_asj_fft_data_ram_fft_120_2 (
	q_b_1,
	q_b_0,
	q_b_7,
	q_b_6,
	q_b_5,
	q_b_4,
	q_b_3,
	q_b_2,
	q_b_9,
	q_b_8,
	q_b_15,
	q_b_14,
	q_b_13,
	q_b_12,
	q_b_11,
	q_b_10,
	ram_in_reg_1_6,
	ram_in_reg_0_6,
	ram_in_reg_7_6,
	ram_in_reg_6_6,
	ram_in_reg_5_6,
	ram_in_reg_4_6,
	ram_in_reg_3_6,
	ram_in_reg_2_6,
	ram_in_reg_1_2,
	ram_in_reg_0_2,
	ram_in_reg_7_2,
	ram_in_reg_6_2,
	ram_in_reg_5_2,
	ram_in_reg_4_2,
	ram_in_reg_3_2,
	ram_in_reg_2_2,
	global_clock_enable,
	wc_vec_6,
	ram_in_reg_0_0,
	ram_in_reg_1_21,
	ram_in_reg_2_0,
	ram_in_reg_3_21,
	ram_in_reg_4_0,
	ram_in_reg_5_21,
	ram_in_reg_6_0,
	rdaddress_c_bus_0,
	rdaddress_c_bus_15,
	rdaddress_c_bus_16,
	rdaddress_c_bus_10,
	rdaddress_c_bus_11,
	rdaddress_c_bus_12,
	rdaddress_c_bus_13,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_1;
output 	q_b_0;
output 	q_b_7;
output 	q_b_6;
output 	q_b_5;
output 	q_b_4;
output 	q_b_3;
output 	q_b_2;
output 	q_b_9;
output 	q_b_8;
output 	q_b_15;
output 	q_b_14;
output 	q_b_13;
output 	q_b_12;
output 	q_b_11;
output 	q_b_10;
input 	ram_in_reg_1_6;
input 	ram_in_reg_0_6;
input 	ram_in_reg_7_6;
input 	ram_in_reg_6_6;
input 	ram_in_reg_5_6;
input 	ram_in_reg_4_6;
input 	ram_in_reg_3_6;
input 	ram_in_reg_2_6;
input 	ram_in_reg_1_2;
input 	ram_in_reg_0_2;
input 	ram_in_reg_7_2;
input 	ram_in_reg_6_2;
input 	ram_in_reg_5_2;
input 	ram_in_reg_4_2;
input 	ram_in_reg_3_2;
input 	ram_in_reg_2_2;
input 	global_clock_enable;
input 	wc_vec_6;
input 	ram_in_reg_0_0;
input 	ram_in_reg_1_21;
input 	ram_in_reg_2_0;
input 	ram_in_reg_3_21;
input 	ram_in_reg_4_0;
input 	ram_in_reg_5_21;
input 	ram_in_reg_6_0;
input 	rdaddress_c_bus_0;
input 	rdaddress_c_bus_15;
input 	rdaddress_c_bus_16;
input 	rdaddress_c_bus_10;
input 	rdaddress_c_bus_11;
input 	rdaddress_c_bus_12;
input 	rdaddress_c_bus_13;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_altsyncram_9 \gen_M4K:altsyncram_component (
	.q_b({q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.data_a({ram_in_reg_7_2,ram_in_reg_6_2,ram_in_reg_5_2,ram_in_reg_4_2,ram_in_reg_3_2,ram_in_reg_2_2,ram_in_reg_1_2,ram_in_reg_0_2,ram_in_reg_7_6,ram_in_reg_6_6,ram_in_reg_5_6,ram_in_reg_4_6,ram_in_reg_3_6,ram_in_reg_2_6,ram_in_reg_1_6,ram_in_reg_0_6}),
	.clocken0(global_clock_enable),
	.wren_a(wc_vec_6),
	.address_a({ram_in_reg_6_0,ram_in_reg_5_21,ram_in_reg_4_0,ram_in_reg_3_21,ram_in_reg_2_0,ram_in_reg_1_21,ram_in_reg_0_0}),
	.address_b({rdaddress_c_bus_13,rdaddress_c_bus_12,rdaddress_c_bus_11,rdaddress_c_bus_10,rdaddress_c_bus_16,rdaddress_c_bus_15,rdaddress_c_bus_0}),
	.clock0(clk));

endmodule

module fft_altsyncram_9 (
	q_b,
	data_a,
	clocken0,
	wren_a,
	address_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	[15:0] data_a;
input 	clocken0;
input 	wren_a;
input 	[6:0] address_a;
input 	[6:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_altsyncram_lmu3_2 auto_generated(
	.q_b({q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.data_a({data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.clocken0(clocken0),
	.wren_a(wren_a),
	.address_a({address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.clock0(clock0));

endmodule

module fft_altsyncram_lmu3_2 (
	q_b,
	data_a,
	clocken0,
	wren_a,
	address_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	[15:0] data_a;
input 	clocken0;
input 	wren_a;
input 	[6:0] address_a;
input 	[6:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

cycloneiii_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "old";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 7;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 127;
defparam ram_block1a1.port_a_logical_ram_depth = 128;
defparam ram_block1a1.port_a_logical_ram_width = 16;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 7;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "clock0";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 127;
defparam ram_block1a1.port_b_logical_ram_depth = 128;
defparam ram_block1a1.port_b_logical_ram_width = 16;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "old";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 7;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 127;
defparam ram_block1a0.port_a_logical_ram_depth = 128;
defparam ram_block1a0.port_a_logical_ram_width = 16;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 7;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "clock0";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 127;
defparam ram_block1a0.port_b_logical_ram_depth = 128;
defparam ram_block1a0.port_b_logical_ram_width = 16;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "old";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 7;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 127;
defparam ram_block1a7.port_a_logical_ram_depth = 128;
defparam ram_block1a7.port_a_logical_ram_width = 16;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 7;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "clock0";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 127;
defparam ram_block1a7.port_b_logical_ram_depth = 128;
defparam ram_block1a7.port_b_logical_ram_width = 16;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "old";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 7;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 127;
defparam ram_block1a6.port_a_logical_ram_depth = 128;
defparam ram_block1a6.port_a_logical_ram_width = 16;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 7;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "clock0";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 127;
defparam ram_block1a6.port_b_logical_ram_depth = 128;
defparam ram_block1a6.port_b_logical_ram_width = 16;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "old";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 7;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 127;
defparam ram_block1a5.port_a_logical_ram_depth = 128;
defparam ram_block1a5.port_a_logical_ram_width = 16;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 7;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "clock0";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 127;
defparam ram_block1a5.port_b_logical_ram_depth = 128;
defparam ram_block1a5.port_b_logical_ram_width = 16;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "old";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 7;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 127;
defparam ram_block1a4.port_a_logical_ram_depth = 128;
defparam ram_block1a4.port_a_logical_ram_width = 16;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 7;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "clock0";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 127;
defparam ram_block1a4.port_b_logical_ram_depth = 128;
defparam ram_block1a4.port_b_logical_ram_width = 16;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "old";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 7;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 127;
defparam ram_block1a3.port_a_logical_ram_depth = 128;
defparam ram_block1a3.port_a_logical_ram_width = 16;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 7;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "clock0";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 127;
defparam ram_block1a3.port_b_logical_ram_depth = 128;
defparam ram_block1a3.port_b_logical_ram_width = 16;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "old";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 7;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 127;
defparam ram_block1a2.port_a_logical_ram_depth = 128;
defparam ram_block1a2.port_a_logical_ram_width = 16;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 7;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "clock0";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 127;
defparam ram_block1a2.port_b_logical_ram_depth = 128;
defparam ram_block1a2.port_b_logical_ram_width = 16;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.clk0_output_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "old";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 7;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 127;
defparam ram_block1a9.port_a_logical_ram_depth = 128;
defparam ram_block1a9.port_a_logical_ram_width = 16;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 7;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "clock0";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 127;
defparam ram_block1a9.port_b_logical_ram_depth = 128;
defparam ram_block1a9.port_b_logical_ram_width = 16;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.clk0_output_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "old";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 7;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 127;
defparam ram_block1a8.port_a_logical_ram_depth = 128;
defparam ram_block1a8.port_a_logical_ram_width = 16;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 7;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "clock0";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 127;
defparam ram_block1a8.port_b_logical_ram_depth = 128;
defparam ram_block1a8.port_b_logical_ram_width = 16;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.clk0_output_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "old";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 7;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 127;
defparam ram_block1a15.port_a_logical_ram_depth = 128;
defparam ram_block1a15.port_a_logical_ram_width = 16;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 7;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "clock0";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 127;
defparam ram_block1a15.port_b_logical_ram_depth = 128;
defparam ram_block1a15.port_b_logical_ram_width = 16;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.clk0_output_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "old";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 7;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 127;
defparam ram_block1a14.port_a_logical_ram_depth = 128;
defparam ram_block1a14.port_a_logical_ram_width = 16;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 7;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "clock0";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 127;
defparam ram_block1a14.port_b_logical_ram_depth = 128;
defparam ram_block1a14.port_b_logical_ram_width = 16;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.clk0_output_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "old";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 7;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 127;
defparam ram_block1a13.port_a_logical_ram_depth = 128;
defparam ram_block1a13.port_a_logical_ram_width = 16;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 7;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "clock0";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 127;
defparam ram_block1a13.port_b_logical_ram_depth = 128;
defparam ram_block1a13.port_b_logical_ram_width = 16;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.clk0_output_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "old";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 7;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 127;
defparam ram_block1a12.port_a_logical_ram_depth = 128;
defparam ram_block1a12.port_a_logical_ram_width = 16;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 7;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "clock0";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 127;
defparam ram_block1a12.port_b_logical_ram_depth = 128;
defparam ram_block1a12.port_b_logical_ram_width = 16;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.clk0_output_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "old";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 7;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 127;
defparam ram_block1a11.port_a_logical_ram_depth = 128;
defparam ram_block1a11.port_a_logical_ram_width = 16;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 7;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "clock0";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 127;
defparam ram_block1a11.port_b_logical_ram_depth = 128;
defparam ram_block1a11.port_b_logical_ram_width = 16;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.clk0_output_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "old";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 7;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 127;
defparam ram_block1a10.port_a_logical_ram_depth = 128;
defparam ram_block1a10.port_a_logical_ram_width = 16;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 7;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "clock0";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 127;
defparam ram_block1a10.port_b_logical_ram_depth = 128;
defparam ram_block1a10.port_b_logical_ram_width = 16;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";

endmodule

module fft_asj_fft_data_ram_fft_120_3 (
	q_b_1,
	q_b_0,
	q_b_7,
	q_b_6,
	q_b_5,
	q_b_4,
	q_b_3,
	q_b_2,
	q_b_9,
	q_b_8,
	q_b_15,
	q_b_14,
	q_b_13,
	q_b_12,
	q_b_11,
	q_b_10,
	ram_in_reg_1_7,
	ram_in_reg_0_7,
	ram_in_reg_7_7,
	ram_in_reg_6_7,
	ram_in_reg_5_7,
	ram_in_reg_4_7,
	ram_in_reg_3_7,
	ram_in_reg_2_7,
	ram_in_reg_1_3,
	ram_in_reg_0_3,
	ram_in_reg_7_3,
	ram_in_reg_6_3,
	ram_in_reg_5_3,
	ram_in_reg_4_3,
	ram_in_reg_3_3,
	ram_in_reg_2_3,
	global_clock_enable,
	wc_vec_6,
	ram_in_reg_6_0,
	rdaddress_c_bus_0,
	rdaddress_c_bus_15,
	rdaddress_c_bus_16,
	rdaddress_c_bus_10,
	rdaddress_c_bus_11,
	rdaddress_c_bus_12,
	ram_in_reg_0_1,
	ram_in_reg_2_1,
	ram_in_reg_4_1,
	rdaddress_c_bus_20,
	ram_in_reg_1_31,
	ram_in_reg_3_31,
	ram_in_reg_5_31,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_1;
output 	q_b_0;
output 	q_b_7;
output 	q_b_6;
output 	q_b_5;
output 	q_b_4;
output 	q_b_3;
output 	q_b_2;
output 	q_b_9;
output 	q_b_8;
output 	q_b_15;
output 	q_b_14;
output 	q_b_13;
output 	q_b_12;
output 	q_b_11;
output 	q_b_10;
input 	ram_in_reg_1_7;
input 	ram_in_reg_0_7;
input 	ram_in_reg_7_7;
input 	ram_in_reg_6_7;
input 	ram_in_reg_5_7;
input 	ram_in_reg_4_7;
input 	ram_in_reg_3_7;
input 	ram_in_reg_2_7;
input 	ram_in_reg_1_3;
input 	ram_in_reg_0_3;
input 	ram_in_reg_7_3;
input 	ram_in_reg_6_3;
input 	ram_in_reg_5_3;
input 	ram_in_reg_4_3;
input 	ram_in_reg_3_3;
input 	ram_in_reg_2_3;
input 	global_clock_enable;
input 	wc_vec_6;
input 	ram_in_reg_6_0;
input 	rdaddress_c_bus_0;
input 	rdaddress_c_bus_15;
input 	rdaddress_c_bus_16;
input 	rdaddress_c_bus_10;
input 	rdaddress_c_bus_11;
input 	rdaddress_c_bus_12;
input 	ram_in_reg_0_1;
input 	ram_in_reg_2_1;
input 	ram_in_reg_4_1;
input 	rdaddress_c_bus_20;
input 	ram_in_reg_1_31;
input 	ram_in_reg_3_31;
input 	ram_in_reg_5_31;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_altsyncram_10 \gen_M4K:altsyncram_component (
	.q_b({q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.data_a({ram_in_reg_7_3,ram_in_reg_6_3,ram_in_reg_5_3,ram_in_reg_4_3,ram_in_reg_3_3,ram_in_reg_2_3,ram_in_reg_1_3,ram_in_reg_0_3,ram_in_reg_7_7,ram_in_reg_6_7,ram_in_reg_5_7,ram_in_reg_4_7,ram_in_reg_3_7,ram_in_reg_2_7,ram_in_reg_1_7,ram_in_reg_0_7}),
	.clocken0(global_clock_enable),
	.wren_a(wc_vec_6),
	.address_a({ram_in_reg_6_0,ram_in_reg_5_31,ram_in_reg_4_1,ram_in_reg_3_31,ram_in_reg_2_1,ram_in_reg_1_31,ram_in_reg_0_1}),
	.address_b({rdaddress_c_bus_20,rdaddress_c_bus_12,rdaddress_c_bus_11,rdaddress_c_bus_10,rdaddress_c_bus_16,rdaddress_c_bus_15,rdaddress_c_bus_0}),
	.clock0(clk));

endmodule

module fft_altsyncram_10 (
	q_b,
	data_a,
	clocken0,
	wren_a,
	address_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	[15:0] data_a;
input 	clocken0;
input 	wren_a;
input 	[6:0] address_a;
input 	[6:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_altsyncram_lmu3_3 auto_generated(
	.q_b({q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.data_a({data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.clocken0(clocken0),
	.wren_a(wren_a),
	.address_a({address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.clock0(clock0));

endmodule

module fft_altsyncram_lmu3_3 (
	q_b,
	data_a,
	clocken0,
	wren_a,
	address_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	[15:0] data_a;
input 	clocken0;
input 	wren_a;
input 	[6:0] address_a;
input 	[6:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

cycloneiii_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "old";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 7;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 127;
defparam ram_block1a1.port_a_logical_ram_depth = 128;
defparam ram_block1a1.port_a_logical_ram_width = 16;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 7;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "clock0";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 127;
defparam ram_block1a1.port_b_logical_ram_depth = 128;
defparam ram_block1a1.port_b_logical_ram_width = 16;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "old";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 7;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 127;
defparam ram_block1a0.port_a_logical_ram_depth = 128;
defparam ram_block1a0.port_a_logical_ram_width = 16;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 7;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "clock0";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 127;
defparam ram_block1a0.port_b_logical_ram_depth = 128;
defparam ram_block1a0.port_b_logical_ram_width = 16;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "old";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 7;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 127;
defparam ram_block1a7.port_a_logical_ram_depth = 128;
defparam ram_block1a7.port_a_logical_ram_width = 16;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 7;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "clock0";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 127;
defparam ram_block1a7.port_b_logical_ram_depth = 128;
defparam ram_block1a7.port_b_logical_ram_width = 16;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "old";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 7;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 127;
defparam ram_block1a6.port_a_logical_ram_depth = 128;
defparam ram_block1a6.port_a_logical_ram_width = 16;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 7;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "clock0";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 127;
defparam ram_block1a6.port_b_logical_ram_depth = 128;
defparam ram_block1a6.port_b_logical_ram_width = 16;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "old";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 7;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 127;
defparam ram_block1a5.port_a_logical_ram_depth = 128;
defparam ram_block1a5.port_a_logical_ram_width = 16;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 7;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "clock0";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 127;
defparam ram_block1a5.port_b_logical_ram_depth = 128;
defparam ram_block1a5.port_b_logical_ram_width = 16;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "old";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 7;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 127;
defparam ram_block1a4.port_a_logical_ram_depth = 128;
defparam ram_block1a4.port_a_logical_ram_width = 16;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 7;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "clock0";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 127;
defparam ram_block1a4.port_b_logical_ram_depth = 128;
defparam ram_block1a4.port_b_logical_ram_width = 16;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "old";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 7;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 127;
defparam ram_block1a3.port_a_logical_ram_depth = 128;
defparam ram_block1a3.port_a_logical_ram_width = 16;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 7;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "clock0";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 127;
defparam ram_block1a3.port_b_logical_ram_depth = 128;
defparam ram_block1a3.port_b_logical_ram_width = 16;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "old";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 7;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 127;
defparam ram_block1a2.port_a_logical_ram_depth = 128;
defparam ram_block1a2.port_a_logical_ram_width = 16;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 7;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "clock0";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 127;
defparam ram_block1a2.port_b_logical_ram_depth = 128;
defparam ram_block1a2.port_b_logical_ram_width = 16;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.clk0_output_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "old";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 7;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 127;
defparam ram_block1a9.port_a_logical_ram_depth = 128;
defparam ram_block1a9.port_a_logical_ram_width = 16;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 7;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "clock0";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 127;
defparam ram_block1a9.port_b_logical_ram_depth = 128;
defparam ram_block1a9.port_b_logical_ram_width = 16;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.clk0_output_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "old";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 7;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 127;
defparam ram_block1a8.port_a_logical_ram_depth = 128;
defparam ram_block1a8.port_a_logical_ram_width = 16;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 7;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "clock0";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 127;
defparam ram_block1a8.port_b_logical_ram_depth = 128;
defparam ram_block1a8.port_b_logical_ram_width = 16;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.clk0_output_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "old";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 7;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 127;
defparam ram_block1a15.port_a_logical_ram_depth = 128;
defparam ram_block1a15.port_a_logical_ram_width = 16;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 7;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "clock0";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 127;
defparam ram_block1a15.port_b_logical_ram_depth = 128;
defparam ram_block1a15.port_b_logical_ram_width = 16;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.clk0_output_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "old";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 7;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 127;
defparam ram_block1a14.port_a_logical_ram_depth = 128;
defparam ram_block1a14.port_a_logical_ram_width = 16;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 7;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "clock0";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 127;
defparam ram_block1a14.port_b_logical_ram_depth = 128;
defparam ram_block1a14.port_b_logical_ram_width = 16;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.clk0_output_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "old";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 7;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 127;
defparam ram_block1a13.port_a_logical_ram_depth = 128;
defparam ram_block1a13.port_a_logical_ram_width = 16;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 7;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "clock0";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 127;
defparam ram_block1a13.port_b_logical_ram_depth = 128;
defparam ram_block1a13.port_b_logical_ram_width = 16;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.clk0_output_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "old";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 7;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 127;
defparam ram_block1a12.port_a_logical_ram_depth = 128;
defparam ram_block1a12.port_a_logical_ram_width = 16;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 7;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "clock0";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 127;
defparam ram_block1a12.port_b_logical_ram_depth = 128;
defparam ram_block1a12.port_b_logical_ram_width = 16;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.clk0_output_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "old";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 7;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 127;
defparam ram_block1a11.port_a_logical_ram_depth = 128;
defparam ram_block1a11.port_a_logical_ram_width = 16;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 7;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "clock0";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 127;
defparam ram_block1a11.port_b_logical_ram_depth = 128;
defparam ram_block1a11.port_b_logical_ram_width = 16;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.clk0_output_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_C|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "old";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 7;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 127;
defparam ram_block1a10.port_a_logical_ram_depth = 128;
defparam ram_block1a10.port_a_logical_ram_width = 16;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 7;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "clock0";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 127;
defparam ram_block1a10.port_b_logical_ram_depth = 128;
defparam ram_block1a10.port_b_logical_ram_width = 16;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";

endmodule

module fft_asj_fft_4dp_ram_fft_120_1 (
	q_b_1,
	q_b_11,
	q_b_12,
	q_b_13,
	q_b_0,
	q_b_01,
	q_b_02,
	q_b_03,
	q_b_7,
	q_b_71,
	q_b_72,
	q_b_73,
	q_b_6,
	q_b_61,
	q_b_62,
	q_b_63,
	q_b_5,
	q_b_51,
	q_b_52,
	q_b_53,
	q_b_4,
	q_b_41,
	q_b_42,
	q_b_43,
	q_b_3,
	q_b_31,
	q_b_32,
	q_b_33,
	q_b_2,
	q_b_21,
	q_b_22,
	q_b_23,
	q_b_9,
	q_b_91,
	q_b_92,
	q_b_93,
	q_b_8,
	q_b_81,
	q_b_82,
	q_b_83,
	q_b_15,
	q_b_151,
	q_b_152,
	q_b_153,
	q_b_14,
	q_b_141,
	q_b_142,
	q_b_143,
	q_b_131,
	q_b_132,
	q_b_133,
	q_b_134,
	q_b_121,
	q_b_122,
	q_b_123,
	q_b_124,
	q_b_111,
	q_b_112,
	q_b_113,
	q_b_114,
	q_b_10,
	q_b_101,
	q_b_102,
	q_b_103,
	ram_in_reg_1_6,
	ram_in_reg_1_5,
	ram_in_reg_1_4,
	ram_in_reg_1_7,
	ram_in_reg_0_6,
	ram_in_reg_0_5,
	ram_in_reg_0_4,
	ram_in_reg_0_7,
	ram_in_reg_7_6,
	ram_in_reg_7_5,
	ram_in_reg_7_4,
	ram_in_reg_7_7,
	ram_in_reg_6_6,
	ram_in_reg_6_5,
	ram_in_reg_6_4,
	ram_in_reg_6_7,
	ram_in_reg_5_6,
	ram_in_reg_5_5,
	ram_in_reg_5_4,
	ram_in_reg_5_7,
	ram_in_reg_4_6,
	ram_in_reg_4_5,
	ram_in_reg_4_4,
	ram_in_reg_4_7,
	ram_in_reg_3_6,
	ram_in_reg_3_5,
	ram_in_reg_3_4,
	ram_in_reg_3_7,
	ram_in_reg_2_6,
	ram_in_reg_2_5,
	ram_in_reg_2_4,
	ram_in_reg_2_7,
	ram_in_reg_1_2,
	ram_in_reg_1_1,
	ram_in_reg_1_0,
	ram_in_reg_1_3,
	ram_in_reg_0_2,
	ram_in_reg_0_1,
	ram_in_reg_0_0,
	ram_in_reg_0_3,
	ram_in_reg_7_2,
	ram_in_reg_7_1,
	ram_in_reg_7_0,
	ram_in_reg_7_3,
	ram_in_reg_6_2,
	ram_in_reg_6_1,
	ram_in_reg_6_0,
	ram_in_reg_6_3,
	ram_in_reg_5_2,
	ram_in_reg_5_1,
	ram_in_reg_5_0,
	ram_in_reg_5_3,
	ram_in_reg_4_2,
	ram_in_reg_4_1,
	ram_in_reg_4_0,
	ram_in_reg_4_3,
	ram_in_reg_3_2,
	ram_in_reg_3_1,
	ram_in_reg_3_0,
	ram_in_reg_3_3,
	ram_in_reg_2_2,
	ram_in_reg_2_1,
	ram_in_reg_2_0,
	ram_in_reg_2_3,
	global_clock_enable,
	ram_in_reg_0_01,
	ram_in_reg_1_21,
	ram_in_reg_2_01,
	ram_in_reg_3_21,
	ram_in_reg_4_01,
	ram_in_reg_5_21,
	ram_in_reg_6_01,
	rdaddress_c_bus_0,
	rdaddress_c_bus_15,
	rdaddress_c_bus_16,
	rdaddress_c_bus_10,
	rdaddress_c_bus_11,
	rdaddress_c_bus_12,
	rdaddress_c_bus_13,
	wd_vec_6,
	ram_in_reg_0_11,
	ram_in_reg_1_11,
	ram_in_reg_2_11,
	ram_in_reg_3_11,
	ram_in_reg_4_11,
	ram_in_reg_5_11,
	rdaddress_c_bus_20,
	ram_in_reg_1_01,
	ram_in_reg_3_01,
	ram_in_reg_5_01,
	ram_in_reg_1_31,
	ram_in_reg_3_31,
	ram_in_reg_5_31,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_1;
output 	q_b_11;
output 	q_b_12;
output 	q_b_13;
output 	q_b_0;
output 	q_b_01;
output 	q_b_02;
output 	q_b_03;
output 	q_b_7;
output 	q_b_71;
output 	q_b_72;
output 	q_b_73;
output 	q_b_6;
output 	q_b_61;
output 	q_b_62;
output 	q_b_63;
output 	q_b_5;
output 	q_b_51;
output 	q_b_52;
output 	q_b_53;
output 	q_b_4;
output 	q_b_41;
output 	q_b_42;
output 	q_b_43;
output 	q_b_3;
output 	q_b_31;
output 	q_b_32;
output 	q_b_33;
output 	q_b_2;
output 	q_b_21;
output 	q_b_22;
output 	q_b_23;
output 	q_b_9;
output 	q_b_91;
output 	q_b_92;
output 	q_b_93;
output 	q_b_8;
output 	q_b_81;
output 	q_b_82;
output 	q_b_83;
output 	q_b_15;
output 	q_b_151;
output 	q_b_152;
output 	q_b_153;
output 	q_b_14;
output 	q_b_141;
output 	q_b_142;
output 	q_b_143;
output 	q_b_131;
output 	q_b_132;
output 	q_b_133;
output 	q_b_134;
output 	q_b_121;
output 	q_b_122;
output 	q_b_123;
output 	q_b_124;
output 	q_b_111;
output 	q_b_112;
output 	q_b_113;
output 	q_b_114;
output 	q_b_10;
output 	q_b_101;
output 	q_b_102;
output 	q_b_103;
input 	ram_in_reg_1_6;
input 	ram_in_reg_1_5;
input 	ram_in_reg_1_4;
input 	ram_in_reg_1_7;
input 	ram_in_reg_0_6;
input 	ram_in_reg_0_5;
input 	ram_in_reg_0_4;
input 	ram_in_reg_0_7;
input 	ram_in_reg_7_6;
input 	ram_in_reg_7_5;
input 	ram_in_reg_7_4;
input 	ram_in_reg_7_7;
input 	ram_in_reg_6_6;
input 	ram_in_reg_6_5;
input 	ram_in_reg_6_4;
input 	ram_in_reg_6_7;
input 	ram_in_reg_5_6;
input 	ram_in_reg_5_5;
input 	ram_in_reg_5_4;
input 	ram_in_reg_5_7;
input 	ram_in_reg_4_6;
input 	ram_in_reg_4_5;
input 	ram_in_reg_4_4;
input 	ram_in_reg_4_7;
input 	ram_in_reg_3_6;
input 	ram_in_reg_3_5;
input 	ram_in_reg_3_4;
input 	ram_in_reg_3_7;
input 	ram_in_reg_2_6;
input 	ram_in_reg_2_5;
input 	ram_in_reg_2_4;
input 	ram_in_reg_2_7;
input 	ram_in_reg_1_2;
input 	ram_in_reg_1_1;
input 	ram_in_reg_1_0;
input 	ram_in_reg_1_3;
input 	ram_in_reg_0_2;
input 	ram_in_reg_0_1;
input 	ram_in_reg_0_0;
input 	ram_in_reg_0_3;
input 	ram_in_reg_7_2;
input 	ram_in_reg_7_1;
input 	ram_in_reg_7_0;
input 	ram_in_reg_7_3;
input 	ram_in_reg_6_2;
input 	ram_in_reg_6_1;
input 	ram_in_reg_6_0;
input 	ram_in_reg_6_3;
input 	ram_in_reg_5_2;
input 	ram_in_reg_5_1;
input 	ram_in_reg_5_0;
input 	ram_in_reg_5_3;
input 	ram_in_reg_4_2;
input 	ram_in_reg_4_1;
input 	ram_in_reg_4_0;
input 	ram_in_reg_4_3;
input 	ram_in_reg_3_2;
input 	ram_in_reg_3_1;
input 	ram_in_reg_3_0;
input 	ram_in_reg_3_3;
input 	ram_in_reg_2_2;
input 	ram_in_reg_2_1;
input 	ram_in_reg_2_0;
input 	ram_in_reg_2_3;
input 	global_clock_enable;
input 	ram_in_reg_0_01;
input 	ram_in_reg_1_21;
input 	ram_in_reg_2_01;
input 	ram_in_reg_3_21;
input 	ram_in_reg_4_01;
input 	ram_in_reg_5_21;
input 	ram_in_reg_6_01;
input 	rdaddress_c_bus_0;
input 	rdaddress_c_bus_15;
input 	rdaddress_c_bus_16;
input 	rdaddress_c_bus_10;
input 	rdaddress_c_bus_11;
input 	rdaddress_c_bus_12;
input 	rdaddress_c_bus_13;
input 	wd_vec_6;
input 	ram_in_reg_0_11;
input 	ram_in_reg_1_11;
input 	ram_in_reg_2_11;
input 	ram_in_reg_3_11;
input 	ram_in_reg_4_11;
input 	ram_in_reg_5_11;
input 	rdaddress_c_bus_20;
input 	ram_in_reg_1_01;
input 	ram_in_reg_3_01;
input 	ram_in_reg_5_01;
input 	ram_in_reg_1_31;
input 	ram_in_reg_3_31;
input 	ram_in_reg_5_31;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_asj_fft_data_ram_fft_120_7 \gen_rams:3:dat_A (
	.q_b_1(q_b_13),
	.q_b_0(q_b_03),
	.q_b_7(q_b_73),
	.q_b_6(q_b_63),
	.q_b_5(q_b_53),
	.q_b_4(q_b_43),
	.q_b_3(q_b_33),
	.q_b_2(q_b_23),
	.q_b_9(q_b_93),
	.q_b_8(q_b_83),
	.q_b_15(q_b_153),
	.q_b_14(q_b_143),
	.q_b_13(q_b_134),
	.q_b_12(q_b_124),
	.q_b_11(q_b_114),
	.q_b_10(q_b_103),
	.ram_in_reg_1_7(ram_in_reg_1_7),
	.ram_in_reg_0_7(ram_in_reg_0_7),
	.ram_in_reg_7_7(ram_in_reg_7_7),
	.ram_in_reg_6_7(ram_in_reg_6_7),
	.ram_in_reg_5_7(ram_in_reg_5_7),
	.ram_in_reg_4_7(ram_in_reg_4_7),
	.ram_in_reg_3_7(ram_in_reg_3_7),
	.ram_in_reg_2_7(ram_in_reg_2_7),
	.ram_in_reg_1_3(ram_in_reg_1_3),
	.ram_in_reg_0_3(ram_in_reg_0_3),
	.ram_in_reg_7_3(ram_in_reg_7_3),
	.ram_in_reg_6_3(ram_in_reg_6_3),
	.ram_in_reg_5_3(ram_in_reg_5_3),
	.ram_in_reg_4_3(ram_in_reg_4_3),
	.ram_in_reg_3_3(ram_in_reg_3_3),
	.ram_in_reg_2_3(ram_in_reg_2_3),
	.global_clock_enable(global_clock_enable),
	.ram_in_reg_6_0(ram_in_reg_6_01),
	.rdaddress_c_bus_0(rdaddress_c_bus_0),
	.rdaddress_c_bus_15(rdaddress_c_bus_15),
	.rdaddress_c_bus_16(rdaddress_c_bus_16),
	.rdaddress_c_bus_10(rdaddress_c_bus_10),
	.rdaddress_c_bus_11(rdaddress_c_bus_11),
	.rdaddress_c_bus_12(rdaddress_c_bus_12),
	.wd_vec_6(wd_vec_6),
	.ram_in_reg_0_1(ram_in_reg_0_11),
	.ram_in_reg_2_1(ram_in_reg_2_11),
	.ram_in_reg_4_1(ram_in_reg_4_11),
	.rdaddress_c_bus_20(rdaddress_c_bus_20),
	.ram_in_reg_1_31(ram_in_reg_1_31),
	.ram_in_reg_3_31(ram_in_reg_3_31),
	.ram_in_reg_5_31(ram_in_reg_5_31),
	.clk(clk));

fft_asj_fft_data_ram_fft_120_6 \gen_rams:2:dat_A (
	.q_b_1(q_b_1),
	.q_b_0(q_b_0),
	.q_b_7(q_b_7),
	.q_b_6(q_b_6),
	.q_b_5(q_b_5),
	.q_b_4(q_b_4),
	.q_b_3(q_b_3),
	.q_b_2(q_b_2),
	.q_b_9(q_b_9),
	.q_b_8(q_b_8),
	.q_b_15(q_b_15),
	.q_b_14(q_b_14),
	.q_b_13(q_b_131),
	.q_b_12(q_b_121),
	.q_b_11(q_b_111),
	.q_b_10(q_b_10),
	.ram_in_reg_1_6(ram_in_reg_1_6),
	.ram_in_reg_0_6(ram_in_reg_0_6),
	.ram_in_reg_7_6(ram_in_reg_7_6),
	.ram_in_reg_6_6(ram_in_reg_6_6),
	.ram_in_reg_5_6(ram_in_reg_5_6),
	.ram_in_reg_4_6(ram_in_reg_4_6),
	.ram_in_reg_3_6(ram_in_reg_3_6),
	.ram_in_reg_2_6(ram_in_reg_2_6),
	.ram_in_reg_1_2(ram_in_reg_1_2),
	.ram_in_reg_0_2(ram_in_reg_0_2),
	.ram_in_reg_7_2(ram_in_reg_7_2),
	.ram_in_reg_6_2(ram_in_reg_6_2),
	.ram_in_reg_5_2(ram_in_reg_5_2),
	.ram_in_reg_4_2(ram_in_reg_4_2),
	.ram_in_reg_3_2(ram_in_reg_3_2),
	.ram_in_reg_2_2(ram_in_reg_2_2),
	.global_clock_enable(global_clock_enable),
	.ram_in_reg_0_0(ram_in_reg_0_01),
	.ram_in_reg_1_21(ram_in_reg_1_21),
	.ram_in_reg_2_0(ram_in_reg_2_01),
	.ram_in_reg_3_21(ram_in_reg_3_21),
	.ram_in_reg_4_0(ram_in_reg_4_01),
	.ram_in_reg_5_21(ram_in_reg_5_21),
	.ram_in_reg_6_0(ram_in_reg_6_01),
	.rdaddress_c_bus_0(rdaddress_c_bus_0),
	.rdaddress_c_bus_15(rdaddress_c_bus_15),
	.rdaddress_c_bus_16(rdaddress_c_bus_16),
	.rdaddress_c_bus_10(rdaddress_c_bus_10),
	.rdaddress_c_bus_11(rdaddress_c_bus_11),
	.rdaddress_c_bus_12(rdaddress_c_bus_12),
	.rdaddress_c_bus_13(rdaddress_c_bus_13),
	.wd_vec_6(wd_vec_6),
	.clk(clk));

fft_asj_fft_data_ram_fft_120_5 \gen_rams:1:dat_A (
	.q_b_1(q_b_11),
	.q_b_0(q_b_01),
	.q_b_7(q_b_71),
	.q_b_6(q_b_61),
	.q_b_5(q_b_51),
	.q_b_4(q_b_41),
	.q_b_3(q_b_31),
	.q_b_2(q_b_21),
	.q_b_9(q_b_91),
	.q_b_8(q_b_81),
	.q_b_15(q_b_151),
	.q_b_14(q_b_141),
	.q_b_13(q_b_132),
	.q_b_12(q_b_122),
	.q_b_11(q_b_112),
	.q_b_10(q_b_101),
	.ram_in_reg_1_5(ram_in_reg_1_5),
	.ram_in_reg_0_5(ram_in_reg_0_5),
	.ram_in_reg_7_5(ram_in_reg_7_5),
	.ram_in_reg_6_5(ram_in_reg_6_5),
	.ram_in_reg_5_5(ram_in_reg_5_5),
	.ram_in_reg_4_5(ram_in_reg_4_5),
	.ram_in_reg_3_5(ram_in_reg_3_5),
	.ram_in_reg_2_5(ram_in_reg_2_5),
	.ram_in_reg_1_1(ram_in_reg_1_1),
	.ram_in_reg_0_1(ram_in_reg_0_1),
	.ram_in_reg_7_1(ram_in_reg_7_1),
	.ram_in_reg_6_1(ram_in_reg_6_1),
	.ram_in_reg_5_1(ram_in_reg_5_1),
	.ram_in_reg_4_1(ram_in_reg_4_1),
	.ram_in_reg_3_1(ram_in_reg_3_1),
	.ram_in_reg_2_1(ram_in_reg_2_1),
	.global_clock_enable(global_clock_enable),
	.ram_in_reg_6_0(ram_in_reg_6_01),
	.rdaddress_c_bus_0(rdaddress_c_bus_0),
	.rdaddress_c_bus_15(rdaddress_c_bus_15),
	.rdaddress_c_bus_16(rdaddress_c_bus_16),
	.rdaddress_c_bus_10(rdaddress_c_bus_10),
	.rdaddress_c_bus_11(rdaddress_c_bus_11),
	.rdaddress_c_bus_12(rdaddress_c_bus_12),
	.wd_vec_6(wd_vec_6),
	.ram_in_reg_0_11(ram_in_reg_0_11),
	.ram_in_reg_1_11(ram_in_reg_1_11),
	.ram_in_reg_2_11(ram_in_reg_2_11),
	.ram_in_reg_3_11(ram_in_reg_3_11),
	.ram_in_reg_4_11(ram_in_reg_4_11),
	.ram_in_reg_5_11(ram_in_reg_5_11),
	.rdaddress_c_bus_20(rdaddress_c_bus_20),
	.clk(clk));

fft_asj_fft_data_ram_fft_120_4 \gen_rams:0:dat_A (
	.q_b_1(q_b_12),
	.q_b_0(q_b_02),
	.q_b_7(q_b_72),
	.q_b_6(q_b_62),
	.q_b_5(q_b_52),
	.q_b_4(q_b_42),
	.q_b_3(q_b_32),
	.q_b_2(q_b_22),
	.q_b_9(q_b_92),
	.q_b_8(q_b_82),
	.q_b_15(q_b_152),
	.q_b_14(q_b_142),
	.q_b_13(q_b_133),
	.q_b_12(q_b_123),
	.q_b_11(q_b_113),
	.q_b_10(q_b_102),
	.ram_in_reg_1_4(ram_in_reg_1_4),
	.ram_in_reg_0_4(ram_in_reg_0_4),
	.ram_in_reg_7_4(ram_in_reg_7_4),
	.ram_in_reg_6_4(ram_in_reg_6_4),
	.ram_in_reg_5_4(ram_in_reg_5_4),
	.ram_in_reg_4_4(ram_in_reg_4_4),
	.ram_in_reg_3_4(ram_in_reg_3_4),
	.ram_in_reg_2_4(ram_in_reg_2_4),
	.ram_in_reg_1_0(ram_in_reg_1_0),
	.ram_in_reg_0_0(ram_in_reg_0_0),
	.ram_in_reg_7_0(ram_in_reg_7_0),
	.ram_in_reg_6_0(ram_in_reg_6_0),
	.ram_in_reg_5_0(ram_in_reg_5_0),
	.ram_in_reg_4_0(ram_in_reg_4_0),
	.ram_in_reg_3_0(ram_in_reg_3_0),
	.ram_in_reg_2_0(ram_in_reg_2_0),
	.global_clock_enable(global_clock_enable),
	.ram_in_reg_0_01(ram_in_reg_0_01),
	.ram_in_reg_2_01(ram_in_reg_2_01),
	.ram_in_reg_4_01(ram_in_reg_4_01),
	.ram_in_reg_6_01(ram_in_reg_6_01),
	.rdaddress_c_bus_0(rdaddress_c_bus_0),
	.rdaddress_c_bus_15(rdaddress_c_bus_15),
	.rdaddress_c_bus_16(rdaddress_c_bus_16),
	.rdaddress_c_bus_10(rdaddress_c_bus_10),
	.rdaddress_c_bus_11(rdaddress_c_bus_11),
	.rdaddress_c_bus_12(rdaddress_c_bus_12),
	.rdaddress_c_bus_13(rdaddress_c_bus_13),
	.wd_vec_6(wd_vec_6),
	.ram_in_reg_1_01(ram_in_reg_1_01),
	.ram_in_reg_3_01(ram_in_reg_3_01),
	.ram_in_reg_5_01(ram_in_reg_5_01),
	.clk(clk));

endmodule

module fft_asj_fft_data_ram_fft_120_4 (
	q_b_1,
	q_b_0,
	q_b_7,
	q_b_6,
	q_b_5,
	q_b_4,
	q_b_3,
	q_b_2,
	q_b_9,
	q_b_8,
	q_b_15,
	q_b_14,
	q_b_13,
	q_b_12,
	q_b_11,
	q_b_10,
	ram_in_reg_1_4,
	ram_in_reg_0_4,
	ram_in_reg_7_4,
	ram_in_reg_6_4,
	ram_in_reg_5_4,
	ram_in_reg_4_4,
	ram_in_reg_3_4,
	ram_in_reg_2_4,
	ram_in_reg_1_0,
	ram_in_reg_0_0,
	ram_in_reg_7_0,
	ram_in_reg_6_0,
	ram_in_reg_5_0,
	ram_in_reg_4_0,
	ram_in_reg_3_0,
	ram_in_reg_2_0,
	global_clock_enable,
	ram_in_reg_0_01,
	ram_in_reg_2_01,
	ram_in_reg_4_01,
	ram_in_reg_6_01,
	rdaddress_c_bus_0,
	rdaddress_c_bus_15,
	rdaddress_c_bus_16,
	rdaddress_c_bus_10,
	rdaddress_c_bus_11,
	rdaddress_c_bus_12,
	rdaddress_c_bus_13,
	wd_vec_6,
	ram_in_reg_1_01,
	ram_in_reg_3_01,
	ram_in_reg_5_01,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_1;
output 	q_b_0;
output 	q_b_7;
output 	q_b_6;
output 	q_b_5;
output 	q_b_4;
output 	q_b_3;
output 	q_b_2;
output 	q_b_9;
output 	q_b_8;
output 	q_b_15;
output 	q_b_14;
output 	q_b_13;
output 	q_b_12;
output 	q_b_11;
output 	q_b_10;
input 	ram_in_reg_1_4;
input 	ram_in_reg_0_4;
input 	ram_in_reg_7_4;
input 	ram_in_reg_6_4;
input 	ram_in_reg_5_4;
input 	ram_in_reg_4_4;
input 	ram_in_reg_3_4;
input 	ram_in_reg_2_4;
input 	ram_in_reg_1_0;
input 	ram_in_reg_0_0;
input 	ram_in_reg_7_0;
input 	ram_in_reg_6_0;
input 	ram_in_reg_5_0;
input 	ram_in_reg_4_0;
input 	ram_in_reg_3_0;
input 	ram_in_reg_2_0;
input 	global_clock_enable;
input 	ram_in_reg_0_01;
input 	ram_in_reg_2_01;
input 	ram_in_reg_4_01;
input 	ram_in_reg_6_01;
input 	rdaddress_c_bus_0;
input 	rdaddress_c_bus_15;
input 	rdaddress_c_bus_16;
input 	rdaddress_c_bus_10;
input 	rdaddress_c_bus_11;
input 	rdaddress_c_bus_12;
input 	rdaddress_c_bus_13;
input 	wd_vec_6;
input 	ram_in_reg_1_01;
input 	ram_in_reg_3_01;
input 	ram_in_reg_5_01;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_altsyncram_11 \gen_M4K:altsyncram_component (
	.q_b({q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.data_a({ram_in_reg_7_0,ram_in_reg_6_0,ram_in_reg_5_0,ram_in_reg_4_0,ram_in_reg_3_0,ram_in_reg_2_0,ram_in_reg_1_0,ram_in_reg_0_0,ram_in_reg_7_4,ram_in_reg_6_4,ram_in_reg_5_4,ram_in_reg_4_4,ram_in_reg_3_4,ram_in_reg_2_4,ram_in_reg_1_4,ram_in_reg_0_4}),
	.clocken0(global_clock_enable),
	.address_a({ram_in_reg_6_01,ram_in_reg_5_01,ram_in_reg_4_01,ram_in_reg_3_01,ram_in_reg_2_01,ram_in_reg_1_01,ram_in_reg_0_01}),
	.address_b({rdaddress_c_bus_13,rdaddress_c_bus_12,rdaddress_c_bus_11,rdaddress_c_bus_10,rdaddress_c_bus_16,rdaddress_c_bus_15,rdaddress_c_bus_0}),
	.wren_a(wd_vec_6),
	.clock0(clk));

endmodule

module fft_altsyncram_11 (
	q_b,
	data_a,
	clocken0,
	address_a,
	address_b,
	wren_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	[15:0] data_a;
input 	clocken0;
input 	[6:0] address_a;
input 	[6:0] address_b;
input 	wren_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_altsyncram_lmu3_4 auto_generated(
	.q_b({q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.data_a({data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.clocken0(clocken0),
	.address_a({address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.wren_a(wren_a),
	.clock0(clock0));

endmodule

module fft_altsyncram_lmu3_4 (
	q_b,
	data_a,
	clocken0,
	address_a,
	address_b,
	wren_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	[15:0] data_a;
input 	clocken0;
input 	[6:0] address_a;
input 	[6:0] address_b;
input 	wren_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

cycloneiii_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "old";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 7;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 127;
defparam ram_block1a1.port_a_logical_ram_depth = 128;
defparam ram_block1a1.port_a_logical_ram_width = 16;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 7;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "clock0";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 127;
defparam ram_block1a1.port_b_logical_ram_depth = 128;
defparam ram_block1a1.port_b_logical_ram_width = 16;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "old";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 7;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 127;
defparam ram_block1a0.port_a_logical_ram_depth = 128;
defparam ram_block1a0.port_a_logical_ram_width = 16;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 7;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "clock0";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 127;
defparam ram_block1a0.port_b_logical_ram_depth = 128;
defparam ram_block1a0.port_b_logical_ram_width = 16;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "old";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 7;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 127;
defparam ram_block1a7.port_a_logical_ram_depth = 128;
defparam ram_block1a7.port_a_logical_ram_width = 16;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 7;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "clock0";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 127;
defparam ram_block1a7.port_b_logical_ram_depth = 128;
defparam ram_block1a7.port_b_logical_ram_width = 16;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "old";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 7;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 127;
defparam ram_block1a6.port_a_logical_ram_depth = 128;
defparam ram_block1a6.port_a_logical_ram_width = 16;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 7;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "clock0";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 127;
defparam ram_block1a6.port_b_logical_ram_depth = 128;
defparam ram_block1a6.port_b_logical_ram_width = 16;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "old";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 7;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 127;
defparam ram_block1a5.port_a_logical_ram_depth = 128;
defparam ram_block1a5.port_a_logical_ram_width = 16;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 7;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "clock0";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 127;
defparam ram_block1a5.port_b_logical_ram_depth = 128;
defparam ram_block1a5.port_b_logical_ram_width = 16;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "old";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 7;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 127;
defparam ram_block1a4.port_a_logical_ram_depth = 128;
defparam ram_block1a4.port_a_logical_ram_width = 16;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 7;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "clock0";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 127;
defparam ram_block1a4.port_b_logical_ram_depth = 128;
defparam ram_block1a4.port_b_logical_ram_width = 16;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "old";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 7;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 127;
defparam ram_block1a3.port_a_logical_ram_depth = 128;
defparam ram_block1a3.port_a_logical_ram_width = 16;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 7;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "clock0";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 127;
defparam ram_block1a3.port_b_logical_ram_depth = 128;
defparam ram_block1a3.port_b_logical_ram_width = 16;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "old";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 7;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 127;
defparam ram_block1a2.port_a_logical_ram_depth = 128;
defparam ram_block1a2.port_a_logical_ram_width = 16;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 7;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "clock0";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 127;
defparam ram_block1a2.port_b_logical_ram_depth = 128;
defparam ram_block1a2.port_b_logical_ram_width = 16;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.clk0_output_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "old";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 7;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 127;
defparam ram_block1a9.port_a_logical_ram_depth = 128;
defparam ram_block1a9.port_a_logical_ram_width = 16;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 7;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "clock0";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 127;
defparam ram_block1a9.port_b_logical_ram_depth = 128;
defparam ram_block1a9.port_b_logical_ram_width = 16;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.clk0_output_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "old";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 7;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 127;
defparam ram_block1a8.port_a_logical_ram_depth = 128;
defparam ram_block1a8.port_a_logical_ram_width = 16;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 7;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "clock0";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 127;
defparam ram_block1a8.port_b_logical_ram_depth = 128;
defparam ram_block1a8.port_b_logical_ram_width = 16;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.clk0_output_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "old";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 7;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 127;
defparam ram_block1a15.port_a_logical_ram_depth = 128;
defparam ram_block1a15.port_a_logical_ram_width = 16;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 7;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "clock0";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 127;
defparam ram_block1a15.port_b_logical_ram_depth = 128;
defparam ram_block1a15.port_b_logical_ram_width = 16;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.clk0_output_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "old";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 7;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 127;
defparam ram_block1a14.port_a_logical_ram_depth = 128;
defparam ram_block1a14.port_a_logical_ram_width = 16;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 7;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "clock0";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 127;
defparam ram_block1a14.port_b_logical_ram_depth = 128;
defparam ram_block1a14.port_b_logical_ram_width = 16;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.clk0_output_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "old";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 7;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 127;
defparam ram_block1a13.port_a_logical_ram_depth = 128;
defparam ram_block1a13.port_a_logical_ram_width = 16;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 7;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "clock0";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 127;
defparam ram_block1a13.port_b_logical_ram_depth = 128;
defparam ram_block1a13.port_b_logical_ram_width = 16;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.clk0_output_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "old";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 7;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 127;
defparam ram_block1a12.port_a_logical_ram_depth = 128;
defparam ram_block1a12.port_a_logical_ram_width = 16;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 7;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "clock0";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 127;
defparam ram_block1a12.port_b_logical_ram_depth = 128;
defparam ram_block1a12.port_b_logical_ram_width = 16;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.clk0_output_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "old";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 7;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 127;
defparam ram_block1a11.port_a_logical_ram_depth = 128;
defparam ram_block1a11.port_a_logical_ram_width = 16;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 7;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "clock0";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 127;
defparam ram_block1a11.port_b_logical_ram_depth = 128;
defparam ram_block1a11.port_b_logical_ram_width = 16;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.clk0_output_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "old";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 7;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 127;
defparam ram_block1a10.port_a_logical_ram_depth = 128;
defparam ram_block1a10.port_a_logical_ram_width = 16;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 7;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "clock0";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 127;
defparam ram_block1a10.port_b_logical_ram_depth = 128;
defparam ram_block1a10.port_b_logical_ram_width = 16;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";

endmodule

module fft_asj_fft_data_ram_fft_120_5 (
	q_b_1,
	q_b_0,
	q_b_7,
	q_b_6,
	q_b_5,
	q_b_4,
	q_b_3,
	q_b_2,
	q_b_9,
	q_b_8,
	q_b_15,
	q_b_14,
	q_b_13,
	q_b_12,
	q_b_11,
	q_b_10,
	ram_in_reg_1_5,
	ram_in_reg_0_5,
	ram_in_reg_7_5,
	ram_in_reg_6_5,
	ram_in_reg_5_5,
	ram_in_reg_4_5,
	ram_in_reg_3_5,
	ram_in_reg_2_5,
	ram_in_reg_1_1,
	ram_in_reg_0_1,
	ram_in_reg_7_1,
	ram_in_reg_6_1,
	ram_in_reg_5_1,
	ram_in_reg_4_1,
	ram_in_reg_3_1,
	ram_in_reg_2_1,
	global_clock_enable,
	ram_in_reg_6_0,
	rdaddress_c_bus_0,
	rdaddress_c_bus_15,
	rdaddress_c_bus_16,
	rdaddress_c_bus_10,
	rdaddress_c_bus_11,
	rdaddress_c_bus_12,
	wd_vec_6,
	ram_in_reg_0_11,
	ram_in_reg_1_11,
	ram_in_reg_2_11,
	ram_in_reg_3_11,
	ram_in_reg_4_11,
	ram_in_reg_5_11,
	rdaddress_c_bus_20,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_1;
output 	q_b_0;
output 	q_b_7;
output 	q_b_6;
output 	q_b_5;
output 	q_b_4;
output 	q_b_3;
output 	q_b_2;
output 	q_b_9;
output 	q_b_8;
output 	q_b_15;
output 	q_b_14;
output 	q_b_13;
output 	q_b_12;
output 	q_b_11;
output 	q_b_10;
input 	ram_in_reg_1_5;
input 	ram_in_reg_0_5;
input 	ram_in_reg_7_5;
input 	ram_in_reg_6_5;
input 	ram_in_reg_5_5;
input 	ram_in_reg_4_5;
input 	ram_in_reg_3_5;
input 	ram_in_reg_2_5;
input 	ram_in_reg_1_1;
input 	ram_in_reg_0_1;
input 	ram_in_reg_7_1;
input 	ram_in_reg_6_1;
input 	ram_in_reg_5_1;
input 	ram_in_reg_4_1;
input 	ram_in_reg_3_1;
input 	ram_in_reg_2_1;
input 	global_clock_enable;
input 	ram_in_reg_6_0;
input 	rdaddress_c_bus_0;
input 	rdaddress_c_bus_15;
input 	rdaddress_c_bus_16;
input 	rdaddress_c_bus_10;
input 	rdaddress_c_bus_11;
input 	rdaddress_c_bus_12;
input 	wd_vec_6;
input 	ram_in_reg_0_11;
input 	ram_in_reg_1_11;
input 	ram_in_reg_2_11;
input 	ram_in_reg_3_11;
input 	ram_in_reg_4_11;
input 	ram_in_reg_5_11;
input 	rdaddress_c_bus_20;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_altsyncram_12 \gen_M4K:altsyncram_component (
	.q_b({q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.data_a({ram_in_reg_7_1,ram_in_reg_6_1,ram_in_reg_5_1,ram_in_reg_4_1,ram_in_reg_3_1,ram_in_reg_2_1,ram_in_reg_1_1,ram_in_reg_0_1,ram_in_reg_7_5,ram_in_reg_6_5,ram_in_reg_5_5,ram_in_reg_4_5,ram_in_reg_3_5,ram_in_reg_2_5,ram_in_reg_1_5,ram_in_reg_0_5}),
	.clocken0(global_clock_enable),
	.address_a({ram_in_reg_6_0,ram_in_reg_5_11,ram_in_reg_4_11,ram_in_reg_3_11,ram_in_reg_2_11,ram_in_reg_1_11,ram_in_reg_0_11}),
	.address_b({rdaddress_c_bus_20,rdaddress_c_bus_12,rdaddress_c_bus_11,rdaddress_c_bus_10,rdaddress_c_bus_16,rdaddress_c_bus_15,rdaddress_c_bus_0}),
	.wren_a(wd_vec_6),
	.clock0(clk));

endmodule

module fft_altsyncram_12 (
	q_b,
	data_a,
	clocken0,
	address_a,
	address_b,
	wren_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	[15:0] data_a;
input 	clocken0;
input 	[6:0] address_a;
input 	[6:0] address_b;
input 	wren_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_altsyncram_lmu3_5 auto_generated(
	.q_b({q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.data_a({data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.clocken0(clocken0),
	.address_a({address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.wren_a(wren_a),
	.clock0(clock0));

endmodule

module fft_altsyncram_lmu3_5 (
	q_b,
	data_a,
	clocken0,
	address_a,
	address_b,
	wren_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	[15:0] data_a;
input 	clocken0;
input 	[6:0] address_a;
input 	[6:0] address_b;
input 	wren_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

cycloneiii_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "old";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 7;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 127;
defparam ram_block1a1.port_a_logical_ram_depth = 128;
defparam ram_block1a1.port_a_logical_ram_width = 16;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 7;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "clock0";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 127;
defparam ram_block1a1.port_b_logical_ram_depth = 128;
defparam ram_block1a1.port_b_logical_ram_width = 16;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "old";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 7;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 127;
defparam ram_block1a0.port_a_logical_ram_depth = 128;
defparam ram_block1a0.port_a_logical_ram_width = 16;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 7;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "clock0";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 127;
defparam ram_block1a0.port_b_logical_ram_depth = 128;
defparam ram_block1a0.port_b_logical_ram_width = 16;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "old";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 7;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 127;
defparam ram_block1a7.port_a_logical_ram_depth = 128;
defparam ram_block1a7.port_a_logical_ram_width = 16;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 7;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "clock0";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 127;
defparam ram_block1a7.port_b_logical_ram_depth = 128;
defparam ram_block1a7.port_b_logical_ram_width = 16;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "old";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 7;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 127;
defparam ram_block1a6.port_a_logical_ram_depth = 128;
defparam ram_block1a6.port_a_logical_ram_width = 16;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 7;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "clock0";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 127;
defparam ram_block1a6.port_b_logical_ram_depth = 128;
defparam ram_block1a6.port_b_logical_ram_width = 16;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "old";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 7;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 127;
defparam ram_block1a5.port_a_logical_ram_depth = 128;
defparam ram_block1a5.port_a_logical_ram_width = 16;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 7;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "clock0";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 127;
defparam ram_block1a5.port_b_logical_ram_depth = 128;
defparam ram_block1a5.port_b_logical_ram_width = 16;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "old";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 7;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 127;
defparam ram_block1a4.port_a_logical_ram_depth = 128;
defparam ram_block1a4.port_a_logical_ram_width = 16;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 7;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "clock0";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 127;
defparam ram_block1a4.port_b_logical_ram_depth = 128;
defparam ram_block1a4.port_b_logical_ram_width = 16;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "old";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 7;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 127;
defparam ram_block1a3.port_a_logical_ram_depth = 128;
defparam ram_block1a3.port_a_logical_ram_width = 16;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 7;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "clock0";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 127;
defparam ram_block1a3.port_b_logical_ram_depth = 128;
defparam ram_block1a3.port_b_logical_ram_width = 16;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "old";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 7;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 127;
defparam ram_block1a2.port_a_logical_ram_depth = 128;
defparam ram_block1a2.port_a_logical_ram_width = 16;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 7;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "clock0";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 127;
defparam ram_block1a2.port_b_logical_ram_depth = 128;
defparam ram_block1a2.port_b_logical_ram_width = 16;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.clk0_output_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "old";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 7;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 127;
defparam ram_block1a9.port_a_logical_ram_depth = 128;
defparam ram_block1a9.port_a_logical_ram_width = 16;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 7;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "clock0";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 127;
defparam ram_block1a9.port_b_logical_ram_depth = 128;
defparam ram_block1a9.port_b_logical_ram_width = 16;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.clk0_output_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "old";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 7;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 127;
defparam ram_block1a8.port_a_logical_ram_depth = 128;
defparam ram_block1a8.port_a_logical_ram_width = 16;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 7;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "clock0";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 127;
defparam ram_block1a8.port_b_logical_ram_depth = 128;
defparam ram_block1a8.port_b_logical_ram_width = 16;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.clk0_output_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "old";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 7;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 127;
defparam ram_block1a15.port_a_logical_ram_depth = 128;
defparam ram_block1a15.port_a_logical_ram_width = 16;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 7;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "clock0";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 127;
defparam ram_block1a15.port_b_logical_ram_depth = 128;
defparam ram_block1a15.port_b_logical_ram_width = 16;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.clk0_output_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "old";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 7;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 127;
defparam ram_block1a14.port_a_logical_ram_depth = 128;
defparam ram_block1a14.port_a_logical_ram_width = 16;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 7;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "clock0";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 127;
defparam ram_block1a14.port_b_logical_ram_depth = 128;
defparam ram_block1a14.port_b_logical_ram_width = 16;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.clk0_output_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "old";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 7;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 127;
defparam ram_block1a13.port_a_logical_ram_depth = 128;
defparam ram_block1a13.port_a_logical_ram_width = 16;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 7;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "clock0";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 127;
defparam ram_block1a13.port_b_logical_ram_depth = 128;
defparam ram_block1a13.port_b_logical_ram_width = 16;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.clk0_output_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "old";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 7;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 127;
defparam ram_block1a12.port_a_logical_ram_depth = 128;
defparam ram_block1a12.port_a_logical_ram_width = 16;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 7;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "clock0";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 127;
defparam ram_block1a12.port_b_logical_ram_depth = 128;
defparam ram_block1a12.port_b_logical_ram_width = 16;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.clk0_output_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "old";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 7;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 127;
defparam ram_block1a11.port_a_logical_ram_depth = 128;
defparam ram_block1a11.port_a_logical_ram_width = 16;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 7;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "clock0";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 127;
defparam ram_block1a11.port_b_logical_ram_depth = 128;
defparam ram_block1a11.port_b_logical_ram_width = 16;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.clk0_output_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "old";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 7;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 127;
defparam ram_block1a10.port_a_logical_ram_depth = 128;
defparam ram_block1a10.port_a_logical_ram_width = 16;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 7;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "clock0";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 127;
defparam ram_block1a10.port_b_logical_ram_depth = 128;
defparam ram_block1a10.port_b_logical_ram_width = 16;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";

endmodule

module fft_asj_fft_data_ram_fft_120_6 (
	q_b_1,
	q_b_0,
	q_b_7,
	q_b_6,
	q_b_5,
	q_b_4,
	q_b_3,
	q_b_2,
	q_b_9,
	q_b_8,
	q_b_15,
	q_b_14,
	q_b_13,
	q_b_12,
	q_b_11,
	q_b_10,
	ram_in_reg_1_6,
	ram_in_reg_0_6,
	ram_in_reg_7_6,
	ram_in_reg_6_6,
	ram_in_reg_5_6,
	ram_in_reg_4_6,
	ram_in_reg_3_6,
	ram_in_reg_2_6,
	ram_in_reg_1_2,
	ram_in_reg_0_2,
	ram_in_reg_7_2,
	ram_in_reg_6_2,
	ram_in_reg_5_2,
	ram_in_reg_4_2,
	ram_in_reg_3_2,
	ram_in_reg_2_2,
	global_clock_enable,
	ram_in_reg_0_0,
	ram_in_reg_1_21,
	ram_in_reg_2_0,
	ram_in_reg_3_21,
	ram_in_reg_4_0,
	ram_in_reg_5_21,
	ram_in_reg_6_0,
	rdaddress_c_bus_0,
	rdaddress_c_bus_15,
	rdaddress_c_bus_16,
	rdaddress_c_bus_10,
	rdaddress_c_bus_11,
	rdaddress_c_bus_12,
	rdaddress_c_bus_13,
	wd_vec_6,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_1;
output 	q_b_0;
output 	q_b_7;
output 	q_b_6;
output 	q_b_5;
output 	q_b_4;
output 	q_b_3;
output 	q_b_2;
output 	q_b_9;
output 	q_b_8;
output 	q_b_15;
output 	q_b_14;
output 	q_b_13;
output 	q_b_12;
output 	q_b_11;
output 	q_b_10;
input 	ram_in_reg_1_6;
input 	ram_in_reg_0_6;
input 	ram_in_reg_7_6;
input 	ram_in_reg_6_6;
input 	ram_in_reg_5_6;
input 	ram_in_reg_4_6;
input 	ram_in_reg_3_6;
input 	ram_in_reg_2_6;
input 	ram_in_reg_1_2;
input 	ram_in_reg_0_2;
input 	ram_in_reg_7_2;
input 	ram_in_reg_6_2;
input 	ram_in_reg_5_2;
input 	ram_in_reg_4_2;
input 	ram_in_reg_3_2;
input 	ram_in_reg_2_2;
input 	global_clock_enable;
input 	ram_in_reg_0_0;
input 	ram_in_reg_1_21;
input 	ram_in_reg_2_0;
input 	ram_in_reg_3_21;
input 	ram_in_reg_4_0;
input 	ram_in_reg_5_21;
input 	ram_in_reg_6_0;
input 	rdaddress_c_bus_0;
input 	rdaddress_c_bus_15;
input 	rdaddress_c_bus_16;
input 	rdaddress_c_bus_10;
input 	rdaddress_c_bus_11;
input 	rdaddress_c_bus_12;
input 	rdaddress_c_bus_13;
input 	wd_vec_6;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_altsyncram_13 \gen_M4K:altsyncram_component (
	.q_b({q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.data_a({ram_in_reg_7_2,ram_in_reg_6_2,ram_in_reg_5_2,ram_in_reg_4_2,ram_in_reg_3_2,ram_in_reg_2_2,ram_in_reg_1_2,ram_in_reg_0_2,ram_in_reg_7_6,ram_in_reg_6_6,ram_in_reg_5_6,ram_in_reg_4_6,ram_in_reg_3_6,ram_in_reg_2_6,ram_in_reg_1_6,ram_in_reg_0_6}),
	.clocken0(global_clock_enable),
	.address_a({ram_in_reg_6_0,ram_in_reg_5_21,ram_in_reg_4_0,ram_in_reg_3_21,ram_in_reg_2_0,ram_in_reg_1_21,ram_in_reg_0_0}),
	.address_b({rdaddress_c_bus_13,rdaddress_c_bus_12,rdaddress_c_bus_11,rdaddress_c_bus_10,rdaddress_c_bus_16,rdaddress_c_bus_15,rdaddress_c_bus_0}),
	.wren_a(wd_vec_6),
	.clock0(clk));

endmodule

module fft_altsyncram_13 (
	q_b,
	data_a,
	clocken0,
	address_a,
	address_b,
	wren_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	[15:0] data_a;
input 	clocken0;
input 	[6:0] address_a;
input 	[6:0] address_b;
input 	wren_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_altsyncram_lmu3_6 auto_generated(
	.q_b({q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.data_a({data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.clocken0(clocken0),
	.address_a({address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.wren_a(wren_a),
	.clock0(clock0));

endmodule

module fft_altsyncram_lmu3_6 (
	q_b,
	data_a,
	clocken0,
	address_a,
	address_b,
	wren_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	[15:0] data_a;
input 	clocken0;
input 	[6:0] address_a;
input 	[6:0] address_b;
input 	wren_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

cycloneiii_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "old";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 7;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 127;
defparam ram_block1a1.port_a_logical_ram_depth = 128;
defparam ram_block1a1.port_a_logical_ram_width = 16;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 7;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "clock0";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 127;
defparam ram_block1a1.port_b_logical_ram_depth = 128;
defparam ram_block1a1.port_b_logical_ram_width = 16;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "old";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 7;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 127;
defparam ram_block1a0.port_a_logical_ram_depth = 128;
defparam ram_block1a0.port_a_logical_ram_width = 16;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 7;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "clock0";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 127;
defparam ram_block1a0.port_b_logical_ram_depth = 128;
defparam ram_block1a0.port_b_logical_ram_width = 16;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "old";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 7;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 127;
defparam ram_block1a7.port_a_logical_ram_depth = 128;
defparam ram_block1a7.port_a_logical_ram_width = 16;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 7;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "clock0";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 127;
defparam ram_block1a7.port_b_logical_ram_depth = 128;
defparam ram_block1a7.port_b_logical_ram_width = 16;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "old";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 7;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 127;
defparam ram_block1a6.port_a_logical_ram_depth = 128;
defparam ram_block1a6.port_a_logical_ram_width = 16;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 7;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "clock0";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 127;
defparam ram_block1a6.port_b_logical_ram_depth = 128;
defparam ram_block1a6.port_b_logical_ram_width = 16;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "old";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 7;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 127;
defparam ram_block1a5.port_a_logical_ram_depth = 128;
defparam ram_block1a5.port_a_logical_ram_width = 16;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 7;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "clock0";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 127;
defparam ram_block1a5.port_b_logical_ram_depth = 128;
defparam ram_block1a5.port_b_logical_ram_width = 16;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "old";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 7;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 127;
defparam ram_block1a4.port_a_logical_ram_depth = 128;
defparam ram_block1a4.port_a_logical_ram_width = 16;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 7;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "clock0";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 127;
defparam ram_block1a4.port_b_logical_ram_depth = 128;
defparam ram_block1a4.port_b_logical_ram_width = 16;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "old";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 7;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 127;
defparam ram_block1a3.port_a_logical_ram_depth = 128;
defparam ram_block1a3.port_a_logical_ram_width = 16;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 7;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "clock0";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 127;
defparam ram_block1a3.port_b_logical_ram_depth = 128;
defparam ram_block1a3.port_b_logical_ram_width = 16;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "old";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 7;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 127;
defparam ram_block1a2.port_a_logical_ram_depth = 128;
defparam ram_block1a2.port_a_logical_ram_width = 16;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 7;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "clock0";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 127;
defparam ram_block1a2.port_b_logical_ram_depth = 128;
defparam ram_block1a2.port_b_logical_ram_width = 16;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.clk0_output_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "old";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 7;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 127;
defparam ram_block1a9.port_a_logical_ram_depth = 128;
defparam ram_block1a9.port_a_logical_ram_width = 16;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 7;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "clock0";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 127;
defparam ram_block1a9.port_b_logical_ram_depth = 128;
defparam ram_block1a9.port_b_logical_ram_width = 16;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.clk0_output_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "old";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 7;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 127;
defparam ram_block1a8.port_a_logical_ram_depth = 128;
defparam ram_block1a8.port_a_logical_ram_width = 16;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 7;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "clock0";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 127;
defparam ram_block1a8.port_b_logical_ram_depth = 128;
defparam ram_block1a8.port_b_logical_ram_width = 16;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.clk0_output_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "old";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 7;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 127;
defparam ram_block1a15.port_a_logical_ram_depth = 128;
defparam ram_block1a15.port_a_logical_ram_width = 16;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 7;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "clock0";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 127;
defparam ram_block1a15.port_b_logical_ram_depth = 128;
defparam ram_block1a15.port_b_logical_ram_width = 16;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.clk0_output_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "old";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 7;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 127;
defparam ram_block1a14.port_a_logical_ram_depth = 128;
defparam ram_block1a14.port_a_logical_ram_width = 16;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 7;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "clock0";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 127;
defparam ram_block1a14.port_b_logical_ram_depth = 128;
defparam ram_block1a14.port_b_logical_ram_width = 16;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.clk0_output_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "old";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 7;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 127;
defparam ram_block1a13.port_a_logical_ram_depth = 128;
defparam ram_block1a13.port_a_logical_ram_width = 16;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 7;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "clock0";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 127;
defparam ram_block1a13.port_b_logical_ram_depth = 128;
defparam ram_block1a13.port_b_logical_ram_width = 16;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.clk0_output_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "old";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 7;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 127;
defparam ram_block1a12.port_a_logical_ram_depth = 128;
defparam ram_block1a12.port_a_logical_ram_width = 16;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 7;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "clock0";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 127;
defparam ram_block1a12.port_b_logical_ram_depth = 128;
defparam ram_block1a12.port_b_logical_ram_width = 16;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.clk0_output_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "old";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 7;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 127;
defparam ram_block1a11.port_a_logical_ram_depth = 128;
defparam ram_block1a11.port_a_logical_ram_width = 16;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 7;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "clock0";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 127;
defparam ram_block1a11.port_b_logical_ram_depth = 128;
defparam ram_block1a11.port_b_logical_ram_width = 16;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.clk0_output_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "old";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 7;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 127;
defparam ram_block1a10.port_a_logical_ram_depth = 128;
defparam ram_block1a10.port_a_logical_ram_width = 16;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 7;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "clock0";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 127;
defparam ram_block1a10.port_b_logical_ram_depth = 128;
defparam ram_block1a10.port_b_logical_ram_width = 16;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";

endmodule

module fft_asj_fft_data_ram_fft_120_7 (
	q_b_1,
	q_b_0,
	q_b_7,
	q_b_6,
	q_b_5,
	q_b_4,
	q_b_3,
	q_b_2,
	q_b_9,
	q_b_8,
	q_b_15,
	q_b_14,
	q_b_13,
	q_b_12,
	q_b_11,
	q_b_10,
	ram_in_reg_1_7,
	ram_in_reg_0_7,
	ram_in_reg_7_7,
	ram_in_reg_6_7,
	ram_in_reg_5_7,
	ram_in_reg_4_7,
	ram_in_reg_3_7,
	ram_in_reg_2_7,
	ram_in_reg_1_3,
	ram_in_reg_0_3,
	ram_in_reg_7_3,
	ram_in_reg_6_3,
	ram_in_reg_5_3,
	ram_in_reg_4_3,
	ram_in_reg_3_3,
	ram_in_reg_2_3,
	global_clock_enable,
	ram_in_reg_6_0,
	rdaddress_c_bus_0,
	rdaddress_c_bus_15,
	rdaddress_c_bus_16,
	rdaddress_c_bus_10,
	rdaddress_c_bus_11,
	rdaddress_c_bus_12,
	wd_vec_6,
	ram_in_reg_0_1,
	ram_in_reg_2_1,
	ram_in_reg_4_1,
	rdaddress_c_bus_20,
	ram_in_reg_1_31,
	ram_in_reg_3_31,
	ram_in_reg_5_31,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_1;
output 	q_b_0;
output 	q_b_7;
output 	q_b_6;
output 	q_b_5;
output 	q_b_4;
output 	q_b_3;
output 	q_b_2;
output 	q_b_9;
output 	q_b_8;
output 	q_b_15;
output 	q_b_14;
output 	q_b_13;
output 	q_b_12;
output 	q_b_11;
output 	q_b_10;
input 	ram_in_reg_1_7;
input 	ram_in_reg_0_7;
input 	ram_in_reg_7_7;
input 	ram_in_reg_6_7;
input 	ram_in_reg_5_7;
input 	ram_in_reg_4_7;
input 	ram_in_reg_3_7;
input 	ram_in_reg_2_7;
input 	ram_in_reg_1_3;
input 	ram_in_reg_0_3;
input 	ram_in_reg_7_3;
input 	ram_in_reg_6_3;
input 	ram_in_reg_5_3;
input 	ram_in_reg_4_3;
input 	ram_in_reg_3_3;
input 	ram_in_reg_2_3;
input 	global_clock_enable;
input 	ram_in_reg_6_0;
input 	rdaddress_c_bus_0;
input 	rdaddress_c_bus_15;
input 	rdaddress_c_bus_16;
input 	rdaddress_c_bus_10;
input 	rdaddress_c_bus_11;
input 	rdaddress_c_bus_12;
input 	wd_vec_6;
input 	ram_in_reg_0_1;
input 	ram_in_reg_2_1;
input 	ram_in_reg_4_1;
input 	rdaddress_c_bus_20;
input 	ram_in_reg_1_31;
input 	ram_in_reg_3_31;
input 	ram_in_reg_5_31;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_altsyncram_14 \gen_M4K:altsyncram_component (
	.q_b({q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.data_a({ram_in_reg_7_3,ram_in_reg_6_3,ram_in_reg_5_3,ram_in_reg_4_3,ram_in_reg_3_3,ram_in_reg_2_3,ram_in_reg_1_3,ram_in_reg_0_3,ram_in_reg_7_7,ram_in_reg_6_7,ram_in_reg_5_7,ram_in_reg_4_7,ram_in_reg_3_7,ram_in_reg_2_7,ram_in_reg_1_7,ram_in_reg_0_7}),
	.clocken0(global_clock_enable),
	.address_a({ram_in_reg_6_0,ram_in_reg_5_31,ram_in_reg_4_1,ram_in_reg_3_31,ram_in_reg_2_1,ram_in_reg_1_31,ram_in_reg_0_1}),
	.address_b({rdaddress_c_bus_20,rdaddress_c_bus_12,rdaddress_c_bus_11,rdaddress_c_bus_10,rdaddress_c_bus_16,rdaddress_c_bus_15,rdaddress_c_bus_0}),
	.wren_a(wd_vec_6),
	.clock0(clk));

endmodule

module fft_altsyncram_14 (
	q_b,
	data_a,
	clocken0,
	address_a,
	address_b,
	wren_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	[15:0] data_a;
input 	clocken0;
input 	[6:0] address_a;
input 	[6:0] address_b;
input 	wren_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_altsyncram_lmu3_7 auto_generated(
	.q_b({q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.data_a({data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.clocken0(clocken0),
	.address_a({address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.wren_a(wren_a),
	.clock0(clock0));

endmodule

module fft_altsyncram_lmu3_7 (
	q_b,
	data_a,
	clocken0,
	address_a,
	address_b,
	wren_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	[15:0] data_a;
input 	clocken0;
input 	[6:0] address_a;
input 	[6:0] address_b;
input 	wren_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

cycloneiii_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "old";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 7;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 127;
defparam ram_block1a1.port_a_logical_ram_depth = 128;
defparam ram_block1a1.port_a_logical_ram_width = 16;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 7;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "clock0";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 127;
defparam ram_block1a1.port_b_logical_ram_depth = 128;
defparam ram_block1a1.port_b_logical_ram_width = 16;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "old";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 7;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 127;
defparam ram_block1a0.port_a_logical_ram_depth = 128;
defparam ram_block1a0.port_a_logical_ram_width = 16;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 7;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "clock0";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 127;
defparam ram_block1a0.port_b_logical_ram_depth = 128;
defparam ram_block1a0.port_b_logical_ram_width = 16;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "old";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 7;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 127;
defparam ram_block1a7.port_a_logical_ram_depth = 128;
defparam ram_block1a7.port_a_logical_ram_width = 16;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 7;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "clock0";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 127;
defparam ram_block1a7.port_b_logical_ram_depth = 128;
defparam ram_block1a7.port_b_logical_ram_width = 16;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "old";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 7;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 127;
defparam ram_block1a6.port_a_logical_ram_depth = 128;
defparam ram_block1a6.port_a_logical_ram_width = 16;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 7;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "clock0";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 127;
defparam ram_block1a6.port_b_logical_ram_depth = 128;
defparam ram_block1a6.port_b_logical_ram_width = 16;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "old";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 7;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 127;
defparam ram_block1a5.port_a_logical_ram_depth = 128;
defparam ram_block1a5.port_a_logical_ram_width = 16;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 7;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "clock0";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 127;
defparam ram_block1a5.port_b_logical_ram_depth = 128;
defparam ram_block1a5.port_b_logical_ram_width = 16;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "old";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 7;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 127;
defparam ram_block1a4.port_a_logical_ram_depth = 128;
defparam ram_block1a4.port_a_logical_ram_width = 16;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 7;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "clock0";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 127;
defparam ram_block1a4.port_b_logical_ram_depth = 128;
defparam ram_block1a4.port_b_logical_ram_width = 16;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "old";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 7;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 127;
defparam ram_block1a3.port_a_logical_ram_depth = 128;
defparam ram_block1a3.port_a_logical_ram_width = 16;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 7;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "clock0";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 127;
defparam ram_block1a3.port_b_logical_ram_depth = 128;
defparam ram_block1a3.port_b_logical_ram_width = 16;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "old";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 7;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 127;
defparam ram_block1a2.port_a_logical_ram_depth = 128;
defparam ram_block1a2.port_a_logical_ram_width = 16;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 7;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "clock0";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 127;
defparam ram_block1a2.port_b_logical_ram_depth = 128;
defparam ram_block1a2.port_b_logical_ram_width = 16;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.clk0_output_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "old";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 7;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 127;
defparam ram_block1a9.port_a_logical_ram_depth = 128;
defparam ram_block1a9.port_a_logical_ram_width = 16;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 7;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "clock0";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 127;
defparam ram_block1a9.port_b_logical_ram_depth = 128;
defparam ram_block1a9.port_b_logical_ram_width = 16;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.clk0_output_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "old";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 7;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 127;
defparam ram_block1a8.port_a_logical_ram_depth = 128;
defparam ram_block1a8.port_a_logical_ram_width = 16;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 7;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "clock0";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 127;
defparam ram_block1a8.port_b_logical_ram_depth = 128;
defparam ram_block1a8.port_b_logical_ram_width = 16;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.clk0_output_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "old";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 7;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 127;
defparam ram_block1a15.port_a_logical_ram_depth = 128;
defparam ram_block1a15.port_a_logical_ram_width = 16;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 7;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "clock0";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 127;
defparam ram_block1a15.port_b_logical_ram_depth = 128;
defparam ram_block1a15.port_b_logical_ram_width = 16;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.clk0_output_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "old";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 7;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 127;
defparam ram_block1a14.port_a_logical_ram_depth = 128;
defparam ram_block1a14.port_a_logical_ram_width = 16;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 7;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "clock0";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 127;
defparam ram_block1a14.port_b_logical_ram_depth = 128;
defparam ram_block1a14.port_b_logical_ram_width = 16;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.clk0_output_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "old";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 7;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 127;
defparam ram_block1a13.port_a_logical_ram_depth = 128;
defparam ram_block1a13.port_a_logical_ram_width = 16;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 7;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "clock0";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 127;
defparam ram_block1a13.port_b_logical_ram_depth = 128;
defparam ram_block1a13.port_b_logical_ram_width = 16;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.clk0_output_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "old";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 7;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 127;
defparam ram_block1a12.port_a_logical_ram_depth = 128;
defparam ram_block1a12.port_a_logical_ram_width = 16;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 7;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "clock0";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 127;
defparam ram_block1a12.port_b_logical_ram_depth = 128;
defparam ram_block1a12.port_b_logical_ram_width = 16;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.clk0_output_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "old";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 7;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 127;
defparam ram_block1a11.port_a_logical_ram_depth = 128;
defparam ram_block1a11.port_a_logical_ram_width = 16;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 7;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "clock0";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 127;
defparam ram_block1a11.port_b_logical_ram_depth = 128;
defparam ram_block1a11.port_b_logical_ram_width = 16;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.clk0_output_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:\\gen_M4K_Output:dat_D|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "old";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 7;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 127;
defparam ram_block1a10.port_a_logical_ram_depth = 128;
defparam ram_block1a10.port_a_logical_ram_width = 16;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 7;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "clock0";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 127;
defparam ram_block1a10.port_b_logical_ram_depth = 128;
defparam ram_block1a10.port_b_logical_ram_width = 16;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";

endmodule

module fft_asj_fft_4dp_ram_fft_120_2 (
	q_b_10,
	q_b_101,
	q_b_102,
	q_b_103,
	q_b_14,
	q_b_141,
	q_b_142,
	q_b_143,
	q_b_12,
	q_b_121,
	q_b_122,
	q_b_123,
	q_b_11,
	q_b_111,
	q_b_112,
	q_b_113,
	q_b_13,
	q_b_131,
	q_b_132,
	q_b_133,
	q_b_9,
	q_b_91,
	q_b_92,
	q_b_93,
	q_b_8,
	q_b_81,
	q_b_82,
	q_b_83,
	q_b_15,
	q_b_151,
	q_b_152,
	q_b_153,
	q_b_7,
	q_b_71,
	q_b_72,
	q_b_73,
	q_b_3,
	q_b_31,
	q_b_32,
	q_b_33,
	q_b_5,
	q_b_51,
	q_b_52,
	q_b_53,
	q_b_4,
	q_b_41,
	q_b_42,
	q_b_43,
	q_b_6,
	q_b_61,
	q_b_62,
	q_b_63,
	q_b_2,
	q_b_21,
	q_b_22,
	q_b_23,
	q_b_1,
	q_b_16,
	q_b_17,
	q_b_18,
	q_b_0,
	q_b_01,
	q_b_02,
	q_b_03,
	wren_a_0,
	wren_a_1,
	wren_a_2,
	wren_a_3,
	global_clock_enable,
	a_ram_data_in_bus_58,
	wraddress_a_bus_21,
	wraddress_a_bus_22,
	wraddress_a_bus_23,
	wraddress_a_bus_24,
	wraddress_a_bus_11,
	wraddress_a_bus_26,
	wraddress_a_bus_13,
	rdaddress_a_bus_21,
	rdaddress_a_bus_22,
	rdaddress_a_bus_23,
	rdaddress_a_bus_24,
	rdaddress_a_bus_11,
	rdaddress_a_bus_26,
	rdaddress_a_bus_13,
	a_ram_data_in_bus_42,
	wraddress_a_bus_0,
	wraddress_a_bus_15,
	wraddress_a_bus_16,
	wraddress_a_bus_17,
	wraddress_a_bus_18,
	wraddress_a_bus_19,
	rdaddress_a_bus_0,
	rdaddress_a_bus_15,
	rdaddress_a_bus_16,
	rdaddress_a_bus_17,
	rdaddress_a_bus_18,
	rdaddress_a_bus_19,
	a_ram_data_in_bus_26,
	wraddress_a_bus_8,
	wraddress_a_bus_10,
	wraddress_a_bus_12,
	rdaddress_a_bus_8,
	rdaddress_a_bus_10,
	rdaddress_a_bus_12,
	a_ram_data_in_bus_10,
	wraddress_a_bus_1,
	wraddress_a_bus_3,
	wraddress_a_bus_5,
	rdaddress_a_bus_1,
	rdaddress_a_bus_3,
	rdaddress_a_bus_5,
	a_ram_data_in_bus_62,
	a_ram_data_in_bus_46,
	a_ram_data_in_bus_30,
	a_ram_data_in_bus_14,
	a_ram_data_in_bus_60,
	a_ram_data_in_bus_44,
	a_ram_data_in_bus_28,
	a_ram_data_in_bus_12,
	a_ram_data_in_bus_59,
	a_ram_data_in_bus_43,
	a_ram_data_in_bus_27,
	a_ram_data_in_bus_11,
	a_ram_data_in_bus_61,
	a_ram_data_in_bus_45,
	a_ram_data_in_bus_29,
	a_ram_data_in_bus_13,
	a_ram_data_in_bus_57,
	a_ram_data_in_bus_41,
	a_ram_data_in_bus_25,
	a_ram_data_in_bus_9,
	a_ram_data_in_bus_56,
	a_ram_data_in_bus_40,
	a_ram_data_in_bus_24,
	a_ram_data_in_bus_8,
	a_ram_data_in_bus_63,
	a_ram_data_in_bus_47,
	a_ram_data_in_bus_31,
	a_ram_data_in_bus_15,
	a_ram_data_in_bus_55,
	a_ram_data_in_bus_39,
	a_ram_data_in_bus_23,
	a_ram_data_in_bus_7,
	a_ram_data_in_bus_51,
	a_ram_data_in_bus_35,
	a_ram_data_in_bus_19,
	a_ram_data_in_bus_3,
	a_ram_data_in_bus_53,
	a_ram_data_in_bus_37,
	a_ram_data_in_bus_21,
	a_ram_data_in_bus_5,
	a_ram_data_in_bus_52,
	a_ram_data_in_bus_36,
	a_ram_data_in_bus_20,
	a_ram_data_in_bus_4,
	a_ram_data_in_bus_54,
	a_ram_data_in_bus_38,
	a_ram_data_in_bus_22,
	a_ram_data_in_bus_6,
	a_ram_data_in_bus_50,
	a_ram_data_in_bus_34,
	a_ram_data_in_bus_18,
	a_ram_data_in_bus_2,
	a_ram_data_in_bus_49,
	a_ram_data_in_bus_33,
	a_ram_data_in_bus_17,
	a_ram_data_in_bus_1,
	a_ram_data_in_bus_48,
	a_ram_data_in_bus_32,
	a_ram_data_in_bus_16,
	a_ram_data_in_bus_0,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_10;
output 	q_b_101;
output 	q_b_102;
output 	q_b_103;
output 	q_b_14;
output 	q_b_141;
output 	q_b_142;
output 	q_b_143;
output 	q_b_12;
output 	q_b_121;
output 	q_b_122;
output 	q_b_123;
output 	q_b_11;
output 	q_b_111;
output 	q_b_112;
output 	q_b_113;
output 	q_b_13;
output 	q_b_131;
output 	q_b_132;
output 	q_b_133;
output 	q_b_9;
output 	q_b_91;
output 	q_b_92;
output 	q_b_93;
output 	q_b_8;
output 	q_b_81;
output 	q_b_82;
output 	q_b_83;
output 	q_b_15;
output 	q_b_151;
output 	q_b_152;
output 	q_b_153;
output 	q_b_7;
output 	q_b_71;
output 	q_b_72;
output 	q_b_73;
output 	q_b_3;
output 	q_b_31;
output 	q_b_32;
output 	q_b_33;
output 	q_b_5;
output 	q_b_51;
output 	q_b_52;
output 	q_b_53;
output 	q_b_4;
output 	q_b_41;
output 	q_b_42;
output 	q_b_43;
output 	q_b_6;
output 	q_b_61;
output 	q_b_62;
output 	q_b_63;
output 	q_b_2;
output 	q_b_21;
output 	q_b_22;
output 	q_b_23;
output 	q_b_1;
output 	q_b_16;
output 	q_b_17;
output 	q_b_18;
output 	q_b_0;
output 	q_b_01;
output 	q_b_02;
output 	q_b_03;
input 	wren_a_0;
input 	wren_a_1;
input 	wren_a_2;
input 	wren_a_3;
input 	global_clock_enable;
input 	a_ram_data_in_bus_58;
input 	wraddress_a_bus_21;
input 	wraddress_a_bus_22;
input 	wraddress_a_bus_23;
input 	wraddress_a_bus_24;
input 	wraddress_a_bus_11;
input 	wraddress_a_bus_26;
input 	wraddress_a_bus_13;
input 	rdaddress_a_bus_21;
input 	rdaddress_a_bus_22;
input 	rdaddress_a_bus_23;
input 	rdaddress_a_bus_24;
input 	rdaddress_a_bus_11;
input 	rdaddress_a_bus_26;
input 	rdaddress_a_bus_13;
input 	a_ram_data_in_bus_42;
input 	wraddress_a_bus_0;
input 	wraddress_a_bus_15;
input 	wraddress_a_bus_16;
input 	wraddress_a_bus_17;
input 	wraddress_a_bus_18;
input 	wraddress_a_bus_19;
input 	rdaddress_a_bus_0;
input 	rdaddress_a_bus_15;
input 	rdaddress_a_bus_16;
input 	rdaddress_a_bus_17;
input 	rdaddress_a_bus_18;
input 	rdaddress_a_bus_19;
input 	a_ram_data_in_bus_26;
input 	wraddress_a_bus_8;
input 	wraddress_a_bus_10;
input 	wraddress_a_bus_12;
input 	rdaddress_a_bus_8;
input 	rdaddress_a_bus_10;
input 	rdaddress_a_bus_12;
input 	a_ram_data_in_bus_10;
input 	wraddress_a_bus_1;
input 	wraddress_a_bus_3;
input 	wraddress_a_bus_5;
input 	rdaddress_a_bus_1;
input 	rdaddress_a_bus_3;
input 	rdaddress_a_bus_5;
input 	a_ram_data_in_bus_62;
input 	a_ram_data_in_bus_46;
input 	a_ram_data_in_bus_30;
input 	a_ram_data_in_bus_14;
input 	a_ram_data_in_bus_60;
input 	a_ram_data_in_bus_44;
input 	a_ram_data_in_bus_28;
input 	a_ram_data_in_bus_12;
input 	a_ram_data_in_bus_59;
input 	a_ram_data_in_bus_43;
input 	a_ram_data_in_bus_27;
input 	a_ram_data_in_bus_11;
input 	a_ram_data_in_bus_61;
input 	a_ram_data_in_bus_45;
input 	a_ram_data_in_bus_29;
input 	a_ram_data_in_bus_13;
input 	a_ram_data_in_bus_57;
input 	a_ram_data_in_bus_41;
input 	a_ram_data_in_bus_25;
input 	a_ram_data_in_bus_9;
input 	a_ram_data_in_bus_56;
input 	a_ram_data_in_bus_40;
input 	a_ram_data_in_bus_24;
input 	a_ram_data_in_bus_8;
input 	a_ram_data_in_bus_63;
input 	a_ram_data_in_bus_47;
input 	a_ram_data_in_bus_31;
input 	a_ram_data_in_bus_15;
input 	a_ram_data_in_bus_55;
input 	a_ram_data_in_bus_39;
input 	a_ram_data_in_bus_23;
input 	a_ram_data_in_bus_7;
input 	a_ram_data_in_bus_51;
input 	a_ram_data_in_bus_35;
input 	a_ram_data_in_bus_19;
input 	a_ram_data_in_bus_3;
input 	a_ram_data_in_bus_53;
input 	a_ram_data_in_bus_37;
input 	a_ram_data_in_bus_21;
input 	a_ram_data_in_bus_5;
input 	a_ram_data_in_bus_52;
input 	a_ram_data_in_bus_36;
input 	a_ram_data_in_bus_20;
input 	a_ram_data_in_bus_4;
input 	a_ram_data_in_bus_54;
input 	a_ram_data_in_bus_38;
input 	a_ram_data_in_bus_22;
input 	a_ram_data_in_bus_6;
input 	a_ram_data_in_bus_50;
input 	a_ram_data_in_bus_34;
input 	a_ram_data_in_bus_18;
input 	a_ram_data_in_bus_2;
input 	a_ram_data_in_bus_49;
input 	a_ram_data_in_bus_33;
input 	a_ram_data_in_bus_17;
input 	a_ram_data_in_bus_1;
input 	a_ram_data_in_bus_48;
input 	a_ram_data_in_bus_32;
input 	a_ram_data_in_bus_16;
input 	a_ram_data_in_bus_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_asj_fft_data_ram_fft_120_11 \gen_rams:3:dat_A (
	.q_b_10(q_b_103),
	.q_b_14(q_b_143),
	.q_b_12(q_b_123),
	.q_b_11(q_b_113),
	.q_b_13(q_b_133),
	.q_b_9(q_b_93),
	.q_b_8(q_b_83),
	.q_b_15(q_b_153),
	.q_b_7(q_b_73),
	.q_b_3(q_b_33),
	.q_b_5(q_b_53),
	.q_b_4(q_b_43),
	.q_b_6(q_b_63),
	.q_b_2(q_b_23),
	.q_b_1(q_b_18),
	.q_b_0(q_b_03),
	.wren_a_3(wren_a_3),
	.global_clock_enable(global_clock_enable),
	.wraddress_a_bus_13(wraddress_a_bus_13),
	.rdaddress_a_bus_13(rdaddress_a_bus_13),
	.wraddress_a_bus_0(wraddress_a_bus_0),
	.wraddress_a_bus_16(wraddress_a_bus_16),
	.wraddress_a_bus_18(wraddress_a_bus_18),
	.rdaddress_a_bus_0(rdaddress_a_bus_0),
	.rdaddress_a_bus_16(rdaddress_a_bus_16),
	.rdaddress_a_bus_18(rdaddress_a_bus_18),
	.a_ram_data_in_bus_10(a_ram_data_in_bus_10),
	.wraddress_a_bus_1(wraddress_a_bus_1),
	.wraddress_a_bus_3(wraddress_a_bus_3),
	.wraddress_a_bus_5(wraddress_a_bus_5),
	.rdaddress_a_bus_1(rdaddress_a_bus_1),
	.rdaddress_a_bus_3(rdaddress_a_bus_3),
	.rdaddress_a_bus_5(rdaddress_a_bus_5),
	.a_ram_data_in_bus_14(a_ram_data_in_bus_14),
	.a_ram_data_in_bus_12(a_ram_data_in_bus_12),
	.a_ram_data_in_bus_11(a_ram_data_in_bus_11),
	.a_ram_data_in_bus_13(a_ram_data_in_bus_13),
	.a_ram_data_in_bus_9(a_ram_data_in_bus_9),
	.a_ram_data_in_bus_8(a_ram_data_in_bus_8),
	.a_ram_data_in_bus_15(a_ram_data_in_bus_15),
	.a_ram_data_in_bus_7(a_ram_data_in_bus_7),
	.a_ram_data_in_bus_3(a_ram_data_in_bus_3),
	.a_ram_data_in_bus_5(a_ram_data_in_bus_5),
	.a_ram_data_in_bus_4(a_ram_data_in_bus_4),
	.a_ram_data_in_bus_6(a_ram_data_in_bus_6),
	.a_ram_data_in_bus_2(a_ram_data_in_bus_2),
	.a_ram_data_in_bus_1(a_ram_data_in_bus_1),
	.a_ram_data_in_bus_0(a_ram_data_in_bus_0),
	.clk(clk));

fft_asj_fft_data_ram_fft_120_10 \gen_rams:2:dat_A (
	.q_b_10(q_b_102),
	.q_b_14(q_b_142),
	.q_b_12(q_b_122),
	.q_b_11(q_b_112),
	.q_b_13(q_b_132),
	.q_b_9(q_b_92),
	.q_b_8(q_b_82),
	.q_b_15(q_b_152),
	.q_b_7(q_b_72),
	.q_b_3(q_b_32),
	.q_b_5(q_b_52),
	.q_b_4(q_b_42),
	.q_b_6(q_b_62),
	.q_b_2(q_b_22),
	.q_b_1(q_b_17),
	.q_b_0(q_b_02),
	.wren_a_2(wren_a_2),
	.global_clock_enable(global_clock_enable),
	.wraddress_a_bus_21(wraddress_a_bus_21),
	.wraddress_a_bus_23(wraddress_a_bus_23),
	.wraddress_a_bus_11(wraddress_a_bus_11),
	.wraddress_a_bus_13(wraddress_a_bus_13),
	.rdaddress_a_bus_21(rdaddress_a_bus_21),
	.rdaddress_a_bus_23(rdaddress_a_bus_23),
	.rdaddress_a_bus_11(rdaddress_a_bus_11),
	.rdaddress_a_bus_13(rdaddress_a_bus_13),
	.a_ram_data_in_bus_26(a_ram_data_in_bus_26),
	.wraddress_a_bus_8(wraddress_a_bus_8),
	.wraddress_a_bus_10(wraddress_a_bus_10),
	.wraddress_a_bus_12(wraddress_a_bus_12),
	.rdaddress_a_bus_8(rdaddress_a_bus_8),
	.rdaddress_a_bus_10(rdaddress_a_bus_10),
	.rdaddress_a_bus_12(rdaddress_a_bus_12),
	.a_ram_data_in_bus_30(a_ram_data_in_bus_30),
	.a_ram_data_in_bus_28(a_ram_data_in_bus_28),
	.a_ram_data_in_bus_27(a_ram_data_in_bus_27),
	.a_ram_data_in_bus_29(a_ram_data_in_bus_29),
	.a_ram_data_in_bus_25(a_ram_data_in_bus_25),
	.a_ram_data_in_bus_24(a_ram_data_in_bus_24),
	.a_ram_data_in_bus_31(a_ram_data_in_bus_31),
	.a_ram_data_in_bus_23(a_ram_data_in_bus_23),
	.a_ram_data_in_bus_19(a_ram_data_in_bus_19),
	.a_ram_data_in_bus_21(a_ram_data_in_bus_21),
	.a_ram_data_in_bus_20(a_ram_data_in_bus_20),
	.a_ram_data_in_bus_22(a_ram_data_in_bus_22),
	.a_ram_data_in_bus_18(a_ram_data_in_bus_18),
	.a_ram_data_in_bus_17(a_ram_data_in_bus_17),
	.a_ram_data_in_bus_16(a_ram_data_in_bus_16),
	.clk(clk));

fft_asj_fft_data_ram_fft_120_9 \gen_rams:1:dat_A (
	.q_b_10(q_b_101),
	.q_b_14(q_b_141),
	.q_b_12(q_b_121),
	.q_b_11(q_b_111),
	.q_b_13(q_b_131),
	.q_b_9(q_b_91),
	.q_b_8(q_b_81),
	.q_b_15(q_b_151),
	.q_b_7(q_b_71),
	.q_b_3(q_b_31),
	.q_b_5(q_b_51),
	.q_b_4(q_b_41),
	.q_b_6(q_b_61),
	.q_b_2(q_b_21),
	.q_b_1(q_b_16),
	.q_b_0(q_b_01),
	.wren_a_1(wren_a_1),
	.global_clock_enable(global_clock_enable),
	.wraddress_a_bus_13(wraddress_a_bus_13),
	.rdaddress_a_bus_13(rdaddress_a_bus_13),
	.a_ram_data_in_bus_42(a_ram_data_in_bus_42),
	.wraddress_a_bus_0(wraddress_a_bus_0),
	.wraddress_a_bus_15(wraddress_a_bus_15),
	.wraddress_a_bus_16(wraddress_a_bus_16),
	.wraddress_a_bus_17(wraddress_a_bus_17),
	.wraddress_a_bus_18(wraddress_a_bus_18),
	.wraddress_a_bus_19(wraddress_a_bus_19),
	.rdaddress_a_bus_0(rdaddress_a_bus_0),
	.rdaddress_a_bus_15(rdaddress_a_bus_15),
	.rdaddress_a_bus_16(rdaddress_a_bus_16),
	.rdaddress_a_bus_17(rdaddress_a_bus_17),
	.rdaddress_a_bus_18(rdaddress_a_bus_18),
	.rdaddress_a_bus_19(rdaddress_a_bus_19),
	.a_ram_data_in_bus_46(a_ram_data_in_bus_46),
	.a_ram_data_in_bus_44(a_ram_data_in_bus_44),
	.a_ram_data_in_bus_43(a_ram_data_in_bus_43),
	.a_ram_data_in_bus_45(a_ram_data_in_bus_45),
	.a_ram_data_in_bus_41(a_ram_data_in_bus_41),
	.a_ram_data_in_bus_40(a_ram_data_in_bus_40),
	.a_ram_data_in_bus_47(a_ram_data_in_bus_47),
	.a_ram_data_in_bus_39(a_ram_data_in_bus_39),
	.a_ram_data_in_bus_35(a_ram_data_in_bus_35),
	.a_ram_data_in_bus_37(a_ram_data_in_bus_37),
	.a_ram_data_in_bus_36(a_ram_data_in_bus_36),
	.a_ram_data_in_bus_38(a_ram_data_in_bus_38),
	.a_ram_data_in_bus_34(a_ram_data_in_bus_34),
	.a_ram_data_in_bus_33(a_ram_data_in_bus_33),
	.a_ram_data_in_bus_32(a_ram_data_in_bus_32),
	.clk(clk));

fft_asj_fft_data_ram_fft_120_8 \gen_rams:0:dat_A (
	.q_b_10(q_b_10),
	.q_b_14(q_b_14),
	.q_b_12(q_b_12),
	.q_b_11(q_b_11),
	.q_b_13(q_b_13),
	.q_b_9(q_b_9),
	.q_b_8(q_b_8),
	.q_b_15(q_b_15),
	.q_b_7(q_b_7),
	.q_b_3(q_b_3),
	.q_b_5(q_b_5),
	.q_b_4(q_b_4),
	.q_b_6(q_b_6),
	.q_b_2(q_b_2),
	.q_b_1(q_b_1),
	.q_b_0(q_b_0),
	.wren_a_0(wren_a_0),
	.global_clock_enable(global_clock_enable),
	.a_ram_data_in_bus_58(a_ram_data_in_bus_58),
	.wraddress_a_bus_21(wraddress_a_bus_21),
	.wraddress_a_bus_22(wraddress_a_bus_22),
	.wraddress_a_bus_23(wraddress_a_bus_23),
	.wraddress_a_bus_24(wraddress_a_bus_24),
	.wraddress_a_bus_11(wraddress_a_bus_11),
	.wraddress_a_bus_26(wraddress_a_bus_26),
	.wraddress_a_bus_13(wraddress_a_bus_13),
	.rdaddress_a_bus_21(rdaddress_a_bus_21),
	.rdaddress_a_bus_22(rdaddress_a_bus_22),
	.rdaddress_a_bus_23(rdaddress_a_bus_23),
	.rdaddress_a_bus_24(rdaddress_a_bus_24),
	.rdaddress_a_bus_11(rdaddress_a_bus_11),
	.rdaddress_a_bus_26(rdaddress_a_bus_26),
	.rdaddress_a_bus_13(rdaddress_a_bus_13),
	.a_ram_data_in_bus_62(a_ram_data_in_bus_62),
	.a_ram_data_in_bus_60(a_ram_data_in_bus_60),
	.a_ram_data_in_bus_59(a_ram_data_in_bus_59),
	.a_ram_data_in_bus_61(a_ram_data_in_bus_61),
	.a_ram_data_in_bus_57(a_ram_data_in_bus_57),
	.a_ram_data_in_bus_56(a_ram_data_in_bus_56),
	.a_ram_data_in_bus_63(a_ram_data_in_bus_63),
	.a_ram_data_in_bus_55(a_ram_data_in_bus_55),
	.a_ram_data_in_bus_51(a_ram_data_in_bus_51),
	.a_ram_data_in_bus_53(a_ram_data_in_bus_53),
	.a_ram_data_in_bus_52(a_ram_data_in_bus_52),
	.a_ram_data_in_bus_54(a_ram_data_in_bus_54),
	.a_ram_data_in_bus_50(a_ram_data_in_bus_50),
	.a_ram_data_in_bus_49(a_ram_data_in_bus_49),
	.a_ram_data_in_bus_48(a_ram_data_in_bus_48),
	.clk(clk));

endmodule

module fft_asj_fft_data_ram_fft_120_8 (
	q_b_10,
	q_b_14,
	q_b_12,
	q_b_11,
	q_b_13,
	q_b_9,
	q_b_8,
	q_b_15,
	q_b_7,
	q_b_3,
	q_b_5,
	q_b_4,
	q_b_6,
	q_b_2,
	q_b_1,
	q_b_0,
	wren_a_0,
	global_clock_enable,
	a_ram_data_in_bus_58,
	wraddress_a_bus_21,
	wraddress_a_bus_22,
	wraddress_a_bus_23,
	wraddress_a_bus_24,
	wraddress_a_bus_11,
	wraddress_a_bus_26,
	wraddress_a_bus_13,
	rdaddress_a_bus_21,
	rdaddress_a_bus_22,
	rdaddress_a_bus_23,
	rdaddress_a_bus_24,
	rdaddress_a_bus_11,
	rdaddress_a_bus_26,
	rdaddress_a_bus_13,
	a_ram_data_in_bus_62,
	a_ram_data_in_bus_60,
	a_ram_data_in_bus_59,
	a_ram_data_in_bus_61,
	a_ram_data_in_bus_57,
	a_ram_data_in_bus_56,
	a_ram_data_in_bus_63,
	a_ram_data_in_bus_55,
	a_ram_data_in_bus_51,
	a_ram_data_in_bus_53,
	a_ram_data_in_bus_52,
	a_ram_data_in_bus_54,
	a_ram_data_in_bus_50,
	a_ram_data_in_bus_49,
	a_ram_data_in_bus_48,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_10;
output 	q_b_14;
output 	q_b_12;
output 	q_b_11;
output 	q_b_13;
output 	q_b_9;
output 	q_b_8;
output 	q_b_15;
output 	q_b_7;
output 	q_b_3;
output 	q_b_5;
output 	q_b_4;
output 	q_b_6;
output 	q_b_2;
output 	q_b_1;
output 	q_b_0;
input 	wren_a_0;
input 	global_clock_enable;
input 	a_ram_data_in_bus_58;
input 	wraddress_a_bus_21;
input 	wraddress_a_bus_22;
input 	wraddress_a_bus_23;
input 	wraddress_a_bus_24;
input 	wraddress_a_bus_11;
input 	wraddress_a_bus_26;
input 	wraddress_a_bus_13;
input 	rdaddress_a_bus_21;
input 	rdaddress_a_bus_22;
input 	rdaddress_a_bus_23;
input 	rdaddress_a_bus_24;
input 	rdaddress_a_bus_11;
input 	rdaddress_a_bus_26;
input 	rdaddress_a_bus_13;
input 	a_ram_data_in_bus_62;
input 	a_ram_data_in_bus_60;
input 	a_ram_data_in_bus_59;
input 	a_ram_data_in_bus_61;
input 	a_ram_data_in_bus_57;
input 	a_ram_data_in_bus_56;
input 	a_ram_data_in_bus_63;
input 	a_ram_data_in_bus_55;
input 	a_ram_data_in_bus_51;
input 	a_ram_data_in_bus_53;
input 	a_ram_data_in_bus_52;
input 	a_ram_data_in_bus_54;
input 	a_ram_data_in_bus_50;
input 	a_ram_data_in_bus_49;
input 	a_ram_data_in_bus_48;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_altsyncram_15 \gen_M4K:altsyncram_component (
	.q_b({q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.wren_a(wren_a_0),
	.clocken0(global_clock_enable),
	.data_a({a_ram_data_in_bus_63,a_ram_data_in_bus_62,a_ram_data_in_bus_61,a_ram_data_in_bus_60,a_ram_data_in_bus_59,a_ram_data_in_bus_58,a_ram_data_in_bus_57,a_ram_data_in_bus_56,a_ram_data_in_bus_55,a_ram_data_in_bus_54,a_ram_data_in_bus_53,a_ram_data_in_bus_52,
a_ram_data_in_bus_51,a_ram_data_in_bus_50,a_ram_data_in_bus_49,a_ram_data_in_bus_48}),
	.address_a({wraddress_a_bus_13,wraddress_a_bus_26,wraddress_a_bus_11,wraddress_a_bus_24,wraddress_a_bus_23,wraddress_a_bus_22,wraddress_a_bus_21}),
	.address_b({rdaddress_a_bus_13,rdaddress_a_bus_26,rdaddress_a_bus_11,rdaddress_a_bus_24,rdaddress_a_bus_23,rdaddress_a_bus_22,rdaddress_a_bus_21}),
	.clock0(clk));

endmodule

module fft_altsyncram_15 (
	q_b,
	wren_a,
	clocken0,
	data_a,
	address_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	wren_a;
input 	clocken0;
input 	[15:0] data_a;
input 	[6:0] address_a;
input 	[6:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_altsyncram_lmu3_8 auto_generated(
	.q_b({q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.wren_a(wren_a),
	.clocken0(clocken0),
	.data_a({data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_a({address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.clock0(clock0));

endmodule

module fft_altsyncram_lmu3_8 (
	q_b,
	wren_a,
	clocken0,
	data_a,
	address_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	wren_a;
input 	clocken0;
input 	[15:0] data_a;
input 	[6:0] address_a;
input 	[6:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

cycloneiii_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.clk0_output_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "old";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 7;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 127;
defparam ram_block1a10.port_a_logical_ram_depth = 128;
defparam ram_block1a10.port_a_logical_ram_width = 16;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 7;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "clock0";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 127;
defparam ram_block1a10.port_b_logical_ram_depth = 128;
defparam ram_block1a10.port_b_logical_ram_width = 16;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.clk0_output_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "old";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 7;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 127;
defparam ram_block1a14.port_a_logical_ram_depth = 128;
defparam ram_block1a14.port_a_logical_ram_width = 16;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 7;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "clock0";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 127;
defparam ram_block1a14.port_b_logical_ram_depth = 128;
defparam ram_block1a14.port_b_logical_ram_width = 16;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.clk0_output_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "old";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 7;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 127;
defparam ram_block1a12.port_a_logical_ram_depth = 128;
defparam ram_block1a12.port_a_logical_ram_width = 16;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 7;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "clock0";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 127;
defparam ram_block1a12.port_b_logical_ram_depth = 128;
defparam ram_block1a12.port_b_logical_ram_width = 16;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.clk0_output_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "old";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 7;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 127;
defparam ram_block1a11.port_a_logical_ram_depth = 128;
defparam ram_block1a11.port_a_logical_ram_width = 16;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 7;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "clock0";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 127;
defparam ram_block1a11.port_b_logical_ram_depth = 128;
defparam ram_block1a11.port_b_logical_ram_width = 16;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.clk0_output_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "old";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 7;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 127;
defparam ram_block1a13.port_a_logical_ram_depth = 128;
defparam ram_block1a13.port_a_logical_ram_width = 16;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 7;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "clock0";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 127;
defparam ram_block1a13.port_b_logical_ram_depth = 128;
defparam ram_block1a13.port_b_logical_ram_width = 16;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.clk0_output_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "old";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 7;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 127;
defparam ram_block1a9.port_a_logical_ram_depth = 128;
defparam ram_block1a9.port_a_logical_ram_width = 16;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 7;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "clock0";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 127;
defparam ram_block1a9.port_b_logical_ram_depth = 128;
defparam ram_block1a9.port_b_logical_ram_width = 16;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.clk0_output_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "old";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 7;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 127;
defparam ram_block1a8.port_a_logical_ram_depth = 128;
defparam ram_block1a8.port_a_logical_ram_width = 16;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 7;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "clock0";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 127;
defparam ram_block1a8.port_b_logical_ram_depth = 128;
defparam ram_block1a8.port_b_logical_ram_width = 16;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.clk0_output_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "old";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 7;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 127;
defparam ram_block1a15.port_a_logical_ram_depth = 128;
defparam ram_block1a15.port_a_logical_ram_width = 16;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 7;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "clock0";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 127;
defparam ram_block1a15.port_b_logical_ram_depth = 128;
defparam ram_block1a15.port_b_logical_ram_width = 16;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "old";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 7;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 127;
defparam ram_block1a7.port_a_logical_ram_depth = 128;
defparam ram_block1a7.port_a_logical_ram_width = 16;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 7;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "clock0";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 127;
defparam ram_block1a7.port_b_logical_ram_depth = 128;
defparam ram_block1a7.port_b_logical_ram_width = 16;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "old";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 7;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 127;
defparam ram_block1a3.port_a_logical_ram_depth = 128;
defparam ram_block1a3.port_a_logical_ram_width = 16;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 7;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "clock0";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 127;
defparam ram_block1a3.port_b_logical_ram_depth = 128;
defparam ram_block1a3.port_b_logical_ram_width = 16;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "old";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 7;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 127;
defparam ram_block1a5.port_a_logical_ram_depth = 128;
defparam ram_block1a5.port_a_logical_ram_width = 16;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 7;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "clock0";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 127;
defparam ram_block1a5.port_b_logical_ram_depth = 128;
defparam ram_block1a5.port_b_logical_ram_width = 16;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "old";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 7;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 127;
defparam ram_block1a4.port_a_logical_ram_depth = 128;
defparam ram_block1a4.port_a_logical_ram_width = 16;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 7;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "clock0";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 127;
defparam ram_block1a4.port_b_logical_ram_depth = 128;
defparam ram_block1a4.port_b_logical_ram_width = 16;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "old";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 7;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 127;
defparam ram_block1a6.port_a_logical_ram_depth = 128;
defparam ram_block1a6.port_a_logical_ram_width = 16;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 7;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "clock0";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 127;
defparam ram_block1a6.port_b_logical_ram_depth = 128;
defparam ram_block1a6.port_b_logical_ram_width = 16;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "old";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 7;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 127;
defparam ram_block1a2.port_a_logical_ram_depth = 128;
defparam ram_block1a2.port_a_logical_ram_width = 16;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 7;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "clock0";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 127;
defparam ram_block1a2.port_b_logical_ram_depth = 128;
defparam ram_block1a2.port_b_logical_ram_width = 16;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "old";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 7;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 127;
defparam ram_block1a1.port_a_logical_ram_depth = 128;
defparam ram_block1a1.port_a_logical_ram_width = 16;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 7;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "clock0";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 127;
defparam ram_block1a1.port_b_logical_ram_depth = 128;
defparam ram_block1a1.port_b_logical_ram_width = 16;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "old";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 7;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 127;
defparam ram_block1a0.port_a_logical_ram_depth = 128;
defparam ram_block1a0.port_a_logical_ram_width = 16;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 7;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "clock0";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 127;
defparam ram_block1a0.port_b_logical_ram_depth = 128;
defparam ram_block1a0.port_b_logical_ram_width = 16;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";

endmodule

module fft_asj_fft_data_ram_fft_120_9 (
	q_b_10,
	q_b_14,
	q_b_12,
	q_b_11,
	q_b_13,
	q_b_9,
	q_b_8,
	q_b_15,
	q_b_7,
	q_b_3,
	q_b_5,
	q_b_4,
	q_b_6,
	q_b_2,
	q_b_1,
	q_b_0,
	wren_a_1,
	global_clock_enable,
	wraddress_a_bus_13,
	rdaddress_a_bus_13,
	a_ram_data_in_bus_42,
	wraddress_a_bus_0,
	wraddress_a_bus_15,
	wraddress_a_bus_16,
	wraddress_a_bus_17,
	wraddress_a_bus_18,
	wraddress_a_bus_19,
	rdaddress_a_bus_0,
	rdaddress_a_bus_15,
	rdaddress_a_bus_16,
	rdaddress_a_bus_17,
	rdaddress_a_bus_18,
	rdaddress_a_bus_19,
	a_ram_data_in_bus_46,
	a_ram_data_in_bus_44,
	a_ram_data_in_bus_43,
	a_ram_data_in_bus_45,
	a_ram_data_in_bus_41,
	a_ram_data_in_bus_40,
	a_ram_data_in_bus_47,
	a_ram_data_in_bus_39,
	a_ram_data_in_bus_35,
	a_ram_data_in_bus_37,
	a_ram_data_in_bus_36,
	a_ram_data_in_bus_38,
	a_ram_data_in_bus_34,
	a_ram_data_in_bus_33,
	a_ram_data_in_bus_32,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_10;
output 	q_b_14;
output 	q_b_12;
output 	q_b_11;
output 	q_b_13;
output 	q_b_9;
output 	q_b_8;
output 	q_b_15;
output 	q_b_7;
output 	q_b_3;
output 	q_b_5;
output 	q_b_4;
output 	q_b_6;
output 	q_b_2;
output 	q_b_1;
output 	q_b_0;
input 	wren_a_1;
input 	global_clock_enable;
input 	wraddress_a_bus_13;
input 	rdaddress_a_bus_13;
input 	a_ram_data_in_bus_42;
input 	wraddress_a_bus_0;
input 	wraddress_a_bus_15;
input 	wraddress_a_bus_16;
input 	wraddress_a_bus_17;
input 	wraddress_a_bus_18;
input 	wraddress_a_bus_19;
input 	rdaddress_a_bus_0;
input 	rdaddress_a_bus_15;
input 	rdaddress_a_bus_16;
input 	rdaddress_a_bus_17;
input 	rdaddress_a_bus_18;
input 	rdaddress_a_bus_19;
input 	a_ram_data_in_bus_46;
input 	a_ram_data_in_bus_44;
input 	a_ram_data_in_bus_43;
input 	a_ram_data_in_bus_45;
input 	a_ram_data_in_bus_41;
input 	a_ram_data_in_bus_40;
input 	a_ram_data_in_bus_47;
input 	a_ram_data_in_bus_39;
input 	a_ram_data_in_bus_35;
input 	a_ram_data_in_bus_37;
input 	a_ram_data_in_bus_36;
input 	a_ram_data_in_bus_38;
input 	a_ram_data_in_bus_34;
input 	a_ram_data_in_bus_33;
input 	a_ram_data_in_bus_32;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_altsyncram_16 \gen_M4K:altsyncram_component (
	.q_b({q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.wren_a(wren_a_1),
	.clocken0(global_clock_enable),
	.address_a({wraddress_a_bus_13,wraddress_a_bus_19,wraddress_a_bus_18,wraddress_a_bus_17,wraddress_a_bus_16,wraddress_a_bus_15,wraddress_a_bus_0}),
	.address_b({rdaddress_a_bus_13,rdaddress_a_bus_19,rdaddress_a_bus_18,rdaddress_a_bus_17,rdaddress_a_bus_16,rdaddress_a_bus_15,rdaddress_a_bus_0}),
	.data_a({a_ram_data_in_bus_47,a_ram_data_in_bus_46,a_ram_data_in_bus_45,a_ram_data_in_bus_44,a_ram_data_in_bus_43,a_ram_data_in_bus_42,a_ram_data_in_bus_41,a_ram_data_in_bus_40,a_ram_data_in_bus_39,a_ram_data_in_bus_38,a_ram_data_in_bus_37,a_ram_data_in_bus_36,
a_ram_data_in_bus_35,a_ram_data_in_bus_34,a_ram_data_in_bus_33,a_ram_data_in_bus_32}),
	.clock0(clk));

endmodule

module fft_altsyncram_16 (
	q_b,
	wren_a,
	clocken0,
	address_a,
	address_b,
	data_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	wren_a;
input 	clocken0;
input 	[6:0] address_a;
input 	[6:0] address_b;
input 	[15:0] data_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_altsyncram_lmu3_9 auto_generated(
	.q_b({q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.wren_a(wren_a),
	.clocken0(clocken0),
	.address_a({address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.data_a({data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.clock0(clock0));

endmodule

module fft_altsyncram_lmu3_9 (
	q_b,
	wren_a,
	clocken0,
	address_a,
	address_b,
	data_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	wren_a;
input 	clocken0;
input 	[6:0] address_a;
input 	[6:0] address_b;
input 	[15:0] data_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

cycloneiii_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.clk0_output_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "old";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 7;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 127;
defparam ram_block1a10.port_a_logical_ram_depth = 128;
defparam ram_block1a10.port_a_logical_ram_width = 16;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 7;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "clock0";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 127;
defparam ram_block1a10.port_b_logical_ram_depth = 128;
defparam ram_block1a10.port_b_logical_ram_width = 16;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.clk0_output_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "old";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 7;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 127;
defparam ram_block1a14.port_a_logical_ram_depth = 128;
defparam ram_block1a14.port_a_logical_ram_width = 16;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 7;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "clock0";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 127;
defparam ram_block1a14.port_b_logical_ram_depth = 128;
defparam ram_block1a14.port_b_logical_ram_width = 16;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.clk0_output_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "old";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 7;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 127;
defparam ram_block1a12.port_a_logical_ram_depth = 128;
defparam ram_block1a12.port_a_logical_ram_width = 16;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 7;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "clock0";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 127;
defparam ram_block1a12.port_b_logical_ram_depth = 128;
defparam ram_block1a12.port_b_logical_ram_width = 16;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.clk0_output_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "old";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 7;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 127;
defparam ram_block1a11.port_a_logical_ram_depth = 128;
defparam ram_block1a11.port_a_logical_ram_width = 16;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 7;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "clock0";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 127;
defparam ram_block1a11.port_b_logical_ram_depth = 128;
defparam ram_block1a11.port_b_logical_ram_width = 16;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.clk0_output_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "old";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 7;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 127;
defparam ram_block1a13.port_a_logical_ram_depth = 128;
defparam ram_block1a13.port_a_logical_ram_width = 16;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 7;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "clock0";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 127;
defparam ram_block1a13.port_b_logical_ram_depth = 128;
defparam ram_block1a13.port_b_logical_ram_width = 16;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.clk0_output_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "old";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 7;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 127;
defparam ram_block1a9.port_a_logical_ram_depth = 128;
defparam ram_block1a9.port_a_logical_ram_width = 16;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 7;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "clock0";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 127;
defparam ram_block1a9.port_b_logical_ram_depth = 128;
defparam ram_block1a9.port_b_logical_ram_width = 16;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.clk0_output_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "old";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 7;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 127;
defparam ram_block1a8.port_a_logical_ram_depth = 128;
defparam ram_block1a8.port_a_logical_ram_width = 16;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 7;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "clock0";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 127;
defparam ram_block1a8.port_b_logical_ram_depth = 128;
defparam ram_block1a8.port_b_logical_ram_width = 16;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.clk0_output_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "old";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 7;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 127;
defparam ram_block1a15.port_a_logical_ram_depth = 128;
defparam ram_block1a15.port_a_logical_ram_width = 16;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 7;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "clock0";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 127;
defparam ram_block1a15.port_b_logical_ram_depth = 128;
defparam ram_block1a15.port_b_logical_ram_width = 16;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "old";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 7;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 127;
defparam ram_block1a7.port_a_logical_ram_depth = 128;
defparam ram_block1a7.port_a_logical_ram_width = 16;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 7;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "clock0";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 127;
defparam ram_block1a7.port_b_logical_ram_depth = 128;
defparam ram_block1a7.port_b_logical_ram_width = 16;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "old";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 7;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 127;
defparam ram_block1a3.port_a_logical_ram_depth = 128;
defparam ram_block1a3.port_a_logical_ram_width = 16;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 7;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "clock0";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 127;
defparam ram_block1a3.port_b_logical_ram_depth = 128;
defparam ram_block1a3.port_b_logical_ram_width = 16;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "old";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 7;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 127;
defparam ram_block1a5.port_a_logical_ram_depth = 128;
defparam ram_block1a5.port_a_logical_ram_width = 16;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 7;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "clock0";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 127;
defparam ram_block1a5.port_b_logical_ram_depth = 128;
defparam ram_block1a5.port_b_logical_ram_width = 16;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "old";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 7;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 127;
defparam ram_block1a4.port_a_logical_ram_depth = 128;
defparam ram_block1a4.port_a_logical_ram_width = 16;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 7;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "clock0";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 127;
defparam ram_block1a4.port_b_logical_ram_depth = 128;
defparam ram_block1a4.port_b_logical_ram_width = 16;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "old";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 7;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 127;
defparam ram_block1a6.port_a_logical_ram_depth = 128;
defparam ram_block1a6.port_a_logical_ram_width = 16;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 7;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "clock0";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 127;
defparam ram_block1a6.port_b_logical_ram_depth = 128;
defparam ram_block1a6.port_b_logical_ram_width = 16;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "old";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 7;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 127;
defparam ram_block1a2.port_a_logical_ram_depth = 128;
defparam ram_block1a2.port_a_logical_ram_width = 16;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 7;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "clock0";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 127;
defparam ram_block1a2.port_b_logical_ram_depth = 128;
defparam ram_block1a2.port_b_logical_ram_width = 16;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "old";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 7;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 127;
defparam ram_block1a1.port_a_logical_ram_depth = 128;
defparam ram_block1a1.port_a_logical_ram_width = 16;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 7;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "clock0";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 127;
defparam ram_block1a1.port_b_logical_ram_depth = 128;
defparam ram_block1a1.port_b_logical_ram_width = 16;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "old";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 7;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 127;
defparam ram_block1a0.port_a_logical_ram_depth = 128;
defparam ram_block1a0.port_a_logical_ram_width = 16;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 7;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "clock0";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 127;
defparam ram_block1a0.port_b_logical_ram_depth = 128;
defparam ram_block1a0.port_b_logical_ram_width = 16;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";

endmodule

module fft_asj_fft_data_ram_fft_120_10 (
	q_b_10,
	q_b_14,
	q_b_12,
	q_b_11,
	q_b_13,
	q_b_9,
	q_b_8,
	q_b_15,
	q_b_7,
	q_b_3,
	q_b_5,
	q_b_4,
	q_b_6,
	q_b_2,
	q_b_1,
	q_b_0,
	wren_a_2,
	global_clock_enable,
	wraddress_a_bus_21,
	wraddress_a_bus_23,
	wraddress_a_bus_11,
	wraddress_a_bus_13,
	rdaddress_a_bus_21,
	rdaddress_a_bus_23,
	rdaddress_a_bus_11,
	rdaddress_a_bus_13,
	a_ram_data_in_bus_26,
	wraddress_a_bus_8,
	wraddress_a_bus_10,
	wraddress_a_bus_12,
	rdaddress_a_bus_8,
	rdaddress_a_bus_10,
	rdaddress_a_bus_12,
	a_ram_data_in_bus_30,
	a_ram_data_in_bus_28,
	a_ram_data_in_bus_27,
	a_ram_data_in_bus_29,
	a_ram_data_in_bus_25,
	a_ram_data_in_bus_24,
	a_ram_data_in_bus_31,
	a_ram_data_in_bus_23,
	a_ram_data_in_bus_19,
	a_ram_data_in_bus_21,
	a_ram_data_in_bus_20,
	a_ram_data_in_bus_22,
	a_ram_data_in_bus_18,
	a_ram_data_in_bus_17,
	a_ram_data_in_bus_16,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_10;
output 	q_b_14;
output 	q_b_12;
output 	q_b_11;
output 	q_b_13;
output 	q_b_9;
output 	q_b_8;
output 	q_b_15;
output 	q_b_7;
output 	q_b_3;
output 	q_b_5;
output 	q_b_4;
output 	q_b_6;
output 	q_b_2;
output 	q_b_1;
output 	q_b_0;
input 	wren_a_2;
input 	global_clock_enable;
input 	wraddress_a_bus_21;
input 	wraddress_a_bus_23;
input 	wraddress_a_bus_11;
input 	wraddress_a_bus_13;
input 	rdaddress_a_bus_21;
input 	rdaddress_a_bus_23;
input 	rdaddress_a_bus_11;
input 	rdaddress_a_bus_13;
input 	a_ram_data_in_bus_26;
input 	wraddress_a_bus_8;
input 	wraddress_a_bus_10;
input 	wraddress_a_bus_12;
input 	rdaddress_a_bus_8;
input 	rdaddress_a_bus_10;
input 	rdaddress_a_bus_12;
input 	a_ram_data_in_bus_30;
input 	a_ram_data_in_bus_28;
input 	a_ram_data_in_bus_27;
input 	a_ram_data_in_bus_29;
input 	a_ram_data_in_bus_25;
input 	a_ram_data_in_bus_24;
input 	a_ram_data_in_bus_31;
input 	a_ram_data_in_bus_23;
input 	a_ram_data_in_bus_19;
input 	a_ram_data_in_bus_21;
input 	a_ram_data_in_bus_20;
input 	a_ram_data_in_bus_22;
input 	a_ram_data_in_bus_18;
input 	a_ram_data_in_bus_17;
input 	a_ram_data_in_bus_16;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_altsyncram_17 \gen_M4K:altsyncram_component (
	.q_b({q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.wren_a(wren_a_2),
	.clocken0(global_clock_enable),
	.address_a({wraddress_a_bus_13,wraddress_a_bus_12,wraddress_a_bus_11,wraddress_a_bus_10,wraddress_a_bus_23,wraddress_a_bus_8,wraddress_a_bus_21}),
	.address_b({rdaddress_a_bus_13,rdaddress_a_bus_12,rdaddress_a_bus_11,rdaddress_a_bus_10,rdaddress_a_bus_23,rdaddress_a_bus_8,rdaddress_a_bus_21}),
	.data_a({a_ram_data_in_bus_31,a_ram_data_in_bus_30,a_ram_data_in_bus_29,a_ram_data_in_bus_28,a_ram_data_in_bus_27,a_ram_data_in_bus_26,a_ram_data_in_bus_25,a_ram_data_in_bus_24,a_ram_data_in_bus_23,a_ram_data_in_bus_22,a_ram_data_in_bus_21,a_ram_data_in_bus_20,
a_ram_data_in_bus_19,a_ram_data_in_bus_18,a_ram_data_in_bus_17,a_ram_data_in_bus_16}),
	.clock0(clk));

endmodule

module fft_altsyncram_17 (
	q_b,
	wren_a,
	clocken0,
	address_a,
	address_b,
	data_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	wren_a;
input 	clocken0;
input 	[6:0] address_a;
input 	[6:0] address_b;
input 	[15:0] data_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_altsyncram_lmu3_10 auto_generated(
	.q_b({q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.wren_a(wren_a),
	.clocken0(clocken0),
	.address_a({address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.data_a({data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.clock0(clock0));

endmodule

module fft_altsyncram_lmu3_10 (
	q_b,
	wren_a,
	clocken0,
	address_a,
	address_b,
	data_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	wren_a;
input 	clocken0;
input 	[6:0] address_a;
input 	[6:0] address_b;
input 	[15:0] data_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

cycloneiii_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.clk0_output_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "old";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 7;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 127;
defparam ram_block1a10.port_a_logical_ram_depth = 128;
defparam ram_block1a10.port_a_logical_ram_width = 16;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 7;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "clock0";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 127;
defparam ram_block1a10.port_b_logical_ram_depth = 128;
defparam ram_block1a10.port_b_logical_ram_width = 16;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.clk0_output_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "old";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 7;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 127;
defparam ram_block1a14.port_a_logical_ram_depth = 128;
defparam ram_block1a14.port_a_logical_ram_width = 16;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 7;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "clock0";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 127;
defparam ram_block1a14.port_b_logical_ram_depth = 128;
defparam ram_block1a14.port_b_logical_ram_width = 16;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.clk0_output_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "old";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 7;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 127;
defparam ram_block1a12.port_a_logical_ram_depth = 128;
defparam ram_block1a12.port_a_logical_ram_width = 16;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 7;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "clock0";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 127;
defparam ram_block1a12.port_b_logical_ram_depth = 128;
defparam ram_block1a12.port_b_logical_ram_width = 16;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.clk0_output_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "old";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 7;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 127;
defparam ram_block1a11.port_a_logical_ram_depth = 128;
defparam ram_block1a11.port_a_logical_ram_width = 16;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 7;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "clock0";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 127;
defparam ram_block1a11.port_b_logical_ram_depth = 128;
defparam ram_block1a11.port_b_logical_ram_width = 16;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.clk0_output_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "old";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 7;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 127;
defparam ram_block1a13.port_a_logical_ram_depth = 128;
defparam ram_block1a13.port_a_logical_ram_width = 16;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 7;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "clock0";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 127;
defparam ram_block1a13.port_b_logical_ram_depth = 128;
defparam ram_block1a13.port_b_logical_ram_width = 16;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.clk0_output_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "old";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 7;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 127;
defparam ram_block1a9.port_a_logical_ram_depth = 128;
defparam ram_block1a9.port_a_logical_ram_width = 16;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 7;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "clock0";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 127;
defparam ram_block1a9.port_b_logical_ram_depth = 128;
defparam ram_block1a9.port_b_logical_ram_width = 16;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.clk0_output_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "old";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 7;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 127;
defparam ram_block1a8.port_a_logical_ram_depth = 128;
defparam ram_block1a8.port_a_logical_ram_width = 16;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 7;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "clock0";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 127;
defparam ram_block1a8.port_b_logical_ram_depth = 128;
defparam ram_block1a8.port_b_logical_ram_width = 16;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.clk0_output_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "old";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 7;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 127;
defparam ram_block1a15.port_a_logical_ram_depth = 128;
defparam ram_block1a15.port_a_logical_ram_width = 16;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 7;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "clock0";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 127;
defparam ram_block1a15.port_b_logical_ram_depth = 128;
defparam ram_block1a15.port_b_logical_ram_width = 16;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "old";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 7;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 127;
defparam ram_block1a7.port_a_logical_ram_depth = 128;
defparam ram_block1a7.port_a_logical_ram_width = 16;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 7;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "clock0";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 127;
defparam ram_block1a7.port_b_logical_ram_depth = 128;
defparam ram_block1a7.port_b_logical_ram_width = 16;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "old";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 7;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 127;
defparam ram_block1a3.port_a_logical_ram_depth = 128;
defparam ram_block1a3.port_a_logical_ram_width = 16;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 7;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "clock0";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 127;
defparam ram_block1a3.port_b_logical_ram_depth = 128;
defparam ram_block1a3.port_b_logical_ram_width = 16;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "old";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 7;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 127;
defparam ram_block1a5.port_a_logical_ram_depth = 128;
defparam ram_block1a5.port_a_logical_ram_width = 16;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 7;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "clock0";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 127;
defparam ram_block1a5.port_b_logical_ram_depth = 128;
defparam ram_block1a5.port_b_logical_ram_width = 16;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "old";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 7;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 127;
defparam ram_block1a4.port_a_logical_ram_depth = 128;
defparam ram_block1a4.port_a_logical_ram_width = 16;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 7;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "clock0";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 127;
defparam ram_block1a4.port_b_logical_ram_depth = 128;
defparam ram_block1a4.port_b_logical_ram_width = 16;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "old";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 7;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 127;
defparam ram_block1a6.port_a_logical_ram_depth = 128;
defparam ram_block1a6.port_a_logical_ram_width = 16;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 7;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "clock0";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 127;
defparam ram_block1a6.port_b_logical_ram_depth = 128;
defparam ram_block1a6.port_b_logical_ram_width = 16;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "old";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 7;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 127;
defparam ram_block1a2.port_a_logical_ram_depth = 128;
defparam ram_block1a2.port_a_logical_ram_width = 16;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 7;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "clock0";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 127;
defparam ram_block1a2.port_b_logical_ram_depth = 128;
defparam ram_block1a2.port_b_logical_ram_width = 16;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "old";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 7;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 127;
defparam ram_block1a1.port_a_logical_ram_depth = 128;
defparam ram_block1a1.port_a_logical_ram_width = 16;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 7;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "clock0";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 127;
defparam ram_block1a1.port_b_logical_ram_depth = 128;
defparam ram_block1a1.port_b_logical_ram_width = 16;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "old";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 7;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 127;
defparam ram_block1a0.port_a_logical_ram_depth = 128;
defparam ram_block1a0.port_a_logical_ram_width = 16;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 7;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "clock0";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 127;
defparam ram_block1a0.port_b_logical_ram_depth = 128;
defparam ram_block1a0.port_b_logical_ram_width = 16;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";

endmodule

module fft_asj_fft_data_ram_fft_120_11 (
	q_b_10,
	q_b_14,
	q_b_12,
	q_b_11,
	q_b_13,
	q_b_9,
	q_b_8,
	q_b_15,
	q_b_7,
	q_b_3,
	q_b_5,
	q_b_4,
	q_b_6,
	q_b_2,
	q_b_1,
	q_b_0,
	wren_a_3,
	global_clock_enable,
	wraddress_a_bus_13,
	rdaddress_a_bus_13,
	wraddress_a_bus_0,
	wraddress_a_bus_16,
	wraddress_a_bus_18,
	rdaddress_a_bus_0,
	rdaddress_a_bus_16,
	rdaddress_a_bus_18,
	a_ram_data_in_bus_10,
	wraddress_a_bus_1,
	wraddress_a_bus_3,
	wraddress_a_bus_5,
	rdaddress_a_bus_1,
	rdaddress_a_bus_3,
	rdaddress_a_bus_5,
	a_ram_data_in_bus_14,
	a_ram_data_in_bus_12,
	a_ram_data_in_bus_11,
	a_ram_data_in_bus_13,
	a_ram_data_in_bus_9,
	a_ram_data_in_bus_8,
	a_ram_data_in_bus_15,
	a_ram_data_in_bus_7,
	a_ram_data_in_bus_3,
	a_ram_data_in_bus_5,
	a_ram_data_in_bus_4,
	a_ram_data_in_bus_6,
	a_ram_data_in_bus_2,
	a_ram_data_in_bus_1,
	a_ram_data_in_bus_0,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_10;
output 	q_b_14;
output 	q_b_12;
output 	q_b_11;
output 	q_b_13;
output 	q_b_9;
output 	q_b_8;
output 	q_b_15;
output 	q_b_7;
output 	q_b_3;
output 	q_b_5;
output 	q_b_4;
output 	q_b_6;
output 	q_b_2;
output 	q_b_1;
output 	q_b_0;
input 	wren_a_3;
input 	global_clock_enable;
input 	wraddress_a_bus_13;
input 	rdaddress_a_bus_13;
input 	wraddress_a_bus_0;
input 	wraddress_a_bus_16;
input 	wraddress_a_bus_18;
input 	rdaddress_a_bus_0;
input 	rdaddress_a_bus_16;
input 	rdaddress_a_bus_18;
input 	a_ram_data_in_bus_10;
input 	wraddress_a_bus_1;
input 	wraddress_a_bus_3;
input 	wraddress_a_bus_5;
input 	rdaddress_a_bus_1;
input 	rdaddress_a_bus_3;
input 	rdaddress_a_bus_5;
input 	a_ram_data_in_bus_14;
input 	a_ram_data_in_bus_12;
input 	a_ram_data_in_bus_11;
input 	a_ram_data_in_bus_13;
input 	a_ram_data_in_bus_9;
input 	a_ram_data_in_bus_8;
input 	a_ram_data_in_bus_15;
input 	a_ram_data_in_bus_7;
input 	a_ram_data_in_bus_3;
input 	a_ram_data_in_bus_5;
input 	a_ram_data_in_bus_4;
input 	a_ram_data_in_bus_6;
input 	a_ram_data_in_bus_2;
input 	a_ram_data_in_bus_1;
input 	a_ram_data_in_bus_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_altsyncram_18 \gen_M4K:altsyncram_component (
	.q_b({q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.wren_a(wren_a_3),
	.clocken0(global_clock_enable),
	.address_a({wraddress_a_bus_13,wraddress_a_bus_5,wraddress_a_bus_18,wraddress_a_bus_3,wraddress_a_bus_16,wraddress_a_bus_1,wraddress_a_bus_0}),
	.address_b({rdaddress_a_bus_13,rdaddress_a_bus_5,rdaddress_a_bus_18,rdaddress_a_bus_3,rdaddress_a_bus_16,rdaddress_a_bus_1,rdaddress_a_bus_0}),
	.data_a({a_ram_data_in_bus_15,a_ram_data_in_bus_14,a_ram_data_in_bus_13,a_ram_data_in_bus_12,a_ram_data_in_bus_11,a_ram_data_in_bus_10,a_ram_data_in_bus_9,a_ram_data_in_bus_8,a_ram_data_in_bus_7,a_ram_data_in_bus_6,a_ram_data_in_bus_5,a_ram_data_in_bus_4,a_ram_data_in_bus_3,
a_ram_data_in_bus_2,a_ram_data_in_bus_1,a_ram_data_in_bus_0}),
	.clock0(clk));

endmodule

module fft_altsyncram_18 (
	q_b,
	wren_a,
	clocken0,
	address_a,
	address_b,
	data_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	wren_a;
input 	clocken0;
input 	[6:0] address_a;
input 	[6:0] address_b;
input 	[15:0] data_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_altsyncram_lmu3_11 auto_generated(
	.q_b({q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.wren_a(wren_a),
	.clocken0(clocken0),
	.address_a({address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.data_a({data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.clock0(clock0));

endmodule

module fft_altsyncram_lmu3_11 (
	q_b,
	wren_a,
	clocken0,
	address_a,
	address_b,
	data_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	wren_a;
input 	clocken0;
input 	[6:0] address_a;
input 	[6:0] address_b;
input 	[15:0] data_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

cycloneiii_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.clk0_output_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "old";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 7;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 127;
defparam ram_block1a10.port_a_logical_ram_depth = 128;
defparam ram_block1a10.port_a_logical_ram_width = 16;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 7;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "clock0";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 127;
defparam ram_block1a10.port_b_logical_ram_depth = 128;
defparam ram_block1a10.port_b_logical_ram_width = 16;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.clk0_output_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "old";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 7;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 127;
defparam ram_block1a14.port_a_logical_ram_depth = 128;
defparam ram_block1a14.port_a_logical_ram_width = 16;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 7;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "clock0";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 127;
defparam ram_block1a14.port_b_logical_ram_depth = 128;
defparam ram_block1a14.port_b_logical_ram_width = 16;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.clk0_output_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "old";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 7;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 127;
defparam ram_block1a12.port_a_logical_ram_depth = 128;
defparam ram_block1a12.port_a_logical_ram_width = 16;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 7;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "clock0";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 127;
defparam ram_block1a12.port_b_logical_ram_depth = 128;
defparam ram_block1a12.port_b_logical_ram_width = 16;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.clk0_output_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "old";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 7;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 127;
defparam ram_block1a11.port_a_logical_ram_depth = 128;
defparam ram_block1a11.port_a_logical_ram_width = 16;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 7;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "clock0";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 127;
defparam ram_block1a11.port_b_logical_ram_depth = 128;
defparam ram_block1a11.port_b_logical_ram_width = 16;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.clk0_output_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "old";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 7;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 127;
defparam ram_block1a13.port_a_logical_ram_depth = 128;
defparam ram_block1a13.port_a_logical_ram_width = 16;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 7;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "clock0";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 127;
defparam ram_block1a13.port_b_logical_ram_depth = 128;
defparam ram_block1a13.port_b_logical_ram_width = 16;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.clk0_output_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "old";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 7;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 127;
defparam ram_block1a9.port_a_logical_ram_depth = 128;
defparam ram_block1a9.port_a_logical_ram_width = 16;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 7;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "clock0";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 127;
defparam ram_block1a9.port_b_logical_ram_depth = 128;
defparam ram_block1a9.port_b_logical_ram_width = 16;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.clk0_output_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "old";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 7;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 127;
defparam ram_block1a8.port_a_logical_ram_depth = 128;
defparam ram_block1a8.port_a_logical_ram_width = 16;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 7;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "clock0";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 127;
defparam ram_block1a8.port_b_logical_ram_depth = 128;
defparam ram_block1a8.port_b_logical_ram_width = 16;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.clk0_output_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "old";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 7;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 127;
defparam ram_block1a15.port_a_logical_ram_depth = 128;
defparam ram_block1a15.port_a_logical_ram_width = 16;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 7;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "clock0";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 127;
defparam ram_block1a15.port_b_logical_ram_depth = 128;
defparam ram_block1a15.port_b_logical_ram_width = 16;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "old";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 7;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 127;
defparam ram_block1a7.port_a_logical_ram_depth = 128;
defparam ram_block1a7.port_a_logical_ram_width = 16;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 7;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "clock0";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 127;
defparam ram_block1a7.port_b_logical_ram_depth = 128;
defparam ram_block1a7.port_b_logical_ram_width = 16;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "old";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 7;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 127;
defparam ram_block1a3.port_a_logical_ram_depth = 128;
defparam ram_block1a3.port_a_logical_ram_width = 16;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 7;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "clock0";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 127;
defparam ram_block1a3.port_b_logical_ram_depth = 128;
defparam ram_block1a3.port_b_logical_ram_width = 16;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "old";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 7;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 127;
defparam ram_block1a5.port_a_logical_ram_depth = 128;
defparam ram_block1a5.port_a_logical_ram_width = 16;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 7;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "clock0";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 127;
defparam ram_block1a5.port_b_logical_ram_depth = 128;
defparam ram_block1a5.port_b_logical_ram_width = 16;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "old";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 7;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 127;
defparam ram_block1a4.port_a_logical_ram_depth = 128;
defparam ram_block1a4.port_a_logical_ram_width = 16;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 7;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "clock0";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 127;
defparam ram_block1a4.port_b_logical_ram_depth = 128;
defparam ram_block1a4.port_b_logical_ram_width = 16;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "old";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 7;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 127;
defparam ram_block1a6.port_a_logical_ram_depth = 128;
defparam ram_block1a6.port_a_logical_ram_width = 16;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 7;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "clock0";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 127;
defparam ram_block1a6.port_b_logical_ram_depth = 128;
defparam ram_block1a6.port_b_logical_ram_width = 16;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "old";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 7;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 127;
defparam ram_block1a2.port_a_logical_ram_depth = 128;
defparam ram_block1a2.port_a_logical_ram_width = 16;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 7;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "clock0";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 127;
defparam ram_block1a2.port_b_logical_ram_depth = 128;
defparam ram_block1a2.port_b_logical_ram_width = 16;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "old";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 7;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 127;
defparam ram_block1a1.port_a_logical_ram_depth = 128;
defparam ram_block1a1.port_a_logical_ram_width = 16;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 7;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "clock0";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 127;
defparam ram_block1a1.port_b_logical_ram_depth = 128;
defparam ram_block1a1.port_b_logical_ram_width = 16;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_A|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "old";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 7;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 127;
defparam ram_block1a0.port_a_logical_ram_depth = 128;
defparam ram_block1a0.port_a_logical_ram_width = 16;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 7;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "clock0";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 127;
defparam ram_block1a0.port_b_logical_ram_depth = 128;
defparam ram_block1a0.port_b_logical_ram_width = 16;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";

endmodule

module fft_asj_fft_4dp_ram_fft_120_3 (
	q_b_10,
	q_b_101,
	q_b_102,
	q_b_103,
	q_b_14,
	q_b_141,
	q_b_142,
	q_b_143,
	q_b_12,
	q_b_121,
	q_b_122,
	q_b_123,
	q_b_11,
	q_b_111,
	q_b_112,
	q_b_113,
	q_b_13,
	q_b_131,
	q_b_132,
	q_b_133,
	q_b_9,
	q_b_91,
	q_b_92,
	q_b_93,
	q_b_8,
	q_b_81,
	q_b_82,
	q_b_83,
	q_b_15,
	q_b_151,
	q_b_152,
	q_b_153,
	q_b_7,
	q_b_71,
	q_b_72,
	q_b_73,
	q_b_3,
	q_b_31,
	q_b_32,
	q_b_33,
	q_b_5,
	q_b_51,
	q_b_52,
	q_b_53,
	q_b_4,
	q_b_41,
	q_b_42,
	q_b_43,
	q_b_6,
	q_b_61,
	q_b_62,
	q_b_63,
	q_b_2,
	q_b_21,
	q_b_22,
	q_b_23,
	q_b_1,
	q_b_16,
	q_b_17,
	q_b_18,
	q_b_0,
	q_b_01,
	q_b_02,
	q_b_03,
	wren_b_0,
	wren_b_1,
	wren_b_2,
	wren_b_3,
	global_clock_enable,
	b_ram_data_in_bus_58,
	wraddress_b_bus_21,
	wraddress_b_bus_22,
	wraddress_b_bus_23,
	wraddress_b_bus_24,
	wraddress_b_bus_11,
	wraddress_b_bus_26,
	wraddress_b_bus_13,
	rdaddress_b_bus_21,
	rdaddress_b_bus_22,
	rdaddress_b_bus_23,
	rdaddress_b_bus_24,
	rdaddress_b_bus_11,
	rdaddress_b_bus_26,
	rdaddress_b_bus_13,
	b_ram_data_in_bus_42,
	wraddress_b_bus_0,
	wraddress_b_bus_15,
	wraddress_b_bus_16,
	wraddress_b_bus_17,
	wraddress_b_bus_18,
	wraddress_b_bus_19,
	rdaddress_b_bus_0,
	rdaddress_b_bus_15,
	rdaddress_b_bus_16,
	rdaddress_b_bus_17,
	rdaddress_b_bus_18,
	rdaddress_b_bus_19,
	b_ram_data_in_bus_26,
	wraddress_b_bus_8,
	wraddress_b_bus_10,
	wraddress_b_bus_12,
	rdaddress_b_bus_8,
	rdaddress_b_bus_10,
	rdaddress_b_bus_12,
	b_ram_data_in_bus_10,
	wraddress_b_bus_1,
	wraddress_b_bus_3,
	wraddress_b_bus_5,
	rdaddress_b_bus_1,
	rdaddress_b_bus_3,
	rdaddress_b_bus_5,
	b_ram_data_in_bus_62,
	b_ram_data_in_bus_46,
	b_ram_data_in_bus_30,
	b_ram_data_in_bus_14,
	b_ram_data_in_bus_60,
	b_ram_data_in_bus_44,
	b_ram_data_in_bus_28,
	b_ram_data_in_bus_12,
	b_ram_data_in_bus_59,
	b_ram_data_in_bus_43,
	b_ram_data_in_bus_27,
	b_ram_data_in_bus_11,
	b_ram_data_in_bus_61,
	b_ram_data_in_bus_45,
	b_ram_data_in_bus_29,
	b_ram_data_in_bus_13,
	b_ram_data_in_bus_57,
	b_ram_data_in_bus_41,
	b_ram_data_in_bus_25,
	b_ram_data_in_bus_9,
	b_ram_data_in_bus_56,
	b_ram_data_in_bus_40,
	b_ram_data_in_bus_24,
	b_ram_data_in_bus_8,
	b_ram_data_in_bus_63,
	b_ram_data_in_bus_47,
	b_ram_data_in_bus_31,
	b_ram_data_in_bus_15,
	b_ram_data_in_bus_55,
	b_ram_data_in_bus_39,
	b_ram_data_in_bus_23,
	b_ram_data_in_bus_7,
	b_ram_data_in_bus_51,
	b_ram_data_in_bus_35,
	b_ram_data_in_bus_19,
	b_ram_data_in_bus_3,
	b_ram_data_in_bus_53,
	b_ram_data_in_bus_37,
	b_ram_data_in_bus_21,
	b_ram_data_in_bus_5,
	b_ram_data_in_bus_52,
	b_ram_data_in_bus_36,
	b_ram_data_in_bus_20,
	b_ram_data_in_bus_4,
	b_ram_data_in_bus_54,
	b_ram_data_in_bus_38,
	b_ram_data_in_bus_22,
	b_ram_data_in_bus_6,
	b_ram_data_in_bus_50,
	b_ram_data_in_bus_34,
	b_ram_data_in_bus_18,
	b_ram_data_in_bus_2,
	b_ram_data_in_bus_49,
	b_ram_data_in_bus_33,
	b_ram_data_in_bus_17,
	b_ram_data_in_bus_1,
	b_ram_data_in_bus_48,
	b_ram_data_in_bus_32,
	b_ram_data_in_bus_16,
	b_ram_data_in_bus_0,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_10;
output 	q_b_101;
output 	q_b_102;
output 	q_b_103;
output 	q_b_14;
output 	q_b_141;
output 	q_b_142;
output 	q_b_143;
output 	q_b_12;
output 	q_b_121;
output 	q_b_122;
output 	q_b_123;
output 	q_b_11;
output 	q_b_111;
output 	q_b_112;
output 	q_b_113;
output 	q_b_13;
output 	q_b_131;
output 	q_b_132;
output 	q_b_133;
output 	q_b_9;
output 	q_b_91;
output 	q_b_92;
output 	q_b_93;
output 	q_b_8;
output 	q_b_81;
output 	q_b_82;
output 	q_b_83;
output 	q_b_15;
output 	q_b_151;
output 	q_b_152;
output 	q_b_153;
output 	q_b_7;
output 	q_b_71;
output 	q_b_72;
output 	q_b_73;
output 	q_b_3;
output 	q_b_31;
output 	q_b_32;
output 	q_b_33;
output 	q_b_5;
output 	q_b_51;
output 	q_b_52;
output 	q_b_53;
output 	q_b_4;
output 	q_b_41;
output 	q_b_42;
output 	q_b_43;
output 	q_b_6;
output 	q_b_61;
output 	q_b_62;
output 	q_b_63;
output 	q_b_2;
output 	q_b_21;
output 	q_b_22;
output 	q_b_23;
output 	q_b_1;
output 	q_b_16;
output 	q_b_17;
output 	q_b_18;
output 	q_b_0;
output 	q_b_01;
output 	q_b_02;
output 	q_b_03;
input 	wren_b_0;
input 	wren_b_1;
input 	wren_b_2;
input 	wren_b_3;
input 	global_clock_enable;
input 	b_ram_data_in_bus_58;
input 	wraddress_b_bus_21;
input 	wraddress_b_bus_22;
input 	wraddress_b_bus_23;
input 	wraddress_b_bus_24;
input 	wraddress_b_bus_11;
input 	wraddress_b_bus_26;
input 	wraddress_b_bus_13;
input 	rdaddress_b_bus_21;
input 	rdaddress_b_bus_22;
input 	rdaddress_b_bus_23;
input 	rdaddress_b_bus_24;
input 	rdaddress_b_bus_11;
input 	rdaddress_b_bus_26;
input 	rdaddress_b_bus_13;
input 	b_ram_data_in_bus_42;
input 	wraddress_b_bus_0;
input 	wraddress_b_bus_15;
input 	wraddress_b_bus_16;
input 	wraddress_b_bus_17;
input 	wraddress_b_bus_18;
input 	wraddress_b_bus_19;
input 	rdaddress_b_bus_0;
input 	rdaddress_b_bus_15;
input 	rdaddress_b_bus_16;
input 	rdaddress_b_bus_17;
input 	rdaddress_b_bus_18;
input 	rdaddress_b_bus_19;
input 	b_ram_data_in_bus_26;
input 	wraddress_b_bus_8;
input 	wraddress_b_bus_10;
input 	wraddress_b_bus_12;
input 	rdaddress_b_bus_8;
input 	rdaddress_b_bus_10;
input 	rdaddress_b_bus_12;
input 	b_ram_data_in_bus_10;
input 	wraddress_b_bus_1;
input 	wraddress_b_bus_3;
input 	wraddress_b_bus_5;
input 	rdaddress_b_bus_1;
input 	rdaddress_b_bus_3;
input 	rdaddress_b_bus_5;
input 	b_ram_data_in_bus_62;
input 	b_ram_data_in_bus_46;
input 	b_ram_data_in_bus_30;
input 	b_ram_data_in_bus_14;
input 	b_ram_data_in_bus_60;
input 	b_ram_data_in_bus_44;
input 	b_ram_data_in_bus_28;
input 	b_ram_data_in_bus_12;
input 	b_ram_data_in_bus_59;
input 	b_ram_data_in_bus_43;
input 	b_ram_data_in_bus_27;
input 	b_ram_data_in_bus_11;
input 	b_ram_data_in_bus_61;
input 	b_ram_data_in_bus_45;
input 	b_ram_data_in_bus_29;
input 	b_ram_data_in_bus_13;
input 	b_ram_data_in_bus_57;
input 	b_ram_data_in_bus_41;
input 	b_ram_data_in_bus_25;
input 	b_ram_data_in_bus_9;
input 	b_ram_data_in_bus_56;
input 	b_ram_data_in_bus_40;
input 	b_ram_data_in_bus_24;
input 	b_ram_data_in_bus_8;
input 	b_ram_data_in_bus_63;
input 	b_ram_data_in_bus_47;
input 	b_ram_data_in_bus_31;
input 	b_ram_data_in_bus_15;
input 	b_ram_data_in_bus_55;
input 	b_ram_data_in_bus_39;
input 	b_ram_data_in_bus_23;
input 	b_ram_data_in_bus_7;
input 	b_ram_data_in_bus_51;
input 	b_ram_data_in_bus_35;
input 	b_ram_data_in_bus_19;
input 	b_ram_data_in_bus_3;
input 	b_ram_data_in_bus_53;
input 	b_ram_data_in_bus_37;
input 	b_ram_data_in_bus_21;
input 	b_ram_data_in_bus_5;
input 	b_ram_data_in_bus_52;
input 	b_ram_data_in_bus_36;
input 	b_ram_data_in_bus_20;
input 	b_ram_data_in_bus_4;
input 	b_ram_data_in_bus_54;
input 	b_ram_data_in_bus_38;
input 	b_ram_data_in_bus_22;
input 	b_ram_data_in_bus_6;
input 	b_ram_data_in_bus_50;
input 	b_ram_data_in_bus_34;
input 	b_ram_data_in_bus_18;
input 	b_ram_data_in_bus_2;
input 	b_ram_data_in_bus_49;
input 	b_ram_data_in_bus_33;
input 	b_ram_data_in_bus_17;
input 	b_ram_data_in_bus_1;
input 	b_ram_data_in_bus_48;
input 	b_ram_data_in_bus_32;
input 	b_ram_data_in_bus_16;
input 	b_ram_data_in_bus_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_asj_fft_data_ram_fft_120_15 \gen_rams:3:dat_A (
	.q_b_10(q_b_103),
	.q_b_14(q_b_143),
	.q_b_12(q_b_123),
	.q_b_11(q_b_113),
	.q_b_13(q_b_133),
	.q_b_9(q_b_93),
	.q_b_8(q_b_83),
	.q_b_15(q_b_153),
	.q_b_7(q_b_73),
	.q_b_3(q_b_33),
	.q_b_5(q_b_53),
	.q_b_4(q_b_43),
	.q_b_6(q_b_63),
	.q_b_2(q_b_23),
	.q_b_1(q_b_18),
	.q_b_0(q_b_03),
	.wren_b_3(wren_b_3),
	.global_clock_enable(global_clock_enable),
	.wraddress_b_bus_13(wraddress_b_bus_13),
	.rdaddress_b_bus_13(rdaddress_b_bus_13),
	.wraddress_b_bus_0(wraddress_b_bus_0),
	.wraddress_b_bus_16(wraddress_b_bus_16),
	.wraddress_b_bus_18(wraddress_b_bus_18),
	.rdaddress_b_bus_0(rdaddress_b_bus_0),
	.rdaddress_b_bus_16(rdaddress_b_bus_16),
	.rdaddress_b_bus_18(rdaddress_b_bus_18),
	.b_ram_data_in_bus_10(b_ram_data_in_bus_10),
	.wraddress_b_bus_1(wraddress_b_bus_1),
	.wraddress_b_bus_3(wraddress_b_bus_3),
	.wraddress_b_bus_5(wraddress_b_bus_5),
	.rdaddress_b_bus_1(rdaddress_b_bus_1),
	.rdaddress_b_bus_3(rdaddress_b_bus_3),
	.rdaddress_b_bus_5(rdaddress_b_bus_5),
	.b_ram_data_in_bus_14(b_ram_data_in_bus_14),
	.b_ram_data_in_bus_12(b_ram_data_in_bus_12),
	.b_ram_data_in_bus_11(b_ram_data_in_bus_11),
	.b_ram_data_in_bus_13(b_ram_data_in_bus_13),
	.b_ram_data_in_bus_9(b_ram_data_in_bus_9),
	.b_ram_data_in_bus_8(b_ram_data_in_bus_8),
	.b_ram_data_in_bus_15(b_ram_data_in_bus_15),
	.b_ram_data_in_bus_7(b_ram_data_in_bus_7),
	.b_ram_data_in_bus_3(b_ram_data_in_bus_3),
	.b_ram_data_in_bus_5(b_ram_data_in_bus_5),
	.b_ram_data_in_bus_4(b_ram_data_in_bus_4),
	.b_ram_data_in_bus_6(b_ram_data_in_bus_6),
	.b_ram_data_in_bus_2(b_ram_data_in_bus_2),
	.b_ram_data_in_bus_1(b_ram_data_in_bus_1),
	.b_ram_data_in_bus_0(b_ram_data_in_bus_0),
	.clk(clk));

fft_asj_fft_data_ram_fft_120_14 \gen_rams:2:dat_A (
	.q_b_10(q_b_102),
	.q_b_14(q_b_142),
	.q_b_12(q_b_122),
	.q_b_11(q_b_112),
	.q_b_13(q_b_132),
	.q_b_9(q_b_92),
	.q_b_8(q_b_82),
	.q_b_15(q_b_152),
	.q_b_7(q_b_72),
	.q_b_3(q_b_32),
	.q_b_5(q_b_52),
	.q_b_4(q_b_42),
	.q_b_6(q_b_62),
	.q_b_2(q_b_22),
	.q_b_1(q_b_17),
	.q_b_0(q_b_02),
	.wren_b_2(wren_b_2),
	.global_clock_enable(global_clock_enable),
	.wraddress_b_bus_21(wraddress_b_bus_21),
	.wraddress_b_bus_23(wraddress_b_bus_23),
	.wraddress_b_bus_11(wraddress_b_bus_11),
	.wraddress_b_bus_13(wraddress_b_bus_13),
	.rdaddress_b_bus_21(rdaddress_b_bus_21),
	.rdaddress_b_bus_23(rdaddress_b_bus_23),
	.rdaddress_b_bus_11(rdaddress_b_bus_11),
	.rdaddress_b_bus_13(rdaddress_b_bus_13),
	.b_ram_data_in_bus_26(b_ram_data_in_bus_26),
	.wraddress_b_bus_8(wraddress_b_bus_8),
	.wraddress_b_bus_10(wraddress_b_bus_10),
	.wraddress_b_bus_12(wraddress_b_bus_12),
	.rdaddress_b_bus_8(rdaddress_b_bus_8),
	.rdaddress_b_bus_10(rdaddress_b_bus_10),
	.rdaddress_b_bus_12(rdaddress_b_bus_12),
	.b_ram_data_in_bus_30(b_ram_data_in_bus_30),
	.b_ram_data_in_bus_28(b_ram_data_in_bus_28),
	.b_ram_data_in_bus_27(b_ram_data_in_bus_27),
	.b_ram_data_in_bus_29(b_ram_data_in_bus_29),
	.b_ram_data_in_bus_25(b_ram_data_in_bus_25),
	.b_ram_data_in_bus_24(b_ram_data_in_bus_24),
	.b_ram_data_in_bus_31(b_ram_data_in_bus_31),
	.b_ram_data_in_bus_23(b_ram_data_in_bus_23),
	.b_ram_data_in_bus_19(b_ram_data_in_bus_19),
	.b_ram_data_in_bus_21(b_ram_data_in_bus_21),
	.b_ram_data_in_bus_20(b_ram_data_in_bus_20),
	.b_ram_data_in_bus_22(b_ram_data_in_bus_22),
	.b_ram_data_in_bus_18(b_ram_data_in_bus_18),
	.b_ram_data_in_bus_17(b_ram_data_in_bus_17),
	.b_ram_data_in_bus_16(b_ram_data_in_bus_16),
	.clk(clk));

fft_asj_fft_data_ram_fft_120_13 \gen_rams:1:dat_A (
	.q_b_10(q_b_101),
	.q_b_14(q_b_141),
	.q_b_12(q_b_121),
	.q_b_11(q_b_111),
	.q_b_13(q_b_131),
	.q_b_9(q_b_91),
	.q_b_8(q_b_81),
	.q_b_15(q_b_151),
	.q_b_7(q_b_71),
	.q_b_3(q_b_31),
	.q_b_5(q_b_51),
	.q_b_4(q_b_41),
	.q_b_6(q_b_61),
	.q_b_2(q_b_21),
	.q_b_1(q_b_16),
	.q_b_0(q_b_01),
	.wren_b_1(wren_b_1),
	.global_clock_enable(global_clock_enable),
	.wraddress_b_bus_13(wraddress_b_bus_13),
	.rdaddress_b_bus_13(rdaddress_b_bus_13),
	.b_ram_data_in_bus_42(b_ram_data_in_bus_42),
	.wraddress_b_bus_0(wraddress_b_bus_0),
	.wraddress_b_bus_15(wraddress_b_bus_15),
	.wraddress_b_bus_16(wraddress_b_bus_16),
	.wraddress_b_bus_17(wraddress_b_bus_17),
	.wraddress_b_bus_18(wraddress_b_bus_18),
	.wraddress_b_bus_19(wraddress_b_bus_19),
	.rdaddress_b_bus_0(rdaddress_b_bus_0),
	.rdaddress_b_bus_15(rdaddress_b_bus_15),
	.rdaddress_b_bus_16(rdaddress_b_bus_16),
	.rdaddress_b_bus_17(rdaddress_b_bus_17),
	.rdaddress_b_bus_18(rdaddress_b_bus_18),
	.rdaddress_b_bus_19(rdaddress_b_bus_19),
	.b_ram_data_in_bus_46(b_ram_data_in_bus_46),
	.b_ram_data_in_bus_44(b_ram_data_in_bus_44),
	.b_ram_data_in_bus_43(b_ram_data_in_bus_43),
	.b_ram_data_in_bus_45(b_ram_data_in_bus_45),
	.b_ram_data_in_bus_41(b_ram_data_in_bus_41),
	.b_ram_data_in_bus_40(b_ram_data_in_bus_40),
	.b_ram_data_in_bus_47(b_ram_data_in_bus_47),
	.b_ram_data_in_bus_39(b_ram_data_in_bus_39),
	.b_ram_data_in_bus_35(b_ram_data_in_bus_35),
	.b_ram_data_in_bus_37(b_ram_data_in_bus_37),
	.b_ram_data_in_bus_36(b_ram_data_in_bus_36),
	.b_ram_data_in_bus_38(b_ram_data_in_bus_38),
	.b_ram_data_in_bus_34(b_ram_data_in_bus_34),
	.b_ram_data_in_bus_33(b_ram_data_in_bus_33),
	.b_ram_data_in_bus_32(b_ram_data_in_bus_32),
	.clk(clk));

fft_asj_fft_data_ram_fft_120_12 \gen_rams:0:dat_A (
	.q_b_10(q_b_10),
	.q_b_14(q_b_14),
	.q_b_12(q_b_12),
	.q_b_11(q_b_11),
	.q_b_13(q_b_13),
	.q_b_9(q_b_9),
	.q_b_8(q_b_8),
	.q_b_15(q_b_15),
	.q_b_7(q_b_7),
	.q_b_3(q_b_3),
	.q_b_5(q_b_5),
	.q_b_4(q_b_4),
	.q_b_6(q_b_6),
	.q_b_2(q_b_2),
	.q_b_1(q_b_1),
	.q_b_0(q_b_0),
	.wren_b_0(wren_b_0),
	.global_clock_enable(global_clock_enable),
	.b_ram_data_in_bus_58(b_ram_data_in_bus_58),
	.wraddress_b_bus_21(wraddress_b_bus_21),
	.wraddress_b_bus_22(wraddress_b_bus_22),
	.wraddress_b_bus_23(wraddress_b_bus_23),
	.wraddress_b_bus_24(wraddress_b_bus_24),
	.wraddress_b_bus_11(wraddress_b_bus_11),
	.wraddress_b_bus_26(wraddress_b_bus_26),
	.wraddress_b_bus_13(wraddress_b_bus_13),
	.rdaddress_b_bus_21(rdaddress_b_bus_21),
	.rdaddress_b_bus_22(rdaddress_b_bus_22),
	.rdaddress_b_bus_23(rdaddress_b_bus_23),
	.rdaddress_b_bus_24(rdaddress_b_bus_24),
	.rdaddress_b_bus_11(rdaddress_b_bus_11),
	.rdaddress_b_bus_26(rdaddress_b_bus_26),
	.rdaddress_b_bus_13(rdaddress_b_bus_13),
	.b_ram_data_in_bus_62(b_ram_data_in_bus_62),
	.b_ram_data_in_bus_60(b_ram_data_in_bus_60),
	.b_ram_data_in_bus_59(b_ram_data_in_bus_59),
	.b_ram_data_in_bus_61(b_ram_data_in_bus_61),
	.b_ram_data_in_bus_57(b_ram_data_in_bus_57),
	.b_ram_data_in_bus_56(b_ram_data_in_bus_56),
	.b_ram_data_in_bus_63(b_ram_data_in_bus_63),
	.b_ram_data_in_bus_55(b_ram_data_in_bus_55),
	.b_ram_data_in_bus_51(b_ram_data_in_bus_51),
	.b_ram_data_in_bus_53(b_ram_data_in_bus_53),
	.b_ram_data_in_bus_52(b_ram_data_in_bus_52),
	.b_ram_data_in_bus_54(b_ram_data_in_bus_54),
	.b_ram_data_in_bus_50(b_ram_data_in_bus_50),
	.b_ram_data_in_bus_49(b_ram_data_in_bus_49),
	.b_ram_data_in_bus_48(b_ram_data_in_bus_48),
	.clk(clk));

endmodule

module fft_asj_fft_data_ram_fft_120_12 (
	q_b_10,
	q_b_14,
	q_b_12,
	q_b_11,
	q_b_13,
	q_b_9,
	q_b_8,
	q_b_15,
	q_b_7,
	q_b_3,
	q_b_5,
	q_b_4,
	q_b_6,
	q_b_2,
	q_b_1,
	q_b_0,
	wren_b_0,
	global_clock_enable,
	b_ram_data_in_bus_58,
	wraddress_b_bus_21,
	wraddress_b_bus_22,
	wraddress_b_bus_23,
	wraddress_b_bus_24,
	wraddress_b_bus_11,
	wraddress_b_bus_26,
	wraddress_b_bus_13,
	rdaddress_b_bus_21,
	rdaddress_b_bus_22,
	rdaddress_b_bus_23,
	rdaddress_b_bus_24,
	rdaddress_b_bus_11,
	rdaddress_b_bus_26,
	rdaddress_b_bus_13,
	b_ram_data_in_bus_62,
	b_ram_data_in_bus_60,
	b_ram_data_in_bus_59,
	b_ram_data_in_bus_61,
	b_ram_data_in_bus_57,
	b_ram_data_in_bus_56,
	b_ram_data_in_bus_63,
	b_ram_data_in_bus_55,
	b_ram_data_in_bus_51,
	b_ram_data_in_bus_53,
	b_ram_data_in_bus_52,
	b_ram_data_in_bus_54,
	b_ram_data_in_bus_50,
	b_ram_data_in_bus_49,
	b_ram_data_in_bus_48,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_10;
output 	q_b_14;
output 	q_b_12;
output 	q_b_11;
output 	q_b_13;
output 	q_b_9;
output 	q_b_8;
output 	q_b_15;
output 	q_b_7;
output 	q_b_3;
output 	q_b_5;
output 	q_b_4;
output 	q_b_6;
output 	q_b_2;
output 	q_b_1;
output 	q_b_0;
input 	wren_b_0;
input 	global_clock_enable;
input 	b_ram_data_in_bus_58;
input 	wraddress_b_bus_21;
input 	wraddress_b_bus_22;
input 	wraddress_b_bus_23;
input 	wraddress_b_bus_24;
input 	wraddress_b_bus_11;
input 	wraddress_b_bus_26;
input 	wraddress_b_bus_13;
input 	rdaddress_b_bus_21;
input 	rdaddress_b_bus_22;
input 	rdaddress_b_bus_23;
input 	rdaddress_b_bus_24;
input 	rdaddress_b_bus_11;
input 	rdaddress_b_bus_26;
input 	rdaddress_b_bus_13;
input 	b_ram_data_in_bus_62;
input 	b_ram_data_in_bus_60;
input 	b_ram_data_in_bus_59;
input 	b_ram_data_in_bus_61;
input 	b_ram_data_in_bus_57;
input 	b_ram_data_in_bus_56;
input 	b_ram_data_in_bus_63;
input 	b_ram_data_in_bus_55;
input 	b_ram_data_in_bus_51;
input 	b_ram_data_in_bus_53;
input 	b_ram_data_in_bus_52;
input 	b_ram_data_in_bus_54;
input 	b_ram_data_in_bus_50;
input 	b_ram_data_in_bus_49;
input 	b_ram_data_in_bus_48;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_altsyncram_19 \gen_M4K:altsyncram_component (
	.q_b({q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.wren_a(wren_b_0),
	.clocken0(global_clock_enable),
	.data_a({b_ram_data_in_bus_63,b_ram_data_in_bus_62,b_ram_data_in_bus_61,b_ram_data_in_bus_60,b_ram_data_in_bus_59,b_ram_data_in_bus_58,b_ram_data_in_bus_57,b_ram_data_in_bus_56,b_ram_data_in_bus_55,b_ram_data_in_bus_54,b_ram_data_in_bus_53,b_ram_data_in_bus_52,
b_ram_data_in_bus_51,b_ram_data_in_bus_50,b_ram_data_in_bus_49,b_ram_data_in_bus_48}),
	.address_a({wraddress_b_bus_13,wraddress_b_bus_26,wraddress_b_bus_11,wraddress_b_bus_24,wraddress_b_bus_23,wraddress_b_bus_22,wraddress_b_bus_21}),
	.address_b({rdaddress_b_bus_13,rdaddress_b_bus_26,rdaddress_b_bus_11,rdaddress_b_bus_24,rdaddress_b_bus_23,rdaddress_b_bus_22,rdaddress_b_bus_21}),
	.clock0(clk));

endmodule

module fft_altsyncram_19 (
	q_b,
	wren_a,
	clocken0,
	data_a,
	address_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	wren_a;
input 	clocken0;
input 	[15:0] data_a;
input 	[6:0] address_a;
input 	[6:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_altsyncram_lmu3_12 auto_generated(
	.q_b({q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.wren_a(wren_a),
	.clocken0(clocken0),
	.data_a({data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_a({address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.clock0(clock0));

endmodule

module fft_altsyncram_lmu3_12 (
	q_b,
	wren_a,
	clocken0,
	data_a,
	address_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	wren_a;
input 	clocken0;
input 	[15:0] data_a;
input 	[6:0] address_a;
input 	[6:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

cycloneiii_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.clk0_output_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "old";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 7;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 127;
defparam ram_block1a10.port_a_logical_ram_depth = 128;
defparam ram_block1a10.port_a_logical_ram_width = 16;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 7;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "clock0";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 127;
defparam ram_block1a10.port_b_logical_ram_depth = 128;
defparam ram_block1a10.port_b_logical_ram_width = 16;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.clk0_output_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "old";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 7;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 127;
defparam ram_block1a14.port_a_logical_ram_depth = 128;
defparam ram_block1a14.port_a_logical_ram_width = 16;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 7;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "clock0";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 127;
defparam ram_block1a14.port_b_logical_ram_depth = 128;
defparam ram_block1a14.port_b_logical_ram_width = 16;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.clk0_output_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "old";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 7;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 127;
defparam ram_block1a12.port_a_logical_ram_depth = 128;
defparam ram_block1a12.port_a_logical_ram_width = 16;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 7;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "clock0";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 127;
defparam ram_block1a12.port_b_logical_ram_depth = 128;
defparam ram_block1a12.port_b_logical_ram_width = 16;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.clk0_output_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "old";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 7;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 127;
defparam ram_block1a11.port_a_logical_ram_depth = 128;
defparam ram_block1a11.port_a_logical_ram_width = 16;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 7;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "clock0";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 127;
defparam ram_block1a11.port_b_logical_ram_depth = 128;
defparam ram_block1a11.port_b_logical_ram_width = 16;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.clk0_output_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "old";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 7;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 127;
defparam ram_block1a13.port_a_logical_ram_depth = 128;
defparam ram_block1a13.port_a_logical_ram_width = 16;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 7;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "clock0";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 127;
defparam ram_block1a13.port_b_logical_ram_depth = 128;
defparam ram_block1a13.port_b_logical_ram_width = 16;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.clk0_output_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "old";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 7;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 127;
defparam ram_block1a9.port_a_logical_ram_depth = 128;
defparam ram_block1a9.port_a_logical_ram_width = 16;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 7;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "clock0";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 127;
defparam ram_block1a9.port_b_logical_ram_depth = 128;
defparam ram_block1a9.port_b_logical_ram_width = 16;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.clk0_output_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "old";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 7;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 127;
defparam ram_block1a8.port_a_logical_ram_depth = 128;
defparam ram_block1a8.port_a_logical_ram_width = 16;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 7;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "clock0";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 127;
defparam ram_block1a8.port_b_logical_ram_depth = 128;
defparam ram_block1a8.port_b_logical_ram_width = 16;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.clk0_output_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "old";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 7;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 127;
defparam ram_block1a15.port_a_logical_ram_depth = 128;
defparam ram_block1a15.port_a_logical_ram_width = 16;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 7;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "clock0";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 127;
defparam ram_block1a15.port_b_logical_ram_depth = 128;
defparam ram_block1a15.port_b_logical_ram_width = 16;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "old";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 7;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 127;
defparam ram_block1a7.port_a_logical_ram_depth = 128;
defparam ram_block1a7.port_a_logical_ram_width = 16;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 7;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "clock0";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 127;
defparam ram_block1a7.port_b_logical_ram_depth = 128;
defparam ram_block1a7.port_b_logical_ram_width = 16;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "old";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 7;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 127;
defparam ram_block1a3.port_a_logical_ram_depth = 128;
defparam ram_block1a3.port_a_logical_ram_width = 16;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 7;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "clock0";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 127;
defparam ram_block1a3.port_b_logical_ram_depth = 128;
defparam ram_block1a3.port_b_logical_ram_width = 16;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "old";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 7;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 127;
defparam ram_block1a5.port_a_logical_ram_depth = 128;
defparam ram_block1a5.port_a_logical_ram_width = 16;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 7;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "clock0";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 127;
defparam ram_block1a5.port_b_logical_ram_depth = 128;
defparam ram_block1a5.port_b_logical_ram_width = 16;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "old";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 7;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 127;
defparam ram_block1a4.port_a_logical_ram_depth = 128;
defparam ram_block1a4.port_a_logical_ram_width = 16;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 7;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "clock0";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 127;
defparam ram_block1a4.port_b_logical_ram_depth = 128;
defparam ram_block1a4.port_b_logical_ram_width = 16;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "old";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 7;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 127;
defparam ram_block1a6.port_a_logical_ram_depth = 128;
defparam ram_block1a6.port_a_logical_ram_width = 16;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 7;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "clock0";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 127;
defparam ram_block1a6.port_b_logical_ram_depth = 128;
defparam ram_block1a6.port_b_logical_ram_width = 16;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "old";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 7;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 127;
defparam ram_block1a2.port_a_logical_ram_depth = 128;
defparam ram_block1a2.port_a_logical_ram_width = 16;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 7;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "clock0";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 127;
defparam ram_block1a2.port_b_logical_ram_depth = 128;
defparam ram_block1a2.port_b_logical_ram_width = 16;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "old";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 7;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 127;
defparam ram_block1a1.port_a_logical_ram_depth = 128;
defparam ram_block1a1.port_a_logical_ram_width = 16;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 7;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "clock0";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 127;
defparam ram_block1a1.port_b_logical_ram_depth = 128;
defparam ram_block1a1.port_b_logical_ram_width = 16;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:0:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "old";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 7;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 127;
defparam ram_block1a0.port_a_logical_ram_depth = 128;
defparam ram_block1a0.port_a_logical_ram_width = 16;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 7;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "clock0";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 127;
defparam ram_block1a0.port_b_logical_ram_depth = 128;
defparam ram_block1a0.port_b_logical_ram_width = 16;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";

endmodule

module fft_asj_fft_data_ram_fft_120_13 (
	q_b_10,
	q_b_14,
	q_b_12,
	q_b_11,
	q_b_13,
	q_b_9,
	q_b_8,
	q_b_15,
	q_b_7,
	q_b_3,
	q_b_5,
	q_b_4,
	q_b_6,
	q_b_2,
	q_b_1,
	q_b_0,
	wren_b_1,
	global_clock_enable,
	wraddress_b_bus_13,
	rdaddress_b_bus_13,
	b_ram_data_in_bus_42,
	wraddress_b_bus_0,
	wraddress_b_bus_15,
	wraddress_b_bus_16,
	wraddress_b_bus_17,
	wraddress_b_bus_18,
	wraddress_b_bus_19,
	rdaddress_b_bus_0,
	rdaddress_b_bus_15,
	rdaddress_b_bus_16,
	rdaddress_b_bus_17,
	rdaddress_b_bus_18,
	rdaddress_b_bus_19,
	b_ram_data_in_bus_46,
	b_ram_data_in_bus_44,
	b_ram_data_in_bus_43,
	b_ram_data_in_bus_45,
	b_ram_data_in_bus_41,
	b_ram_data_in_bus_40,
	b_ram_data_in_bus_47,
	b_ram_data_in_bus_39,
	b_ram_data_in_bus_35,
	b_ram_data_in_bus_37,
	b_ram_data_in_bus_36,
	b_ram_data_in_bus_38,
	b_ram_data_in_bus_34,
	b_ram_data_in_bus_33,
	b_ram_data_in_bus_32,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_10;
output 	q_b_14;
output 	q_b_12;
output 	q_b_11;
output 	q_b_13;
output 	q_b_9;
output 	q_b_8;
output 	q_b_15;
output 	q_b_7;
output 	q_b_3;
output 	q_b_5;
output 	q_b_4;
output 	q_b_6;
output 	q_b_2;
output 	q_b_1;
output 	q_b_0;
input 	wren_b_1;
input 	global_clock_enable;
input 	wraddress_b_bus_13;
input 	rdaddress_b_bus_13;
input 	b_ram_data_in_bus_42;
input 	wraddress_b_bus_0;
input 	wraddress_b_bus_15;
input 	wraddress_b_bus_16;
input 	wraddress_b_bus_17;
input 	wraddress_b_bus_18;
input 	wraddress_b_bus_19;
input 	rdaddress_b_bus_0;
input 	rdaddress_b_bus_15;
input 	rdaddress_b_bus_16;
input 	rdaddress_b_bus_17;
input 	rdaddress_b_bus_18;
input 	rdaddress_b_bus_19;
input 	b_ram_data_in_bus_46;
input 	b_ram_data_in_bus_44;
input 	b_ram_data_in_bus_43;
input 	b_ram_data_in_bus_45;
input 	b_ram_data_in_bus_41;
input 	b_ram_data_in_bus_40;
input 	b_ram_data_in_bus_47;
input 	b_ram_data_in_bus_39;
input 	b_ram_data_in_bus_35;
input 	b_ram_data_in_bus_37;
input 	b_ram_data_in_bus_36;
input 	b_ram_data_in_bus_38;
input 	b_ram_data_in_bus_34;
input 	b_ram_data_in_bus_33;
input 	b_ram_data_in_bus_32;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_altsyncram_20 \gen_M4K:altsyncram_component (
	.q_b({q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.wren_a(wren_b_1),
	.clocken0(global_clock_enable),
	.address_a({wraddress_b_bus_13,wraddress_b_bus_19,wraddress_b_bus_18,wraddress_b_bus_17,wraddress_b_bus_16,wraddress_b_bus_15,wraddress_b_bus_0}),
	.address_b({rdaddress_b_bus_13,rdaddress_b_bus_19,rdaddress_b_bus_18,rdaddress_b_bus_17,rdaddress_b_bus_16,rdaddress_b_bus_15,rdaddress_b_bus_0}),
	.data_a({b_ram_data_in_bus_47,b_ram_data_in_bus_46,b_ram_data_in_bus_45,b_ram_data_in_bus_44,b_ram_data_in_bus_43,b_ram_data_in_bus_42,b_ram_data_in_bus_41,b_ram_data_in_bus_40,b_ram_data_in_bus_39,b_ram_data_in_bus_38,b_ram_data_in_bus_37,b_ram_data_in_bus_36,
b_ram_data_in_bus_35,b_ram_data_in_bus_34,b_ram_data_in_bus_33,b_ram_data_in_bus_32}),
	.clock0(clk));

endmodule

module fft_altsyncram_20 (
	q_b,
	wren_a,
	clocken0,
	address_a,
	address_b,
	data_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	wren_a;
input 	clocken0;
input 	[6:0] address_a;
input 	[6:0] address_b;
input 	[15:0] data_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_altsyncram_lmu3_13 auto_generated(
	.q_b({q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.wren_a(wren_a),
	.clocken0(clocken0),
	.address_a({address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.data_a({data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.clock0(clock0));

endmodule

module fft_altsyncram_lmu3_13 (
	q_b,
	wren_a,
	clocken0,
	address_a,
	address_b,
	data_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	wren_a;
input 	clocken0;
input 	[6:0] address_a;
input 	[6:0] address_b;
input 	[15:0] data_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

cycloneiii_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.clk0_output_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "old";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 7;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 127;
defparam ram_block1a10.port_a_logical_ram_depth = 128;
defparam ram_block1a10.port_a_logical_ram_width = 16;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 7;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "clock0";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 127;
defparam ram_block1a10.port_b_logical_ram_depth = 128;
defparam ram_block1a10.port_b_logical_ram_width = 16;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.clk0_output_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "old";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 7;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 127;
defparam ram_block1a14.port_a_logical_ram_depth = 128;
defparam ram_block1a14.port_a_logical_ram_width = 16;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 7;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "clock0";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 127;
defparam ram_block1a14.port_b_logical_ram_depth = 128;
defparam ram_block1a14.port_b_logical_ram_width = 16;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.clk0_output_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "old";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 7;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 127;
defparam ram_block1a12.port_a_logical_ram_depth = 128;
defparam ram_block1a12.port_a_logical_ram_width = 16;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 7;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "clock0";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 127;
defparam ram_block1a12.port_b_logical_ram_depth = 128;
defparam ram_block1a12.port_b_logical_ram_width = 16;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.clk0_output_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "old";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 7;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 127;
defparam ram_block1a11.port_a_logical_ram_depth = 128;
defparam ram_block1a11.port_a_logical_ram_width = 16;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 7;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "clock0";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 127;
defparam ram_block1a11.port_b_logical_ram_depth = 128;
defparam ram_block1a11.port_b_logical_ram_width = 16;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.clk0_output_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "old";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 7;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 127;
defparam ram_block1a13.port_a_logical_ram_depth = 128;
defparam ram_block1a13.port_a_logical_ram_width = 16;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 7;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "clock0";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 127;
defparam ram_block1a13.port_b_logical_ram_depth = 128;
defparam ram_block1a13.port_b_logical_ram_width = 16;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.clk0_output_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "old";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 7;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 127;
defparam ram_block1a9.port_a_logical_ram_depth = 128;
defparam ram_block1a9.port_a_logical_ram_width = 16;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 7;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "clock0";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 127;
defparam ram_block1a9.port_b_logical_ram_depth = 128;
defparam ram_block1a9.port_b_logical_ram_width = 16;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.clk0_output_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "old";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 7;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 127;
defparam ram_block1a8.port_a_logical_ram_depth = 128;
defparam ram_block1a8.port_a_logical_ram_width = 16;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 7;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "clock0";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 127;
defparam ram_block1a8.port_b_logical_ram_depth = 128;
defparam ram_block1a8.port_b_logical_ram_width = 16;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.clk0_output_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "old";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 7;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 127;
defparam ram_block1a15.port_a_logical_ram_depth = 128;
defparam ram_block1a15.port_a_logical_ram_width = 16;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 7;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "clock0";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 127;
defparam ram_block1a15.port_b_logical_ram_depth = 128;
defparam ram_block1a15.port_b_logical_ram_width = 16;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "old";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 7;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 127;
defparam ram_block1a7.port_a_logical_ram_depth = 128;
defparam ram_block1a7.port_a_logical_ram_width = 16;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 7;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "clock0";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 127;
defparam ram_block1a7.port_b_logical_ram_depth = 128;
defparam ram_block1a7.port_b_logical_ram_width = 16;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "old";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 7;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 127;
defparam ram_block1a3.port_a_logical_ram_depth = 128;
defparam ram_block1a3.port_a_logical_ram_width = 16;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 7;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "clock0";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 127;
defparam ram_block1a3.port_b_logical_ram_depth = 128;
defparam ram_block1a3.port_b_logical_ram_width = 16;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "old";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 7;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 127;
defparam ram_block1a5.port_a_logical_ram_depth = 128;
defparam ram_block1a5.port_a_logical_ram_width = 16;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 7;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "clock0";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 127;
defparam ram_block1a5.port_b_logical_ram_depth = 128;
defparam ram_block1a5.port_b_logical_ram_width = 16;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "old";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 7;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 127;
defparam ram_block1a4.port_a_logical_ram_depth = 128;
defparam ram_block1a4.port_a_logical_ram_width = 16;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 7;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "clock0";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 127;
defparam ram_block1a4.port_b_logical_ram_depth = 128;
defparam ram_block1a4.port_b_logical_ram_width = 16;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "old";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 7;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 127;
defparam ram_block1a6.port_a_logical_ram_depth = 128;
defparam ram_block1a6.port_a_logical_ram_width = 16;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 7;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "clock0";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 127;
defparam ram_block1a6.port_b_logical_ram_depth = 128;
defparam ram_block1a6.port_b_logical_ram_width = 16;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "old";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 7;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 127;
defparam ram_block1a2.port_a_logical_ram_depth = 128;
defparam ram_block1a2.port_a_logical_ram_width = 16;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 7;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "clock0";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 127;
defparam ram_block1a2.port_b_logical_ram_depth = 128;
defparam ram_block1a2.port_b_logical_ram_width = 16;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "old";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 7;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 127;
defparam ram_block1a1.port_a_logical_ram_depth = 128;
defparam ram_block1a1.port_a_logical_ram_width = 16;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 7;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "clock0";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 127;
defparam ram_block1a1.port_b_logical_ram_depth = 128;
defparam ram_block1a1.port_b_logical_ram_width = 16;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:1:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "old";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 7;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 127;
defparam ram_block1a0.port_a_logical_ram_depth = 128;
defparam ram_block1a0.port_a_logical_ram_width = 16;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 7;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "clock0";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 127;
defparam ram_block1a0.port_b_logical_ram_depth = 128;
defparam ram_block1a0.port_b_logical_ram_width = 16;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";

endmodule

module fft_asj_fft_data_ram_fft_120_14 (
	q_b_10,
	q_b_14,
	q_b_12,
	q_b_11,
	q_b_13,
	q_b_9,
	q_b_8,
	q_b_15,
	q_b_7,
	q_b_3,
	q_b_5,
	q_b_4,
	q_b_6,
	q_b_2,
	q_b_1,
	q_b_0,
	wren_b_2,
	global_clock_enable,
	wraddress_b_bus_21,
	wraddress_b_bus_23,
	wraddress_b_bus_11,
	wraddress_b_bus_13,
	rdaddress_b_bus_21,
	rdaddress_b_bus_23,
	rdaddress_b_bus_11,
	rdaddress_b_bus_13,
	b_ram_data_in_bus_26,
	wraddress_b_bus_8,
	wraddress_b_bus_10,
	wraddress_b_bus_12,
	rdaddress_b_bus_8,
	rdaddress_b_bus_10,
	rdaddress_b_bus_12,
	b_ram_data_in_bus_30,
	b_ram_data_in_bus_28,
	b_ram_data_in_bus_27,
	b_ram_data_in_bus_29,
	b_ram_data_in_bus_25,
	b_ram_data_in_bus_24,
	b_ram_data_in_bus_31,
	b_ram_data_in_bus_23,
	b_ram_data_in_bus_19,
	b_ram_data_in_bus_21,
	b_ram_data_in_bus_20,
	b_ram_data_in_bus_22,
	b_ram_data_in_bus_18,
	b_ram_data_in_bus_17,
	b_ram_data_in_bus_16,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_10;
output 	q_b_14;
output 	q_b_12;
output 	q_b_11;
output 	q_b_13;
output 	q_b_9;
output 	q_b_8;
output 	q_b_15;
output 	q_b_7;
output 	q_b_3;
output 	q_b_5;
output 	q_b_4;
output 	q_b_6;
output 	q_b_2;
output 	q_b_1;
output 	q_b_0;
input 	wren_b_2;
input 	global_clock_enable;
input 	wraddress_b_bus_21;
input 	wraddress_b_bus_23;
input 	wraddress_b_bus_11;
input 	wraddress_b_bus_13;
input 	rdaddress_b_bus_21;
input 	rdaddress_b_bus_23;
input 	rdaddress_b_bus_11;
input 	rdaddress_b_bus_13;
input 	b_ram_data_in_bus_26;
input 	wraddress_b_bus_8;
input 	wraddress_b_bus_10;
input 	wraddress_b_bus_12;
input 	rdaddress_b_bus_8;
input 	rdaddress_b_bus_10;
input 	rdaddress_b_bus_12;
input 	b_ram_data_in_bus_30;
input 	b_ram_data_in_bus_28;
input 	b_ram_data_in_bus_27;
input 	b_ram_data_in_bus_29;
input 	b_ram_data_in_bus_25;
input 	b_ram_data_in_bus_24;
input 	b_ram_data_in_bus_31;
input 	b_ram_data_in_bus_23;
input 	b_ram_data_in_bus_19;
input 	b_ram_data_in_bus_21;
input 	b_ram_data_in_bus_20;
input 	b_ram_data_in_bus_22;
input 	b_ram_data_in_bus_18;
input 	b_ram_data_in_bus_17;
input 	b_ram_data_in_bus_16;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_altsyncram_21 \gen_M4K:altsyncram_component (
	.q_b({q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.wren_a(wren_b_2),
	.clocken0(global_clock_enable),
	.address_a({wraddress_b_bus_13,wraddress_b_bus_12,wraddress_b_bus_11,wraddress_b_bus_10,wraddress_b_bus_23,wraddress_b_bus_8,wraddress_b_bus_21}),
	.address_b({rdaddress_b_bus_13,rdaddress_b_bus_12,rdaddress_b_bus_11,rdaddress_b_bus_10,rdaddress_b_bus_23,rdaddress_b_bus_8,rdaddress_b_bus_21}),
	.data_a({b_ram_data_in_bus_31,b_ram_data_in_bus_30,b_ram_data_in_bus_29,b_ram_data_in_bus_28,b_ram_data_in_bus_27,b_ram_data_in_bus_26,b_ram_data_in_bus_25,b_ram_data_in_bus_24,b_ram_data_in_bus_23,b_ram_data_in_bus_22,b_ram_data_in_bus_21,b_ram_data_in_bus_20,
b_ram_data_in_bus_19,b_ram_data_in_bus_18,b_ram_data_in_bus_17,b_ram_data_in_bus_16}),
	.clock0(clk));

endmodule

module fft_altsyncram_21 (
	q_b,
	wren_a,
	clocken0,
	address_a,
	address_b,
	data_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	wren_a;
input 	clocken0;
input 	[6:0] address_a;
input 	[6:0] address_b;
input 	[15:0] data_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_altsyncram_lmu3_14 auto_generated(
	.q_b({q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.wren_a(wren_a),
	.clocken0(clocken0),
	.address_a({address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.data_a({data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.clock0(clock0));

endmodule

module fft_altsyncram_lmu3_14 (
	q_b,
	wren_a,
	clocken0,
	address_a,
	address_b,
	data_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	wren_a;
input 	clocken0;
input 	[6:0] address_a;
input 	[6:0] address_b;
input 	[15:0] data_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

cycloneiii_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.clk0_output_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "old";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 7;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 127;
defparam ram_block1a10.port_a_logical_ram_depth = 128;
defparam ram_block1a10.port_a_logical_ram_width = 16;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 7;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "clock0";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 127;
defparam ram_block1a10.port_b_logical_ram_depth = 128;
defparam ram_block1a10.port_b_logical_ram_width = 16;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.clk0_output_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "old";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 7;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 127;
defparam ram_block1a14.port_a_logical_ram_depth = 128;
defparam ram_block1a14.port_a_logical_ram_width = 16;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 7;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "clock0";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 127;
defparam ram_block1a14.port_b_logical_ram_depth = 128;
defparam ram_block1a14.port_b_logical_ram_width = 16;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.clk0_output_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "old";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 7;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 127;
defparam ram_block1a12.port_a_logical_ram_depth = 128;
defparam ram_block1a12.port_a_logical_ram_width = 16;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 7;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "clock0";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 127;
defparam ram_block1a12.port_b_logical_ram_depth = 128;
defparam ram_block1a12.port_b_logical_ram_width = 16;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.clk0_output_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "old";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 7;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 127;
defparam ram_block1a11.port_a_logical_ram_depth = 128;
defparam ram_block1a11.port_a_logical_ram_width = 16;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 7;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "clock0";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 127;
defparam ram_block1a11.port_b_logical_ram_depth = 128;
defparam ram_block1a11.port_b_logical_ram_width = 16;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.clk0_output_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "old";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 7;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 127;
defparam ram_block1a13.port_a_logical_ram_depth = 128;
defparam ram_block1a13.port_a_logical_ram_width = 16;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 7;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "clock0";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 127;
defparam ram_block1a13.port_b_logical_ram_depth = 128;
defparam ram_block1a13.port_b_logical_ram_width = 16;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.clk0_output_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "old";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 7;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 127;
defparam ram_block1a9.port_a_logical_ram_depth = 128;
defparam ram_block1a9.port_a_logical_ram_width = 16;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 7;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "clock0";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 127;
defparam ram_block1a9.port_b_logical_ram_depth = 128;
defparam ram_block1a9.port_b_logical_ram_width = 16;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.clk0_output_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "old";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 7;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 127;
defparam ram_block1a8.port_a_logical_ram_depth = 128;
defparam ram_block1a8.port_a_logical_ram_width = 16;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 7;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "clock0";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 127;
defparam ram_block1a8.port_b_logical_ram_depth = 128;
defparam ram_block1a8.port_b_logical_ram_width = 16;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.clk0_output_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "old";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 7;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 127;
defparam ram_block1a15.port_a_logical_ram_depth = 128;
defparam ram_block1a15.port_a_logical_ram_width = 16;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 7;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "clock0";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 127;
defparam ram_block1a15.port_b_logical_ram_depth = 128;
defparam ram_block1a15.port_b_logical_ram_width = 16;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "old";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 7;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 127;
defparam ram_block1a7.port_a_logical_ram_depth = 128;
defparam ram_block1a7.port_a_logical_ram_width = 16;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 7;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "clock0";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 127;
defparam ram_block1a7.port_b_logical_ram_depth = 128;
defparam ram_block1a7.port_b_logical_ram_width = 16;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "old";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 7;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 127;
defparam ram_block1a3.port_a_logical_ram_depth = 128;
defparam ram_block1a3.port_a_logical_ram_width = 16;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 7;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "clock0";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 127;
defparam ram_block1a3.port_b_logical_ram_depth = 128;
defparam ram_block1a3.port_b_logical_ram_width = 16;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "old";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 7;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 127;
defparam ram_block1a5.port_a_logical_ram_depth = 128;
defparam ram_block1a5.port_a_logical_ram_width = 16;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 7;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "clock0";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 127;
defparam ram_block1a5.port_b_logical_ram_depth = 128;
defparam ram_block1a5.port_b_logical_ram_width = 16;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "old";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 7;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 127;
defparam ram_block1a4.port_a_logical_ram_depth = 128;
defparam ram_block1a4.port_a_logical_ram_width = 16;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 7;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "clock0";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 127;
defparam ram_block1a4.port_b_logical_ram_depth = 128;
defparam ram_block1a4.port_b_logical_ram_width = 16;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "old";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 7;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 127;
defparam ram_block1a6.port_a_logical_ram_depth = 128;
defparam ram_block1a6.port_a_logical_ram_width = 16;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 7;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "clock0";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 127;
defparam ram_block1a6.port_b_logical_ram_depth = 128;
defparam ram_block1a6.port_b_logical_ram_width = 16;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "old";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 7;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 127;
defparam ram_block1a2.port_a_logical_ram_depth = 128;
defparam ram_block1a2.port_a_logical_ram_width = 16;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 7;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "clock0";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 127;
defparam ram_block1a2.port_b_logical_ram_depth = 128;
defparam ram_block1a2.port_b_logical_ram_width = 16;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "old";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 7;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 127;
defparam ram_block1a1.port_a_logical_ram_depth = 128;
defparam ram_block1a1.port_a_logical_ram_width = 16;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 7;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "clock0";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 127;
defparam ram_block1a1.port_b_logical_ram_depth = 128;
defparam ram_block1a1.port_b_logical_ram_width = 16;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:2:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "old";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 7;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 127;
defparam ram_block1a0.port_a_logical_ram_depth = 128;
defparam ram_block1a0.port_a_logical_ram_width = 16;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 7;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "clock0";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 127;
defparam ram_block1a0.port_b_logical_ram_depth = 128;
defparam ram_block1a0.port_b_logical_ram_width = 16;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";

endmodule

module fft_asj_fft_data_ram_fft_120_15 (
	q_b_10,
	q_b_14,
	q_b_12,
	q_b_11,
	q_b_13,
	q_b_9,
	q_b_8,
	q_b_15,
	q_b_7,
	q_b_3,
	q_b_5,
	q_b_4,
	q_b_6,
	q_b_2,
	q_b_1,
	q_b_0,
	wren_b_3,
	global_clock_enable,
	wraddress_b_bus_13,
	rdaddress_b_bus_13,
	wraddress_b_bus_0,
	wraddress_b_bus_16,
	wraddress_b_bus_18,
	rdaddress_b_bus_0,
	rdaddress_b_bus_16,
	rdaddress_b_bus_18,
	b_ram_data_in_bus_10,
	wraddress_b_bus_1,
	wraddress_b_bus_3,
	wraddress_b_bus_5,
	rdaddress_b_bus_1,
	rdaddress_b_bus_3,
	rdaddress_b_bus_5,
	b_ram_data_in_bus_14,
	b_ram_data_in_bus_12,
	b_ram_data_in_bus_11,
	b_ram_data_in_bus_13,
	b_ram_data_in_bus_9,
	b_ram_data_in_bus_8,
	b_ram_data_in_bus_15,
	b_ram_data_in_bus_7,
	b_ram_data_in_bus_3,
	b_ram_data_in_bus_5,
	b_ram_data_in_bus_4,
	b_ram_data_in_bus_6,
	b_ram_data_in_bus_2,
	b_ram_data_in_bus_1,
	b_ram_data_in_bus_0,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_10;
output 	q_b_14;
output 	q_b_12;
output 	q_b_11;
output 	q_b_13;
output 	q_b_9;
output 	q_b_8;
output 	q_b_15;
output 	q_b_7;
output 	q_b_3;
output 	q_b_5;
output 	q_b_4;
output 	q_b_6;
output 	q_b_2;
output 	q_b_1;
output 	q_b_0;
input 	wren_b_3;
input 	global_clock_enable;
input 	wraddress_b_bus_13;
input 	rdaddress_b_bus_13;
input 	wraddress_b_bus_0;
input 	wraddress_b_bus_16;
input 	wraddress_b_bus_18;
input 	rdaddress_b_bus_0;
input 	rdaddress_b_bus_16;
input 	rdaddress_b_bus_18;
input 	b_ram_data_in_bus_10;
input 	wraddress_b_bus_1;
input 	wraddress_b_bus_3;
input 	wraddress_b_bus_5;
input 	rdaddress_b_bus_1;
input 	rdaddress_b_bus_3;
input 	rdaddress_b_bus_5;
input 	b_ram_data_in_bus_14;
input 	b_ram_data_in_bus_12;
input 	b_ram_data_in_bus_11;
input 	b_ram_data_in_bus_13;
input 	b_ram_data_in_bus_9;
input 	b_ram_data_in_bus_8;
input 	b_ram_data_in_bus_15;
input 	b_ram_data_in_bus_7;
input 	b_ram_data_in_bus_3;
input 	b_ram_data_in_bus_5;
input 	b_ram_data_in_bus_4;
input 	b_ram_data_in_bus_6;
input 	b_ram_data_in_bus_2;
input 	b_ram_data_in_bus_1;
input 	b_ram_data_in_bus_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_altsyncram_22 \gen_M4K:altsyncram_component (
	.q_b({q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.wren_a(wren_b_3),
	.clocken0(global_clock_enable),
	.address_a({wraddress_b_bus_13,wraddress_b_bus_5,wraddress_b_bus_18,wraddress_b_bus_3,wraddress_b_bus_16,wraddress_b_bus_1,wraddress_b_bus_0}),
	.address_b({rdaddress_b_bus_13,rdaddress_b_bus_5,rdaddress_b_bus_18,rdaddress_b_bus_3,rdaddress_b_bus_16,rdaddress_b_bus_1,rdaddress_b_bus_0}),
	.data_a({b_ram_data_in_bus_15,b_ram_data_in_bus_14,b_ram_data_in_bus_13,b_ram_data_in_bus_12,b_ram_data_in_bus_11,b_ram_data_in_bus_10,b_ram_data_in_bus_9,b_ram_data_in_bus_8,b_ram_data_in_bus_7,b_ram_data_in_bus_6,b_ram_data_in_bus_5,b_ram_data_in_bus_4,b_ram_data_in_bus_3,
b_ram_data_in_bus_2,b_ram_data_in_bus_1,b_ram_data_in_bus_0}),
	.clock0(clk));

endmodule

module fft_altsyncram_22 (
	q_b,
	wren_a,
	clocken0,
	address_a,
	address_b,
	data_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	wren_a;
input 	clocken0;
input 	[6:0] address_a;
input 	[6:0] address_b;
input 	[15:0] data_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_altsyncram_lmu3_15 auto_generated(
	.q_b({q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.wren_a(wren_a),
	.clocken0(clocken0),
	.address_a({address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.data_a({data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.clock0(clock0));

endmodule

module fft_altsyncram_lmu3_15 (
	q_b,
	wren_a,
	clocken0,
	address_a,
	address_b,
	data_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	wren_a;
input 	clocken0;
input 	[6:0] address_a;
input 	[6:0] address_b;
input 	[15:0] data_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

cycloneiii_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.clk0_output_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "old";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 7;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 127;
defparam ram_block1a10.port_a_logical_ram_depth = 128;
defparam ram_block1a10.port_a_logical_ram_width = 16;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 7;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "clock0";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 127;
defparam ram_block1a10.port_b_logical_ram_depth = 128;
defparam ram_block1a10.port_b_logical_ram_width = 16;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.clk0_output_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "old";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 7;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 127;
defparam ram_block1a14.port_a_logical_ram_depth = 128;
defparam ram_block1a14.port_a_logical_ram_width = 16;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 7;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "clock0";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 127;
defparam ram_block1a14.port_b_logical_ram_depth = 128;
defparam ram_block1a14.port_b_logical_ram_width = 16;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.clk0_output_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "old";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 7;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 127;
defparam ram_block1a12.port_a_logical_ram_depth = 128;
defparam ram_block1a12.port_a_logical_ram_width = 16;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 7;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "clock0";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 127;
defparam ram_block1a12.port_b_logical_ram_depth = 128;
defparam ram_block1a12.port_b_logical_ram_width = 16;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.clk0_output_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "old";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 7;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 127;
defparam ram_block1a11.port_a_logical_ram_depth = 128;
defparam ram_block1a11.port_a_logical_ram_width = 16;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 7;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "clock0";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 127;
defparam ram_block1a11.port_b_logical_ram_depth = 128;
defparam ram_block1a11.port_b_logical_ram_width = 16;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.clk0_output_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "old";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 7;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 127;
defparam ram_block1a13.port_a_logical_ram_depth = 128;
defparam ram_block1a13.port_a_logical_ram_width = 16;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 7;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "clock0";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 127;
defparam ram_block1a13.port_b_logical_ram_depth = 128;
defparam ram_block1a13.port_b_logical_ram_width = 16;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.clk0_output_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "old";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 7;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 127;
defparam ram_block1a9.port_a_logical_ram_depth = 128;
defparam ram_block1a9.port_a_logical_ram_width = 16;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 7;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "clock0";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 127;
defparam ram_block1a9.port_b_logical_ram_depth = 128;
defparam ram_block1a9.port_b_logical_ram_width = 16;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.clk0_output_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "old";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 7;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 127;
defparam ram_block1a8.port_a_logical_ram_depth = 128;
defparam ram_block1a8.port_a_logical_ram_width = 16;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 7;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "clock0";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 127;
defparam ram_block1a8.port_b_logical_ram_depth = 128;
defparam ram_block1a8.port_b_logical_ram_width = 16;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.clk0_output_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "old";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 7;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 127;
defparam ram_block1a15.port_a_logical_ram_depth = 128;
defparam ram_block1a15.port_a_logical_ram_width = 16;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 7;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "clock0";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 127;
defparam ram_block1a15.port_b_logical_ram_depth = 128;
defparam ram_block1a15.port_b_logical_ram_width = 16;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "old";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 7;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 127;
defparam ram_block1a7.port_a_logical_ram_depth = 128;
defparam ram_block1a7.port_a_logical_ram_width = 16;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 7;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "clock0";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 127;
defparam ram_block1a7.port_b_logical_ram_depth = 128;
defparam ram_block1a7.port_b_logical_ram_width = 16;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "old";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 7;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 127;
defparam ram_block1a3.port_a_logical_ram_depth = 128;
defparam ram_block1a3.port_a_logical_ram_width = 16;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 7;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "clock0";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 127;
defparam ram_block1a3.port_b_logical_ram_depth = 128;
defparam ram_block1a3.port_b_logical_ram_width = 16;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "old";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 7;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 127;
defparam ram_block1a5.port_a_logical_ram_depth = 128;
defparam ram_block1a5.port_a_logical_ram_width = 16;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 7;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "clock0";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 127;
defparam ram_block1a5.port_b_logical_ram_depth = 128;
defparam ram_block1a5.port_b_logical_ram_width = 16;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "old";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 7;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 127;
defparam ram_block1a4.port_a_logical_ram_depth = 128;
defparam ram_block1a4.port_a_logical_ram_width = 16;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 7;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "clock0";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 127;
defparam ram_block1a4.port_b_logical_ram_depth = 128;
defparam ram_block1a4.port_b_logical_ram_width = 16;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "old";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 7;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 127;
defparam ram_block1a6.port_a_logical_ram_depth = 128;
defparam ram_block1a6.port_a_logical_ram_width = 16;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 7;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "clock0";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 127;
defparam ram_block1a6.port_b_logical_ram_depth = 128;
defparam ram_block1a6.port_b_logical_ram_width = 16;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "old";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 7;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 127;
defparam ram_block1a2.port_a_logical_ram_depth = 128;
defparam ram_block1a2.port_a_logical_ram_width = 16;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 7;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "clock0";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 127;
defparam ram_block1a2.port_b_logical_ram_depth = 128;
defparam ram_block1a2.port_b_logical_ram_width = 16;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "old";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 7;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 127;
defparam ram_block1a1.port_a_logical_ram_depth = 128;
defparam ram_block1a1.port_a_logical_ram_width = 16;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 7;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "clock0";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 127;
defparam ram_block1a1.port_b_logical_ram_depth = 128;
defparam ram_block1a1.port_b_logical_ram_width = 16;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|asj_fft_4dp_ram_fft_120:dat_B|asj_fft_data_ram_fft_120:\\gen_rams:3:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_lmu3:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "old";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 7;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 127;
defparam ram_block1a0.port_a_logical_ram_depth = 128;
defparam ram_block1a0.port_a_logical_ram_width = 16;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 7;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "clock0";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 127;
defparam ram_block1a0.port_b_logical_ram_depth = 128;
defparam ram_block1a0.port_b_logical_ram_width = 16;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";

endmodule

module fft_asj_fft_bfp_ctrl_fft_120 (
	source_valid_ctrl_sop,
	stall_reg,
	source_stall_int_d,
	global_clock_enable,
	blk_exp_0,
	blk_exp_1,
	blk_exp_2,
	blk_exp_3,
	blk_exp_4,
	blk_exp_5,
	tdl_arr_4,
	slb_last_0,
	slb_last_1,
	slb_last_2,
	slb_i_0,
	slb_i_1,
	slb_i_2,
	slb_i_3,
	Mux2,
	tdl_arr_11,
	Mux1,
	en_slb,
	GND_port,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	source_valid_ctrl_sop;
input 	stall_reg;
input 	source_stall_int_d;
input 	global_clock_enable;
output 	blk_exp_0;
output 	blk_exp_1;
output 	blk_exp_2;
output 	blk_exp_3;
output 	blk_exp_4;
output 	blk_exp_5;
input 	tdl_arr_4;
output 	slb_last_0;
output 	slb_last_1;
output 	slb_last_2;
input 	slb_i_0;
input 	slb_i_1;
input 	slb_i_2;
input 	slb_i_3;
input 	Mux2;
input 	tdl_arr_11;
input 	Mux1;
input 	en_slb;
input 	GND_port;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \gen_quad_str_ctrl:gen_se_bfp:gen_4bit_accum:gen_cont:delay_next_pass2|tdl_arr[0]~q ;
wire \gen_quad_str_ctrl:gen_se_bfp:gen_4bit_accum:gen_cont:delay_next_pass|tdl_arr[10]~q ;
wire \blk_exp_acc[0]~6_combout ;
wire \blk_exp_acc[5]~8_combout ;
wire \blk_exp_acc[0]~9_combout ;
wire \blk_exp_acc[0]~10_combout ;
wire \blk_exp_acc[0]~q ;
wire \blk_exp~0_combout ;
wire \blk_exp[0]~1_combout ;
wire \blk_exp_acc[0]~7 ;
wire \blk_exp_acc[1]~11_combout ;
wire \blk_exp_acc[1]~q ;
wire \blk_exp~2_combout ;
wire \blk_exp_acc[1]~12 ;
wire \blk_exp_acc[2]~13_combout ;
wire \blk_exp_acc[2]~q ;
wire \blk_exp~3_combout ;
wire \blk_exp_acc[2]~14 ;
wire \blk_exp_acc[3]~15_combout ;
wire \blk_exp_acc[3]~q ;
wire \blk_exp~4_combout ;
wire \blk_exp_acc[3]~16 ;
wire \blk_exp_acc[4]~17_combout ;
wire \blk_exp_acc[4]~q ;
wire \blk_exp~5_combout ;
wire \blk_exp_acc[4]~18 ;
wire \blk_exp_acc[5]~19_combout ;
wire \blk_exp_acc[5]~q ;
wire \blk_exp~6_combout ;
wire \slb_last~8_combout ;
wire \slb_last[2]~4_combout ;
wire \slb_last[2]~5_combout ;
wire \slb_last~9_combout ;
wire \slb_last~6_combout ;
wire \slb_last~7_combout ;


fft_asj_fft_tdl_bit_rst_fft_120_1 \gen_quad_str_ctrl:gen_se_bfp:gen_4bit_accum:gen_cont:delay_next_pass2 (
	.global_clock_enable(global_clock_enable),
	.tdl_arr_0(\gen_quad_str_ctrl:gen_se_bfp:gen_4bit_accum:gen_cont:delay_next_pass2|tdl_arr[0]~q ),
	.tdl_arr_10(\gen_quad_str_ctrl:gen_se_bfp:gen_4bit_accum:gen_cont:delay_next_pass|tdl_arr[10]~q ),
	.clk(clk),
	.reset_n(reset_n));

fft_asj_fft_tdl_bit_rst_fft_120 \gen_quad_str_ctrl:gen_se_bfp:gen_4bit_accum:gen_cont:delay_next_pass (
	.global_clock_enable(global_clock_enable),
	.tdl_arr_10(\gen_quad_str_ctrl:gen_se_bfp:gen_4bit_accum:gen_cont:delay_next_pass|tdl_arr[10]~q ),
	.en_slb(en_slb),
	.clk(clk),
	.reset_n(reset_n));

dffeas \blk_exp[0] (
	.clk(clk),
	.d(\blk_exp~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\blk_exp[0]~1_combout ),
	.q(blk_exp_0),
	.prn(vcc));
defparam \blk_exp[0] .is_wysiwyg = "true";
defparam \blk_exp[0] .power_up = "low";

dffeas \blk_exp[1] (
	.clk(clk),
	.d(\blk_exp~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\blk_exp[0]~1_combout ),
	.q(blk_exp_1),
	.prn(vcc));
defparam \blk_exp[1] .is_wysiwyg = "true";
defparam \blk_exp[1] .power_up = "low";

dffeas \blk_exp[2] (
	.clk(clk),
	.d(\blk_exp~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\blk_exp[0]~1_combout ),
	.q(blk_exp_2),
	.prn(vcc));
defparam \blk_exp[2] .is_wysiwyg = "true";
defparam \blk_exp[2] .power_up = "low";

dffeas \blk_exp[3] (
	.clk(clk),
	.d(\blk_exp~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\blk_exp[0]~1_combout ),
	.q(blk_exp_3),
	.prn(vcc));
defparam \blk_exp[3] .is_wysiwyg = "true";
defparam \blk_exp[3] .power_up = "low";

dffeas \blk_exp[4] (
	.clk(clk),
	.d(\blk_exp~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\blk_exp[0]~1_combout ),
	.q(blk_exp_4),
	.prn(vcc));
defparam \blk_exp[4] .is_wysiwyg = "true";
defparam \blk_exp[4] .power_up = "low";

dffeas \blk_exp[5] (
	.clk(clk),
	.d(\blk_exp~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\blk_exp[0]~1_combout ),
	.q(blk_exp_5),
	.prn(vcc));
defparam \blk_exp[5] .is_wysiwyg = "true";
defparam \blk_exp[5] .power_up = "low";

dffeas \slb_last[0] (
	.clk(clk),
	.d(\slb_last~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\slb_last[2]~5_combout ),
	.q(slb_last_0),
	.prn(vcc));
defparam \slb_last[0] .is_wysiwyg = "true";
defparam \slb_last[0] .power_up = "low";

dffeas \slb_last[1] (
	.clk(clk),
	.d(\slb_last~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\slb_last[2]~5_combout ),
	.q(slb_last_1),
	.prn(vcc));
defparam \slb_last[1] .is_wysiwyg = "true";
defparam \slb_last[1] .power_up = "low";

dffeas \slb_last[2] (
	.clk(clk),
	.d(\slb_last~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\slb_last[2]~5_combout ),
	.q(slb_last_2),
	.prn(vcc));
defparam \slb_last[2] .is_wysiwyg = "true";
defparam \slb_last[2] .power_up = "low";

cycloneiii_lcell_comb \blk_exp_acc[0]~6 (
	.dataa(\blk_exp_acc[0]~q ),
	.datab(slb_last_0),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\blk_exp_acc[0]~6_combout ),
	.cout(\blk_exp_acc[0]~7 ));
defparam \blk_exp_acc[0]~6 .lut_mask = 16'h66EE;
defparam \blk_exp_acc[0]~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \blk_exp_acc[5]~8 (
	.dataa(reset_n),
	.datab(\gen_quad_str_ctrl:gen_se_bfp:gen_4bit_accum:gen_cont:delay_next_pass2|tdl_arr[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\blk_exp_acc[5]~8_combout ),
	.cout());
defparam \blk_exp_acc[5]~8 .lut_mask = 16'h7777;
defparam \blk_exp_acc[5]~8 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \blk_exp_acc[0]~9 (
	.dataa(\gen_quad_str_ctrl:gen_se_bfp:gen_4bit_accum:gen_cont:delay_next_pass2|tdl_arr[0]~q ),
	.datab(tdl_arr_4),
	.datac(reset_n),
	.datad(gnd),
	.cin(gnd),
	.combout(\blk_exp_acc[0]~9_combout ),
	.cout());
defparam \blk_exp_acc[0]~9 .lut_mask = 16'hEFEF;
defparam \blk_exp_acc[0]~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \blk_exp_acc[0]~10 (
	.dataa(source_stall_int_d),
	.datab(source_valid_ctrl_sop),
	.datac(stall_reg),
	.datad(\blk_exp_acc[0]~9_combout ),
	.cin(gnd),
	.combout(\blk_exp_acc[0]~10_combout ),
	.cout());
defparam \blk_exp_acc[0]~10 .lut_mask = 16'hF7D5;
defparam \blk_exp_acc[0]~10 .sum_lutc_input = "datac";

dffeas \blk_exp_acc[0] (
	.clk(clk),
	.d(\blk_exp_acc[0]~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\blk_exp_acc[5]~8_combout ),
	.ena(\blk_exp_acc[0]~10_combout ),
	.q(\blk_exp_acc[0]~q ),
	.prn(vcc));
defparam \blk_exp_acc[0] .is_wysiwyg = "true";
defparam \blk_exp_acc[0] .power_up = "low";

cycloneiii_lcell_comb \blk_exp~0 (
	.dataa(reset_n),
	.datab(\blk_exp_acc[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\blk_exp~0_combout ),
	.cout());
defparam \blk_exp~0 .lut_mask = 16'hEEEE;
defparam \blk_exp~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \blk_exp[0]~1 (
	.dataa(global_clock_enable),
	.datab(reset_n),
	.datac(\gen_quad_str_ctrl:gen_se_bfp:gen_4bit_accum:gen_cont:delay_next_pass2|tdl_arr[0]~q ),
	.datad(tdl_arr_4),
	.cin(gnd),
	.combout(\blk_exp[0]~1_combout ),
	.cout());
defparam \blk_exp[0]~1 .lut_mask = 16'hFFBF;
defparam \blk_exp[0]~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \blk_exp_acc[1]~11 (
	.dataa(\blk_exp_acc[1]~q ),
	.datab(slb_last_1),
	.datac(gnd),
	.datad(vcc),
	.cin(\blk_exp_acc[0]~7 ),
	.combout(\blk_exp_acc[1]~11_combout ),
	.cout(\blk_exp_acc[1]~12 ));
defparam \blk_exp_acc[1]~11 .lut_mask = 16'h967F;
defparam \blk_exp_acc[1]~11 .sum_lutc_input = "cin";

dffeas \blk_exp_acc[1] (
	.clk(clk),
	.d(\blk_exp_acc[1]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\blk_exp_acc[5]~8_combout ),
	.ena(\blk_exp_acc[0]~10_combout ),
	.q(\blk_exp_acc[1]~q ),
	.prn(vcc));
defparam \blk_exp_acc[1] .is_wysiwyg = "true";
defparam \blk_exp_acc[1] .power_up = "low";

cycloneiii_lcell_comb \blk_exp~2 (
	.dataa(reset_n),
	.datab(\blk_exp_acc[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\blk_exp~2_combout ),
	.cout());
defparam \blk_exp~2 .lut_mask = 16'hEEEE;
defparam \blk_exp~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \blk_exp_acc[2]~13 (
	.dataa(\blk_exp_acc[2]~q ),
	.datab(slb_last_2),
	.datac(gnd),
	.datad(vcc),
	.cin(\blk_exp_acc[1]~12 ),
	.combout(\blk_exp_acc[2]~13_combout ),
	.cout(\blk_exp_acc[2]~14 ));
defparam \blk_exp_acc[2]~13 .lut_mask = 16'h96EF;
defparam \blk_exp_acc[2]~13 .sum_lutc_input = "cin";

dffeas \blk_exp_acc[2] (
	.clk(clk),
	.d(\blk_exp_acc[2]~13_combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\blk_exp_acc[5]~8_combout ),
	.ena(\blk_exp_acc[0]~10_combout ),
	.q(\blk_exp_acc[2]~q ),
	.prn(vcc));
defparam \blk_exp_acc[2] .is_wysiwyg = "true";
defparam \blk_exp_acc[2] .power_up = "low";

cycloneiii_lcell_comb \blk_exp~3 (
	.dataa(reset_n),
	.datab(\blk_exp_acc[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\blk_exp~3_combout ),
	.cout());
defparam \blk_exp~3 .lut_mask = 16'hEEEE;
defparam \blk_exp~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \blk_exp_acc[3]~15 (
	.dataa(\blk_exp_acc[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\blk_exp_acc[2]~14 ),
	.combout(\blk_exp_acc[3]~15_combout ),
	.cout(\blk_exp_acc[3]~16 ));
defparam \blk_exp_acc[3]~15 .lut_mask = 16'h5A5F;
defparam \blk_exp_acc[3]~15 .sum_lutc_input = "cin";

dffeas \blk_exp_acc[3] (
	.clk(clk),
	.d(\blk_exp_acc[3]~15_combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\blk_exp_acc[5]~8_combout ),
	.ena(\blk_exp_acc[0]~10_combout ),
	.q(\blk_exp_acc[3]~q ),
	.prn(vcc));
defparam \blk_exp_acc[3] .is_wysiwyg = "true";
defparam \blk_exp_acc[3] .power_up = "low";

cycloneiii_lcell_comb \blk_exp~4 (
	.dataa(reset_n),
	.datab(\blk_exp_acc[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\blk_exp~4_combout ),
	.cout());
defparam \blk_exp~4 .lut_mask = 16'hEEEE;
defparam \blk_exp~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \blk_exp_acc[4]~17 (
	.dataa(\blk_exp_acc[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\blk_exp_acc[3]~16 ),
	.combout(\blk_exp_acc[4]~17_combout ),
	.cout(\blk_exp_acc[4]~18 ));
defparam \blk_exp_acc[4]~17 .lut_mask = 16'h5AAF;
defparam \blk_exp_acc[4]~17 .sum_lutc_input = "cin";

dffeas \blk_exp_acc[4] (
	.clk(clk),
	.d(\blk_exp_acc[4]~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\blk_exp_acc[5]~8_combout ),
	.ena(\blk_exp_acc[0]~10_combout ),
	.q(\blk_exp_acc[4]~q ),
	.prn(vcc));
defparam \blk_exp_acc[4] .is_wysiwyg = "true";
defparam \blk_exp_acc[4] .power_up = "low";

cycloneiii_lcell_comb \blk_exp~5 (
	.dataa(reset_n),
	.datab(\blk_exp_acc[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\blk_exp~5_combout ),
	.cout());
defparam \blk_exp~5 .lut_mask = 16'hEEEE;
defparam \blk_exp~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \blk_exp_acc[5]~19 (
	.dataa(\blk_exp_acc[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\blk_exp_acc[4]~18 ),
	.combout(\blk_exp_acc[5]~19_combout ),
	.cout());
defparam \blk_exp_acc[5]~19 .lut_mask = 16'h5A5A;
defparam \blk_exp_acc[5]~19 .sum_lutc_input = "cin";

dffeas \blk_exp_acc[5] (
	.clk(clk),
	.d(\blk_exp_acc[5]~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\blk_exp_acc[5]~8_combout ),
	.ena(\blk_exp_acc[0]~10_combout ),
	.q(\blk_exp_acc[5]~q ),
	.prn(vcc));
defparam \blk_exp_acc[5] .is_wysiwyg = "true";
defparam \blk_exp_acc[5] .power_up = "low";

cycloneiii_lcell_comb \blk_exp~6 (
	.dataa(reset_n),
	.datab(\blk_exp_acc[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\blk_exp~6_combout ),
	.cout());
defparam \blk_exp~6 .lut_mask = 16'hEEEE;
defparam \blk_exp~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \slb_last~8 (
	.dataa(reset_n),
	.datab(\gen_quad_str_ctrl:gen_se_bfp:gen_4bit_accum:gen_cont:delay_next_pass|tdl_arr[10]~q ),
	.datac(Mux2),
	.datad(gnd),
	.cin(gnd),
	.combout(\slb_last~8_combout ),
	.cout());
defparam \slb_last~8 .lut_mask = 16'hFEFE;
defparam \slb_last~8 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \slb_last[2]~4 (
	.dataa(\gen_quad_str_ctrl:gen_se_bfp:gen_4bit_accum:gen_cont:delay_next_pass|tdl_arr[10]~q ),
	.datab(tdl_arr_11),
	.datac(reset_n),
	.datad(gnd),
	.cin(gnd),
	.combout(\slb_last[2]~4_combout ),
	.cout());
defparam \slb_last[2]~4 .lut_mask = 16'hEFEF;
defparam \slb_last[2]~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \slb_last[2]~5 (
	.dataa(source_stall_int_d),
	.datab(source_valid_ctrl_sop),
	.datac(stall_reg),
	.datad(\slb_last[2]~4_combout ),
	.cin(gnd),
	.combout(\slb_last[2]~5_combout ),
	.cout());
defparam \slb_last[2]~5 .lut_mask = 16'hF7D5;
defparam \slb_last[2]~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \slb_last~9 (
	.dataa(reset_n),
	.datab(\gen_quad_str_ctrl:gen_se_bfp:gen_4bit_accum:gen_cont:delay_next_pass|tdl_arr[10]~q ),
	.datac(Mux1),
	.datad(gnd),
	.cin(gnd),
	.combout(\slb_last~9_combout ),
	.cout());
defparam \slb_last~9 .lut_mask = 16'hFEFE;
defparam \slb_last~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \slb_last~6 (
	.dataa(reset_n),
	.datab(\gen_quad_str_ctrl:gen_se_bfp:gen_4bit_accum:gen_cont:delay_next_pass|tdl_arr[10]~q ),
	.datac(slb_i_2),
	.datad(slb_i_3),
	.cin(gnd),
	.combout(\slb_last~6_combout ),
	.cout());
defparam \slb_last~6 .lut_mask = 16'hEFFF;
defparam \slb_last~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \slb_last~7 (
	.dataa(\slb_last~6_combout ),
	.datab(gnd),
	.datac(slb_i_0),
	.datad(slb_i_1),
	.cin(gnd),
	.combout(\slb_last~7_combout ),
	.cout());
defparam \slb_last~7 .lut_mask = 16'hAFFF;
defparam \slb_last~7 .sum_lutc_input = "datac";

endmodule

module fft_asj_fft_tdl_bit_rst_fft_120 (
	global_clock_enable,
	tdl_arr_10,
	en_slb,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	global_clock_enable;
output 	tdl_arr_10;
input 	en_slb;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \tdl_arr~10_combout ;
wire \tdl_arr[0]~q ;
wire \tdl_arr~9_combout ;
wire \tdl_arr[1]~q ;
wire \tdl_arr~8_combout ;
wire \tdl_arr[2]~q ;
wire \tdl_arr~7_combout ;
wire \tdl_arr[3]~q ;
wire \tdl_arr~6_combout ;
wire \tdl_arr[4]~q ;
wire \tdl_arr~5_combout ;
wire \tdl_arr[5]~q ;
wire \tdl_arr~4_combout ;
wire \tdl_arr[6]~q ;
wire \tdl_arr~3_combout ;
wire \tdl_arr[7]~q ;
wire \tdl_arr~2_combout ;
wire \tdl_arr[8]~q ;
wire \tdl_arr~1_combout ;
wire \tdl_arr[9]~q ;
wire \tdl_arr~0_combout ;


dffeas \tdl_arr[10] (
	.clk(clk),
	.d(\tdl_arr~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_10),
	.prn(vcc));
defparam \tdl_arr[10] .is_wysiwyg = "true";
defparam \tdl_arr[10] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~10 (
	.dataa(reset_n),
	.datab(en_slb),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~10_combout ),
	.cout());
defparam \tdl_arr~10 .lut_mask = 16'hEEEE;
defparam \tdl_arr~10 .sum_lutc_input = "datac";

dffeas \tdl_arr[0] (
	.clk(clk),
	.d(\tdl_arr~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0]~q ),
	.prn(vcc));
defparam \tdl_arr[0] .is_wysiwyg = "true";
defparam \tdl_arr[0] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~9 (
	.dataa(reset_n),
	.datab(\tdl_arr[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~9_combout ),
	.cout());
defparam \tdl_arr~9 .lut_mask = 16'hEEEE;
defparam \tdl_arr~9 .sum_lutc_input = "datac";

dffeas \tdl_arr[1] (
	.clk(clk),
	.d(\tdl_arr~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[1]~q ),
	.prn(vcc));
defparam \tdl_arr[1] .is_wysiwyg = "true";
defparam \tdl_arr[1] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~8 (
	.dataa(reset_n),
	.datab(\tdl_arr[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~8_combout ),
	.cout());
defparam \tdl_arr~8 .lut_mask = 16'hEEEE;
defparam \tdl_arr~8 .sum_lutc_input = "datac";

dffeas \tdl_arr[2] (
	.clk(clk),
	.d(\tdl_arr~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[2]~q ),
	.prn(vcc));
defparam \tdl_arr[2] .is_wysiwyg = "true";
defparam \tdl_arr[2] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~7 (
	.dataa(reset_n),
	.datab(\tdl_arr[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~7_combout ),
	.cout());
defparam \tdl_arr~7 .lut_mask = 16'hEEEE;
defparam \tdl_arr~7 .sum_lutc_input = "datac";

dffeas \tdl_arr[3] (
	.clk(clk),
	.d(\tdl_arr~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[3]~q ),
	.prn(vcc));
defparam \tdl_arr[3] .is_wysiwyg = "true";
defparam \tdl_arr[3] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~6 (
	.dataa(reset_n),
	.datab(\tdl_arr[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~6_combout ),
	.cout());
defparam \tdl_arr~6 .lut_mask = 16'hEEEE;
defparam \tdl_arr~6 .sum_lutc_input = "datac";

dffeas \tdl_arr[4] (
	.clk(clk),
	.d(\tdl_arr~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[4]~q ),
	.prn(vcc));
defparam \tdl_arr[4] .is_wysiwyg = "true";
defparam \tdl_arr[4] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~5 (
	.dataa(reset_n),
	.datab(\tdl_arr[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~5_combout ),
	.cout());
defparam \tdl_arr~5 .lut_mask = 16'hEEEE;
defparam \tdl_arr~5 .sum_lutc_input = "datac";

dffeas \tdl_arr[5] (
	.clk(clk),
	.d(\tdl_arr~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[5]~q ),
	.prn(vcc));
defparam \tdl_arr[5] .is_wysiwyg = "true";
defparam \tdl_arr[5] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~4 (
	.dataa(reset_n),
	.datab(\tdl_arr[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~4_combout ),
	.cout());
defparam \tdl_arr~4 .lut_mask = 16'hEEEE;
defparam \tdl_arr~4 .sum_lutc_input = "datac";

dffeas \tdl_arr[6] (
	.clk(clk),
	.d(\tdl_arr~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[6]~q ),
	.prn(vcc));
defparam \tdl_arr[6] .is_wysiwyg = "true";
defparam \tdl_arr[6] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~3 (
	.dataa(reset_n),
	.datab(\tdl_arr[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~3_combout ),
	.cout());
defparam \tdl_arr~3 .lut_mask = 16'hEEEE;
defparam \tdl_arr~3 .sum_lutc_input = "datac";

dffeas \tdl_arr[7] (
	.clk(clk),
	.d(\tdl_arr~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[7]~q ),
	.prn(vcc));
defparam \tdl_arr[7] .is_wysiwyg = "true";
defparam \tdl_arr[7] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~2 (
	.dataa(reset_n),
	.datab(\tdl_arr[7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~2_combout ),
	.cout());
defparam \tdl_arr~2 .lut_mask = 16'hEEEE;
defparam \tdl_arr~2 .sum_lutc_input = "datac";

dffeas \tdl_arr[8] (
	.clk(clk),
	.d(\tdl_arr~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[8]~q ),
	.prn(vcc));
defparam \tdl_arr[8] .is_wysiwyg = "true";
defparam \tdl_arr[8] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~1 (
	.dataa(reset_n),
	.datab(\tdl_arr[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~1_combout ),
	.cout());
defparam \tdl_arr~1 .lut_mask = 16'hEEEE;
defparam \tdl_arr~1 .sum_lutc_input = "datac";

dffeas \tdl_arr[9] (
	.clk(clk),
	.d(\tdl_arr~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[9]~q ),
	.prn(vcc));
defparam \tdl_arr[9] .is_wysiwyg = "true";
defparam \tdl_arr[9] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~0 (
	.dataa(reset_n),
	.datab(\tdl_arr[9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~0_combout ),
	.cout());
defparam \tdl_arr~0 .lut_mask = 16'hEEEE;
defparam \tdl_arr~0 .sum_lutc_input = "datac";

endmodule

module fft_asj_fft_tdl_bit_rst_fft_120_1 (
	global_clock_enable,
	tdl_arr_0,
	tdl_arr_10,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	global_clock_enable;
output 	tdl_arr_0;
input 	tdl_arr_10;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \tdl_arr~0_combout ;


dffeas \tdl_arr[0] (
	.clk(clk),
	.d(\tdl_arr~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_0),
	.prn(vcc));
defparam \tdl_arr[0] .is_wysiwyg = "true";
defparam \tdl_arr[0] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~0 (
	.dataa(reset_n),
	.datab(tdl_arr_10),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~0_combout ),
	.cout());
defparam \tdl_arr~0 .lut_mask = 16'hEEEE;
defparam \tdl_arr~0 .sum_lutc_input = "datac";

endmodule

module fft_asj_fft_cnt_ctrl_fft_120 (
	ram_in_reg_1_6,
	ram_in_reg_1_5,
	ram_in_reg_1_4,
	ram_in_reg_1_7,
	ram_in_reg_0_6,
	ram_in_reg_0_5,
	ram_in_reg_0_4,
	ram_in_reg_0_7,
	ram_in_reg_7_6,
	ram_in_reg_7_5,
	ram_in_reg_7_4,
	ram_in_reg_7_7,
	ram_in_reg_6_6,
	ram_in_reg_6_5,
	ram_in_reg_6_4,
	ram_in_reg_6_7,
	ram_in_reg_5_6,
	ram_in_reg_5_5,
	ram_in_reg_5_4,
	ram_in_reg_5_7,
	ram_in_reg_4_6,
	ram_in_reg_4_5,
	ram_in_reg_4_4,
	ram_in_reg_4_7,
	ram_in_reg_3_6,
	ram_in_reg_3_5,
	ram_in_reg_3_4,
	ram_in_reg_3_7,
	ram_in_reg_2_6,
	ram_in_reg_2_5,
	ram_in_reg_2_4,
	ram_in_reg_2_7,
	ram_in_reg_1_2,
	ram_in_reg_1_1,
	ram_in_reg_1_0,
	ram_in_reg_1_3,
	ram_in_reg_0_2,
	ram_in_reg_0_1,
	ram_in_reg_0_0,
	ram_in_reg_0_3,
	ram_in_reg_7_2,
	ram_in_reg_7_1,
	ram_in_reg_7_0,
	ram_in_reg_7_3,
	ram_in_reg_6_2,
	ram_in_reg_6_1,
	ram_in_reg_6_0,
	ram_in_reg_6_3,
	ram_in_reg_5_2,
	ram_in_reg_5_1,
	ram_in_reg_5_0,
	ram_in_reg_5_3,
	ram_in_reg_4_2,
	ram_in_reg_4_1,
	ram_in_reg_4_0,
	ram_in_reg_4_3,
	ram_in_reg_3_2,
	ram_in_reg_3_1,
	ram_in_reg_3_0,
	ram_in_reg_3_3,
	ram_in_reg_2_2,
	ram_in_reg_2_1,
	ram_in_reg_2_0,
	ram_in_reg_2_3,
	q_b_10,
	q_b_101,
	q_b_102,
	q_b_103,
	q_b_104,
	q_b_105,
	q_b_106,
	q_b_107,
	q_b_14,
	q_b_141,
	q_b_142,
	q_b_143,
	q_b_144,
	q_b_145,
	q_b_146,
	q_b_147,
	q_b_12,
	q_b_121,
	q_b_122,
	q_b_123,
	q_b_124,
	q_b_125,
	q_b_126,
	q_b_127,
	q_b_11,
	q_b_111,
	q_b_112,
	q_b_113,
	q_b_114,
	q_b_115,
	q_b_116,
	q_b_117,
	q_b_13,
	q_b_131,
	q_b_132,
	q_b_133,
	q_b_134,
	q_b_135,
	q_b_136,
	q_b_137,
	q_b_9,
	q_b_91,
	q_b_92,
	q_b_93,
	q_b_94,
	q_b_95,
	q_b_96,
	q_b_97,
	q_b_8,
	q_b_81,
	q_b_82,
	q_b_83,
	q_b_84,
	q_b_85,
	q_b_86,
	q_b_87,
	q_b_15,
	q_b_151,
	q_b_152,
	q_b_153,
	q_b_154,
	q_b_155,
	q_b_156,
	q_b_157,
	q_b_7,
	q_b_71,
	q_b_72,
	q_b_73,
	q_b_74,
	q_b_75,
	q_b_76,
	q_b_77,
	q_b_3,
	q_b_31,
	q_b_32,
	q_b_33,
	q_b_34,
	q_b_35,
	q_b_36,
	q_b_37,
	q_b_5,
	q_b_51,
	q_b_52,
	q_b_53,
	q_b_54,
	q_b_55,
	q_b_56,
	q_b_57,
	q_b_4,
	q_b_41,
	q_b_42,
	q_b_43,
	q_b_44,
	q_b_45,
	q_b_46,
	q_b_47,
	q_b_6,
	q_b_61,
	q_b_62,
	q_b_63,
	q_b_64,
	q_b_65,
	q_b_66,
	q_b_67,
	q_b_2,
	q_b_21,
	q_b_22,
	q_b_23,
	q_b_24,
	q_b_25,
	q_b_26,
	q_b_27,
	q_b_1,
	q_b_16,
	q_b_17,
	q_b_18,
	q_b_19,
	q_b_110,
	q_b_118,
	q_b_119,
	q_b_0,
	q_b_01,
	q_b_02,
	q_b_03,
	q_b_04,
	q_b_05,
	q_b_06,
	q_b_07,
	global_clock_enable,
	ram_in_reg_0_01,
	ram_in_reg_1_21,
	ram_in_reg_2_01,
	ram_in_reg_3_21,
	ram_in_reg_4_01,
	ram_in_reg_5_21,
	ram_in_reg_6_01,
	ram_in_reg_0_11,
	ram_in_reg_1_11,
	ram_in_reg_2_11,
	ram_in_reg_3_11,
	ram_in_reg_4_11,
	ram_in_reg_5_11,
	ram_in_reg_1_01,
	ram_in_reg_3_01,
	ram_in_reg_5_01,
	ram_in_reg_1_31,
	ram_in_reg_3_31,
	ram_in_reg_5_31,
	ram_data_out0_10,
	ram_data_out1_10,
	ram_data_out2_10,
	ram_data_out3_10,
	ram_data_out0_14,
	ram_data_out1_14,
	ram_data_out2_14,
	ram_data_out3_14,
	ram_data_out0_12,
	ram_data_out1_12,
	ram_data_out2_12,
	ram_data_out3_12,
	ram_data_out0_11,
	ram_data_out1_11,
	ram_data_out2_11,
	ram_data_out3_11,
	ram_data_out0_13,
	ram_data_out1_13,
	ram_data_out2_13,
	ram_data_out3_13,
	ram_data_out0_9,
	ram_data_out1_9,
	ram_data_out2_9,
	ram_data_out3_9,
	ram_data_out0_8,
	ram_data_out1_8,
	ram_data_out2_8,
	ram_data_out3_8,
	ram_data_out0_15,
	ram_data_out1_15,
	ram_data_out2_15,
	ram_data_out3_15,
	ram_data_out0_7,
	ram_data_out1_7,
	ram_data_out2_7,
	ram_data_out3_7,
	ram_data_out0_3,
	ram_data_out1_3,
	ram_data_out2_3,
	ram_data_out3_3,
	ram_data_out0_5,
	ram_data_out1_5,
	ram_data_out2_5,
	ram_data_out3_5,
	ram_data_out0_4,
	ram_data_out1_4,
	ram_data_out2_4,
	ram_data_out3_4,
	ram_data_out0_6,
	ram_data_out1_6,
	ram_data_out2_6,
	ram_data_out3_6,
	ram_data_out0_2,
	ram_data_out1_2,
	ram_data_out2_2,
	ram_data_out3_2,
	ram_data_out0_1,
	ram_data_out1_1,
	ram_data_out2_1,
	ram_data_out3_1,
	ram_data_out0_0,
	ram_data_out1_0,
	ram_data_out2_0,
	ram_data_out3_0,
	data_rdy_vec_10,
	ram_a_not_b_vec_10,
	b_ram_data_in_bus_58,
	wraddress_b_bus_21,
	wraddress_b_bus_22,
	wraddress_b_bus_23,
	wraddress_b_bus_24,
	wraddress_b_bus_11,
	wraddress_b_bus_26,
	wraddress_b_bus_13,
	rdaddress_b_bus_21,
	rdaddress_b_bus_22,
	rdaddress_b_bus_23,
	rdaddress_b_bus_24,
	rdaddress_b_bus_11,
	rdaddress_b_bus_26,
	rdaddress_b_bus_13,
	a_ram_data_in_bus_58,
	wraddress_a_bus_21,
	wraddress_a_bus_22,
	wraddress_a_bus_23,
	wraddress_a_bus_24,
	wraddress_a_bus_11,
	wraddress_a_bus_26,
	wraddress_a_bus_13,
	rdaddress_a_bus_21,
	rdaddress_a_bus_22,
	rdaddress_a_bus_23,
	rdaddress_a_bus_24,
	rdaddress_a_bus_11,
	rdaddress_a_bus_26,
	rdaddress_a_bus_13,
	b_ram_data_in_bus_42,
	wraddress_b_bus_0,
	wraddress_b_bus_15,
	wraddress_b_bus_16,
	wraddress_b_bus_17,
	wraddress_b_bus_18,
	wraddress_b_bus_19,
	rdaddress_b_bus_0,
	rdaddress_b_bus_15,
	rdaddress_b_bus_16,
	rdaddress_b_bus_17,
	rdaddress_b_bus_18,
	rdaddress_b_bus_19,
	a_ram_data_in_bus_42,
	wraddress_a_bus_0,
	wraddress_a_bus_15,
	wraddress_a_bus_16,
	wraddress_a_bus_17,
	wraddress_a_bus_18,
	wraddress_a_bus_19,
	rdaddress_a_bus_0,
	rdaddress_a_bus_15,
	rdaddress_a_bus_16,
	rdaddress_a_bus_17,
	rdaddress_a_bus_18,
	rdaddress_a_bus_19,
	b_ram_data_in_bus_26,
	wraddress_b_bus_8,
	wraddress_b_bus_10,
	wraddress_b_bus_12,
	rdaddress_b_bus_8,
	rdaddress_b_bus_10,
	rdaddress_b_bus_12,
	a_ram_data_in_bus_26,
	wraddress_a_bus_8,
	wraddress_a_bus_10,
	wraddress_a_bus_12,
	rdaddress_a_bus_8,
	rdaddress_a_bus_10,
	rdaddress_a_bus_12,
	b_ram_data_in_bus_10,
	wraddress_b_bus_1,
	wraddress_b_bus_3,
	wraddress_b_bus_5,
	rdaddress_b_bus_1,
	rdaddress_b_bus_3,
	rdaddress_b_bus_5,
	a_ram_data_in_bus_10,
	wraddress_a_bus_1,
	wraddress_a_bus_3,
	wraddress_a_bus_5,
	rdaddress_a_bus_1,
	rdaddress_a_bus_3,
	rdaddress_a_bus_5,
	b_ram_data_in_bus_62,
	a_ram_data_in_bus_62,
	b_ram_data_in_bus_46,
	a_ram_data_in_bus_46,
	b_ram_data_in_bus_30,
	a_ram_data_in_bus_30,
	b_ram_data_in_bus_14,
	a_ram_data_in_bus_14,
	b_ram_data_in_bus_60,
	a_ram_data_in_bus_60,
	b_ram_data_in_bus_44,
	a_ram_data_in_bus_44,
	b_ram_data_in_bus_28,
	a_ram_data_in_bus_28,
	b_ram_data_in_bus_12,
	a_ram_data_in_bus_12,
	b_ram_data_in_bus_59,
	a_ram_data_in_bus_59,
	b_ram_data_in_bus_43,
	a_ram_data_in_bus_43,
	b_ram_data_in_bus_27,
	a_ram_data_in_bus_27,
	b_ram_data_in_bus_11,
	a_ram_data_in_bus_11,
	b_ram_data_in_bus_61,
	a_ram_data_in_bus_61,
	b_ram_data_in_bus_45,
	a_ram_data_in_bus_45,
	b_ram_data_in_bus_29,
	a_ram_data_in_bus_29,
	b_ram_data_in_bus_13,
	a_ram_data_in_bus_13,
	b_ram_data_in_bus_57,
	a_ram_data_in_bus_57,
	b_ram_data_in_bus_41,
	a_ram_data_in_bus_41,
	b_ram_data_in_bus_25,
	a_ram_data_in_bus_25,
	b_ram_data_in_bus_9,
	a_ram_data_in_bus_9,
	b_ram_data_in_bus_56,
	a_ram_data_in_bus_56,
	b_ram_data_in_bus_40,
	a_ram_data_in_bus_40,
	b_ram_data_in_bus_24,
	a_ram_data_in_bus_24,
	b_ram_data_in_bus_8,
	a_ram_data_in_bus_8,
	b_ram_data_in_bus_63,
	a_ram_data_in_bus_63,
	b_ram_data_in_bus_47,
	a_ram_data_in_bus_47,
	b_ram_data_in_bus_31,
	a_ram_data_in_bus_31,
	b_ram_data_in_bus_15,
	a_ram_data_in_bus_15,
	b_ram_data_in_bus_55,
	a_ram_data_in_bus_55,
	b_ram_data_in_bus_39,
	a_ram_data_in_bus_39,
	b_ram_data_in_bus_23,
	a_ram_data_in_bus_23,
	b_ram_data_in_bus_7,
	a_ram_data_in_bus_7,
	b_ram_data_in_bus_51,
	a_ram_data_in_bus_51,
	b_ram_data_in_bus_35,
	a_ram_data_in_bus_35,
	b_ram_data_in_bus_19,
	a_ram_data_in_bus_19,
	b_ram_data_in_bus_3,
	a_ram_data_in_bus_3,
	b_ram_data_in_bus_53,
	a_ram_data_in_bus_53,
	b_ram_data_in_bus_37,
	a_ram_data_in_bus_37,
	b_ram_data_in_bus_21,
	a_ram_data_in_bus_21,
	b_ram_data_in_bus_5,
	a_ram_data_in_bus_5,
	b_ram_data_in_bus_52,
	a_ram_data_in_bus_52,
	b_ram_data_in_bus_36,
	a_ram_data_in_bus_36,
	b_ram_data_in_bus_20,
	a_ram_data_in_bus_20,
	b_ram_data_in_bus_4,
	a_ram_data_in_bus_4,
	b_ram_data_in_bus_54,
	a_ram_data_in_bus_54,
	b_ram_data_in_bus_38,
	a_ram_data_in_bus_38,
	b_ram_data_in_bus_22,
	a_ram_data_in_bus_22,
	b_ram_data_in_bus_6,
	a_ram_data_in_bus_6,
	b_ram_data_in_bus_50,
	a_ram_data_in_bus_50,
	b_ram_data_in_bus_34,
	a_ram_data_in_bus_34,
	b_ram_data_in_bus_18,
	a_ram_data_in_bus_18,
	b_ram_data_in_bus_2,
	a_ram_data_in_bus_2,
	b_ram_data_in_bus_49,
	a_ram_data_in_bus_49,
	b_ram_data_in_bus_33,
	a_ram_data_in_bus_33,
	b_ram_data_in_bus_17,
	a_ram_data_in_bus_17,
	b_ram_data_in_bus_1,
	a_ram_data_in_bus_1,
	b_ram_data_in_bus_48,
	a_ram_data_in_bus_48,
	b_ram_data_in_bus_32,
	a_ram_data_in_bus_32,
	b_ram_data_in_bus_16,
	a_ram_data_in_bus_16,
	b_ram_data_in_bus_0,
	a_ram_data_in_bus_0,
	ram_a_not_b_vec_1,
	data_in_r_2,
	wr_address_i_int_0,
	wr_address_i_int_1,
	wr_address_i_int_2,
	wr_address_i_int_3,
	wr_address_i_int_4,
	wr_address_i_int_5,
	wr_address_i_int_6,
	ram_a_not_b_vec_7,
	ram_in_reg_0_02,
	ram_in_reg_1_02,
	ram_in_reg_2_02,
	ram_in_reg_3_02,
	ram_in_reg_4_02,
	ram_in_reg_5_02,
	tdl_arr_6_1,
	ram_in_reg_0_12,
	ram_in_reg_1_12,
	ram_in_reg_2_12,
	ram_in_reg_3_12,
	ram_in_reg_4_12,
	ram_in_reg_5_12,
	ram_in_reg_1_22,
	ram_in_reg_3_22,
	ram_in_reg_5_22,
	ram_in_reg_1_32,
	ram_in_reg_3_32,
	ram_in_reg_5_32,
	data_in_r_6,
	data_in_r_4,
	data_in_r_3,
	data_in_r_5,
	data_in_r_1,
	data_in_r_0,
	data_in_r_7,
	data_in_i_7,
	data_in_i_3,
	data_in_i_5,
	data_in_i_4,
	data_in_i_6,
	data_in_i_2,
	data_in_i_1,
	data_in_i_0,
	clk)/* synthesis synthesis_greybox=1 */;
input 	ram_in_reg_1_6;
input 	ram_in_reg_1_5;
input 	ram_in_reg_1_4;
input 	ram_in_reg_1_7;
input 	ram_in_reg_0_6;
input 	ram_in_reg_0_5;
input 	ram_in_reg_0_4;
input 	ram_in_reg_0_7;
input 	ram_in_reg_7_6;
input 	ram_in_reg_7_5;
input 	ram_in_reg_7_4;
input 	ram_in_reg_7_7;
input 	ram_in_reg_6_6;
input 	ram_in_reg_6_5;
input 	ram_in_reg_6_4;
input 	ram_in_reg_6_7;
input 	ram_in_reg_5_6;
input 	ram_in_reg_5_5;
input 	ram_in_reg_5_4;
input 	ram_in_reg_5_7;
input 	ram_in_reg_4_6;
input 	ram_in_reg_4_5;
input 	ram_in_reg_4_4;
input 	ram_in_reg_4_7;
input 	ram_in_reg_3_6;
input 	ram_in_reg_3_5;
input 	ram_in_reg_3_4;
input 	ram_in_reg_3_7;
input 	ram_in_reg_2_6;
input 	ram_in_reg_2_5;
input 	ram_in_reg_2_4;
input 	ram_in_reg_2_7;
input 	ram_in_reg_1_2;
input 	ram_in_reg_1_1;
input 	ram_in_reg_1_0;
input 	ram_in_reg_1_3;
input 	ram_in_reg_0_2;
input 	ram_in_reg_0_1;
input 	ram_in_reg_0_0;
input 	ram_in_reg_0_3;
input 	ram_in_reg_7_2;
input 	ram_in_reg_7_1;
input 	ram_in_reg_7_0;
input 	ram_in_reg_7_3;
input 	ram_in_reg_6_2;
input 	ram_in_reg_6_1;
input 	ram_in_reg_6_0;
input 	ram_in_reg_6_3;
input 	ram_in_reg_5_2;
input 	ram_in_reg_5_1;
input 	ram_in_reg_5_0;
input 	ram_in_reg_5_3;
input 	ram_in_reg_4_2;
input 	ram_in_reg_4_1;
input 	ram_in_reg_4_0;
input 	ram_in_reg_4_3;
input 	ram_in_reg_3_2;
input 	ram_in_reg_3_1;
input 	ram_in_reg_3_0;
input 	ram_in_reg_3_3;
input 	ram_in_reg_2_2;
input 	ram_in_reg_2_1;
input 	ram_in_reg_2_0;
input 	ram_in_reg_2_3;
input 	q_b_10;
input 	q_b_101;
input 	q_b_102;
input 	q_b_103;
input 	q_b_104;
input 	q_b_105;
input 	q_b_106;
input 	q_b_107;
input 	q_b_14;
input 	q_b_141;
input 	q_b_142;
input 	q_b_143;
input 	q_b_144;
input 	q_b_145;
input 	q_b_146;
input 	q_b_147;
input 	q_b_12;
input 	q_b_121;
input 	q_b_122;
input 	q_b_123;
input 	q_b_124;
input 	q_b_125;
input 	q_b_126;
input 	q_b_127;
input 	q_b_11;
input 	q_b_111;
input 	q_b_112;
input 	q_b_113;
input 	q_b_114;
input 	q_b_115;
input 	q_b_116;
input 	q_b_117;
input 	q_b_13;
input 	q_b_131;
input 	q_b_132;
input 	q_b_133;
input 	q_b_134;
input 	q_b_135;
input 	q_b_136;
input 	q_b_137;
input 	q_b_9;
input 	q_b_91;
input 	q_b_92;
input 	q_b_93;
input 	q_b_94;
input 	q_b_95;
input 	q_b_96;
input 	q_b_97;
input 	q_b_8;
input 	q_b_81;
input 	q_b_82;
input 	q_b_83;
input 	q_b_84;
input 	q_b_85;
input 	q_b_86;
input 	q_b_87;
input 	q_b_15;
input 	q_b_151;
input 	q_b_152;
input 	q_b_153;
input 	q_b_154;
input 	q_b_155;
input 	q_b_156;
input 	q_b_157;
input 	q_b_7;
input 	q_b_71;
input 	q_b_72;
input 	q_b_73;
input 	q_b_74;
input 	q_b_75;
input 	q_b_76;
input 	q_b_77;
input 	q_b_3;
input 	q_b_31;
input 	q_b_32;
input 	q_b_33;
input 	q_b_34;
input 	q_b_35;
input 	q_b_36;
input 	q_b_37;
input 	q_b_5;
input 	q_b_51;
input 	q_b_52;
input 	q_b_53;
input 	q_b_54;
input 	q_b_55;
input 	q_b_56;
input 	q_b_57;
input 	q_b_4;
input 	q_b_41;
input 	q_b_42;
input 	q_b_43;
input 	q_b_44;
input 	q_b_45;
input 	q_b_46;
input 	q_b_47;
input 	q_b_6;
input 	q_b_61;
input 	q_b_62;
input 	q_b_63;
input 	q_b_64;
input 	q_b_65;
input 	q_b_66;
input 	q_b_67;
input 	q_b_2;
input 	q_b_21;
input 	q_b_22;
input 	q_b_23;
input 	q_b_24;
input 	q_b_25;
input 	q_b_26;
input 	q_b_27;
input 	q_b_1;
input 	q_b_16;
input 	q_b_17;
input 	q_b_18;
input 	q_b_19;
input 	q_b_110;
input 	q_b_118;
input 	q_b_119;
input 	q_b_0;
input 	q_b_01;
input 	q_b_02;
input 	q_b_03;
input 	q_b_04;
input 	q_b_05;
input 	q_b_06;
input 	q_b_07;
input 	global_clock_enable;
input 	ram_in_reg_0_01;
input 	ram_in_reg_1_21;
input 	ram_in_reg_2_01;
input 	ram_in_reg_3_21;
input 	ram_in_reg_4_01;
input 	ram_in_reg_5_21;
input 	ram_in_reg_6_01;
input 	ram_in_reg_0_11;
input 	ram_in_reg_1_11;
input 	ram_in_reg_2_11;
input 	ram_in_reg_3_11;
input 	ram_in_reg_4_11;
input 	ram_in_reg_5_11;
input 	ram_in_reg_1_01;
input 	ram_in_reg_3_01;
input 	ram_in_reg_5_01;
input 	ram_in_reg_1_31;
input 	ram_in_reg_3_31;
input 	ram_in_reg_5_31;
output 	ram_data_out0_10;
output 	ram_data_out1_10;
output 	ram_data_out2_10;
output 	ram_data_out3_10;
output 	ram_data_out0_14;
output 	ram_data_out1_14;
output 	ram_data_out2_14;
output 	ram_data_out3_14;
output 	ram_data_out0_12;
output 	ram_data_out1_12;
output 	ram_data_out2_12;
output 	ram_data_out3_12;
output 	ram_data_out0_11;
output 	ram_data_out1_11;
output 	ram_data_out2_11;
output 	ram_data_out3_11;
output 	ram_data_out0_13;
output 	ram_data_out1_13;
output 	ram_data_out2_13;
output 	ram_data_out3_13;
output 	ram_data_out0_9;
output 	ram_data_out1_9;
output 	ram_data_out2_9;
output 	ram_data_out3_9;
output 	ram_data_out0_8;
output 	ram_data_out1_8;
output 	ram_data_out2_8;
output 	ram_data_out3_8;
output 	ram_data_out0_15;
output 	ram_data_out1_15;
output 	ram_data_out2_15;
output 	ram_data_out3_15;
output 	ram_data_out0_7;
output 	ram_data_out1_7;
output 	ram_data_out2_7;
output 	ram_data_out3_7;
output 	ram_data_out0_3;
output 	ram_data_out1_3;
output 	ram_data_out2_3;
output 	ram_data_out3_3;
output 	ram_data_out0_5;
output 	ram_data_out1_5;
output 	ram_data_out2_5;
output 	ram_data_out3_5;
output 	ram_data_out0_4;
output 	ram_data_out1_4;
output 	ram_data_out2_4;
output 	ram_data_out3_4;
output 	ram_data_out0_6;
output 	ram_data_out1_6;
output 	ram_data_out2_6;
output 	ram_data_out3_6;
output 	ram_data_out0_2;
output 	ram_data_out1_2;
output 	ram_data_out2_2;
output 	ram_data_out3_2;
output 	ram_data_out0_1;
output 	ram_data_out1_1;
output 	ram_data_out2_1;
output 	ram_data_out3_1;
output 	ram_data_out0_0;
output 	ram_data_out1_0;
output 	ram_data_out2_0;
output 	ram_data_out3_0;
input 	data_rdy_vec_10;
input 	ram_a_not_b_vec_10;
output 	b_ram_data_in_bus_58;
output 	wraddress_b_bus_21;
output 	wraddress_b_bus_22;
output 	wraddress_b_bus_23;
output 	wraddress_b_bus_24;
output 	wraddress_b_bus_11;
output 	wraddress_b_bus_26;
output 	wraddress_b_bus_13;
output 	rdaddress_b_bus_21;
output 	rdaddress_b_bus_22;
output 	rdaddress_b_bus_23;
output 	rdaddress_b_bus_24;
output 	rdaddress_b_bus_11;
output 	rdaddress_b_bus_26;
output 	rdaddress_b_bus_13;
output 	a_ram_data_in_bus_58;
output 	wraddress_a_bus_21;
output 	wraddress_a_bus_22;
output 	wraddress_a_bus_23;
output 	wraddress_a_bus_24;
output 	wraddress_a_bus_11;
output 	wraddress_a_bus_26;
output 	wraddress_a_bus_13;
output 	rdaddress_a_bus_21;
output 	rdaddress_a_bus_22;
output 	rdaddress_a_bus_23;
output 	rdaddress_a_bus_24;
output 	rdaddress_a_bus_11;
output 	rdaddress_a_bus_26;
output 	rdaddress_a_bus_13;
output 	b_ram_data_in_bus_42;
output 	wraddress_b_bus_0;
output 	wraddress_b_bus_15;
output 	wraddress_b_bus_16;
output 	wraddress_b_bus_17;
output 	wraddress_b_bus_18;
output 	wraddress_b_bus_19;
output 	rdaddress_b_bus_0;
output 	rdaddress_b_bus_15;
output 	rdaddress_b_bus_16;
output 	rdaddress_b_bus_17;
output 	rdaddress_b_bus_18;
output 	rdaddress_b_bus_19;
output 	a_ram_data_in_bus_42;
output 	wraddress_a_bus_0;
output 	wraddress_a_bus_15;
output 	wraddress_a_bus_16;
output 	wraddress_a_bus_17;
output 	wraddress_a_bus_18;
output 	wraddress_a_bus_19;
output 	rdaddress_a_bus_0;
output 	rdaddress_a_bus_15;
output 	rdaddress_a_bus_16;
output 	rdaddress_a_bus_17;
output 	rdaddress_a_bus_18;
output 	rdaddress_a_bus_19;
output 	b_ram_data_in_bus_26;
output 	wraddress_b_bus_8;
output 	wraddress_b_bus_10;
output 	wraddress_b_bus_12;
output 	rdaddress_b_bus_8;
output 	rdaddress_b_bus_10;
output 	rdaddress_b_bus_12;
output 	a_ram_data_in_bus_26;
output 	wraddress_a_bus_8;
output 	wraddress_a_bus_10;
output 	wraddress_a_bus_12;
output 	rdaddress_a_bus_8;
output 	rdaddress_a_bus_10;
output 	rdaddress_a_bus_12;
output 	b_ram_data_in_bus_10;
output 	wraddress_b_bus_1;
output 	wraddress_b_bus_3;
output 	wraddress_b_bus_5;
output 	rdaddress_b_bus_1;
output 	rdaddress_b_bus_3;
output 	rdaddress_b_bus_5;
output 	a_ram_data_in_bus_10;
output 	wraddress_a_bus_1;
output 	wraddress_a_bus_3;
output 	wraddress_a_bus_5;
output 	rdaddress_a_bus_1;
output 	rdaddress_a_bus_3;
output 	rdaddress_a_bus_5;
output 	b_ram_data_in_bus_62;
output 	a_ram_data_in_bus_62;
output 	b_ram_data_in_bus_46;
output 	a_ram_data_in_bus_46;
output 	b_ram_data_in_bus_30;
output 	a_ram_data_in_bus_30;
output 	b_ram_data_in_bus_14;
output 	a_ram_data_in_bus_14;
output 	b_ram_data_in_bus_60;
output 	a_ram_data_in_bus_60;
output 	b_ram_data_in_bus_44;
output 	a_ram_data_in_bus_44;
output 	b_ram_data_in_bus_28;
output 	a_ram_data_in_bus_28;
output 	b_ram_data_in_bus_12;
output 	a_ram_data_in_bus_12;
output 	b_ram_data_in_bus_59;
output 	a_ram_data_in_bus_59;
output 	b_ram_data_in_bus_43;
output 	a_ram_data_in_bus_43;
output 	b_ram_data_in_bus_27;
output 	a_ram_data_in_bus_27;
output 	b_ram_data_in_bus_11;
output 	a_ram_data_in_bus_11;
output 	b_ram_data_in_bus_61;
output 	a_ram_data_in_bus_61;
output 	b_ram_data_in_bus_45;
output 	a_ram_data_in_bus_45;
output 	b_ram_data_in_bus_29;
output 	a_ram_data_in_bus_29;
output 	b_ram_data_in_bus_13;
output 	a_ram_data_in_bus_13;
output 	b_ram_data_in_bus_57;
output 	a_ram_data_in_bus_57;
output 	b_ram_data_in_bus_41;
output 	a_ram_data_in_bus_41;
output 	b_ram_data_in_bus_25;
output 	a_ram_data_in_bus_25;
output 	b_ram_data_in_bus_9;
output 	a_ram_data_in_bus_9;
output 	b_ram_data_in_bus_56;
output 	a_ram_data_in_bus_56;
output 	b_ram_data_in_bus_40;
output 	a_ram_data_in_bus_40;
output 	b_ram_data_in_bus_24;
output 	a_ram_data_in_bus_24;
output 	b_ram_data_in_bus_8;
output 	a_ram_data_in_bus_8;
output 	b_ram_data_in_bus_63;
output 	a_ram_data_in_bus_63;
output 	b_ram_data_in_bus_47;
output 	a_ram_data_in_bus_47;
output 	b_ram_data_in_bus_31;
output 	a_ram_data_in_bus_31;
output 	b_ram_data_in_bus_15;
output 	a_ram_data_in_bus_15;
output 	b_ram_data_in_bus_55;
output 	a_ram_data_in_bus_55;
output 	b_ram_data_in_bus_39;
output 	a_ram_data_in_bus_39;
output 	b_ram_data_in_bus_23;
output 	a_ram_data_in_bus_23;
output 	b_ram_data_in_bus_7;
output 	a_ram_data_in_bus_7;
output 	b_ram_data_in_bus_51;
output 	a_ram_data_in_bus_51;
output 	b_ram_data_in_bus_35;
output 	a_ram_data_in_bus_35;
output 	b_ram_data_in_bus_19;
output 	a_ram_data_in_bus_19;
output 	b_ram_data_in_bus_3;
output 	a_ram_data_in_bus_3;
output 	b_ram_data_in_bus_53;
output 	a_ram_data_in_bus_53;
output 	b_ram_data_in_bus_37;
output 	a_ram_data_in_bus_37;
output 	b_ram_data_in_bus_21;
output 	a_ram_data_in_bus_21;
output 	b_ram_data_in_bus_5;
output 	a_ram_data_in_bus_5;
output 	b_ram_data_in_bus_52;
output 	a_ram_data_in_bus_52;
output 	b_ram_data_in_bus_36;
output 	a_ram_data_in_bus_36;
output 	b_ram_data_in_bus_20;
output 	a_ram_data_in_bus_20;
output 	b_ram_data_in_bus_4;
output 	a_ram_data_in_bus_4;
output 	b_ram_data_in_bus_54;
output 	a_ram_data_in_bus_54;
output 	b_ram_data_in_bus_38;
output 	a_ram_data_in_bus_38;
output 	b_ram_data_in_bus_22;
output 	a_ram_data_in_bus_22;
output 	b_ram_data_in_bus_6;
output 	a_ram_data_in_bus_6;
output 	b_ram_data_in_bus_50;
output 	a_ram_data_in_bus_50;
output 	b_ram_data_in_bus_34;
output 	a_ram_data_in_bus_34;
output 	b_ram_data_in_bus_18;
output 	a_ram_data_in_bus_18;
output 	b_ram_data_in_bus_2;
output 	a_ram_data_in_bus_2;
output 	b_ram_data_in_bus_49;
output 	a_ram_data_in_bus_49;
output 	b_ram_data_in_bus_33;
output 	a_ram_data_in_bus_33;
output 	b_ram_data_in_bus_17;
output 	a_ram_data_in_bus_17;
output 	b_ram_data_in_bus_1;
output 	a_ram_data_in_bus_1;
output 	b_ram_data_in_bus_48;
output 	a_ram_data_in_bus_48;
output 	b_ram_data_in_bus_32;
output 	a_ram_data_in_bus_32;
output 	b_ram_data_in_bus_16;
output 	a_ram_data_in_bus_16;
output 	b_ram_data_in_bus_0;
output 	a_ram_data_in_bus_0;
input 	ram_a_not_b_vec_1;
input 	data_in_r_2;
input 	wr_address_i_int_0;
input 	wr_address_i_int_1;
input 	wr_address_i_int_2;
input 	wr_address_i_int_3;
input 	wr_address_i_int_4;
input 	wr_address_i_int_5;
input 	wr_address_i_int_6;
input 	ram_a_not_b_vec_7;
input 	ram_in_reg_0_02;
input 	ram_in_reg_1_02;
input 	ram_in_reg_2_02;
input 	ram_in_reg_3_02;
input 	ram_in_reg_4_02;
input 	ram_in_reg_5_02;
input 	tdl_arr_6_1;
input 	ram_in_reg_0_12;
input 	ram_in_reg_1_12;
input 	ram_in_reg_2_12;
input 	ram_in_reg_3_12;
input 	ram_in_reg_4_12;
input 	ram_in_reg_5_12;
input 	ram_in_reg_1_22;
input 	ram_in_reg_3_22;
input 	ram_in_reg_5_22;
input 	ram_in_reg_1_32;
input 	ram_in_reg_3_32;
input 	ram_in_reg_5_32;
input 	data_in_r_6;
input 	data_in_r_4;
input 	data_in_r_3;
input 	data_in_r_5;
input 	data_in_r_1;
input 	data_in_r_0;
input 	data_in_r_7;
input 	data_in_i_7;
input 	data_in_i_3;
input 	data_in_i_5;
input 	data_in_i_4;
input 	data_in_i_6;
input 	data_in_i_2;
input 	data_in_i_1;
input 	data_in_i_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ram_data_out0~0_combout ;
wire \ram_data_out1~0_combout ;
wire \ram_data_out2~0_combout ;
wire \ram_data_out3~0_combout ;
wire \ram_data_out0~1_combout ;
wire \ram_data_out1~1_combout ;
wire \ram_data_out2~1_combout ;
wire \ram_data_out3~1_combout ;
wire \ram_data_out0~2_combout ;
wire \ram_data_out1~2_combout ;
wire \ram_data_out2~2_combout ;
wire \ram_data_out3~2_combout ;
wire \ram_data_out0~3_combout ;
wire \ram_data_out1~3_combout ;
wire \ram_data_out2~3_combout ;
wire \ram_data_out3~3_combout ;
wire \ram_data_out0~4_combout ;
wire \ram_data_out1~4_combout ;
wire \ram_data_out2~4_combout ;
wire \ram_data_out3~4_combout ;
wire \ram_data_out0~5_combout ;
wire \ram_data_out1~5_combout ;
wire \ram_data_out2~5_combout ;
wire \ram_data_out3~5_combout ;
wire \ram_data_out0~6_combout ;
wire \ram_data_out1~6_combout ;
wire \ram_data_out2~6_combout ;
wire \ram_data_out3~6_combout ;
wire \ram_data_out0~7_combout ;
wire \ram_data_out1~7_combout ;
wire \ram_data_out2~7_combout ;
wire \ram_data_out3~7_combout ;
wire \ram_data_out0~8_combout ;
wire \ram_data_out1~8_combout ;
wire \ram_data_out2~8_combout ;
wire \ram_data_out3~8_combout ;
wire \ram_data_out0~9_combout ;
wire \ram_data_out1~9_combout ;
wire \ram_data_out2~9_combout ;
wire \ram_data_out3~9_combout ;
wire \ram_data_out0~10_combout ;
wire \ram_data_out1~10_combout ;
wire \ram_data_out2~10_combout ;
wire \ram_data_out3~10_combout ;
wire \ram_data_out0~11_combout ;
wire \ram_data_out1~11_combout ;
wire \ram_data_out2~11_combout ;
wire \ram_data_out3~11_combout ;
wire \ram_data_out0~12_combout ;
wire \ram_data_out1~12_combout ;
wire \ram_data_out2~12_combout ;
wire \ram_data_out3~12_combout ;
wire \ram_data_out0~13_combout ;
wire \ram_data_out1~13_combout ;
wire \ram_data_out2~13_combout ;
wire \ram_data_out3~13_combout ;
wire \ram_data_out0~14_combout ;
wire \ram_data_out1~14_combout ;
wire \ram_data_out2~14_combout ;
wire \ram_data_out3~14_combout ;
wire \ram_data_out0~15_combout ;
wire \ram_data_out1~15_combout ;
wire \ram_data_out2~15_combout ;
wire \ram_data_out3~15_combout ;
wire \b_ram_data_in_bus~0_combout ;
wire \wraddress_b_bus~0_combout ;
wire \wraddress_b_bus~1_combout ;
wire \wraddress_b_bus~2_combout ;
wire \wraddress_b_bus~3_combout ;
wire \wraddress_b_bus~4_combout ;
wire \wraddress_b_bus~5_combout ;
wire \wraddress_b_bus~6_combout ;
wire \rdaddress_b_bus~0_combout ;
wire \rdaddress_b_bus~1_combout ;
wire \rdaddress_b_bus~2_combout ;
wire \rdaddress_b_bus~3_combout ;
wire \rdaddress_b_bus~4_combout ;
wire \rdaddress_b_bus~5_combout ;
wire \rdaddress_b_bus~6_combout ;
wire \a_ram_data_in_bus~0_combout ;
wire \wraddress_a_bus~0_combout ;
wire \wraddress_a_bus~1_combout ;
wire \wraddress_a_bus~2_combout ;
wire \wraddress_a_bus~3_combout ;
wire \wraddress_a_bus~4_combout ;
wire \wraddress_a_bus~5_combout ;
wire \wraddress_a_bus~6_combout ;
wire \rdaddress_a_bus~0_combout ;
wire \rdaddress_a_bus~1_combout ;
wire \rdaddress_a_bus~2_combout ;
wire \rdaddress_a_bus~3_combout ;
wire \rdaddress_a_bus~4_combout ;
wire \rdaddress_a_bus~5_combout ;
wire \rdaddress_a_bus~6_combout ;
wire \b_ram_data_in_bus~1_combout ;
wire \wraddress_b_bus~7_combout ;
wire \wraddress_b_bus~8_combout ;
wire \wraddress_b_bus~9_combout ;
wire \wraddress_b_bus~10_combout ;
wire \wraddress_b_bus~11_combout ;
wire \wraddress_b_bus~12_combout ;
wire \rdaddress_b_bus~7_combout ;
wire \rdaddress_b_bus~8_combout ;
wire \rdaddress_b_bus~9_combout ;
wire \rdaddress_b_bus~10_combout ;
wire \rdaddress_b_bus~11_combout ;
wire \rdaddress_b_bus~12_combout ;
wire \a_ram_data_in_bus~1_combout ;
wire \wraddress_a_bus~7_combout ;
wire \wraddress_a_bus~8_combout ;
wire \wraddress_a_bus~9_combout ;
wire \wraddress_a_bus~10_combout ;
wire \wraddress_a_bus~11_combout ;
wire \wraddress_a_bus~12_combout ;
wire \rdaddress_a_bus~7_combout ;
wire \rdaddress_a_bus~8_combout ;
wire \rdaddress_a_bus~9_combout ;
wire \rdaddress_a_bus~10_combout ;
wire \rdaddress_a_bus~11_combout ;
wire \rdaddress_a_bus~12_combout ;
wire \b_ram_data_in_bus~2_combout ;
wire \wraddress_b_bus~13_combout ;
wire \wraddress_b_bus~14_combout ;
wire \wraddress_b_bus~15_combout ;
wire \rdaddress_b_bus~13_combout ;
wire \rdaddress_b_bus~14_combout ;
wire \rdaddress_b_bus~15_combout ;
wire \a_ram_data_in_bus~2_combout ;
wire \wraddress_a_bus~13_combout ;
wire \wraddress_a_bus~14_combout ;
wire \wraddress_a_bus~15_combout ;
wire \rdaddress_a_bus~13_combout ;
wire \rdaddress_a_bus~14_combout ;
wire \rdaddress_a_bus~15_combout ;
wire \b_ram_data_in_bus~3_combout ;
wire \wraddress_b_bus~16_combout ;
wire \wraddress_b_bus~17_combout ;
wire \wraddress_b_bus~18_combout ;
wire \rdaddress_b_bus~16_combout ;
wire \rdaddress_b_bus~17_combout ;
wire \rdaddress_b_bus~18_combout ;
wire \a_ram_data_in_bus~3_combout ;
wire \wraddress_a_bus~16_combout ;
wire \wraddress_a_bus~17_combout ;
wire \wraddress_a_bus~18_combout ;
wire \rdaddress_a_bus~16_combout ;
wire \rdaddress_a_bus~17_combout ;
wire \rdaddress_a_bus~18_combout ;
wire \b_ram_data_in_bus~4_combout ;
wire \a_ram_data_in_bus~4_combout ;
wire \b_ram_data_in_bus~5_combout ;
wire \a_ram_data_in_bus~5_combout ;
wire \b_ram_data_in_bus~6_combout ;
wire \a_ram_data_in_bus~6_combout ;
wire \b_ram_data_in_bus~7_combout ;
wire \a_ram_data_in_bus~7_combout ;
wire \b_ram_data_in_bus~8_combout ;
wire \a_ram_data_in_bus~8_combout ;
wire \b_ram_data_in_bus~9_combout ;
wire \a_ram_data_in_bus~9_combout ;
wire \b_ram_data_in_bus~10_combout ;
wire \a_ram_data_in_bus~10_combout ;
wire \b_ram_data_in_bus~11_combout ;
wire \a_ram_data_in_bus~11_combout ;
wire \b_ram_data_in_bus~12_combout ;
wire \a_ram_data_in_bus~12_combout ;
wire \b_ram_data_in_bus~13_combout ;
wire \a_ram_data_in_bus~13_combout ;
wire \b_ram_data_in_bus~14_combout ;
wire \a_ram_data_in_bus~14_combout ;
wire \b_ram_data_in_bus~15_combout ;
wire \a_ram_data_in_bus~15_combout ;
wire \b_ram_data_in_bus~16_combout ;
wire \a_ram_data_in_bus~16_combout ;
wire \b_ram_data_in_bus~17_combout ;
wire \a_ram_data_in_bus~17_combout ;
wire \b_ram_data_in_bus~18_combout ;
wire \a_ram_data_in_bus~18_combout ;
wire \b_ram_data_in_bus~19_combout ;
wire \a_ram_data_in_bus~19_combout ;
wire \b_ram_data_in_bus~20_combout ;
wire \a_ram_data_in_bus~20_combout ;
wire \b_ram_data_in_bus~21_combout ;
wire \a_ram_data_in_bus~21_combout ;
wire \b_ram_data_in_bus~22_combout ;
wire \a_ram_data_in_bus~22_combout ;
wire \b_ram_data_in_bus~23_combout ;
wire \a_ram_data_in_bus~23_combout ;
wire \b_ram_data_in_bus~24_combout ;
wire \a_ram_data_in_bus~24_combout ;
wire \b_ram_data_in_bus~25_combout ;
wire \a_ram_data_in_bus~25_combout ;
wire \b_ram_data_in_bus~26_combout ;
wire \a_ram_data_in_bus~26_combout ;
wire \b_ram_data_in_bus~27_combout ;
wire \a_ram_data_in_bus~27_combout ;
wire \b_ram_data_in_bus~28_combout ;
wire \a_ram_data_in_bus~28_combout ;
wire \b_ram_data_in_bus~29_combout ;
wire \a_ram_data_in_bus~29_combout ;
wire \b_ram_data_in_bus~30_combout ;
wire \a_ram_data_in_bus~30_combout ;
wire \b_ram_data_in_bus~31_combout ;
wire \a_ram_data_in_bus~31_combout ;
wire \b_ram_data_in_bus~32_combout ;
wire \a_ram_data_in_bus~32_combout ;
wire \b_ram_data_in_bus~33_combout ;
wire \a_ram_data_in_bus~33_combout ;
wire \b_ram_data_in_bus~34_combout ;
wire \a_ram_data_in_bus~34_combout ;
wire \b_ram_data_in_bus~35_combout ;
wire \a_ram_data_in_bus~35_combout ;
wire \b_ram_data_in_bus~36_combout ;
wire \a_ram_data_in_bus~36_combout ;
wire \b_ram_data_in_bus~37_combout ;
wire \a_ram_data_in_bus~37_combout ;
wire \b_ram_data_in_bus~38_combout ;
wire \a_ram_data_in_bus~38_combout ;
wire \b_ram_data_in_bus~39_combout ;
wire \a_ram_data_in_bus~39_combout ;
wire \b_ram_data_in_bus~40_combout ;
wire \a_ram_data_in_bus~40_combout ;
wire \b_ram_data_in_bus~41_combout ;
wire \a_ram_data_in_bus~41_combout ;
wire \b_ram_data_in_bus~42_combout ;
wire \a_ram_data_in_bus~42_combout ;
wire \b_ram_data_in_bus~43_combout ;
wire \a_ram_data_in_bus~43_combout ;
wire \b_ram_data_in_bus~44_combout ;
wire \a_ram_data_in_bus~44_combout ;
wire \b_ram_data_in_bus~45_combout ;
wire \a_ram_data_in_bus~45_combout ;
wire \b_ram_data_in_bus~46_combout ;
wire \a_ram_data_in_bus~46_combout ;
wire \b_ram_data_in_bus~47_combout ;
wire \a_ram_data_in_bus~47_combout ;
wire \b_ram_data_in_bus~48_combout ;
wire \a_ram_data_in_bus~48_combout ;
wire \b_ram_data_in_bus~49_combout ;
wire \a_ram_data_in_bus~49_combout ;
wire \b_ram_data_in_bus~50_combout ;
wire \a_ram_data_in_bus~50_combout ;
wire \b_ram_data_in_bus~51_combout ;
wire \a_ram_data_in_bus~51_combout ;
wire \b_ram_data_in_bus~52_combout ;
wire \a_ram_data_in_bus~52_combout ;
wire \b_ram_data_in_bus~53_combout ;
wire \a_ram_data_in_bus~53_combout ;
wire \b_ram_data_in_bus~54_combout ;
wire \a_ram_data_in_bus~54_combout ;
wire \b_ram_data_in_bus~55_combout ;
wire \a_ram_data_in_bus~55_combout ;
wire \b_ram_data_in_bus~56_combout ;
wire \a_ram_data_in_bus~56_combout ;
wire \b_ram_data_in_bus~57_combout ;
wire \a_ram_data_in_bus~57_combout ;
wire \b_ram_data_in_bus~58_combout ;
wire \a_ram_data_in_bus~58_combout ;
wire \b_ram_data_in_bus~59_combout ;
wire \a_ram_data_in_bus~59_combout ;
wire \b_ram_data_in_bus~60_combout ;
wire \a_ram_data_in_bus~60_combout ;
wire \b_ram_data_in_bus~61_combout ;
wire \a_ram_data_in_bus~61_combout ;
wire \b_ram_data_in_bus~62_combout ;
wire \a_ram_data_in_bus~62_combout ;
wire \b_ram_data_in_bus~63_combout ;
wire \a_ram_data_in_bus~63_combout ;


dffeas \ram_data_out0[10] (
	.clk(clk),
	.d(\ram_data_out0~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out0_10),
	.prn(vcc));
defparam \ram_data_out0[10] .is_wysiwyg = "true";
defparam \ram_data_out0[10] .power_up = "low";

dffeas \ram_data_out1[10] (
	.clk(clk),
	.d(\ram_data_out1~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out1_10),
	.prn(vcc));
defparam \ram_data_out1[10] .is_wysiwyg = "true";
defparam \ram_data_out1[10] .power_up = "low";

dffeas \ram_data_out2[10] (
	.clk(clk),
	.d(\ram_data_out2~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out2_10),
	.prn(vcc));
defparam \ram_data_out2[10] .is_wysiwyg = "true";
defparam \ram_data_out2[10] .power_up = "low";

dffeas \ram_data_out3[10] (
	.clk(clk),
	.d(\ram_data_out3~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out3_10),
	.prn(vcc));
defparam \ram_data_out3[10] .is_wysiwyg = "true";
defparam \ram_data_out3[10] .power_up = "low";

dffeas \ram_data_out0[14] (
	.clk(clk),
	.d(\ram_data_out0~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out0_14),
	.prn(vcc));
defparam \ram_data_out0[14] .is_wysiwyg = "true";
defparam \ram_data_out0[14] .power_up = "low";

dffeas \ram_data_out1[14] (
	.clk(clk),
	.d(\ram_data_out1~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out1_14),
	.prn(vcc));
defparam \ram_data_out1[14] .is_wysiwyg = "true";
defparam \ram_data_out1[14] .power_up = "low";

dffeas \ram_data_out2[14] (
	.clk(clk),
	.d(\ram_data_out2~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out2_14),
	.prn(vcc));
defparam \ram_data_out2[14] .is_wysiwyg = "true";
defparam \ram_data_out2[14] .power_up = "low";

dffeas \ram_data_out3[14] (
	.clk(clk),
	.d(\ram_data_out3~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out3_14),
	.prn(vcc));
defparam \ram_data_out3[14] .is_wysiwyg = "true";
defparam \ram_data_out3[14] .power_up = "low";

dffeas \ram_data_out0[12] (
	.clk(clk),
	.d(\ram_data_out0~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out0_12),
	.prn(vcc));
defparam \ram_data_out0[12] .is_wysiwyg = "true";
defparam \ram_data_out0[12] .power_up = "low";

dffeas \ram_data_out1[12] (
	.clk(clk),
	.d(\ram_data_out1~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out1_12),
	.prn(vcc));
defparam \ram_data_out1[12] .is_wysiwyg = "true";
defparam \ram_data_out1[12] .power_up = "low";

dffeas \ram_data_out2[12] (
	.clk(clk),
	.d(\ram_data_out2~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out2_12),
	.prn(vcc));
defparam \ram_data_out2[12] .is_wysiwyg = "true";
defparam \ram_data_out2[12] .power_up = "low";

dffeas \ram_data_out3[12] (
	.clk(clk),
	.d(\ram_data_out3~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out3_12),
	.prn(vcc));
defparam \ram_data_out3[12] .is_wysiwyg = "true";
defparam \ram_data_out3[12] .power_up = "low";

dffeas \ram_data_out0[11] (
	.clk(clk),
	.d(\ram_data_out0~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out0_11),
	.prn(vcc));
defparam \ram_data_out0[11] .is_wysiwyg = "true";
defparam \ram_data_out0[11] .power_up = "low";

dffeas \ram_data_out1[11] (
	.clk(clk),
	.d(\ram_data_out1~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out1_11),
	.prn(vcc));
defparam \ram_data_out1[11] .is_wysiwyg = "true";
defparam \ram_data_out1[11] .power_up = "low";

dffeas \ram_data_out2[11] (
	.clk(clk),
	.d(\ram_data_out2~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out2_11),
	.prn(vcc));
defparam \ram_data_out2[11] .is_wysiwyg = "true";
defparam \ram_data_out2[11] .power_up = "low";

dffeas \ram_data_out3[11] (
	.clk(clk),
	.d(\ram_data_out3~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out3_11),
	.prn(vcc));
defparam \ram_data_out3[11] .is_wysiwyg = "true";
defparam \ram_data_out3[11] .power_up = "low";

dffeas \ram_data_out0[13] (
	.clk(clk),
	.d(\ram_data_out0~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out0_13),
	.prn(vcc));
defparam \ram_data_out0[13] .is_wysiwyg = "true";
defparam \ram_data_out0[13] .power_up = "low";

dffeas \ram_data_out1[13] (
	.clk(clk),
	.d(\ram_data_out1~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out1_13),
	.prn(vcc));
defparam \ram_data_out1[13] .is_wysiwyg = "true";
defparam \ram_data_out1[13] .power_up = "low";

dffeas \ram_data_out2[13] (
	.clk(clk),
	.d(\ram_data_out2~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out2_13),
	.prn(vcc));
defparam \ram_data_out2[13] .is_wysiwyg = "true";
defparam \ram_data_out2[13] .power_up = "low";

dffeas \ram_data_out3[13] (
	.clk(clk),
	.d(\ram_data_out3~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out3_13),
	.prn(vcc));
defparam \ram_data_out3[13] .is_wysiwyg = "true";
defparam \ram_data_out3[13] .power_up = "low";

dffeas \ram_data_out0[9] (
	.clk(clk),
	.d(\ram_data_out0~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out0_9),
	.prn(vcc));
defparam \ram_data_out0[9] .is_wysiwyg = "true";
defparam \ram_data_out0[9] .power_up = "low";

dffeas \ram_data_out1[9] (
	.clk(clk),
	.d(\ram_data_out1~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out1_9),
	.prn(vcc));
defparam \ram_data_out1[9] .is_wysiwyg = "true";
defparam \ram_data_out1[9] .power_up = "low";

dffeas \ram_data_out2[9] (
	.clk(clk),
	.d(\ram_data_out2~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out2_9),
	.prn(vcc));
defparam \ram_data_out2[9] .is_wysiwyg = "true";
defparam \ram_data_out2[9] .power_up = "low";

dffeas \ram_data_out3[9] (
	.clk(clk),
	.d(\ram_data_out3~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out3_9),
	.prn(vcc));
defparam \ram_data_out3[9] .is_wysiwyg = "true";
defparam \ram_data_out3[9] .power_up = "low";

dffeas \ram_data_out0[8] (
	.clk(clk),
	.d(\ram_data_out0~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out0_8),
	.prn(vcc));
defparam \ram_data_out0[8] .is_wysiwyg = "true";
defparam \ram_data_out0[8] .power_up = "low";

dffeas \ram_data_out1[8] (
	.clk(clk),
	.d(\ram_data_out1~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out1_8),
	.prn(vcc));
defparam \ram_data_out1[8] .is_wysiwyg = "true";
defparam \ram_data_out1[8] .power_up = "low";

dffeas \ram_data_out2[8] (
	.clk(clk),
	.d(\ram_data_out2~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out2_8),
	.prn(vcc));
defparam \ram_data_out2[8] .is_wysiwyg = "true";
defparam \ram_data_out2[8] .power_up = "low";

dffeas \ram_data_out3[8] (
	.clk(clk),
	.d(\ram_data_out3~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out3_8),
	.prn(vcc));
defparam \ram_data_out3[8] .is_wysiwyg = "true";
defparam \ram_data_out3[8] .power_up = "low";

dffeas \ram_data_out0[15] (
	.clk(clk),
	.d(\ram_data_out0~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out0_15),
	.prn(vcc));
defparam \ram_data_out0[15] .is_wysiwyg = "true";
defparam \ram_data_out0[15] .power_up = "low";

dffeas \ram_data_out1[15] (
	.clk(clk),
	.d(\ram_data_out1~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out1_15),
	.prn(vcc));
defparam \ram_data_out1[15] .is_wysiwyg = "true";
defparam \ram_data_out1[15] .power_up = "low";

dffeas \ram_data_out2[15] (
	.clk(clk),
	.d(\ram_data_out2~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out2_15),
	.prn(vcc));
defparam \ram_data_out2[15] .is_wysiwyg = "true";
defparam \ram_data_out2[15] .power_up = "low";

dffeas \ram_data_out3[15] (
	.clk(clk),
	.d(\ram_data_out3~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out3_15),
	.prn(vcc));
defparam \ram_data_out3[15] .is_wysiwyg = "true";
defparam \ram_data_out3[15] .power_up = "low";

dffeas \ram_data_out0[7] (
	.clk(clk),
	.d(\ram_data_out0~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out0_7),
	.prn(vcc));
defparam \ram_data_out0[7] .is_wysiwyg = "true";
defparam \ram_data_out0[7] .power_up = "low";

dffeas \ram_data_out1[7] (
	.clk(clk),
	.d(\ram_data_out1~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out1_7),
	.prn(vcc));
defparam \ram_data_out1[7] .is_wysiwyg = "true";
defparam \ram_data_out1[7] .power_up = "low";

dffeas \ram_data_out2[7] (
	.clk(clk),
	.d(\ram_data_out2~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out2_7),
	.prn(vcc));
defparam \ram_data_out2[7] .is_wysiwyg = "true";
defparam \ram_data_out2[7] .power_up = "low";

dffeas \ram_data_out3[7] (
	.clk(clk),
	.d(\ram_data_out3~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out3_7),
	.prn(vcc));
defparam \ram_data_out3[7] .is_wysiwyg = "true";
defparam \ram_data_out3[7] .power_up = "low";

dffeas \ram_data_out0[3] (
	.clk(clk),
	.d(\ram_data_out0~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out0_3),
	.prn(vcc));
defparam \ram_data_out0[3] .is_wysiwyg = "true";
defparam \ram_data_out0[3] .power_up = "low";

dffeas \ram_data_out1[3] (
	.clk(clk),
	.d(\ram_data_out1~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out1_3),
	.prn(vcc));
defparam \ram_data_out1[3] .is_wysiwyg = "true";
defparam \ram_data_out1[3] .power_up = "low";

dffeas \ram_data_out2[3] (
	.clk(clk),
	.d(\ram_data_out2~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out2_3),
	.prn(vcc));
defparam \ram_data_out2[3] .is_wysiwyg = "true";
defparam \ram_data_out2[3] .power_up = "low";

dffeas \ram_data_out3[3] (
	.clk(clk),
	.d(\ram_data_out3~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out3_3),
	.prn(vcc));
defparam \ram_data_out3[3] .is_wysiwyg = "true";
defparam \ram_data_out3[3] .power_up = "low";

dffeas \ram_data_out0[5] (
	.clk(clk),
	.d(\ram_data_out0~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out0_5),
	.prn(vcc));
defparam \ram_data_out0[5] .is_wysiwyg = "true";
defparam \ram_data_out0[5] .power_up = "low";

dffeas \ram_data_out1[5] (
	.clk(clk),
	.d(\ram_data_out1~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out1_5),
	.prn(vcc));
defparam \ram_data_out1[5] .is_wysiwyg = "true";
defparam \ram_data_out1[5] .power_up = "low";

dffeas \ram_data_out2[5] (
	.clk(clk),
	.d(\ram_data_out2~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out2_5),
	.prn(vcc));
defparam \ram_data_out2[5] .is_wysiwyg = "true";
defparam \ram_data_out2[5] .power_up = "low";

dffeas \ram_data_out3[5] (
	.clk(clk),
	.d(\ram_data_out3~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out3_5),
	.prn(vcc));
defparam \ram_data_out3[5] .is_wysiwyg = "true";
defparam \ram_data_out3[5] .power_up = "low";

dffeas \ram_data_out0[4] (
	.clk(clk),
	.d(\ram_data_out0~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out0_4),
	.prn(vcc));
defparam \ram_data_out0[4] .is_wysiwyg = "true";
defparam \ram_data_out0[4] .power_up = "low";

dffeas \ram_data_out1[4] (
	.clk(clk),
	.d(\ram_data_out1~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out1_4),
	.prn(vcc));
defparam \ram_data_out1[4] .is_wysiwyg = "true";
defparam \ram_data_out1[4] .power_up = "low";

dffeas \ram_data_out2[4] (
	.clk(clk),
	.d(\ram_data_out2~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out2_4),
	.prn(vcc));
defparam \ram_data_out2[4] .is_wysiwyg = "true";
defparam \ram_data_out2[4] .power_up = "low";

dffeas \ram_data_out3[4] (
	.clk(clk),
	.d(\ram_data_out3~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out3_4),
	.prn(vcc));
defparam \ram_data_out3[4] .is_wysiwyg = "true";
defparam \ram_data_out3[4] .power_up = "low";

dffeas \ram_data_out0[6] (
	.clk(clk),
	.d(\ram_data_out0~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out0_6),
	.prn(vcc));
defparam \ram_data_out0[6] .is_wysiwyg = "true";
defparam \ram_data_out0[6] .power_up = "low";

dffeas \ram_data_out1[6] (
	.clk(clk),
	.d(\ram_data_out1~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out1_6),
	.prn(vcc));
defparam \ram_data_out1[6] .is_wysiwyg = "true";
defparam \ram_data_out1[6] .power_up = "low";

dffeas \ram_data_out2[6] (
	.clk(clk),
	.d(\ram_data_out2~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out2_6),
	.prn(vcc));
defparam \ram_data_out2[6] .is_wysiwyg = "true";
defparam \ram_data_out2[6] .power_up = "low";

dffeas \ram_data_out3[6] (
	.clk(clk),
	.d(\ram_data_out3~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out3_6),
	.prn(vcc));
defparam \ram_data_out3[6] .is_wysiwyg = "true";
defparam \ram_data_out3[6] .power_up = "low";

dffeas \ram_data_out0[2] (
	.clk(clk),
	.d(\ram_data_out0~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out0_2),
	.prn(vcc));
defparam \ram_data_out0[2] .is_wysiwyg = "true";
defparam \ram_data_out0[2] .power_up = "low";

dffeas \ram_data_out1[2] (
	.clk(clk),
	.d(\ram_data_out1~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out1_2),
	.prn(vcc));
defparam \ram_data_out1[2] .is_wysiwyg = "true";
defparam \ram_data_out1[2] .power_up = "low";

dffeas \ram_data_out2[2] (
	.clk(clk),
	.d(\ram_data_out2~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out2_2),
	.prn(vcc));
defparam \ram_data_out2[2] .is_wysiwyg = "true";
defparam \ram_data_out2[2] .power_up = "low";

dffeas \ram_data_out3[2] (
	.clk(clk),
	.d(\ram_data_out3~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out3_2),
	.prn(vcc));
defparam \ram_data_out3[2] .is_wysiwyg = "true";
defparam \ram_data_out3[2] .power_up = "low";

dffeas \ram_data_out0[1] (
	.clk(clk),
	.d(\ram_data_out0~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out0_1),
	.prn(vcc));
defparam \ram_data_out0[1] .is_wysiwyg = "true";
defparam \ram_data_out0[1] .power_up = "low";

dffeas \ram_data_out1[1] (
	.clk(clk),
	.d(\ram_data_out1~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out1_1),
	.prn(vcc));
defparam \ram_data_out1[1] .is_wysiwyg = "true";
defparam \ram_data_out1[1] .power_up = "low";

dffeas \ram_data_out2[1] (
	.clk(clk),
	.d(\ram_data_out2~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out2_1),
	.prn(vcc));
defparam \ram_data_out2[1] .is_wysiwyg = "true";
defparam \ram_data_out2[1] .power_up = "low";

dffeas \ram_data_out3[1] (
	.clk(clk),
	.d(\ram_data_out3~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out3_1),
	.prn(vcc));
defparam \ram_data_out3[1] .is_wysiwyg = "true";
defparam \ram_data_out3[1] .power_up = "low";

dffeas \ram_data_out0[0] (
	.clk(clk),
	.d(\ram_data_out0~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out0_0),
	.prn(vcc));
defparam \ram_data_out0[0] .is_wysiwyg = "true";
defparam \ram_data_out0[0] .power_up = "low";

dffeas \ram_data_out1[0] (
	.clk(clk),
	.d(\ram_data_out1~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out1_0),
	.prn(vcc));
defparam \ram_data_out1[0] .is_wysiwyg = "true";
defparam \ram_data_out1[0] .power_up = "low";

dffeas \ram_data_out2[0] (
	.clk(clk),
	.d(\ram_data_out2~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out2_0),
	.prn(vcc));
defparam \ram_data_out2[0] .is_wysiwyg = "true";
defparam \ram_data_out2[0] .power_up = "low";

dffeas \ram_data_out3[0] (
	.clk(clk),
	.d(\ram_data_out3~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out3_0),
	.prn(vcc));
defparam \ram_data_out3[0] .is_wysiwyg = "true";
defparam \ram_data_out3[0] .power_up = "low";

dffeas \b_ram_data_in_bus[58] (
	.clk(clk),
	.d(\b_ram_data_in_bus~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_58),
	.prn(vcc));
defparam \b_ram_data_in_bus[58] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[58] .power_up = "low";

dffeas \wraddress_b_bus[21] (
	.clk(clk),
	.d(\wraddress_b_bus~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_b_bus_21),
	.prn(vcc));
defparam \wraddress_b_bus[21] .is_wysiwyg = "true";
defparam \wraddress_b_bus[21] .power_up = "low";

dffeas \wraddress_b_bus[22] (
	.clk(clk),
	.d(\wraddress_b_bus~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_b_bus_22),
	.prn(vcc));
defparam \wraddress_b_bus[22] .is_wysiwyg = "true";
defparam \wraddress_b_bus[22] .power_up = "low";

dffeas \wraddress_b_bus[23] (
	.clk(clk),
	.d(\wraddress_b_bus~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_b_bus_23),
	.prn(vcc));
defparam \wraddress_b_bus[23] .is_wysiwyg = "true";
defparam \wraddress_b_bus[23] .power_up = "low";

dffeas \wraddress_b_bus[24] (
	.clk(clk),
	.d(\wraddress_b_bus~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_b_bus_24),
	.prn(vcc));
defparam \wraddress_b_bus[24] .is_wysiwyg = "true";
defparam \wraddress_b_bus[24] .power_up = "low";

dffeas \wraddress_b_bus[11] (
	.clk(clk),
	.d(\wraddress_b_bus~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_b_bus_11),
	.prn(vcc));
defparam \wraddress_b_bus[11] .is_wysiwyg = "true";
defparam \wraddress_b_bus[11] .power_up = "low";

dffeas \wraddress_b_bus[26] (
	.clk(clk),
	.d(\wraddress_b_bus~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_b_bus_26),
	.prn(vcc));
defparam \wraddress_b_bus[26] .is_wysiwyg = "true";
defparam \wraddress_b_bus[26] .power_up = "low";

dffeas \wraddress_b_bus[13] (
	.clk(clk),
	.d(\wraddress_b_bus~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_b_bus_13),
	.prn(vcc));
defparam \wraddress_b_bus[13] .is_wysiwyg = "true";
defparam \wraddress_b_bus[13] .power_up = "low";

dffeas \rdaddress_b_bus[21] (
	.clk(clk),
	.d(\rdaddress_b_bus~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_b_bus_21),
	.prn(vcc));
defparam \rdaddress_b_bus[21] .is_wysiwyg = "true";
defparam \rdaddress_b_bus[21] .power_up = "low";

dffeas \rdaddress_b_bus[22] (
	.clk(clk),
	.d(\rdaddress_b_bus~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_b_bus_22),
	.prn(vcc));
defparam \rdaddress_b_bus[22] .is_wysiwyg = "true";
defparam \rdaddress_b_bus[22] .power_up = "low";

dffeas \rdaddress_b_bus[23] (
	.clk(clk),
	.d(\rdaddress_b_bus~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_b_bus_23),
	.prn(vcc));
defparam \rdaddress_b_bus[23] .is_wysiwyg = "true";
defparam \rdaddress_b_bus[23] .power_up = "low";

dffeas \rdaddress_b_bus[24] (
	.clk(clk),
	.d(\rdaddress_b_bus~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_b_bus_24),
	.prn(vcc));
defparam \rdaddress_b_bus[24] .is_wysiwyg = "true";
defparam \rdaddress_b_bus[24] .power_up = "low";

dffeas \rdaddress_b_bus[11] (
	.clk(clk),
	.d(\rdaddress_b_bus~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_b_bus_11),
	.prn(vcc));
defparam \rdaddress_b_bus[11] .is_wysiwyg = "true";
defparam \rdaddress_b_bus[11] .power_up = "low";

dffeas \rdaddress_b_bus[26] (
	.clk(clk),
	.d(\rdaddress_b_bus~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_b_bus_26),
	.prn(vcc));
defparam \rdaddress_b_bus[26] .is_wysiwyg = "true";
defparam \rdaddress_b_bus[26] .power_up = "low";

dffeas \rdaddress_b_bus[13] (
	.clk(clk),
	.d(\rdaddress_b_bus~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_b_bus_13),
	.prn(vcc));
defparam \rdaddress_b_bus[13] .is_wysiwyg = "true";
defparam \rdaddress_b_bus[13] .power_up = "low";

dffeas \a_ram_data_in_bus[58] (
	.clk(clk),
	.d(\a_ram_data_in_bus~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_58),
	.prn(vcc));
defparam \a_ram_data_in_bus[58] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[58] .power_up = "low";

dffeas \wraddress_a_bus[21] (
	.clk(clk),
	.d(\wraddress_a_bus~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_a_bus_21),
	.prn(vcc));
defparam \wraddress_a_bus[21] .is_wysiwyg = "true";
defparam \wraddress_a_bus[21] .power_up = "low";

dffeas \wraddress_a_bus[22] (
	.clk(clk),
	.d(\wraddress_a_bus~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_a_bus_22),
	.prn(vcc));
defparam \wraddress_a_bus[22] .is_wysiwyg = "true";
defparam \wraddress_a_bus[22] .power_up = "low";

dffeas \wraddress_a_bus[23] (
	.clk(clk),
	.d(\wraddress_a_bus~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_a_bus_23),
	.prn(vcc));
defparam \wraddress_a_bus[23] .is_wysiwyg = "true";
defparam \wraddress_a_bus[23] .power_up = "low";

dffeas \wraddress_a_bus[24] (
	.clk(clk),
	.d(\wraddress_a_bus~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_a_bus_24),
	.prn(vcc));
defparam \wraddress_a_bus[24] .is_wysiwyg = "true";
defparam \wraddress_a_bus[24] .power_up = "low";

dffeas \wraddress_a_bus[11] (
	.clk(clk),
	.d(\wraddress_a_bus~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_a_bus_11),
	.prn(vcc));
defparam \wraddress_a_bus[11] .is_wysiwyg = "true";
defparam \wraddress_a_bus[11] .power_up = "low";

dffeas \wraddress_a_bus[26] (
	.clk(clk),
	.d(\wraddress_a_bus~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_a_bus_26),
	.prn(vcc));
defparam \wraddress_a_bus[26] .is_wysiwyg = "true";
defparam \wraddress_a_bus[26] .power_up = "low";

dffeas \wraddress_a_bus[13] (
	.clk(clk),
	.d(\wraddress_a_bus~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_a_bus_13),
	.prn(vcc));
defparam \wraddress_a_bus[13] .is_wysiwyg = "true";
defparam \wraddress_a_bus[13] .power_up = "low";

dffeas \rdaddress_a_bus[21] (
	.clk(clk),
	.d(\rdaddress_a_bus~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_a_bus_21),
	.prn(vcc));
defparam \rdaddress_a_bus[21] .is_wysiwyg = "true";
defparam \rdaddress_a_bus[21] .power_up = "low";

dffeas \rdaddress_a_bus[22] (
	.clk(clk),
	.d(\rdaddress_a_bus~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_a_bus_22),
	.prn(vcc));
defparam \rdaddress_a_bus[22] .is_wysiwyg = "true";
defparam \rdaddress_a_bus[22] .power_up = "low";

dffeas \rdaddress_a_bus[23] (
	.clk(clk),
	.d(\rdaddress_a_bus~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_a_bus_23),
	.prn(vcc));
defparam \rdaddress_a_bus[23] .is_wysiwyg = "true";
defparam \rdaddress_a_bus[23] .power_up = "low";

dffeas \rdaddress_a_bus[24] (
	.clk(clk),
	.d(\rdaddress_a_bus~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_a_bus_24),
	.prn(vcc));
defparam \rdaddress_a_bus[24] .is_wysiwyg = "true";
defparam \rdaddress_a_bus[24] .power_up = "low";

dffeas \rdaddress_a_bus[11] (
	.clk(clk),
	.d(\rdaddress_a_bus~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_a_bus_11),
	.prn(vcc));
defparam \rdaddress_a_bus[11] .is_wysiwyg = "true";
defparam \rdaddress_a_bus[11] .power_up = "low";

dffeas \rdaddress_a_bus[26] (
	.clk(clk),
	.d(\rdaddress_a_bus~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_a_bus_26),
	.prn(vcc));
defparam \rdaddress_a_bus[26] .is_wysiwyg = "true";
defparam \rdaddress_a_bus[26] .power_up = "low";

dffeas \rdaddress_a_bus[13] (
	.clk(clk),
	.d(\rdaddress_a_bus~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_a_bus_13),
	.prn(vcc));
defparam \rdaddress_a_bus[13] .is_wysiwyg = "true";
defparam \rdaddress_a_bus[13] .power_up = "low";

dffeas \b_ram_data_in_bus[42] (
	.clk(clk),
	.d(\b_ram_data_in_bus~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_42),
	.prn(vcc));
defparam \b_ram_data_in_bus[42] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[42] .power_up = "low";

dffeas \wraddress_b_bus[0] (
	.clk(clk),
	.d(\wraddress_b_bus~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_b_bus_0),
	.prn(vcc));
defparam \wraddress_b_bus[0] .is_wysiwyg = "true";
defparam \wraddress_b_bus[0] .power_up = "low";

dffeas \wraddress_b_bus[15] (
	.clk(clk),
	.d(\wraddress_b_bus~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_b_bus_15),
	.prn(vcc));
defparam \wraddress_b_bus[15] .is_wysiwyg = "true";
defparam \wraddress_b_bus[15] .power_up = "low";

dffeas \wraddress_b_bus[16] (
	.clk(clk),
	.d(\wraddress_b_bus~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_b_bus_16),
	.prn(vcc));
defparam \wraddress_b_bus[16] .is_wysiwyg = "true";
defparam \wraddress_b_bus[16] .power_up = "low";

dffeas \wraddress_b_bus[17] (
	.clk(clk),
	.d(\wraddress_b_bus~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_b_bus_17),
	.prn(vcc));
defparam \wraddress_b_bus[17] .is_wysiwyg = "true";
defparam \wraddress_b_bus[17] .power_up = "low";

dffeas \wraddress_b_bus[18] (
	.clk(clk),
	.d(\wraddress_b_bus~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_b_bus_18),
	.prn(vcc));
defparam \wraddress_b_bus[18] .is_wysiwyg = "true";
defparam \wraddress_b_bus[18] .power_up = "low";

dffeas \wraddress_b_bus[19] (
	.clk(clk),
	.d(\wraddress_b_bus~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_b_bus_19),
	.prn(vcc));
defparam \wraddress_b_bus[19] .is_wysiwyg = "true";
defparam \wraddress_b_bus[19] .power_up = "low";

dffeas \rdaddress_b_bus[0] (
	.clk(clk),
	.d(\rdaddress_b_bus~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_b_bus_0),
	.prn(vcc));
defparam \rdaddress_b_bus[0] .is_wysiwyg = "true";
defparam \rdaddress_b_bus[0] .power_up = "low";

dffeas \rdaddress_b_bus[15] (
	.clk(clk),
	.d(\rdaddress_b_bus~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_b_bus_15),
	.prn(vcc));
defparam \rdaddress_b_bus[15] .is_wysiwyg = "true";
defparam \rdaddress_b_bus[15] .power_up = "low";

dffeas \rdaddress_b_bus[16] (
	.clk(clk),
	.d(\rdaddress_b_bus~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_b_bus_16),
	.prn(vcc));
defparam \rdaddress_b_bus[16] .is_wysiwyg = "true";
defparam \rdaddress_b_bus[16] .power_up = "low";

dffeas \rdaddress_b_bus[17] (
	.clk(clk),
	.d(\rdaddress_b_bus~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_b_bus_17),
	.prn(vcc));
defparam \rdaddress_b_bus[17] .is_wysiwyg = "true";
defparam \rdaddress_b_bus[17] .power_up = "low";

dffeas \rdaddress_b_bus[18] (
	.clk(clk),
	.d(\rdaddress_b_bus~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_b_bus_18),
	.prn(vcc));
defparam \rdaddress_b_bus[18] .is_wysiwyg = "true";
defparam \rdaddress_b_bus[18] .power_up = "low";

dffeas \rdaddress_b_bus[19] (
	.clk(clk),
	.d(\rdaddress_b_bus~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_b_bus_19),
	.prn(vcc));
defparam \rdaddress_b_bus[19] .is_wysiwyg = "true";
defparam \rdaddress_b_bus[19] .power_up = "low";

dffeas \a_ram_data_in_bus[42] (
	.clk(clk),
	.d(\a_ram_data_in_bus~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_42),
	.prn(vcc));
defparam \a_ram_data_in_bus[42] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[42] .power_up = "low";

dffeas \wraddress_a_bus[0] (
	.clk(clk),
	.d(\wraddress_a_bus~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_a_bus_0),
	.prn(vcc));
defparam \wraddress_a_bus[0] .is_wysiwyg = "true";
defparam \wraddress_a_bus[0] .power_up = "low";

dffeas \wraddress_a_bus[15] (
	.clk(clk),
	.d(\wraddress_a_bus~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_a_bus_15),
	.prn(vcc));
defparam \wraddress_a_bus[15] .is_wysiwyg = "true";
defparam \wraddress_a_bus[15] .power_up = "low";

dffeas \wraddress_a_bus[16] (
	.clk(clk),
	.d(\wraddress_a_bus~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_a_bus_16),
	.prn(vcc));
defparam \wraddress_a_bus[16] .is_wysiwyg = "true";
defparam \wraddress_a_bus[16] .power_up = "low";

dffeas \wraddress_a_bus[17] (
	.clk(clk),
	.d(\wraddress_a_bus~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_a_bus_17),
	.prn(vcc));
defparam \wraddress_a_bus[17] .is_wysiwyg = "true";
defparam \wraddress_a_bus[17] .power_up = "low";

dffeas \wraddress_a_bus[18] (
	.clk(clk),
	.d(\wraddress_a_bus~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_a_bus_18),
	.prn(vcc));
defparam \wraddress_a_bus[18] .is_wysiwyg = "true";
defparam \wraddress_a_bus[18] .power_up = "low";

dffeas \wraddress_a_bus[19] (
	.clk(clk),
	.d(\wraddress_a_bus~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_a_bus_19),
	.prn(vcc));
defparam \wraddress_a_bus[19] .is_wysiwyg = "true";
defparam \wraddress_a_bus[19] .power_up = "low";

dffeas \rdaddress_a_bus[0] (
	.clk(clk),
	.d(\rdaddress_a_bus~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_a_bus_0),
	.prn(vcc));
defparam \rdaddress_a_bus[0] .is_wysiwyg = "true";
defparam \rdaddress_a_bus[0] .power_up = "low";

dffeas \rdaddress_a_bus[15] (
	.clk(clk),
	.d(\rdaddress_a_bus~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_a_bus_15),
	.prn(vcc));
defparam \rdaddress_a_bus[15] .is_wysiwyg = "true";
defparam \rdaddress_a_bus[15] .power_up = "low";

dffeas \rdaddress_a_bus[16] (
	.clk(clk),
	.d(\rdaddress_a_bus~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_a_bus_16),
	.prn(vcc));
defparam \rdaddress_a_bus[16] .is_wysiwyg = "true";
defparam \rdaddress_a_bus[16] .power_up = "low";

dffeas \rdaddress_a_bus[17] (
	.clk(clk),
	.d(\rdaddress_a_bus~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_a_bus_17),
	.prn(vcc));
defparam \rdaddress_a_bus[17] .is_wysiwyg = "true";
defparam \rdaddress_a_bus[17] .power_up = "low";

dffeas \rdaddress_a_bus[18] (
	.clk(clk),
	.d(\rdaddress_a_bus~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_a_bus_18),
	.prn(vcc));
defparam \rdaddress_a_bus[18] .is_wysiwyg = "true";
defparam \rdaddress_a_bus[18] .power_up = "low";

dffeas \rdaddress_a_bus[19] (
	.clk(clk),
	.d(\rdaddress_a_bus~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_a_bus_19),
	.prn(vcc));
defparam \rdaddress_a_bus[19] .is_wysiwyg = "true";
defparam \rdaddress_a_bus[19] .power_up = "low";

dffeas \b_ram_data_in_bus[26] (
	.clk(clk),
	.d(\b_ram_data_in_bus~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_26),
	.prn(vcc));
defparam \b_ram_data_in_bus[26] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[26] .power_up = "low";

dffeas \wraddress_b_bus[8] (
	.clk(clk),
	.d(\wraddress_b_bus~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_b_bus_8),
	.prn(vcc));
defparam \wraddress_b_bus[8] .is_wysiwyg = "true";
defparam \wraddress_b_bus[8] .power_up = "low";

dffeas \wraddress_b_bus[10] (
	.clk(clk),
	.d(\wraddress_b_bus~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_b_bus_10),
	.prn(vcc));
defparam \wraddress_b_bus[10] .is_wysiwyg = "true";
defparam \wraddress_b_bus[10] .power_up = "low";

dffeas \wraddress_b_bus[12] (
	.clk(clk),
	.d(\wraddress_b_bus~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_b_bus_12),
	.prn(vcc));
defparam \wraddress_b_bus[12] .is_wysiwyg = "true";
defparam \wraddress_b_bus[12] .power_up = "low";

dffeas \rdaddress_b_bus[8] (
	.clk(clk),
	.d(\rdaddress_b_bus~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_b_bus_8),
	.prn(vcc));
defparam \rdaddress_b_bus[8] .is_wysiwyg = "true";
defparam \rdaddress_b_bus[8] .power_up = "low";

dffeas \rdaddress_b_bus[10] (
	.clk(clk),
	.d(\rdaddress_b_bus~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_b_bus_10),
	.prn(vcc));
defparam \rdaddress_b_bus[10] .is_wysiwyg = "true";
defparam \rdaddress_b_bus[10] .power_up = "low";

dffeas \rdaddress_b_bus[12] (
	.clk(clk),
	.d(\rdaddress_b_bus~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_b_bus_12),
	.prn(vcc));
defparam \rdaddress_b_bus[12] .is_wysiwyg = "true";
defparam \rdaddress_b_bus[12] .power_up = "low";

dffeas \a_ram_data_in_bus[26] (
	.clk(clk),
	.d(\a_ram_data_in_bus~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_26),
	.prn(vcc));
defparam \a_ram_data_in_bus[26] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[26] .power_up = "low";

dffeas \wraddress_a_bus[8] (
	.clk(clk),
	.d(\wraddress_a_bus~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_a_bus_8),
	.prn(vcc));
defparam \wraddress_a_bus[8] .is_wysiwyg = "true";
defparam \wraddress_a_bus[8] .power_up = "low";

dffeas \wraddress_a_bus[10] (
	.clk(clk),
	.d(\wraddress_a_bus~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_a_bus_10),
	.prn(vcc));
defparam \wraddress_a_bus[10] .is_wysiwyg = "true";
defparam \wraddress_a_bus[10] .power_up = "low";

dffeas \wraddress_a_bus[12] (
	.clk(clk),
	.d(\wraddress_a_bus~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_a_bus_12),
	.prn(vcc));
defparam \wraddress_a_bus[12] .is_wysiwyg = "true";
defparam \wraddress_a_bus[12] .power_up = "low";

dffeas \rdaddress_a_bus[8] (
	.clk(clk),
	.d(\rdaddress_a_bus~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_a_bus_8),
	.prn(vcc));
defparam \rdaddress_a_bus[8] .is_wysiwyg = "true";
defparam \rdaddress_a_bus[8] .power_up = "low";

dffeas \rdaddress_a_bus[10] (
	.clk(clk),
	.d(\rdaddress_a_bus~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_a_bus_10),
	.prn(vcc));
defparam \rdaddress_a_bus[10] .is_wysiwyg = "true";
defparam \rdaddress_a_bus[10] .power_up = "low";

dffeas \rdaddress_a_bus[12] (
	.clk(clk),
	.d(\rdaddress_a_bus~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_a_bus_12),
	.prn(vcc));
defparam \rdaddress_a_bus[12] .is_wysiwyg = "true";
defparam \rdaddress_a_bus[12] .power_up = "low";

dffeas \b_ram_data_in_bus[10] (
	.clk(clk),
	.d(\b_ram_data_in_bus~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_10),
	.prn(vcc));
defparam \b_ram_data_in_bus[10] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[10] .power_up = "low";

dffeas \wraddress_b_bus[1] (
	.clk(clk),
	.d(\wraddress_b_bus~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_b_bus_1),
	.prn(vcc));
defparam \wraddress_b_bus[1] .is_wysiwyg = "true";
defparam \wraddress_b_bus[1] .power_up = "low";

dffeas \wraddress_b_bus[3] (
	.clk(clk),
	.d(\wraddress_b_bus~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_b_bus_3),
	.prn(vcc));
defparam \wraddress_b_bus[3] .is_wysiwyg = "true";
defparam \wraddress_b_bus[3] .power_up = "low";

dffeas \wraddress_b_bus[5] (
	.clk(clk),
	.d(\wraddress_b_bus~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_b_bus_5),
	.prn(vcc));
defparam \wraddress_b_bus[5] .is_wysiwyg = "true";
defparam \wraddress_b_bus[5] .power_up = "low";

dffeas \rdaddress_b_bus[1] (
	.clk(clk),
	.d(\rdaddress_b_bus~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_b_bus_1),
	.prn(vcc));
defparam \rdaddress_b_bus[1] .is_wysiwyg = "true";
defparam \rdaddress_b_bus[1] .power_up = "low";

dffeas \rdaddress_b_bus[3] (
	.clk(clk),
	.d(\rdaddress_b_bus~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_b_bus_3),
	.prn(vcc));
defparam \rdaddress_b_bus[3] .is_wysiwyg = "true";
defparam \rdaddress_b_bus[3] .power_up = "low";

dffeas \rdaddress_b_bus[5] (
	.clk(clk),
	.d(\rdaddress_b_bus~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_b_bus_5),
	.prn(vcc));
defparam \rdaddress_b_bus[5] .is_wysiwyg = "true";
defparam \rdaddress_b_bus[5] .power_up = "low";

dffeas \a_ram_data_in_bus[10] (
	.clk(clk),
	.d(\a_ram_data_in_bus~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_10),
	.prn(vcc));
defparam \a_ram_data_in_bus[10] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[10] .power_up = "low";

dffeas \wraddress_a_bus[1] (
	.clk(clk),
	.d(\wraddress_a_bus~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_a_bus_1),
	.prn(vcc));
defparam \wraddress_a_bus[1] .is_wysiwyg = "true";
defparam \wraddress_a_bus[1] .power_up = "low";

dffeas \wraddress_a_bus[3] (
	.clk(clk),
	.d(\wraddress_a_bus~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_a_bus_3),
	.prn(vcc));
defparam \wraddress_a_bus[3] .is_wysiwyg = "true";
defparam \wraddress_a_bus[3] .power_up = "low";

dffeas \wraddress_a_bus[5] (
	.clk(clk),
	.d(\wraddress_a_bus~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_a_bus_5),
	.prn(vcc));
defparam \wraddress_a_bus[5] .is_wysiwyg = "true";
defparam \wraddress_a_bus[5] .power_up = "low";

dffeas \rdaddress_a_bus[1] (
	.clk(clk),
	.d(\rdaddress_a_bus~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_a_bus_1),
	.prn(vcc));
defparam \rdaddress_a_bus[1] .is_wysiwyg = "true";
defparam \rdaddress_a_bus[1] .power_up = "low";

dffeas \rdaddress_a_bus[3] (
	.clk(clk),
	.d(\rdaddress_a_bus~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_a_bus_3),
	.prn(vcc));
defparam \rdaddress_a_bus[3] .is_wysiwyg = "true";
defparam \rdaddress_a_bus[3] .power_up = "low";

dffeas \rdaddress_a_bus[5] (
	.clk(clk),
	.d(\rdaddress_a_bus~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_a_bus_5),
	.prn(vcc));
defparam \rdaddress_a_bus[5] .is_wysiwyg = "true";
defparam \rdaddress_a_bus[5] .power_up = "low";

dffeas \b_ram_data_in_bus[62] (
	.clk(clk),
	.d(\b_ram_data_in_bus~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_62),
	.prn(vcc));
defparam \b_ram_data_in_bus[62] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[62] .power_up = "low";

dffeas \a_ram_data_in_bus[62] (
	.clk(clk),
	.d(\a_ram_data_in_bus~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_62),
	.prn(vcc));
defparam \a_ram_data_in_bus[62] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[62] .power_up = "low";

dffeas \b_ram_data_in_bus[46] (
	.clk(clk),
	.d(\b_ram_data_in_bus~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_46),
	.prn(vcc));
defparam \b_ram_data_in_bus[46] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[46] .power_up = "low";

dffeas \a_ram_data_in_bus[46] (
	.clk(clk),
	.d(\a_ram_data_in_bus~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_46),
	.prn(vcc));
defparam \a_ram_data_in_bus[46] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[46] .power_up = "low";

dffeas \b_ram_data_in_bus[30] (
	.clk(clk),
	.d(\b_ram_data_in_bus~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_30),
	.prn(vcc));
defparam \b_ram_data_in_bus[30] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[30] .power_up = "low";

dffeas \a_ram_data_in_bus[30] (
	.clk(clk),
	.d(\a_ram_data_in_bus~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_30),
	.prn(vcc));
defparam \a_ram_data_in_bus[30] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[30] .power_up = "low";

dffeas \b_ram_data_in_bus[14] (
	.clk(clk),
	.d(\b_ram_data_in_bus~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_14),
	.prn(vcc));
defparam \b_ram_data_in_bus[14] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[14] .power_up = "low";

dffeas \a_ram_data_in_bus[14] (
	.clk(clk),
	.d(\a_ram_data_in_bus~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_14),
	.prn(vcc));
defparam \a_ram_data_in_bus[14] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[14] .power_up = "low";

dffeas \b_ram_data_in_bus[60] (
	.clk(clk),
	.d(\b_ram_data_in_bus~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_60),
	.prn(vcc));
defparam \b_ram_data_in_bus[60] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[60] .power_up = "low";

dffeas \a_ram_data_in_bus[60] (
	.clk(clk),
	.d(\a_ram_data_in_bus~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_60),
	.prn(vcc));
defparam \a_ram_data_in_bus[60] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[60] .power_up = "low";

dffeas \b_ram_data_in_bus[44] (
	.clk(clk),
	.d(\b_ram_data_in_bus~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_44),
	.prn(vcc));
defparam \b_ram_data_in_bus[44] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[44] .power_up = "low";

dffeas \a_ram_data_in_bus[44] (
	.clk(clk),
	.d(\a_ram_data_in_bus~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_44),
	.prn(vcc));
defparam \a_ram_data_in_bus[44] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[44] .power_up = "low";

dffeas \b_ram_data_in_bus[28] (
	.clk(clk),
	.d(\b_ram_data_in_bus~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_28),
	.prn(vcc));
defparam \b_ram_data_in_bus[28] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[28] .power_up = "low";

dffeas \a_ram_data_in_bus[28] (
	.clk(clk),
	.d(\a_ram_data_in_bus~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_28),
	.prn(vcc));
defparam \a_ram_data_in_bus[28] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[28] .power_up = "low";

dffeas \b_ram_data_in_bus[12] (
	.clk(clk),
	.d(\b_ram_data_in_bus~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_12),
	.prn(vcc));
defparam \b_ram_data_in_bus[12] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[12] .power_up = "low";

dffeas \a_ram_data_in_bus[12] (
	.clk(clk),
	.d(\a_ram_data_in_bus~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_12),
	.prn(vcc));
defparam \a_ram_data_in_bus[12] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[12] .power_up = "low";

dffeas \b_ram_data_in_bus[59] (
	.clk(clk),
	.d(\b_ram_data_in_bus~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_59),
	.prn(vcc));
defparam \b_ram_data_in_bus[59] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[59] .power_up = "low";

dffeas \a_ram_data_in_bus[59] (
	.clk(clk),
	.d(\a_ram_data_in_bus~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_59),
	.prn(vcc));
defparam \a_ram_data_in_bus[59] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[59] .power_up = "low";

dffeas \b_ram_data_in_bus[43] (
	.clk(clk),
	.d(\b_ram_data_in_bus~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_43),
	.prn(vcc));
defparam \b_ram_data_in_bus[43] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[43] .power_up = "low";

dffeas \a_ram_data_in_bus[43] (
	.clk(clk),
	.d(\a_ram_data_in_bus~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_43),
	.prn(vcc));
defparam \a_ram_data_in_bus[43] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[43] .power_up = "low";

dffeas \b_ram_data_in_bus[27] (
	.clk(clk),
	.d(\b_ram_data_in_bus~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_27),
	.prn(vcc));
defparam \b_ram_data_in_bus[27] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[27] .power_up = "low";

dffeas \a_ram_data_in_bus[27] (
	.clk(clk),
	.d(\a_ram_data_in_bus~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_27),
	.prn(vcc));
defparam \a_ram_data_in_bus[27] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[27] .power_up = "low";

dffeas \b_ram_data_in_bus[11] (
	.clk(clk),
	.d(\b_ram_data_in_bus~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_11),
	.prn(vcc));
defparam \b_ram_data_in_bus[11] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[11] .power_up = "low";

dffeas \a_ram_data_in_bus[11] (
	.clk(clk),
	.d(\a_ram_data_in_bus~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_11),
	.prn(vcc));
defparam \a_ram_data_in_bus[11] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[11] .power_up = "low";

dffeas \b_ram_data_in_bus[61] (
	.clk(clk),
	.d(\b_ram_data_in_bus~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_61),
	.prn(vcc));
defparam \b_ram_data_in_bus[61] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[61] .power_up = "low";

dffeas \a_ram_data_in_bus[61] (
	.clk(clk),
	.d(\a_ram_data_in_bus~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_61),
	.prn(vcc));
defparam \a_ram_data_in_bus[61] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[61] .power_up = "low";

dffeas \b_ram_data_in_bus[45] (
	.clk(clk),
	.d(\b_ram_data_in_bus~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_45),
	.prn(vcc));
defparam \b_ram_data_in_bus[45] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[45] .power_up = "low";

dffeas \a_ram_data_in_bus[45] (
	.clk(clk),
	.d(\a_ram_data_in_bus~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_45),
	.prn(vcc));
defparam \a_ram_data_in_bus[45] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[45] .power_up = "low";

dffeas \b_ram_data_in_bus[29] (
	.clk(clk),
	.d(\b_ram_data_in_bus~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_29),
	.prn(vcc));
defparam \b_ram_data_in_bus[29] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[29] .power_up = "low";

dffeas \a_ram_data_in_bus[29] (
	.clk(clk),
	.d(\a_ram_data_in_bus~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_29),
	.prn(vcc));
defparam \a_ram_data_in_bus[29] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[29] .power_up = "low";

dffeas \b_ram_data_in_bus[13] (
	.clk(clk),
	.d(\b_ram_data_in_bus~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_13),
	.prn(vcc));
defparam \b_ram_data_in_bus[13] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[13] .power_up = "low";

dffeas \a_ram_data_in_bus[13] (
	.clk(clk),
	.d(\a_ram_data_in_bus~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_13),
	.prn(vcc));
defparam \a_ram_data_in_bus[13] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[13] .power_up = "low";

dffeas \b_ram_data_in_bus[57] (
	.clk(clk),
	.d(\b_ram_data_in_bus~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_57),
	.prn(vcc));
defparam \b_ram_data_in_bus[57] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[57] .power_up = "low";

dffeas \a_ram_data_in_bus[57] (
	.clk(clk),
	.d(\a_ram_data_in_bus~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_57),
	.prn(vcc));
defparam \a_ram_data_in_bus[57] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[57] .power_up = "low";

dffeas \b_ram_data_in_bus[41] (
	.clk(clk),
	.d(\b_ram_data_in_bus~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_41),
	.prn(vcc));
defparam \b_ram_data_in_bus[41] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[41] .power_up = "low";

dffeas \a_ram_data_in_bus[41] (
	.clk(clk),
	.d(\a_ram_data_in_bus~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_41),
	.prn(vcc));
defparam \a_ram_data_in_bus[41] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[41] .power_up = "low";

dffeas \b_ram_data_in_bus[25] (
	.clk(clk),
	.d(\b_ram_data_in_bus~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_25),
	.prn(vcc));
defparam \b_ram_data_in_bus[25] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[25] .power_up = "low";

dffeas \a_ram_data_in_bus[25] (
	.clk(clk),
	.d(\a_ram_data_in_bus~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_25),
	.prn(vcc));
defparam \a_ram_data_in_bus[25] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[25] .power_up = "low";

dffeas \b_ram_data_in_bus[9] (
	.clk(clk),
	.d(\b_ram_data_in_bus~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_9),
	.prn(vcc));
defparam \b_ram_data_in_bus[9] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[9] .power_up = "low";

dffeas \a_ram_data_in_bus[9] (
	.clk(clk),
	.d(\a_ram_data_in_bus~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_9),
	.prn(vcc));
defparam \a_ram_data_in_bus[9] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[9] .power_up = "low";

dffeas \b_ram_data_in_bus[56] (
	.clk(clk),
	.d(\b_ram_data_in_bus~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_56),
	.prn(vcc));
defparam \b_ram_data_in_bus[56] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[56] .power_up = "low";

dffeas \a_ram_data_in_bus[56] (
	.clk(clk),
	.d(\a_ram_data_in_bus~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_56),
	.prn(vcc));
defparam \a_ram_data_in_bus[56] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[56] .power_up = "low";

dffeas \b_ram_data_in_bus[40] (
	.clk(clk),
	.d(\b_ram_data_in_bus~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_40),
	.prn(vcc));
defparam \b_ram_data_in_bus[40] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[40] .power_up = "low";

dffeas \a_ram_data_in_bus[40] (
	.clk(clk),
	.d(\a_ram_data_in_bus~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_40),
	.prn(vcc));
defparam \a_ram_data_in_bus[40] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[40] .power_up = "low";

dffeas \b_ram_data_in_bus[24] (
	.clk(clk),
	.d(\b_ram_data_in_bus~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_24),
	.prn(vcc));
defparam \b_ram_data_in_bus[24] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[24] .power_up = "low";

dffeas \a_ram_data_in_bus[24] (
	.clk(clk),
	.d(\a_ram_data_in_bus~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_24),
	.prn(vcc));
defparam \a_ram_data_in_bus[24] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[24] .power_up = "low";

dffeas \b_ram_data_in_bus[8] (
	.clk(clk),
	.d(\b_ram_data_in_bus~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_8),
	.prn(vcc));
defparam \b_ram_data_in_bus[8] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[8] .power_up = "low";

dffeas \a_ram_data_in_bus[8] (
	.clk(clk),
	.d(\a_ram_data_in_bus~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_8),
	.prn(vcc));
defparam \a_ram_data_in_bus[8] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[8] .power_up = "low";

dffeas \b_ram_data_in_bus[63] (
	.clk(clk),
	.d(\b_ram_data_in_bus~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_63),
	.prn(vcc));
defparam \b_ram_data_in_bus[63] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[63] .power_up = "low";

dffeas \a_ram_data_in_bus[63] (
	.clk(clk),
	.d(\a_ram_data_in_bus~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_63),
	.prn(vcc));
defparam \a_ram_data_in_bus[63] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[63] .power_up = "low";

dffeas \b_ram_data_in_bus[47] (
	.clk(clk),
	.d(\b_ram_data_in_bus~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_47),
	.prn(vcc));
defparam \b_ram_data_in_bus[47] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[47] .power_up = "low";

dffeas \a_ram_data_in_bus[47] (
	.clk(clk),
	.d(\a_ram_data_in_bus~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_47),
	.prn(vcc));
defparam \a_ram_data_in_bus[47] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[47] .power_up = "low";

dffeas \b_ram_data_in_bus[31] (
	.clk(clk),
	.d(\b_ram_data_in_bus~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_31),
	.prn(vcc));
defparam \b_ram_data_in_bus[31] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[31] .power_up = "low";

dffeas \a_ram_data_in_bus[31] (
	.clk(clk),
	.d(\a_ram_data_in_bus~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_31),
	.prn(vcc));
defparam \a_ram_data_in_bus[31] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[31] .power_up = "low";

dffeas \b_ram_data_in_bus[15] (
	.clk(clk),
	.d(\b_ram_data_in_bus~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_15),
	.prn(vcc));
defparam \b_ram_data_in_bus[15] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[15] .power_up = "low";

dffeas \a_ram_data_in_bus[15] (
	.clk(clk),
	.d(\a_ram_data_in_bus~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_15),
	.prn(vcc));
defparam \a_ram_data_in_bus[15] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[15] .power_up = "low";

dffeas \b_ram_data_in_bus[55] (
	.clk(clk),
	.d(\b_ram_data_in_bus~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_55),
	.prn(vcc));
defparam \b_ram_data_in_bus[55] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[55] .power_up = "low";

dffeas \a_ram_data_in_bus[55] (
	.clk(clk),
	.d(\a_ram_data_in_bus~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_55),
	.prn(vcc));
defparam \a_ram_data_in_bus[55] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[55] .power_up = "low";

dffeas \b_ram_data_in_bus[39] (
	.clk(clk),
	.d(\b_ram_data_in_bus~33_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_39),
	.prn(vcc));
defparam \b_ram_data_in_bus[39] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[39] .power_up = "low";

dffeas \a_ram_data_in_bus[39] (
	.clk(clk),
	.d(\a_ram_data_in_bus~33_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_39),
	.prn(vcc));
defparam \a_ram_data_in_bus[39] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[39] .power_up = "low";

dffeas \b_ram_data_in_bus[23] (
	.clk(clk),
	.d(\b_ram_data_in_bus~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_23),
	.prn(vcc));
defparam \b_ram_data_in_bus[23] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[23] .power_up = "low";

dffeas \a_ram_data_in_bus[23] (
	.clk(clk),
	.d(\a_ram_data_in_bus~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_23),
	.prn(vcc));
defparam \a_ram_data_in_bus[23] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[23] .power_up = "low";

dffeas \b_ram_data_in_bus[7] (
	.clk(clk),
	.d(\b_ram_data_in_bus~35_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_7),
	.prn(vcc));
defparam \b_ram_data_in_bus[7] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[7] .power_up = "low";

dffeas \a_ram_data_in_bus[7] (
	.clk(clk),
	.d(\a_ram_data_in_bus~35_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_7),
	.prn(vcc));
defparam \a_ram_data_in_bus[7] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[7] .power_up = "low";

dffeas \b_ram_data_in_bus[51] (
	.clk(clk),
	.d(\b_ram_data_in_bus~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_51),
	.prn(vcc));
defparam \b_ram_data_in_bus[51] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[51] .power_up = "low";

dffeas \a_ram_data_in_bus[51] (
	.clk(clk),
	.d(\a_ram_data_in_bus~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_51),
	.prn(vcc));
defparam \a_ram_data_in_bus[51] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[51] .power_up = "low";

dffeas \b_ram_data_in_bus[35] (
	.clk(clk),
	.d(\b_ram_data_in_bus~37_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_35),
	.prn(vcc));
defparam \b_ram_data_in_bus[35] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[35] .power_up = "low";

dffeas \a_ram_data_in_bus[35] (
	.clk(clk),
	.d(\a_ram_data_in_bus~37_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_35),
	.prn(vcc));
defparam \a_ram_data_in_bus[35] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[35] .power_up = "low";

dffeas \b_ram_data_in_bus[19] (
	.clk(clk),
	.d(\b_ram_data_in_bus~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_19),
	.prn(vcc));
defparam \b_ram_data_in_bus[19] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[19] .power_up = "low";

dffeas \a_ram_data_in_bus[19] (
	.clk(clk),
	.d(\a_ram_data_in_bus~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_19),
	.prn(vcc));
defparam \a_ram_data_in_bus[19] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[19] .power_up = "low";

dffeas \b_ram_data_in_bus[3] (
	.clk(clk),
	.d(\b_ram_data_in_bus~39_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_3),
	.prn(vcc));
defparam \b_ram_data_in_bus[3] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[3] .power_up = "low";

dffeas \a_ram_data_in_bus[3] (
	.clk(clk),
	.d(\a_ram_data_in_bus~39_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_3),
	.prn(vcc));
defparam \a_ram_data_in_bus[3] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[3] .power_up = "low";

dffeas \b_ram_data_in_bus[53] (
	.clk(clk),
	.d(\b_ram_data_in_bus~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_53),
	.prn(vcc));
defparam \b_ram_data_in_bus[53] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[53] .power_up = "low";

dffeas \a_ram_data_in_bus[53] (
	.clk(clk),
	.d(\a_ram_data_in_bus~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_53),
	.prn(vcc));
defparam \a_ram_data_in_bus[53] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[53] .power_up = "low";

dffeas \b_ram_data_in_bus[37] (
	.clk(clk),
	.d(\b_ram_data_in_bus~41_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_37),
	.prn(vcc));
defparam \b_ram_data_in_bus[37] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[37] .power_up = "low";

dffeas \a_ram_data_in_bus[37] (
	.clk(clk),
	.d(\a_ram_data_in_bus~41_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_37),
	.prn(vcc));
defparam \a_ram_data_in_bus[37] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[37] .power_up = "low";

dffeas \b_ram_data_in_bus[21] (
	.clk(clk),
	.d(\b_ram_data_in_bus~42_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_21),
	.prn(vcc));
defparam \b_ram_data_in_bus[21] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[21] .power_up = "low";

dffeas \a_ram_data_in_bus[21] (
	.clk(clk),
	.d(\a_ram_data_in_bus~42_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_21),
	.prn(vcc));
defparam \a_ram_data_in_bus[21] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[21] .power_up = "low";

dffeas \b_ram_data_in_bus[5] (
	.clk(clk),
	.d(\b_ram_data_in_bus~43_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_5),
	.prn(vcc));
defparam \b_ram_data_in_bus[5] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[5] .power_up = "low";

dffeas \a_ram_data_in_bus[5] (
	.clk(clk),
	.d(\a_ram_data_in_bus~43_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_5),
	.prn(vcc));
defparam \a_ram_data_in_bus[5] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[5] .power_up = "low";

dffeas \b_ram_data_in_bus[52] (
	.clk(clk),
	.d(\b_ram_data_in_bus~44_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_52),
	.prn(vcc));
defparam \b_ram_data_in_bus[52] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[52] .power_up = "low";

dffeas \a_ram_data_in_bus[52] (
	.clk(clk),
	.d(\a_ram_data_in_bus~44_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_52),
	.prn(vcc));
defparam \a_ram_data_in_bus[52] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[52] .power_up = "low";

dffeas \b_ram_data_in_bus[36] (
	.clk(clk),
	.d(\b_ram_data_in_bus~45_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_36),
	.prn(vcc));
defparam \b_ram_data_in_bus[36] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[36] .power_up = "low";

dffeas \a_ram_data_in_bus[36] (
	.clk(clk),
	.d(\a_ram_data_in_bus~45_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_36),
	.prn(vcc));
defparam \a_ram_data_in_bus[36] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[36] .power_up = "low";

dffeas \b_ram_data_in_bus[20] (
	.clk(clk),
	.d(\b_ram_data_in_bus~46_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_20),
	.prn(vcc));
defparam \b_ram_data_in_bus[20] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[20] .power_up = "low";

dffeas \a_ram_data_in_bus[20] (
	.clk(clk),
	.d(\a_ram_data_in_bus~46_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_20),
	.prn(vcc));
defparam \a_ram_data_in_bus[20] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[20] .power_up = "low";

dffeas \b_ram_data_in_bus[4] (
	.clk(clk),
	.d(\b_ram_data_in_bus~47_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_4),
	.prn(vcc));
defparam \b_ram_data_in_bus[4] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[4] .power_up = "low";

dffeas \a_ram_data_in_bus[4] (
	.clk(clk),
	.d(\a_ram_data_in_bus~47_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_4),
	.prn(vcc));
defparam \a_ram_data_in_bus[4] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[4] .power_up = "low";

dffeas \b_ram_data_in_bus[54] (
	.clk(clk),
	.d(\b_ram_data_in_bus~48_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_54),
	.prn(vcc));
defparam \b_ram_data_in_bus[54] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[54] .power_up = "low";

dffeas \a_ram_data_in_bus[54] (
	.clk(clk),
	.d(\a_ram_data_in_bus~48_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_54),
	.prn(vcc));
defparam \a_ram_data_in_bus[54] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[54] .power_up = "low";

dffeas \b_ram_data_in_bus[38] (
	.clk(clk),
	.d(\b_ram_data_in_bus~49_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_38),
	.prn(vcc));
defparam \b_ram_data_in_bus[38] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[38] .power_up = "low";

dffeas \a_ram_data_in_bus[38] (
	.clk(clk),
	.d(\a_ram_data_in_bus~49_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_38),
	.prn(vcc));
defparam \a_ram_data_in_bus[38] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[38] .power_up = "low";

dffeas \b_ram_data_in_bus[22] (
	.clk(clk),
	.d(\b_ram_data_in_bus~50_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_22),
	.prn(vcc));
defparam \b_ram_data_in_bus[22] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[22] .power_up = "low";

dffeas \a_ram_data_in_bus[22] (
	.clk(clk),
	.d(\a_ram_data_in_bus~50_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_22),
	.prn(vcc));
defparam \a_ram_data_in_bus[22] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[22] .power_up = "low";

dffeas \b_ram_data_in_bus[6] (
	.clk(clk),
	.d(\b_ram_data_in_bus~51_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_6),
	.prn(vcc));
defparam \b_ram_data_in_bus[6] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[6] .power_up = "low";

dffeas \a_ram_data_in_bus[6] (
	.clk(clk),
	.d(\a_ram_data_in_bus~51_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_6),
	.prn(vcc));
defparam \a_ram_data_in_bus[6] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[6] .power_up = "low";

dffeas \b_ram_data_in_bus[50] (
	.clk(clk),
	.d(\b_ram_data_in_bus~52_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_50),
	.prn(vcc));
defparam \b_ram_data_in_bus[50] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[50] .power_up = "low";

dffeas \a_ram_data_in_bus[50] (
	.clk(clk),
	.d(\a_ram_data_in_bus~52_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_50),
	.prn(vcc));
defparam \a_ram_data_in_bus[50] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[50] .power_up = "low";

dffeas \b_ram_data_in_bus[34] (
	.clk(clk),
	.d(\b_ram_data_in_bus~53_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_34),
	.prn(vcc));
defparam \b_ram_data_in_bus[34] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[34] .power_up = "low";

dffeas \a_ram_data_in_bus[34] (
	.clk(clk),
	.d(\a_ram_data_in_bus~53_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_34),
	.prn(vcc));
defparam \a_ram_data_in_bus[34] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[34] .power_up = "low";

dffeas \b_ram_data_in_bus[18] (
	.clk(clk),
	.d(\b_ram_data_in_bus~54_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_18),
	.prn(vcc));
defparam \b_ram_data_in_bus[18] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[18] .power_up = "low";

dffeas \a_ram_data_in_bus[18] (
	.clk(clk),
	.d(\a_ram_data_in_bus~54_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_18),
	.prn(vcc));
defparam \a_ram_data_in_bus[18] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[18] .power_up = "low";

dffeas \b_ram_data_in_bus[2] (
	.clk(clk),
	.d(\b_ram_data_in_bus~55_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_2),
	.prn(vcc));
defparam \b_ram_data_in_bus[2] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[2] .power_up = "low";

dffeas \a_ram_data_in_bus[2] (
	.clk(clk),
	.d(\a_ram_data_in_bus~55_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_2),
	.prn(vcc));
defparam \a_ram_data_in_bus[2] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[2] .power_up = "low";

dffeas \b_ram_data_in_bus[49] (
	.clk(clk),
	.d(\b_ram_data_in_bus~56_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_49),
	.prn(vcc));
defparam \b_ram_data_in_bus[49] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[49] .power_up = "low";

dffeas \a_ram_data_in_bus[49] (
	.clk(clk),
	.d(\a_ram_data_in_bus~56_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_49),
	.prn(vcc));
defparam \a_ram_data_in_bus[49] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[49] .power_up = "low";

dffeas \b_ram_data_in_bus[33] (
	.clk(clk),
	.d(\b_ram_data_in_bus~57_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_33),
	.prn(vcc));
defparam \b_ram_data_in_bus[33] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[33] .power_up = "low";

dffeas \a_ram_data_in_bus[33] (
	.clk(clk),
	.d(\a_ram_data_in_bus~57_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_33),
	.prn(vcc));
defparam \a_ram_data_in_bus[33] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[33] .power_up = "low";

dffeas \b_ram_data_in_bus[17] (
	.clk(clk),
	.d(\b_ram_data_in_bus~58_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_17),
	.prn(vcc));
defparam \b_ram_data_in_bus[17] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[17] .power_up = "low";

dffeas \a_ram_data_in_bus[17] (
	.clk(clk),
	.d(\a_ram_data_in_bus~58_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_17),
	.prn(vcc));
defparam \a_ram_data_in_bus[17] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[17] .power_up = "low";

dffeas \b_ram_data_in_bus[1] (
	.clk(clk),
	.d(\b_ram_data_in_bus~59_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_1),
	.prn(vcc));
defparam \b_ram_data_in_bus[1] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[1] .power_up = "low";

dffeas \a_ram_data_in_bus[1] (
	.clk(clk),
	.d(\a_ram_data_in_bus~59_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_1),
	.prn(vcc));
defparam \a_ram_data_in_bus[1] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[1] .power_up = "low";

dffeas \b_ram_data_in_bus[48] (
	.clk(clk),
	.d(\b_ram_data_in_bus~60_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_48),
	.prn(vcc));
defparam \b_ram_data_in_bus[48] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[48] .power_up = "low";

dffeas \a_ram_data_in_bus[48] (
	.clk(clk),
	.d(\a_ram_data_in_bus~60_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_48),
	.prn(vcc));
defparam \a_ram_data_in_bus[48] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[48] .power_up = "low";

dffeas \b_ram_data_in_bus[32] (
	.clk(clk),
	.d(\b_ram_data_in_bus~61_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_32),
	.prn(vcc));
defparam \b_ram_data_in_bus[32] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[32] .power_up = "low";

dffeas \a_ram_data_in_bus[32] (
	.clk(clk),
	.d(\a_ram_data_in_bus~61_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_32),
	.prn(vcc));
defparam \a_ram_data_in_bus[32] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[32] .power_up = "low";

dffeas \b_ram_data_in_bus[16] (
	.clk(clk),
	.d(\b_ram_data_in_bus~62_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_16),
	.prn(vcc));
defparam \b_ram_data_in_bus[16] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[16] .power_up = "low";

dffeas \a_ram_data_in_bus[16] (
	.clk(clk),
	.d(\a_ram_data_in_bus~62_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_16),
	.prn(vcc));
defparam \a_ram_data_in_bus[16] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[16] .power_up = "low";

dffeas \b_ram_data_in_bus[0] (
	.clk(clk),
	.d(\b_ram_data_in_bus~63_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(b_ram_data_in_bus_0),
	.prn(vcc));
defparam \b_ram_data_in_bus[0] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[0] .power_up = "low";

dffeas \a_ram_data_in_bus[0] (
	.clk(clk),
	.d(\a_ram_data_in_bus~63_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_0),
	.prn(vcc));
defparam \a_ram_data_in_bus[0] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[0] .power_up = "low";

cycloneiii_lcell_comb \ram_data_out0~0 (
	.dataa(q_b_10),
	.datab(q_b_101),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out0~0_combout ),
	.cout());
defparam \ram_data_out0~0 .lut_mask = 16'hEFFE;
defparam \ram_data_out0~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out1~0 (
	.dataa(q_b_102),
	.datab(q_b_103),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out1~0_combout ),
	.cout());
defparam \ram_data_out1~0 .lut_mask = 16'hEFFE;
defparam \ram_data_out1~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out2~0 (
	.dataa(q_b_104),
	.datab(q_b_105),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out2~0_combout ),
	.cout());
defparam \ram_data_out2~0 .lut_mask = 16'hEFFE;
defparam \ram_data_out2~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out3~0 (
	.dataa(q_b_106),
	.datab(q_b_107),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out3~0_combout ),
	.cout());
defparam \ram_data_out3~0 .lut_mask = 16'hEFFE;
defparam \ram_data_out3~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out0~1 (
	.dataa(q_b_14),
	.datab(q_b_141),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out0~1_combout ),
	.cout());
defparam \ram_data_out0~1 .lut_mask = 16'hEFFE;
defparam \ram_data_out0~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out1~1 (
	.dataa(q_b_142),
	.datab(q_b_143),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out1~1_combout ),
	.cout());
defparam \ram_data_out1~1 .lut_mask = 16'hEFFE;
defparam \ram_data_out1~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out2~1 (
	.dataa(q_b_144),
	.datab(q_b_145),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out2~1_combout ),
	.cout());
defparam \ram_data_out2~1 .lut_mask = 16'hEFFE;
defparam \ram_data_out2~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out3~1 (
	.dataa(q_b_146),
	.datab(q_b_147),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out3~1_combout ),
	.cout());
defparam \ram_data_out3~1 .lut_mask = 16'hEFFE;
defparam \ram_data_out3~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out0~2 (
	.dataa(q_b_12),
	.datab(q_b_121),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out0~2_combout ),
	.cout());
defparam \ram_data_out0~2 .lut_mask = 16'hEFFE;
defparam \ram_data_out0~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out1~2 (
	.dataa(q_b_122),
	.datab(q_b_123),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out1~2_combout ),
	.cout());
defparam \ram_data_out1~2 .lut_mask = 16'hEFFE;
defparam \ram_data_out1~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out2~2 (
	.dataa(q_b_124),
	.datab(q_b_125),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out2~2_combout ),
	.cout());
defparam \ram_data_out2~2 .lut_mask = 16'hEFFE;
defparam \ram_data_out2~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out3~2 (
	.dataa(q_b_126),
	.datab(q_b_127),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out3~2_combout ),
	.cout());
defparam \ram_data_out3~2 .lut_mask = 16'hEFFE;
defparam \ram_data_out3~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out0~3 (
	.dataa(q_b_11),
	.datab(q_b_111),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out0~3_combout ),
	.cout());
defparam \ram_data_out0~3 .lut_mask = 16'hEFFE;
defparam \ram_data_out0~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out1~3 (
	.dataa(q_b_112),
	.datab(q_b_113),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out1~3_combout ),
	.cout());
defparam \ram_data_out1~3 .lut_mask = 16'hEFFE;
defparam \ram_data_out1~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out2~3 (
	.dataa(q_b_114),
	.datab(q_b_115),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out2~3_combout ),
	.cout());
defparam \ram_data_out2~3 .lut_mask = 16'hEFFE;
defparam \ram_data_out2~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out3~3 (
	.dataa(q_b_116),
	.datab(q_b_117),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out3~3_combout ),
	.cout());
defparam \ram_data_out3~3 .lut_mask = 16'hEFFE;
defparam \ram_data_out3~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out0~4 (
	.dataa(q_b_13),
	.datab(q_b_131),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out0~4_combout ),
	.cout());
defparam \ram_data_out0~4 .lut_mask = 16'hEFFE;
defparam \ram_data_out0~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out1~4 (
	.dataa(q_b_132),
	.datab(q_b_133),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out1~4_combout ),
	.cout());
defparam \ram_data_out1~4 .lut_mask = 16'hEFFE;
defparam \ram_data_out1~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out2~4 (
	.dataa(q_b_134),
	.datab(q_b_135),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out2~4_combout ),
	.cout());
defparam \ram_data_out2~4 .lut_mask = 16'hEFFE;
defparam \ram_data_out2~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out3~4 (
	.dataa(q_b_136),
	.datab(q_b_137),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out3~4_combout ),
	.cout());
defparam \ram_data_out3~4 .lut_mask = 16'hEFFE;
defparam \ram_data_out3~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out0~5 (
	.dataa(q_b_9),
	.datab(q_b_91),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out0~5_combout ),
	.cout());
defparam \ram_data_out0~5 .lut_mask = 16'hEFFE;
defparam \ram_data_out0~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out1~5 (
	.dataa(q_b_92),
	.datab(q_b_93),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out1~5_combout ),
	.cout());
defparam \ram_data_out1~5 .lut_mask = 16'hEFFE;
defparam \ram_data_out1~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out2~5 (
	.dataa(q_b_94),
	.datab(q_b_95),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out2~5_combout ),
	.cout());
defparam \ram_data_out2~5 .lut_mask = 16'hEFFE;
defparam \ram_data_out2~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out3~5 (
	.dataa(q_b_96),
	.datab(q_b_97),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out3~5_combout ),
	.cout());
defparam \ram_data_out3~5 .lut_mask = 16'hEFFE;
defparam \ram_data_out3~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out0~6 (
	.dataa(q_b_8),
	.datab(q_b_81),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out0~6_combout ),
	.cout());
defparam \ram_data_out0~6 .lut_mask = 16'hEFFE;
defparam \ram_data_out0~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out1~6 (
	.dataa(q_b_82),
	.datab(q_b_83),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out1~6_combout ),
	.cout());
defparam \ram_data_out1~6 .lut_mask = 16'hEFFE;
defparam \ram_data_out1~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out2~6 (
	.dataa(q_b_84),
	.datab(q_b_85),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out2~6_combout ),
	.cout());
defparam \ram_data_out2~6 .lut_mask = 16'hEFFE;
defparam \ram_data_out2~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out3~6 (
	.dataa(q_b_86),
	.datab(q_b_87),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out3~6_combout ),
	.cout());
defparam \ram_data_out3~6 .lut_mask = 16'hEFFE;
defparam \ram_data_out3~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out0~7 (
	.dataa(q_b_15),
	.datab(q_b_151),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out0~7_combout ),
	.cout());
defparam \ram_data_out0~7 .lut_mask = 16'hEFFE;
defparam \ram_data_out0~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out1~7 (
	.dataa(q_b_152),
	.datab(q_b_153),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out1~7_combout ),
	.cout());
defparam \ram_data_out1~7 .lut_mask = 16'hEFFE;
defparam \ram_data_out1~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out2~7 (
	.dataa(q_b_154),
	.datab(q_b_155),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out2~7_combout ),
	.cout());
defparam \ram_data_out2~7 .lut_mask = 16'hEFFE;
defparam \ram_data_out2~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out3~7 (
	.dataa(q_b_156),
	.datab(q_b_157),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out3~7_combout ),
	.cout());
defparam \ram_data_out3~7 .lut_mask = 16'hEFFE;
defparam \ram_data_out3~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out0~8 (
	.dataa(q_b_7),
	.datab(q_b_71),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out0~8_combout ),
	.cout());
defparam \ram_data_out0~8 .lut_mask = 16'hEFFE;
defparam \ram_data_out0~8 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out1~8 (
	.dataa(q_b_72),
	.datab(q_b_73),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out1~8_combout ),
	.cout());
defparam \ram_data_out1~8 .lut_mask = 16'hEFFE;
defparam \ram_data_out1~8 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out2~8 (
	.dataa(q_b_74),
	.datab(q_b_75),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out2~8_combout ),
	.cout());
defparam \ram_data_out2~8 .lut_mask = 16'hEFFE;
defparam \ram_data_out2~8 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out3~8 (
	.dataa(q_b_76),
	.datab(q_b_77),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out3~8_combout ),
	.cout());
defparam \ram_data_out3~8 .lut_mask = 16'hEFFE;
defparam \ram_data_out3~8 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out0~9 (
	.dataa(q_b_3),
	.datab(q_b_31),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out0~9_combout ),
	.cout());
defparam \ram_data_out0~9 .lut_mask = 16'hEFFE;
defparam \ram_data_out0~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out1~9 (
	.dataa(q_b_32),
	.datab(q_b_33),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out1~9_combout ),
	.cout());
defparam \ram_data_out1~9 .lut_mask = 16'hEFFE;
defparam \ram_data_out1~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out2~9 (
	.dataa(q_b_34),
	.datab(q_b_35),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out2~9_combout ),
	.cout());
defparam \ram_data_out2~9 .lut_mask = 16'hEFFE;
defparam \ram_data_out2~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out3~9 (
	.dataa(q_b_36),
	.datab(q_b_37),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out3~9_combout ),
	.cout());
defparam \ram_data_out3~9 .lut_mask = 16'hEFFE;
defparam \ram_data_out3~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out0~10 (
	.dataa(q_b_5),
	.datab(q_b_51),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out0~10_combout ),
	.cout());
defparam \ram_data_out0~10 .lut_mask = 16'hEFFE;
defparam \ram_data_out0~10 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out1~10 (
	.dataa(q_b_52),
	.datab(q_b_53),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out1~10_combout ),
	.cout());
defparam \ram_data_out1~10 .lut_mask = 16'hEFFE;
defparam \ram_data_out1~10 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out2~10 (
	.dataa(q_b_54),
	.datab(q_b_55),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out2~10_combout ),
	.cout());
defparam \ram_data_out2~10 .lut_mask = 16'hEFFE;
defparam \ram_data_out2~10 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out3~10 (
	.dataa(q_b_56),
	.datab(q_b_57),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out3~10_combout ),
	.cout());
defparam \ram_data_out3~10 .lut_mask = 16'hEFFE;
defparam \ram_data_out3~10 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out0~11 (
	.dataa(q_b_4),
	.datab(q_b_41),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out0~11_combout ),
	.cout());
defparam \ram_data_out0~11 .lut_mask = 16'hEFFE;
defparam \ram_data_out0~11 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out1~11 (
	.dataa(q_b_42),
	.datab(q_b_43),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out1~11_combout ),
	.cout());
defparam \ram_data_out1~11 .lut_mask = 16'hEFFE;
defparam \ram_data_out1~11 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out2~11 (
	.dataa(q_b_44),
	.datab(q_b_45),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out2~11_combout ),
	.cout());
defparam \ram_data_out2~11 .lut_mask = 16'hEFFE;
defparam \ram_data_out2~11 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out3~11 (
	.dataa(q_b_46),
	.datab(q_b_47),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out3~11_combout ),
	.cout());
defparam \ram_data_out3~11 .lut_mask = 16'hEFFE;
defparam \ram_data_out3~11 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out0~12 (
	.dataa(q_b_6),
	.datab(q_b_61),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out0~12_combout ),
	.cout());
defparam \ram_data_out0~12 .lut_mask = 16'hEFFE;
defparam \ram_data_out0~12 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out1~12 (
	.dataa(q_b_62),
	.datab(q_b_63),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out1~12_combout ),
	.cout());
defparam \ram_data_out1~12 .lut_mask = 16'hEFFE;
defparam \ram_data_out1~12 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out2~12 (
	.dataa(q_b_64),
	.datab(q_b_65),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out2~12_combout ),
	.cout());
defparam \ram_data_out2~12 .lut_mask = 16'hEFFE;
defparam \ram_data_out2~12 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out3~12 (
	.dataa(q_b_66),
	.datab(q_b_67),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out3~12_combout ),
	.cout());
defparam \ram_data_out3~12 .lut_mask = 16'hEFFE;
defparam \ram_data_out3~12 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out0~13 (
	.dataa(q_b_2),
	.datab(q_b_21),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out0~13_combout ),
	.cout());
defparam \ram_data_out0~13 .lut_mask = 16'hEFFE;
defparam \ram_data_out0~13 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out1~13 (
	.dataa(q_b_22),
	.datab(q_b_23),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out1~13_combout ),
	.cout());
defparam \ram_data_out1~13 .lut_mask = 16'hEFFE;
defparam \ram_data_out1~13 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out2~13 (
	.dataa(q_b_24),
	.datab(q_b_25),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out2~13_combout ),
	.cout());
defparam \ram_data_out2~13 .lut_mask = 16'hEFFE;
defparam \ram_data_out2~13 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out3~13 (
	.dataa(q_b_26),
	.datab(q_b_27),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out3~13_combout ),
	.cout());
defparam \ram_data_out3~13 .lut_mask = 16'hEFFE;
defparam \ram_data_out3~13 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out0~14 (
	.dataa(q_b_1),
	.datab(q_b_16),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out0~14_combout ),
	.cout());
defparam \ram_data_out0~14 .lut_mask = 16'hEFFE;
defparam \ram_data_out0~14 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out1~14 (
	.dataa(q_b_17),
	.datab(q_b_18),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out1~14_combout ),
	.cout());
defparam \ram_data_out1~14 .lut_mask = 16'hEFFE;
defparam \ram_data_out1~14 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out2~14 (
	.dataa(q_b_19),
	.datab(q_b_110),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out2~14_combout ),
	.cout());
defparam \ram_data_out2~14 .lut_mask = 16'hEFFE;
defparam \ram_data_out2~14 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out3~14 (
	.dataa(q_b_118),
	.datab(q_b_119),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out3~14_combout ),
	.cout());
defparam \ram_data_out3~14 .lut_mask = 16'hEFFE;
defparam \ram_data_out3~14 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out0~15 (
	.dataa(q_b_0),
	.datab(q_b_01),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out0~15_combout ),
	.cout());
defparam \ram_data_out0~15 .lut_mask = 16'hEFFE;
defparam \ram_data_out0~15 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out1~15 (
	.dataa(q_b_02),
	.datab(q_b_03),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out1~15_combout ),
	.cout());
defparam \ram_data_out1~15 .lut_mask = 16'hEFFE;
defparam \ram_data_out1~15 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out2~15 (
	.dataa(q_b_04),
	.datab(q_b_05),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out2~15_combout ),
	.cout());
defparam \ram_data_out2~15 .lut_mask = 16'hEFFE;
defparam \ram_data_out2~15 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_data_out3~15 (
	.dataa(q_b_06),
	.datab(q_b_07),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_10),
	.cin(gnd),
	.combout(\ram_data_out3~15_combout ),
	.cout());
defparam \ram_data_out3~15 .lut_mask = 16'hEFFE;
defparam \ram_data_out3~15 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~0 (
	.dataa(ram_in_reg_2_0),
	.datab(data_in_r_2),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~0_combout ),
	.cout());
defparam \b_ram_data_in_bus~0 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wraddress_b_bus~0 (
	.dataa(ram_in_reg_0_01),
	.datab(wr_address_i_int_0),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\wraddress_b_bus~0_combout ),
	.cout());
defparam \wraddress_b_bus~0 .lut_mask = 16'hAACC;
defparam \wraddress_b_bus~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wraddress_b_bus~1 (
	.dataa(ram_in_reg_1_01),
	.datab(wr_address_i_int_1),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\wraddress_b_bus~1_combout ),
	.cout());
defparam \wraddress_b_bus~1 .lut_mask = 16'hAACC;
defparam \wraddress_b_bus~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wraddress_b_bus~2 (
	.dataa(ram_in_reg_2_01),
	.datab(wr_address_i_int_2),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\wraddress_b_bus~2_combout ),
	.cout());
defparam \wraddress_b_bus~2 .lut_mask = 16'hAACC;
defparam \wraddress_b_bus~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wraddress_b_bus~3 (
	.dataa(ram_in_reg_3_01),
	.datab(wr_address_i_int_3),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\wraddress_b_bus~3_combout ),
	.cout());
defparam \wraddress_b_bus~3 .lut_mask = 16'hAACC;
defparam \wraddress_b_bus~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wraddress_b_bus~4 (
	.dataa(ram_in_reg_4_01),
	.datab(wr_address_i_int_4),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\wraddress_b_bus~4_combout ),
	.cout());
defparam \wraddress_b_bus~4 .lut_mask = 16'hAACC;
defparam \wraddress_b_bus~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wraddress_b_bus~5 (
	.dataa(ram_in_reg_5_01),
	.datab(wr_address_i_int_5),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\wraddress_b_bus~5_combout ),
	.cout());
defparam \wraddress_b_bus~5 .lut_mask = 16'hAACC;
defparam \wraddress_b_bus~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wraddress_b_bus~6 (
	.dataa(ram_in_reg_6_01),
	.datab(wr_address_i_int_6),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\wraddress_b_bus~6_combout ),
	.cout());
defparam \wraddress_b_bus~6 .lut_mask = 16'hAACC;
defparam \wraddress_b_bus~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rdaddress_b_bus~0 (
	.dataa(data_rdy_vec_10),
	.datab(ram_a_not_b_vec_7),
	.datac(ram_in_reg_0_02),
	.datad(gnd),
	.cin(gnd),
	.combout(\rdaddress_b_bus~0_combout ),
	.cout());
defparam \rdaddress_b_bus~0 .lut_mask = 16'hFEFE;
defparam \rdaddress_b_bus~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rdaddress_b_bus~1 (
	.dataa(data_rdy_vec_10),
	.datab(ram_a_not_b_vec_7),
	.datac(ram_in_reg_1_02),
	.datad(gnd),
	.cin(gnd),
	.combout(\rdaddress_b_bus~1_combout ),
	.cout());
defparam \rdaddress_b_bus~1 .lut_mask = 16'hFEFE;
defparam \rdaddress_b_bus~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rdaddress_b_bus~2 (
	.dataa(data_rdy_vec_10),
	.datab(ram_a_not_b_vec_7),
	.datac(ram_in_reg_2_02),
	.datad(gnd),
	.cin(gnd),
	.combout(\rdaddress_b_bus~2_combout ),
	.cout());
defparam \rdaddress_b_bus~2 .lut_mask = 16'hFEFE;
defparam \rdaddress_b_bus~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rdaddress_b_bus~3 (
	.dataa(data_rdy_vec_10),
	.datab(ram_a_not_b_vec_7),
	.datac(ram_in_reg_3_02),
	.datad(gnd),
	.cin(gnd),
	.combout(\rdaddress_b_bus~3_combout ),
	.cout());
defparam \rdaddress_b_bus~3 .lut_mask = 16'hFEFE;
defparam \rdaddress_b_bus~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rdaddress_b_bus~4 (
	.dataa(data_rdy_vec_10),
	.datab(ram_a_not_b_vec_7),
	.datac(ram_in_reg_4_02),
	.datad(gnd),
	.cin(gnd),
	.combout(\rdaddress_b_bus~4_combout ),
	.cout());
defparam \rdaddress_b_bus~4 .lut_mask = 16'hFEFE;
defparam \rdaddress_b_bus~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rdaddress_b_bus~5 (
	.dataa(data_rdy_vec_10),
	.datab(ram_a_not_b_vec_7),
	.datac(ram_in_reg_5_02),
	.datad(gnd),
	.cin(gnd),
	.combout(\rdaddress_b_bus~5_combout ),
	.cout());
defparam \rdaddress_b_bus~5 .lut_mask = 16'hFEFE;
defparam \rdaddress_b_bus~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rdaddress_b_bus~6 (
	.dataa(data_rdy_vec_10),
	.datab(ram_a_not_b_vec_7),
	.datac(tdl_arr_6_1),
	.datad(gnd),
	.cin(gnd),
	.combout(\rdaddress_b_bus~6_combout ),
	.cout());
defparam \rdaddress_b_bus~6 .lut_mask = 16'hFEFE;
defparam \rdaddress_b_bus~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~0 (
	.dataa(data_in_r_2),
	.datab(ram_in_reg_2_0),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~0_combout ),
	.cout());
defparam \a_ram_data_in_bus~0 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wraddress_a_bus~0 (
	.dataa(wr_address_i_int_0),
	.datab(ram_in_reg_0_01),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\wraddress_a_bus~0_combout ),
	.cout());
defparam \wraddress_a_bus~0 .lut_mask = 16'hAACC;
defparam \wraddress_a_bus~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wraddress_a_bus~1 (
	.dataa(wr_address_i_int_1),
	.datab(ram_in_reg_1_01),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\wraddress_a_bus~1_combout ),
	.cout());
defparam \wraddress_a_bus~1 .lut_mask = 16'hAACC;
defparam \wraddress_a_bus~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wraddress_a_bus~2 (
	.dataa(wr_address_i_int_2),
	.datab(ram_in_reg_2_01),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\wraddress_a_bus~2_combout ),
	.cout());
defparam \wraddress_a_bus~2 .lut_mask = 16'hAACC;
defparam \wraddress_a_bus~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wraddress_a_bus~3 (
	.dataa(wr_address_i_int_3),
	.datab(ram_in_reg_3_01),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\wraddress_a_bus~3_combout ),
	.cout());
defparam \wraddress_a_bus~3 .lut_mask = 16'hAACC;
defparam \wraddress_a_bus~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wraddress_a_bus~4 (
	.dataa(wr_address_i_int_4),
	.datab(ram_in_reg_4_01),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\wraddress_a_bus~4_combout ),
	.cout());
defparam \wraddress_a_bus~4 .lut_mask = 16'hAACC;
defparam \wraddress_a_bus~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wraddress_a_bus~5 (
	.dataa(wr_address_i_int_5),
	.datab(ram_in_reg_5_01),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\wraddress_a_bus~5_combout ),
	.cout());
defparam \wraddress_a_bus~5 .lut_mask = 16'hAACC;
defparam \wraddress_a_bus~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wraddress_a_bus~6 (
	.dataa(wr_address_i_int_6),
	.datab(ram_in_reg_6_01),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\wraddress_a_bus~6_combout ),
	.cout());
defparam \wraddress_a_bus~6 .lut_mask = 16'hAACC;
defparam \wraddress_a_bus~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rdaddress_a_bus~0 (
	.dataa(ram_in_reg_0_02),
	.datab(gnd),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_7),
	.cin(gnd),
	.combout(\rdaddress_a_bus~0_combout ),
	.cout());
defparam \rdaddress_a_bus~0 .lut_mask = 16'hAFFF;
defparam \rdaddress_a_bus~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rdaddress_a_bus~1 (
	.dataa(ram_in_reg_1_02),
	.datab(gnd),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_7),
	.cin(gnd),
	.combout(\rdaddress_a_bus~1_combout ),
	.cout());
defparam \rdaddress_a_bus~1 .lut_mask = 16'hAFFF;
defparam \rdaddress_a_bus~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rdaddress_a_bus~2 (
	.dataa(ram_in_reg_2_02),
	.datab(gnd),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_7),
	.cin(gnd),
	.combout(\rdaddress_a_bus~2_combout ),
	.cout());
defparam \rdaddress_a_bus~2 .lut_mask = 16'hAFFF;
defparam \rdaddress_a_bus~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rdaddress_a_bus~3 (
	.dataa(ram_in_reg_3_02),
	.datab(gnd),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_7),
	.cin(gnd),
	.combout(\rdaddress_a_bus~3_combout ),
	.cout());
defparam \rdaddress_a_bus~3 .lut_mask = 16'hAFFF;
defparam \rdaddress_a_bus~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rdaddress_a_bus~4 (
	.dataa(ram_in_reg_4_02),
	.datab(gnd),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_7),
	.cin(gnd),
	.combout(\rdaddress_a_bus~4_combout ),
	.cout());
defparam \rdaddress_a_bus~4 .lut_mask = 16'hAFFF;
defparam \rdaddress_a_bus~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rdaddress_a_bus~5 (
	.dataa(ram_in_reg_5_02),
	.datab(gnd),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_7),
	.cin(gnd),
	.combout(\rdaddress_a_bus~5_combout ),
	.cout());
defparam \rdaddress_a_bus~5 .lut_mask = 16'hAFFF;
defparam \rdaddress_a_bus~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rdaddress_a_bus~6 (
	.dataa(tdl_arr_6_1),
	.datab(gnd),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_7),
	.cin(gnd),
	.combout(\rdaddress_a_bus~6_combout ),
	.cout());
defparam \rdaddress_a_bus~6 .lut_mask = 16'hAFFF;
defparam \rdaddress_a_bus~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~1 (
	.dataa(ram_in_reg_2_1),
	.datab(data_in_r_2),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~1_combout ),
	.cout());
defparam \b_ram_data_in_bus~1 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wraddress_b_bus~7 (
	.dataa(ram_in_reg_0_11),
	.datab(wr_address_i_int_0),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\wraddress_b_bus~7_combout ),
	.cout());
defparam \wraddress_b_bus~7 .lut_mask = 16'hAACC;
defparam \wraddress_b_bus~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wraddress_b_bus~8 (
	.dataa(ram_in_reg_1_11),
	.datab(wr_address_i_int_1),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\wraddress_b_bus~8_combout ),
	.cout());
defparam \wraddress_b_bus~8 .lut_mask = 16'hAACC;
defparam \wraddress_b_bus~8 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wraddress_b_bus~9 (
	.dataa(ram_in_reg_2_11),
	.datab(wr_address_i_int_2),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\wraddress_b_bus~9_combout ),
	.cout());
defparam \wraddress_b_bus~9 .lut_mask = 16'hAACC;
defparam \wraddress_b_bus~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wraddress_b_bus~10 (
	.dataa(ram_in_reg_3_11),
	.datab(wr_address_i_int_3),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\wraddress_b_bus~10_combout ),
	.cout());
defparam \wraddress_b_bus~10 .lut_mask = 16'hAACC;
defparam \wraddress_b_bus~10 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wraddress_b_bus~11 (
	.dataa(ram_in_reg_4_11),
	.datab(wr_address_i_int_4),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\wraddress_b_bus~11_combout ),
	.cout());
defparam \wraddress_b_bus~11 .lut_mask = 16'hAACC;
defparam \wraddress_b_bus~11 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wraddress_b_bus~12 (
	.dataa(ram_in_reg_5_11),
	.datab(wr_address_i_int_5),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\wraddress_b_bus~12_combout ),
	.cout());
defparam \wraddress_b_bus~12 .lut_mask = 16'hAACC;
defparam \wraddress_b_bus~12 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rdaddress_b_bus~7 (
	.dataa(data_rdy_vec_10),
	.datab(ram_a_not_b_vec_7),
	.datac(ram_in_reg_0_12),
	.datad(gnd),
	.cin(gnd),
	.combout(\rdaddress_b_bus~7_combout ),
	.cout());
defparam \rdaddress_b_bus~7 .lut_mask = 16'hFEFE;
defparam \rdaddress_b_bus~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rdaddress_b_bus~8 (
	.dataa(data_rdy_vec_10),
	.datab(ram_a_not_b_vec_7),
	.datac(ram_in_reg_1_12),
	.datad(gnd),
	.cin(gnd),
	.combout(\rdaddress_b_bus~8_combout ),
	.cout());
defparam \rdaddress_b_bus~8 .lut_mask = 16'hFEFE;
defparam \rdaddress_b_bus~8 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rdaddress_b_bus~9 (
	.dataa(data_rdy_vec_10),
	.datab(ram_a_not_b_vec_7),
	.datac(ram_in_reg_2_12),
	.datad(gnd),
	.cin(gnd),
	.combout(\rdaddress_b_bus~9_combout ),
	.cout());
defparam \rdaddress_b_bus~9 .lut_mask = 16'hFEFE;
defparam \rdaddress_b_bus~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rdaddress_b_bus~10 (
	.dataa(data_rdy_vec_10),
	.datab(ram_a_not_b_vec_7),
	.datac(ram_in_reg_3_12),
	.datad(gnd),
	.cin(gnd),
	.combout(\rdaddress_b_bus~10_combout ),
	.cout());
defparam \rdaddress_b_bus~10 .lut_mask = 16'hFEFE;
defparam \rdaddress_b_bus~10 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rdaddress_b_bus~11 (
	.dataa(data_rdy_vec_10),
	.datab(ram_a_not_b_vec_7),
	.datac(ram_in_reg_4_12),
	.datad(gnd),
	.cin(gnd),
	.combout(\rdaddress_b_bus~11_combout ),
	.cout());
defparam \rdaddress_b_bus~11 .lut_mask = 16'hFEFE;
defparam \rdaddress_b_bus~11 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rdaddress_b_bus~12 (
	.dataa(data_rdy_vec_10),
	.datab(ram_a_not_b_vec_7),
	.datac(ram_in_reg_5_12),
	.datad(gnd),
	.cin(gnd),
	.combout(\rdaddress_b_bus~12_combout ),
	.cout());
defparam \rdaddress_b_bus~12 .lut_mask = 16'hFEFE;
defparam \rdaddress_b_bus~12 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~1 (
	.dataa(data_in_r_2),
	.datab(ram_in_reg_2_1),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~1_combout ),
	.cout());
defparam \a_ram_data_in_bus~1 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wraddress_a_bus~7 (
	.dataa(wr_address_i_int_0),
	.datab(ram_in_reg_0_11),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\wraddress_a_bus~7_combout ),
	.cout());
defparam \wraddress_a_bus~7 .lut_mask = 16'hAACC;
defparam \wraddress_a_bus~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wraddress_a_bus~8 (
	.dataa(wr_address_i_int_1),
	.datab(ram_in_reg_1_11),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\wraddress_a_bus~8_combout ),
	.cout());
defparam \wraddress_a_bus~8 .lut_mask = 16'hAACC;
defparam \wraddress_a_bus~8 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wraddress_a_bus~9 (
	.dataa(wr_address_i_int_2),
	.datab(ram_in_reg_2_11),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\wraddress_a_bus~9_combout ),
	.cout());
defparam \wraddress_a_bus~9 .lut_mask = 16'hAACC;
defparam \wraddress_a_bus~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wraddress_a_bus~10 (
	.dataa(wr_address_i_int_3),
	.datab(ram_in_reg_3_11),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\wraddress_a_bus~10_combout ),
	.cout());
defparam \wraddress_a_bus~10 .lut_mask = 16'hAACC;
defparam \wraddress_a_bus~10 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wraddress_a_bus~11 (
	.dataa(wr_address_i_int_4),
	.datab(ram_in_reg_4_11),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\wraddress_a_bus~11_combout ),
	.cout());
defparam \wraddress_a_bus~11 .lut_mask = 16'hAACC;
defparam \wraddress_a_bus~11 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wraddress_a_bus~12 (
	.dataa(wr_address_i_int_5),
	.datab(ram_in_reg_5_11),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\wraddress_a_bus~12_combout ),
	.cout());
defparam \wraddress_a_bus~12 .lut_mask = 16'hAACC;
defparam \wraddress_a_bus~12 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rdaddress_a_bus~7 (
	.dataa(ram_in_reg_0_12),
	.datab(gnd),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_7),
	.cin(gnd),
	.combout(\rdaddress_a_bus~7_combout ),
	.cout());
defparam \rdaddress_a_bus~7 .lut_mask = 16'hAFFF;
defparam \rdaddress_a_bus~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rdaddress_a_bus~8 (
	.dataa(ram_in_reg_1_12),
	.datab(gnd),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_7),
	.cin(gnd),
	.combout(\rdaddress_a_bus~8_combout ),
	.cout());
defparam \rdaddress_a_bus~8 .lut_mask = 16'hAFFF;
defparam \rdaddress_a_bus~8 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rdaddress_a_bus~9 (
	.dataa(ram_in_reg_2_12),
	.datab(gnd),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_7),
	.cin(gnd),
	.combout(\rdaddress_a_bus~9_combout ),
	.cout());
defparam \rdaddress_a_bus~9 .lut_mask = 16'hAFFF;
defparam \rdaddress_a_bus~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rdaddress_a_bus~10 (
	.dataa(ram_in_reg_3_12),
	.datab(gnd),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_7),
	.cin(gnd),
	.combout(\rdaddress_a_bus~10_combout ),
	.cout());
defparam \rdaddress_a_bus~10 .lut_mask = 16'hAFFF;
defparam \rdaddress_a_bus~10 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rdaddress_a_bus~11 (
	.dataa(ram_in_reg_4_12),
	.datab(gnd),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_7),
	.cin(gnd),
	.combout(\rdaddress_a_bus~11_combout ),
	.cout());
defparam \rdaddress_a_bus~11 .lut_mask = 16'hAFFF;
defparam \rdaddress_a_bus~11 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rdaddress_a_bus~12 (
	.dataa(ram_in_reg_5_12),
	.datab(gnd),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_7),
	.cin(gnd),
	.combout(\rdaddress_a_bus~12_combout ),
	.cout());
defparam \rdaddress_a_bus~12 .lut_mask = 16'hAFFF;
defparam \rdaddress_a_bus~12 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~2 (
	.dataa(ram_in_reg_2_2),
	.datab(data_in_r_2),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~2_combout ),
	.cout());
defparam \b_ram_data_in_bus~2 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wraddress_b_bus~13 (
	.dataa(ram_in_reg_1_21),
	.datab(wr_address_i_int_1),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\wraddress_b_bus~13_combout ),
	.cout());
defparam \wraddress_b_bus~13 .lut_mask = 16'hAACC;
defparam \wraddress_b_bus~13 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wraddress_b_bus~14 (
	.dataa(ram_in_reg_3_21),
	.datab(wr_address_i_int_3),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\wraddress_b_bus~14_combout ),
	.cout());
defparam \wraddress_b_bus~14 .lut_mask = 16'hAACC;
defparam \wraddress_b_bus~14 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wraddress_b_bus~15 (
	.dataa(ram_in_reg_5_21),
	.datab(wr_address_i_int_5),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\wraddress_b_bus~15_combout ),
	.cout());
defparam \wraddress_b_bus~15 .lut_mask = 16'hAACC;
defparam \wraddress_b_bus~15 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rdaddress_b_bus~13 (
	.dataa(data_rdy_vec_10),
	.datab(ram_a_not_b_vec_7),
	.datac(ram_in_reg_1_22),
	.datad(gnd),
	.cin(gnd),
	.combout(\rdaddress_b_bus~13_combout ),
	.cout());
defparam \rdaddress_b_bus~13 .lut_mask = 16'hFEFE;
defparam \rdaddress_b_bus~13 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rdaddress_b_bus~14 (
	.dataa(data_rdy_vec_10),
	.datab(ram_a_not_b_vec_7),
	.datac(ram_in_reg_3_22),
	.datad(gnd),
	.cin(gnd),
	.combout(\rdaddress_b_bus~14_combout ),
	.cout());
defparam \rdaddress_b_bus~14 .lut_mask = 16'hFEFE;
defparam \rdaddress_b_bus~14 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rdaddress_b_bus~15 (
	.dataa(data_rdy_vec_10),
	.datab(ram_a_not_b_vec_7),
	.datac(ram_in_reg_5_22),
	.datad(gnd),
	.cin(gnd),
	.combout(\rdaddress_b_bus~15_combout ),
	.cout());
defparam \rdaddress_b_bus~15 .lut_mask = 16'hFEFE;
defparam \rdaddress_b_bus~15 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~2 (
	.dataa(data_in_r_2),
	.datab(ram_in_reg_2_2),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~2_combout ),
	.cout());
defparam \a_ram_data_in_bus~2 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wraddress_a_bus~13 (
	.dataa(wr_address_i_int_1),
	.datab(ram_in_reg_1_21),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\wraddress_a_bus~13_combout ),
	.cout());
defparam \wraddress_a_bus~13 .lut_mask = 16'hAACC;
defparam \wraddress_a_bus~13 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wraddress_a_bus~14 (
	.dataa(wr_address_i_int_3),
	.datab(ram_in_reg_3_21),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\wraddress_a_bus~14_combout ),
	.cout());
defparam \wraddress_a_bus~14 .lut_mask = 16'hAACC;
defparam \wraddress_a_bus~14 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wraddress_a_bus~15 (
	.dataa(wr_address_i_int_5),
	.datab(ram_in_reg_5_21),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\wraddress_a_bus~15_combout ),
	.cout());
defparam \wraddress_a_bus~15 .lut_mask = 16'hAACC;
defparam \wraddress_a_bus~15 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rdaddress_a_bus~13 (
	.dataa(ram_in_reg_1_22),
	.datab(gnd),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_7),
	.cin(gnd),
	.combout(\rdaddress_a_bus~13_combout ),
	.cout());
defparam \rdaddress_a_bus~13 .lut_mask = 16'hAFFF;
defparam \rdaddress_a_bus~13 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rdaddress_a_bus~14 (
	.dataa(ram_in_reg_3_22),
	.datab(gnd),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_7),
	.cin(gnd),
	.combout(\rdaddress_a_bus~14_combout ),
	.cout());
defparam \rdaddress_a_bus~14 .lut_mask = 16'hAFFF;
defparam \rdaddress_a_bus~14 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rdaddress_a_bus~15 (
	.dataa(ram_in_reg_5_22),
	.datab(gnd),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_7),
	.cin(gnd),
	.combout(\rdaddress_a_bus~15_combout ),
	.cout());
defparam \rdaddress_a_bus~15 .lut_mask = 16'hAFFF;
defparam \rdaddress_a_bus~15 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~3 (
	.dataa(ram_in_reg_2_3),
	.datab(data_in_r_2),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~3_combout ),
	.cout());
defparam \b_ram_data_in_bus~3 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wraddress_b_bus~16 (
	.dataa(ram_in_reg_1_31),
	.datab(wr_address_i_int_1),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\wraddress_b_bus~16_combout ),
	.cout());
defparam \wraddress_b_bus~16 .lut_mask = 16'hAACC;
defparam \wraddress_b_bus~16 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wraddress_b_bus~17 (
	.dataa(ram_in_reg_3_31),
	.datab(wr_address_i_int_3),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\wraddress_b_bus~17_combout ),
	.cout());
defparam \wraddress_b_bus~17 .lut_mask = 16'hAACC;
defparam \wraddress_b_bus~17 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wraddress_b_bus~18 (
	.dataa(ram_in_reg_5_31),
	.datab(wr_address_i_int_5),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\wraddress_b_bus~18_combout ),
	.cout());
defparam \wraddress_b_bus~18 .lut_mask = 16'hAACC;
defparam \wraddress_b_bus~18 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rdaddress_b_bus~16 (
	.dataa(data_rdy_vec_10),
	.datab(ram_a_not_b_vec_7),
	.datac(ram_in_reg_1_32),
	.datad(gnd),
	.cin(gnd),
	.combout(\rdaddress_b_bus~16_combout ),
	.cout());
defparam \rdaddress_b_bus~16 .lut_mask = 16'hFEFE;
defparam \rdaddress_b_bus~16 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rdaddress_b_bus~17 (
	.dataa(data_rdy_vec_10),
	.datab(ram_a_not_b_vec_7),
	.datac(ram_in_reg_3_32),
	.datad(gnd),
	.cin(gnd),
	.combout(\rdaddress_b_bus~17_combout ),
	.cout());
defparam \rdaddress_b_bus~17 .lut_mask = 16'hFEFE;
defparam \rdaddress_b_bus~17 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rdaddress_b_bus~18 (
	.dataa(data_rdy_vec_10),
	.datab(ram_a_not_b_vec_7),
	.datac(ram_in_reg_5_32),
	.datad(gnd),
	.cin(gnd),
	.combout(\rdaddress_b_bus~18_combout ),
	.cout());
defparam \rdaddress_b_bus~18 .lut_mask = 16'hFEFE;
defparam \rdaddress_b_bus~18 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~3 (
	.dataa(data_in_r_2),
	.datab(ram_in_reg_2_3),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~3_combout ),
	.cout());
defparam \a_ram_data_in_bus~3 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wraddress_a_bus~16 (
	.dataa(wr_address_i_int_1),
	.datab(ram_in_reg_1_31),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\wraddress_a_bus~16_combout ),
	.cout());
defparam \wraddress_a_bus~16 .lut_mask = 16'hAACC;
defparam \wraddress_a_bus~16 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wraddress_a_bus~17 (
	.dataa(wr_address_i_int_3),
	.datab(ram_in_reg_3_31),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\wraddress_a_bus~17_combout ),
	.cout());
defparam \wraddress_a_bus~17 .lut_mask = 16'hAACC;
defparam \wraddress_a_bus~17 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wraddress_a_bus~18 (
	.dataa(wr_address_i_int_5),
	.datab(ram_in_reg_5_31),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\wraddress_a_bus~18_combout ),
	.cout());
defparam \wraddress_a_bus~18 .lut_mask = 16'hAACC;
defparam \wraddress_a_bus~18 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rdaddress_a_bus~16 (
	.dataa(ram_in_reg_1_32),
	.datab(gnd),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_7),
	.cin(gnd),
	.combout(\rdaddress_a_bus~16_combout ),
	.cout());
defparam \rdaddress_a_bus~16 .lut_mask = 16'hAFFF;
defparam \rdaddress_a_bus~16 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rdaddress_a_bus~17 (
	.dataa(ram_in_reg_3_32),
	.datab(gnd),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_7),
	.cin(gnd),
	.combout(\rdaddress_a_bus~17_combout ),
	.cout());
defparam \rdaddress_a_bus~17 .lut_mask = 16'hAFFF;
defparam \rdaddress_a_bus~17 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rdaddress_a_bus~18 (
	.dataa(ram_in_reg_5_32),
	.datab(gnd),
	.datac(data_rdy_vec_10),
	.datad(ram_a_not_b_vec_7),
	.cin(gnd),
	.combout(\rdaddress_a_bus~18_combout ),
	.cout());
defparam \rdaddress_a_bus~18 .lut_mask = 16'hAFFF;
defparam \rdaddress_a_bus~18 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~4 (
	.dataa(ram_in_reg_6_0),
	.datab(data_in_r_6),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~4_combout ),
	.cout());
defparam \b_ram_data_in_bus~4 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~4 (
	.dataa(data_in_r_6),
	.datab(ram_in_reg_6_0),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~4_combout ),
	.cout());
defparam \a_ram_data_in_bus~4 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~5 (
	.dataa(ram_in_reg_6_1),
	.datab(data_in_r_6),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~5_combout ),
	.cout());
defparam \b_ram_data_in_bus~5 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~5 (
	.dataa(data_in_r_6),
	.datab(ram_in_reg_6_1),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~5_combout ),
	.cout());
defparam \a_ram_data_in_bus~5 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~6 (
	.dataa(ram_in_reg_6_2),
	.datab(data_in_r_6),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~6_combout ),
	.cout());
defparam \b_ram_data_in_bus~6 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~6 (
	.dataa(data_in_r_6),
	.datab(ram_in_reg_6_2),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~6_combout ),
	.cout());
defparam \a_ram_data_in_bus~6 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~7 (
	.dataa(ram_in_reg_6_3),
	.datab(data_in_r_6),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~7_combout ),
	.cout());
defparam \b_ram_data_in_bus~7 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~7 (
	.dataa(data_in_r_6),
	.datab(ram_in_reg_6_3),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~7_combout ),
	.cout());
defparam \a_ram_data_in_bus~7 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~8 (
	.dataa(ram_in_reg_4_0),
	.datab(data_in_r_4),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~8_combout ),
	.cout());
defparam \b_ram_data_in_bus~8 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~8 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~8 (
	.dataa(data_in_r_4),
	.datab(ram_in_reg_4_0),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~8_combout ),
	.cout());
defparam \a_ram_data_in_bus~8 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~8 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~9 (
	.dataa(ram_in_reg_4_1),
	.datab(data_in_r_4),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~9_combout ),
	.cout());
defparam \b_ram_data_in_bus~9 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~9 (
	.dataa(data_in_r_4),
	.datab(ram_in_reg_4_1),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~9_combout ),
	.cout());
defparam \a_ram_data_in_bus~9 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~10 (
	.dataa(ram_in_reg_4_2),
	.datab(data_in_r_4),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~10_combout ),
	.cout());
defparam \b_ram_data_in_bus~10 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~10 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~10 (
	.dataa(data_in_r_4),
	.datab(ram_in_reg_4_2),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~10_combout ),
	.cout());
defparam \a_ram_data_in_bus~10 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~10 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~11 (
	.dataa(ram_in_reg_4_3),
	.datab(data_in_r_4),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~11_combout ),
	.cout());
defparam \b_ram_data_in_bus~11 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~11 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~11 (
	.dataa(data_in_r_4),
	.datab(ram_in_reg_4_3),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~11_combout ),
	.cout());
defparam \a_ram_data_in_bus~11 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~11 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~12 (
	.dataa(ram_in_reg_3_0),
	.datab(data_in_r_3),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~12_combout ),
	.cout());
defparam \b_ram_data_in_bus~12 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~12 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~12 (
	.dataa(data_in_r_3),
	.datab(ram_in_reg_3_0),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~12_combout ),
	.cout());
defparam \a_ram_data_in_bus~12 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~12 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~13 (
	.dataa(ram_in_reg_3_1),
	.datab(data_in_r_3),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~13_combout ),
	.cout());
defparam \b_ram_data_in_bus~13 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~13 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~13 (
	.dataa(data_in_r_3),
	.datab(ram_in_reg_3_1),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~13_combout ),
	.cout());
defparam \a_ram_data_in_bus~13 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~13 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~14 (
	.dataa(ram_in_reg_3_2),
	.datab(data_in_r_3),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~14_combout ),
	.cout());
defparam \b_ram_data_in_bus~14 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~14 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~14 (
	.dataa(data_in_r_3),
	.datab(ram_in_reg_3_2),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~14_combout ),
	.cout());
defparam \a_ram_data_in_bus~14 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~14 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~15 (
	.dataa(ram_in_reg_3_3),
	.datab(data_in_r_3),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~15_combout ),
	.cout());
defparam \b_ram_data_in_bus~15 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~15 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~15 (
	.dataa(data_in_r_3),
	.datab(ram_in_reg_3_3),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~15_combout ),
	.cout());
defparam \a_ram_data_in_bus~15 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~15 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~16 (
	.dataa(ram_in_reg_5_0),
	.datab(data_in_r_5),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~16_combout ),
	.cout());
defparam \b_ram_data_in_bus~16 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~16 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~16 (
	.dataa(data_in_r_5),
	.datab(ram_in_reg_5_0),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~16_combout ),
	.cout());
defparam \a_ram_data_in_bus~16 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~16 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~17 (
	.dataa(ram_in_reg_5_1),
	.datab(data_in_r_5),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~17_combout ),
	.cout());
defparam \b_ram_data_in_bus~17 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~17 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~17 (
	.dataa(data_in_r_5),
	.datab(ram_in_reg_5_1),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~17_combout ),
	.cout());
defparam \a_ram_data_in_bus~17 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~17 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~18 (
	.dataa(ram_in_reg_5_2),
	.datab(data_in_r_5),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~18_combout ),
	.cout());
defparam \b_ram_data_in_bus~18 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~18 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~18 (
	.dataa(data_in_r_5),
	.datab(ram_in_reg_5_2),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~18_combout ),
	.cout());
defparam \a_ram_data_in_bus~18 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~18 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~19 (
	.dataa(ram_in_reg_5_3),
	.datab(data_in_r_5),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~19_combout ),
	.cout());
defparam \b_ram_data_in_bus~19 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~19 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~19 (
	.dataa(data_in_r_5),
	.datab(ram_in_reg_5_3),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~19_combout ),
	.cout());
defparam \a_ram_data_in_bus~19 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~19 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~20 (
	.dataa(ram_in_reg_1_0),
	.datab(data_in_r_1),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~20_combout ),
	.cout());
defparam \b_ram_data_in_bus~20 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~20 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~20 (
	.dataa(data_in_r_1),
	.datab(ram_in_reg_1_0),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~20_combout ),
	.cout());
defparam \a_ram_data_in_bus~20 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~20 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~21 (
	.dataa(ram_in_reg_1_1),
	.datab(data_in_r_1),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~21_combout ),
	.cout());
defparam \b_ram_data_in_bus~21 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~21 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~21 (
	.dataa(data_in_r_1),
	.datab(ram_in_reg_1_1),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~21_combout ),
	.cout());
defparam \a_ram_data_in_bus~21 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~21 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~22 (
	.dataa(ram_in_reg_1_2),
	.datab(data_in_r_1),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~22_combout ),
	.cout());
defparam \b_ram_data_in_bus~22 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~22 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~22 (
	.dataa(data_in_r_1),
	.datab(ram_in_reg_1_2),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~22_combout ),
	.cout());
defparam \a_ram_data_in_bus~22 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~22 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~23 (
	.dataa(ram_in_reg_1_3),
	.datab(data_in_r_1),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~23_combout ),
	.cout());
defparam \b_ram_data_in_bus~23 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~23 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~23 (
	.dataa(data_in_r_1),
	.datab(ram_in_reg_1_3),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~23_combout ),
	.cout());
defparam \a_ram_data_in_bus~23 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~23 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~24 (
	.dataa(ram_in_reg_0_0),
	.datab(data_in_r_0),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~24_combout ),
	.cout());
defparam \b_ram_data_in_bus~24 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~24 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~24 (
	.dataa(data_in_r_0),
	.datab(ram_in_reg_0_0),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~24_combout ),
	.cout());
defparam \a_ram_data_in_bus~24 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~24 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~25 (
	.dataa(ram_in_reg_0_1),
	.datab(data_in_r_0),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~25_combout ),
	.cout());
defparam \b_ram_data_in_bus~25 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~25 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~25 (
	.dataa(data_in_r_0),
	.datab(ram_in_reg_0_1),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~25_combout ),
	.cout());
defparam \a_ram_data_in_bus~25 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~25 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~26 (
	.dataa(ram_in_reg_0_2),
	.datab(data_in_r_0),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~26_combout ),
	.cout());
defparam \b_ram_data_in_bus~26 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~26 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~26 (
	.dataa(data_in_r_0),
	.datab(ram_in_reg_0_2),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~26_combout ),
	.cout());
defparam \a_ram_data_in_bus~26 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~26 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~27 (
	.dataa(ram_in_reg_0_3),
	.datab(data_in_r_0),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~27_combout ),
	.cout());
defparam \b_ram_data_in_bus~27 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~27 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~27 (
	.dataa(data_in_r_0),
	.datab(ram_in_reg_0_3),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~27_combout ),
	.cout());
defparam \a_ram_data_in_bus~27 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~27 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~28 (
	.dataa(ram_in_reg_7_0),
	.datab(data_in_r_7),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~28_combout ),
	.cout());
defparam \b_ram_data_in_bus~28 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~28 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~28 (
	.dataa(data_in_r_7),
	.datab(ram_in_reg_7_0),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~28_combout ),
	.cout());
defparam \a_ram_data_in_bus~28 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~28 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~29 (
	.dataa(ram_in_reg_7_1),
	.datab(data_in_r_7),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~29_combout ),
	.cout());
defparam \b_ram_data_in_bus~29 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~29 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~29 (
	.dataa(data_in_r_7),
	.datab(ram_in_reg_7_1),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~29_combout ),
	.cout());
defparam \a_ram_data_in_bus~29 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~29 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~30 (
	.dataa(ram_in_reg_7_2),
	.datab(data_in_r_7),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~30_combout ),
	.cout());
defparam \b_ram_data_in_bus~30 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~30 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~30 (
	.dataa(data_in_r_7),
	.datab(ram_in_reg_7_2),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~30_combout ),
	.cout());
defparam \a_ram_data_in_bus~30 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~30 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~31 (
	.dataa(ram_in_reg_7_3),
	.datab(data_in_r_7),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~31_combout ),
	.cout());
defparam \b_ram_data_in_bus~31 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~31 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~31 (
	.dataa(data_in_r_7),
	.datab(ram_in_reg_7_3),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~31_combout ),
	.cout());
defparam \a_ram_data_in_bus~31 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~31 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~32 (
	.dataa(ram_in_reg_7_4),
	.datab(data_in_i_7),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~32_combout ),
	.cout());
defparam \b_ram_data_in_bus~32 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~32 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~32 (
	.dataa(data_in_i_7),
	.datab(ram_in_reg_7_4),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~32_combout ),
	.cout());
defparam \a_ram_data_in_bus~32 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~32 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~33 (
	.dataa(ram_in_reg_7_5),
	.datab(data_in_i_7),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~33_combout ),
	.cout());
defparam \b_ram_data_in_bus~33 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~33 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~33 (
	.dataa(data_in_i_7),
	.datab(ram_in_reg_7_5),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~33_combout ),
	.cout());
defparam \a_ram_data_in_bus~33 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~33 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~34 (
	.dataa(ram_in_reg_7_6),
	.datab(data_in_i_7),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~34_combout ),
	.cout());
defparam \b_ram_data_in_bus~34 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~34 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~34 (
	.dataa(data_in_i_7),
	.datab(ram_in_reg_7_6),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~34_combout ),
	.cout());
defparam \a_ram_data_in_bus~34 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~34 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~35 (
	.dataa(ram_in_reg_7_7),
	.datab(data_in_i_7),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~35_combout ),
	.cout());
defparam \b_ram_data_in_bus~35 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~35 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~35 (
	.dataa(data_in_i_7),
	.datab(ram_in_reg_7_7),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~35_combout ),
	.cout());
defparam \a_ram_data_in_bus~35 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~35 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~36 (
	.dataa(ram_in_reg_3_4),
	.datab(data_in_i_3),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~36_combout ),
	.cout());
defparam \b_ram_data_in_bus~36 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~36 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~36 (
	.dataa(data_in_i_3),
	.datab(ram_in_reg_3_4),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~36_combout ),
	.cout());
defparam \a_ram_data_in_bus~36 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~36 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~37 (
	.dataa(ram_in_reg_3_5),
	.datab(data_in_i_3),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~37_combout ),
	.cout());
defparam \b_ram_data_in_bus~37 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~37 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~37 (
	.dataa(data_in_i_3),
	.datab(ram_in_reg_3_5),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~37_combout ),
	.cout());
defparam \a_ram_data_in_bus~37 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~37 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~38 (
	.dataa(ram_in_reg_3_6),
	.datab(data_in_i_3),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~38_combout ),
	.cout());
defparam \b_ram_data_in_bus~38 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~38 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~38 (
	.dataa(data_in_i_3),
	.datab(ram_in_reg_3_6),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~38_combout ),
	.cout());
defparam \a_ram_data_in_bus~38 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~38 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~39 (
	.dataa(ram_in_reg_3_7),
	.datab(data_in_i_3),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~39_combout ),
	.cout());
defparam \b_ram_data_in_bus~39 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~39 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~39 (
	.dataa(data_in_i_3),
	.datab(ram_in_reg_3_7),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~39_combout ),
	.cout());
defparam \a_ram_data_in_bus~39 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~39 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~40 (
	.dataa(ram_in_reg_5_4),
	.datab(data_in_i_5),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~40_combout ),
	.cout());
defparam \b_ram_data_in_bus~40 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~40 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~40 (
	.dataa(data_in_i_5),
	.datab(ram_in_reg_5_4),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~40_combout ),
	.cout());
defparam \a_ram_data_in_bus~40 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~40 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~41 (
	.dataa(ram_in_reg_5_5),
	.datab(data_in_i_5),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~41_combout ),
	.cout());
defparam \b_ram_data_in_bus~41 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~41 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~41 (
	.dataa(data_in_i_5),
	.datab(ram_in_reg_5_5),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~41_combout ),
	.cout());
defparam \a_ram_data_in_bus~41 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~41 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~42 (
	.dataa(ram_in_reg_5_6),
	.datab(data_in_i_5),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~42_combout ),
	.cout());
defparam \b_ram_data_in_bus~42 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~42 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~42 (
	.dataa(data_in_i_5),
	.datab(ram_in_reg_5_6),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~42_combout ),
	.cout());
defparam \a_ram_data_in_bus~42 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~42 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~43 (
	.dataa(ram_in_reg_5_7),
	.datab(data_in_i_5),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~43_combout ),
	.cout());
defparam \b_ram_data_in_bus~43 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~43 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~43 (
	.dataa(data_in_i_5),
	.datab(ram_in_reg_5_7),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~43_combout ),
	.cout());
defparam \a_ram_data_in_bus~43 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~43 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~44 (
	.dataa(ram_in_reg_4_4),
	.datab(data_in_i_4),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~44_combout ),
	.cout());
defparam \b_ram_data_in_bus~44 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~44 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~44 (
	.dataa(data_in_i_4),
	.datab(ram_in_reg_4_4),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~44_combout ),
	.cout());
defparam \a_ram_data_in_bus~44 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~44 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~45 (
	.dataa(ram_in_reg_4_5),
	.datab(data_in_i_4),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~45_combout ),
	.cout());
defparam \b_ram_data_in_bus~45 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~45 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~45 (
	.dataa(data_in_i_4),
	.datab(ram_in_reg_4_5),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~45_combout ),
	.cout());
defparam \a_ram_data_in_bus~45 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~45 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~46 (
	.dataa(ram_in_reg_4_6),
	.datab(data_in_i_4),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~46_combout ),
	.cout());
defparam \b_ram_data_in_bus~46 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~46 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~46 (
	.dataa(data_in_i_4),
	.datab(ram_in_reg_4_6),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~46_combout ),
	.cout());
defparam \a_ram_data_in_bus~46 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~46 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~47 (
	.dataa(ram_in_reg_4_7),
	.datab(data_in_i_4),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~47_combout ),
	.cout());
defparam \b_ram_data_in_bus~47 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~47 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~47 (
	.dataa(data_in_i_4),
	.datab(ram_in_reg_4_7),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~47_combout ),
	.cout());
defparam \a_ram_data_in_bus~47 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~47 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~48 (
	.dataa(ram_in_reg_6_4),
	.datab(data_in_i_6),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~48_combout ),
	.cout());
defparam \b_ram_data_in_bus~48 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~48 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~48 (
	.dataa(data_in_i_6),
	.datab(ram_in_reg_6_4),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~48_combout ),
	.cout());
defparam \a_ram_data_in_bus~48 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~48 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~49 (
	.dataa(ram_in_reg_6_5),
	.datab(data_in_i_6),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~49_combout ),
	.cout());
defparam \b_ram_data_in_bus~49 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~49 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~49 (
	.dataa(data_in_i_6),
	.datab(ram_in_reg_6_5),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~49_combout ),
	.cout());
defparam \a_ram_data_in_bus~49 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~49 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~50 (
	.dataa(ram_in_reg_6_6),
	.datab(data_in_i_6),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~50_combout ),
	.cout());
defparam \b_ram_data_in_bus~50 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~50 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~50 (
	.dataa(data_in_i_6),
	.datab(ram_in_reg_6_6),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~50_combout ),
	.cout());
defparam \a_ram_data_in_bus~50 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~50 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~51 (
	.dataa(ram_in_reg_6_7),
	.datab(data_in_i_6),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~51_combout ),
	.cout());
defparam \b_ram_data_in_bus~51 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~51 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~51 (
	.dataa(data_in_i_6),
	.datab(ram_in_reg_6_7),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~51_combout ),
	.cout());
defparam \a_ram_data_in_bus~51 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~51 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~52 (
	.dataa(ram_in_reg_2_4),
	.datab(data_in_i_2),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~52_combout ),
	.cout());
defparam \b_ram_data_in_bus~52 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~52 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~52 (
	.dataa(data_in_i_2),
	.datab(ram_in_reg_2_4),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~52_combout ),
	.cout());
defparam \a_ram_data_in_bus~52 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~52 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~53 (
	.dataa(ram_in_reg_2_5),
	.datab(data_in_i_2),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~53_combout ),
	.cout());
defparam \b_ram_data_in_bus~53 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~53 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~53 (
	.dataa(data_in_i_2),
	.datab(ram_in_reg_2_5),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~53_combout ),
	.cout());
defparam \a_ram_data_in_bus~53 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~53 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~54 (
	.dataa(ram_in_reg_2_6),
	.datab(data_in_i_2),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~54_combout ),
	.cout());
defparam \b_ram_data_in_bus~54 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~54 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~54 (
	.dataa(data_in_i_2),
	.datab(ram_in_reg_2_6),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~54_combout ),
	.cout());
defparam \a_ram_data_in_bus~54 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~54 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~55 (
	.dataa(ram_in_reg_2_7),
	.datab(data_in_i_2),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~55_combout ),
	.cout());
defparam \b_ram_data_in_bus~55 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~55 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~55 (
	.dataa(data_in_i_2),
	.datab(ram_in_reg_2_7),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~55_combout ),
	.cout());
defparam \a_ram_data_in_bus~55 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~55 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~56 (
	.dataa(ram_in_reg_1_4),
	.datab(data_in_i_1),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~56_combout ),
	.cout());
defparam \b_ram_data_in_bus~56 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~56 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~56 (
	.dataa(data_in_i_1),
	.datab(ram_in_reg_1_4),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~56_combout ),
	.cout());
defparam \a_ram_data_in_bus~56 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~56 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~57 (
	.dataa(ram_in_reg_1_5),
	.datab(data_in_i_1),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~57_combout ),
	.cout());
defparam \b_ram_data_in_bus~57 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~57 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~57 (
	.dataa(data_in_i_1),
	.datab(ram_in_reg_1_5),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~57_combout ),
	.cout());
defparam \a_ram_data_in_bus~57 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~57 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~58 (
	.dataa(ram_in_reg_1_6),
	.datab(data_in_i_1),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~58_combout ),
	.cout());
defparam \b_ram_data_in_bus~58 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~58 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~58 (
	.dataa(data_in_i_1),
	.datab(ram_in_reg_1_6),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~58_combout ),
	.cout());
defparam \a_ram_data_in_bus~58 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~58 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~59 (
	.dataa(ram_in_reg_1_7),
	.datab(data_in_i_1),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~59_combout ),
	.cout());
defparam \b_ram_data_in_bus~59 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~59 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~59 (
	.dataa(data_in_i_1),
	.datab(ram_in_reg_1_7),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~59_combout ),
	.cout());
defparam \a_ram_data_in_bus~59 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~59 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~60 (
	.dataa(ram_in_reg_0_4),
	.datab(data_in_i_0),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~60_combout ),
	.cout());
defparam \b_ram_data_in_bus~60 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~60 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~60 (
	.dataa(data_in_i_0),
	.datab(ram_in_reg_0_4),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~60_combout ),
	.cout());
defparam \a_ram_data_in_bus~60 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~60 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~61 (
	.dataa(ram_in_reg_0_5),
	.datab(data_in_i_0),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~61_combout ),
	.cout());
defparam \b_ram_data_in_bus~61 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~61 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~61 (
	.dataa(data_in_i_0),
	.datab(ram_in_reg_0_5),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~61_combout ),
	.cout());
defparam \a_ram_data_in_bus~61 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~61 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~62 (
	.dataa(ram_in_reg_0_6),
	.datab(data_in_i_0),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~62_combout ),
	.cout());
defparam \b_ram_data_in_bus~62 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~62 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~62 (
	.dataa(data_in_i_0),
	.datab(ram_in_reg_0_6),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~62_combout ),
	.cout());
defparam \a_ram_data_in_bus~62 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~62 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \b_ram_data_in_bus~63 (
	.dataa(ram_in_reg_0_7),
	.datab(data_in_i_0),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\b_ram_data_in_bus~63_combout ),
	.cout());
defparam \b_ram_data_in_bus~63 .lut_mask = 16'hAACC;
defparam \b_ram_data_in_bus~63 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a_ram_data_in_bus~63 (
	.dataa(data_in_i_0),
	.datab(ram_in_reg_0_7),
	.datac(gnd),
	.datad(ram_a_not_b_vec_1),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~63_combout ),
	.cout());
defparam \a_ram_data_in_bus~63 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~63 .sum_lutc_input = "datac";

endmodule

module fft_asj_fft_cxb_addr_fft_120 (
	sw_0,
	global_clock_enable,
	ram_in_reg_0_0,
	ram_in_reg_1_0,
	ram_in_reg_2_0,
	ram_in_reg_3_0,
	ram_in_reg_4_0,
	ram_in_reg_5_0,
	ram_in_reg_6_1,
	rd_addr_b_0,
	rd_addr_b_1,
	rd_addr_b_2,
	rd_addr_b_3,
	rd_addr_b_4,
	rd_addr_b_5,
	rd_addr_b_6,
	clk)/* synthesis synthesis_greybox=1 */;
input 	sw_0;
input 	global_clock_enable;
output 	ram_in_reg_0_0;
output 	ram_in_reg_1_0;
output 	ram_in_reg_2_0;
output 	ram_in_reg_3_0;
output 	ram_in_reg_4_0;
output 	ram_in_reg_5_0;
output 	ram_in_reg_6_1;
input 	rd_addr_b_0;
input 	rd_addr_b_1;
input 	rd_addr_b_2;
input 	rd_addr_b_3;
input 	rd_addr_b_4;
input 	rd_addr_b_5;
input 	rd_addr_b_6;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Mux7~0_combout ;


dffeas \ram_in_reg[0][0] (
	.clk(clk),
	.d(rd_addr_b_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_0_0),
	.prn(vcc));
defparam \ram_in_reg[0][0] .is_wysiwyg = "true";
defparam \ram_in_reg[0][0] .power_up = "low";

dffeas \ram_in_reg[0][1] (
	.clk(clk),
	.d(rd_addr_b_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_1_0),
	.prn(vcc));
defparam \ram_in_reg[0][1] .is_wysiwyg = "true";
defparam \ram_in_reg[0][1] .power_up = "low";

dffeas \ram_in_reg[0][2] (
	.clk(clk),
	.d(rd_addr_b_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_2_0),
	.prn(vcc));
defparam \ram_in_reg[0][2] .is_wysiwyg = "true";
defparam \ram_in_reg[0][2] .power_up = "low";

dffeas \ram_in_reg[0][3] (
	.clk(clk),
	.d(rd_addr_b_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_3_0),
	.prn(vcc));
defparam \ram_in_reg[0][3] .is_wysiwyg = "true";
defparam \ram_in_reg[0][3] .power_up = "low";

dffeas \ram_in_reg[0][4] (
	.clk(clk),
	.d(rd_addr_b_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_4_0),
	.prn(vcc));
defparam \ram_in_reg[0][4] .is_wysiwyg = "true";
defparam \ram_in_reg[0][4] .power_up = "low";

dffeas \ram_in_reg[0][5] (
	.clk(clk),
	.d(rd_addr_b_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_5_0),
	.prn(vcc));
defparam \ram_in_reg[0][5] .is_wysiwyg = "true";
defparam \ram_in_reg[0][5] .power_up = "low";

dffeas \ram_in_reg[1][6] (
	.clk(clk),
	.d(\Mux7~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_6_1),
	.prn(vcc));
defparam \ram_in_reg[1][6] .is_wysiwyg = "true";
defparam \ram_in_reg[1][6] .power_up = "low";

cycloneiii_lcell_comb \Mux7~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(rd_addr_b_6),
	.datad(sw_0),
	.cin(gnd),
	.combout(\Mux7~0_combout ),
	.cout());
defparam \Mux7~0 .lut_mask = 16'h0FF0;
defparam \Mux7~0 .sum_lutc_input = "datac";

endmodule

module fft_asj_fft_cxb_addr_fft_120_1 (
	global_clock_enable,
	ram_in_reg_0_0,
	ram_in_reg_1_2,
	ram_in_reg_2_0,
	ram_in_reg_3_2,
	ram_in_reg_4_0,
	ram_in_reg_5_2,
	ram_in_reg_6_0,
	ram_in_reg_0_1,
	ram_in_reg_1_1,
	ram_in_reg_2_1,
	ram_in_reg_3_1,
	ram_in_reg_4_1,
	ram_in_reg_5_1,
	ram_in_reg_1_0,
	ram_in_reg_3_0,
	ram_in_reg_5_0,
	ram_in_reg_1_3,
	ram_in_reg_3_3,
	ram_in_reg_5_3,
	swa_tdl_0_0,
	swa_tdl_1_0,
	sw_3_in,
	sw_2_in,
	sw_1_in,
	clk)/* synthesis synthesis_greybox=1 */;
input 	global_clock_enable;
output 	ram_in_reg_0_0;
output 	ram_in_reg_1_2;
output 	ram_in_reg_2_0;
output 	ram_in_reg_3_2;
output 	ram_in_reg_4_0;
output 	ram_in_reg_5_2;
output 	ram_in_reg_6_0;
output 	ram_in_reg_0_1;
output 	ram_in_reg_1_1;
output 	ram_in_reg_2_1;
output 	ram_in_reg_3_1;
output 	ram_in_reg_4_1;
output 	ram_in_reg_5_1;
output 	ram_in_reg_1_0;
output 	ram_in_reg_3_0;
output 	ram_in_reg_5_0;
output 	ram_in_reg_1_3;
output 	ram_in_reg_3_3;
output 	ram_in_reg_5_3;
input 	swa_tdl_0_0;
input 	swa_tdl_1_0;
input 	[6:0] sw_3_in;
input 	[6:0] sw_2_in;
input 	[6:0] sw_1_in;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \sw_3_arr[0][0]~q ;
wire \sw_2_arr[0][0]~q ;
wire \Mux6~0_combout ;
wire \sw_3_arr[0][1]~q ;
wire \sw_1_arr[0][1]~q ;
wire \Mux19~0_combout ;
wire \sw_3_arr[0][2]~q ;
wire \sw_2_arr[0][2]~q ;
wire \Mux4~0_combout ;
wire \sw_3_arr[0][3]~q ;
wire \sw_1_arr[0][3]~q ;
wire \Mux17~0_combout ;
wire \sw_3_arr[0][4]~q ;
wire \sw_2_arr[0][4]~q ;
wire \Mux2~0_combout ;
wire \sw_3_arr[0][5]~q ;
wire \sw_1_arr[0][5]~q ;
wire \Mux15~0_combout ;
wire \sw_3_arr[0][6]~q ;
wire \Mux13~0_combout ;
wire \Mux5~0_combout ;
wire \Mux11~0_combout ;
wire \Mux3~0_combout ;
wire \Mux9~0_combout ;
wire \Mux1~0_combout ;
wire \Mux5~1_combout ;
wire \Mux3~1_combout ;
wire \Mux1~1_combout ;
wire \Mux5~2_combout ;
wire \Mux3~2_combout ;
wire \Mux1~2_combout ;


dffeas \ram_in_reg[0][0] (
	.clk(clk),
	.d(\Mux6~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_0_0),
	.prn(vcc));
defparam \ram_in_reg[0][0] .is_wysiwyg = "true";
defparam \ram_in_reg[0][0] .power_up = "low";

dffeas \ram_in_reg[2][1] (
	.clk(clk),
	.d(\Mux19~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_1_2),
	.prn(vcc));
defparam \ram_in_reg[2][1] .is_wysiwyg = "true";
defparam \ram_in_reg[2][1] .power_up = "low";

dffeas \ram_in_reg[0][2] (
	.clk(clk),
	.d(\Mux4~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_2_0),
	.prn(vcc));
defparam \ram_in_reg[0][2] .is_wysiwyg = "true";
defparam \ram_in_reg[0][2] .power_up = "low";

dffeas \ram_in_reg[2][3] (
	.clk(clk),
	.d(\Mux17~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_3_2),
	.prn(vcc));
defparam \ram_in_reg[2][3] .is_wysiwyg = "true";
defparam \ram_in_reg[2][3] .power_up = "low";

dffeas \ram_in_reg[0][4] (
	.clk(clk),
	.d(\Mux2~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_4_0),
	.prn(vcc));
defparam \ram_in_reg[0][4] .is_wysiwyg = "true";
defparam \ram_in_reg[0][4] .power_up = "low";

dffeas \ram_in_reg[2][5] (
	.clk(clk),
	.d(\Mux15~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_5_2),
	.prn(vcc));
defparam \ram_in_reg[2][5] .is_wysiwyg = "true";
defparam \ram_in_reg[2][5] .power_up = "low";

dffeas \ram_in_reg[0][6] (
	.clk(clk),
	.d(\sw_3_arr[0][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_6_0),
	.prn(vcc));
defparam \ram_in_reg[0][6] .is_wysiwyg = "true";
defparam \ram_in_reg[0][6] .power_up = "low";

dffeas \ram_in_reg[1][0] (
	.clk(clk),
	.d(\Mux13~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_0_1),
	.prn(vcc));
defparam \ram_in_reg[1][0] .is_wysiwyg = "true";
defparam \ram_in_reg[1][0] .power_up = "low";

dffeas \ram_in_reg[1][1] (
	.clk(clk),
	.d(\Mux5~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_1_1),
	.prn(vcc));
defparam \ram_in_reg[1][1] .is_wysiwyg = "true";
defparam \ram_in_reg[1][1] .power_up = "low";

dffeas \ram_in_reg[1][2] (
	.clk(clk),
	.d(\Mux11~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_2_1),
	.prn(vcc));
defparam \ram_in_reg[1][2] .is_wysiwyg = "true";
defparam \ram_in_reg[1][2] .power_up = "low";

dffeas \ram_in_reg[1][3] (
	.clk(clk),
	.d(\Mux3~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_3_1),
	.prn(vcc));
defparam \ram_in_reg[1][3] .is_wysiwyg = "true";
defparam \ram_in_reg[1][3] .power_up = "low";

dffeas \ram_in_reg[1][4] (
	.clk(clk),
	.d(\Mux9~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_4_1),
	.prn(vcc));
defparam \ram_in_reg[1][4] .is_wysiwyg = "true";
defparam \ram_in_reg[1][4] .power_up = "low";

dffeas \ram_in_reg[1][5] (
	.clk(clk),
	.d(\Mux1~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_5_1),
	.prn(vcc));
defparam \ram_in_reg[1][5] .is_wysiwyg = "true";
defparam \ram_in_reg[1][5] .power_up = "low";

dffeas \ram_in_reg[0][1] (
	.clk(clk),
	.d(\Mux5~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_1_0),
	.prn(vcc));
defparam \ram_in_reg[0][1] .is_wysiwyg = "true";
defparam \ram_in_reg[0][1] .power_up = "low";

dffeas \ram_in_reg[0][3] (
	.clk(clk),
	.d(\Mux3~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_3_0),
	.prn(vcc));
defparam \ram_in_reg[0][3] .is_wysiwyg = "true";
defparam \ram_in_reg[0][3] .power_up = "low";

dffeas \ram_in_reg[0][5] (
	.clk(clk),
	.d(\Mux1~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_5_0),
	.prn(vcc));
defparam \ram_in_reg[0][5] .is_wysiwyg = "true";
defparam \ram_in_reg[0][5] .power_up = "low";

dffeas \ram_in_reg[3][1] (
	.clk(clk),
	.d(\Mux5~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_1_3),
	.prn(vcc));
defparam \ram_in_reg[3][1] .is_wysiwyg = "true";
defparam \ram_in_reg[3][1] .power_up = "low";

dffeas \ram_in_reg[3][3] (
	.clk(clk),
	.d(\Mux3~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_3_3),
	.prn(vcc));
defparam \ram_in_reg[3][3] .is_wysiwyg = "true";
defparam \ram_in_reg[3][3] .power_up = "low";

dffeas \ram_in_reg[3][5] (
	.clk(clk),
	.d(\Mux1~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_5_3),
	.prn(vcc));
defparam \ram_in_reg[3][5] .is_wysiwyg = "true";
defparam \ram_in_reg[3][5] .power_up = "low";

dffeas \sw_3_arr[0][0] (
	.clk(clk),
	.d(sw_3_in[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sw_3_arr[0][0]~q ),
	.prn(vcc));
defparam \sw_3_arr[0][0] .is_wysiwyg = "true";
defparam \sw_3_arr[0][0] .power_up = "low";

dffeas \sw_2_arr[0][0] (
	.clk(clk),
	.d(sw_2_in[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sw_2_arr[0][0]~q ),
	.prn(vcc));
defparam \sw_2_arr[0][0] .is_wysiwyg = "true";
defparam \sw_2_arr[0][0] .power_up = "low";

cycloneiii_lcell_comb \Mux6~0 (
	.dataa(\sw_3_arr[0][0]~q ),
	.datab(\sw_2_arr[0][0]~q ),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\Mux6~0_combout ),
	.cout());
defparam \Mux6~0 .lut_mask = 16'hAACC;
defparam \Mux6~0 .sum_lutc_input = "datac";

dffeas \sw_3_arr[0][1] (
	.clk(clk),
	.d(sw_3_in[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sw_3_arr[0][1]~q ),
	.prn(vcc));
defparam \sw_3_arr[0][1] .is_wysiwyg = "true";
defparam \sw_3_arr[0][1] .power_up = "low";

dffeas \sw_1_arr[0][1] (
	.clk(clk),
	.d(sw_1_in[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sw_1_arr[0][1]~q ),
	.prn(vcc));
defparam \sw_1_arr[0][1] .is_wysiwyg = "true";
defparam \sw_1_arr[0][1] .power_up = "low";

cycloneiii_lcell_comb \Mux19~0 (
	.dataa(\sw_3_arr[0][1]~q ),
	.datab(\sw_1_arr[0][1]~q ),
	.datac(swa_tdl_0_0),
	.datad(swa_tdl_1_0),
	.cin(gnd),
	.combout(\Mux19~0_combout ),
	.cout());
defparam \Mux19~0 .lut_mask = 16'hEFFE;
defparam \Mux19~0 .sum_lutc_input = "datac";

dffeas \sw_3_arr[0][2] (
	.clk(clk),
	.d(sw_3_in[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sw_3_arr[0][2]~q ),
	.prn(vcc));
defparam \sw_3_arr[0][2] .is_wysiwyg = "true";
defparam \sw_3_arr[0][2] .power_up = "low";

dffeas \sw_2_arr[0][2] (
	.clk(clk),
	.d(sw_2_in[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sw_2_arr[0][2]~q ),
	.prn(vcc));
defparam \sw_2_arr[0][2] .is_wysiwyg = "true";
defparam \sw_2_arr[0][2] .power_up = "low";

cycloneiii_lcell_comb \Mux4~0 (
	.dataa(\sw_3_arr[0][2]~q ),
	.datab(\sw_2_arr[0][2]~q ),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\Mux4~0_combout ),
	.cout());
defparam \Mux4~0 .lut_mask = 16'hAACC;
defparam \Mux4~0 .sum_lutc_input = "datac";

dffeas \sw_3_arr[0][3] (
	.clk(clk),
	.d(sw_3_in[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sw_3_arr[0][3]~q ),
	.prn(vcc));
defparam \sw_3_arr[0][3] .is_wysiwyg = "true";
defparam \sw_3_arr[0][3] .power_up = "low";

dffeas \sw_1_arr[0][3] (
	.clk(clk),
	.d(sw_1_in[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sw_1_arr[0][3]~q ),
	.prn(vcc));
defparam \sw_1_arr[0][3] .is_wysiwyg = "true";
defparam \sw_1_arr[0][3] .power_up = "low";

cycloneiii_lcell_comb \Mux17~0 (
	.dataa(\sw_3_arr[0][3]~q ),
	.datab(\sw_1_arr[0][3]~q ),
	.datac(swa_tdl_0_0),
	.datad(swa_tdl_1_0),
	.cin(gnd),
	.combout(\Mux17~0_combout ),
	.cout());
defparam \Mux17~0 .lut_mask = 16'hEFFE;
defparam \Mux17~0 .sum_lutc_input = "datac";

dffeas \sw_3_arr[0][4] (
	.clk(clk),
	.d(sw_3_in[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sw_3_arr[0][4]~q ),
	.prn(vcc));
defparam \sw_3_arr[0][4] .is_wysiwyg = "true";
defparam \sw_3_arr[0][4] .power_up = "low";

dffeas \sw_2_arr[0][4] (
	.clk(clk),
	.d(sw_2_in[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sw_2_arr[0][4]~q ),
	.prn(vcc));
defparam \sw_2_arr[0][4] .is_wysiwyg = "true";
defparam \sw_2_arr[0][4] .power_up = "low";

cycloneiii_lcell_comb \Mux2~0 (
	.dataa(\sw_3_arr[0][4]~q ),
	.datab(\sw_2_arr[0][4]~q ),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\Mux2~0_combout ),
	.cout());
defparam \Mux2~0 .lut_mask = 16'hAACC;
defparam \Mux2~0 .sum_lutc_input = "datac";

dffeas \sw_3_arr[0][5] (
	.clk(clk),
	.d(sw_3_in[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sw_3_arr[0][5]~q ),
	.prn(vcc));
defparam \sw_3_arr[0][5] .is_wysiwyg = "true";
defparam \sw_3_arr[0][5] .power_up = "low";

dffeas \sw_1_arr[0][5] (
	.clk(clk),
	.d(sw_1_in[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sw_1_arr[0][5]~q ),
	.prn(vcc));
defparam \sw_1_arr[0][5] .is_wysiwyg = "true";
defparam \sw_1_arr[0][5] .power_up = "low";

cycloneiii_lcell_comb \Mux15~0 (
	.dataa(\sw_3_arr[0][5]~q ),
	.datab(\sw_1_arr[0][5]~q ),
	.datac(swa_tdl_0_0),
	.datad(swa_tdl_1_0),
	.cin(gnd),
	.combout(\Mux15~0_combout ),
	.cout());
defparam \Mux15~0 .lut_mask = 16'hEFFE;
defparam \Mux15~0 .sum_lutc_input = "datac";

dffeas \sw_3_arr[0][6] (
	.clk(clk),
	.d(sw_3_in[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sw_3_arr[0][6]~q ),
	.prn(vcc));
defparam \sw_3_arr[0][6] .is_wysiwyg = "true";
defparam \sw_3_arr[0][6] .power_up = "low";

cycloneiii_lcell_comb \Mux13~0 (
	.dataa(\sw_2_arr[0][0]~q ),
	.datab(\sw_3_arr[0][0]~q ),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\Mux13~0_combout ),
	.cout());
defparam \Mux13~0 .lut_mask = 16'hAACC;
defparam \Mux13~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux5~0 (
	.dataa(\sw_3_arr[0][1]~q ),
	.datab(\sw_1_arr[0][1]~q ),
	.datac(gnd),
	.datad(swa_tdl_1_0),
	.cin(gnd),
	.combout(\Mux5~0_combout ),
	.cout());
defparam \Mux5~0 .lut_mask = 16'hAACC;
defparam \Mux5~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux11~0 (
	.dataa(\sw_2_arr[0][2]~q ),
	.datab(\sw_3_arr[0][2]~q ),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\Mux11~0_combout ),
	.cout());
defparam \Mux11~0 .lut_mask = 16'hAACC;
defparam \Mux11~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux3~0 (
	.dataa(\sw_3_arr[0][3]~q ),
	.datab(\sw_1_arr[0][3]~q ),
	.datac(gnd),
	.datad(swa_tdl_1_0),
	.cin(gnd),
	.combout(\Mux3~0_combout ),
	.cout());
defparam \Mux3~0 .lut_mask = 16'hAACC;
defparam \Mux3~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux9~0 (
	.dataa(\sw_2_arr[0][4]~q ),
	.datab(\sw_3_arr[0][4]~q ),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\Mux9~0_combout ),
	.cout());
defparam \Mux9~0 .lut_mask = 16'hAACC;
defparam \Mux9~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux1~0 (
	.dataa(\sw_3_arr[0][5]~q ),
	.datab(\sw_1_arr[0][5]~q ),
	.datac(gnd),
	.datad(swa_tdl_1_0),
	.cin(gnd),
	.combout(\Mux1~0_combout ),
	.cout());
defparam \Mux1~0 .lut_mask = 16'hAACC;
defparam \Mux1~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux5~1 (
	.dataa(\sw_1_arr[0][1]~q ),
	.datab(\sw_3_arr[0][1]~q ),
	.datac(swa_tdl_0_0),
	.datad(swa_tdl_1_0),
	.cin(gnd),
	.combout(\Mux5~1_combout ),
	.cout());
defparam \Mux5~1 .lut_mask = 16'hEFFE;
defparam \Mux5~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux3~1 (
	.dataa(\sw_1_arr[0][3]~q ),
	.datab(\sw_3_arr[0][3]~q ),
	.datac(swa_tdl_0_0),
	.datad(swa_tdl_1_0),
	.cin(gnd),
	.combout(\Mux3~1_combout ),
	.cout());
defparam \Mux3~1 .lut_mask = 16'hEFFE;
defparam \Mux3~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux1~1 (
	.dataa(\sw_1_arr[0][5]~q ),
	.datab(\sw_3_arr[0][5]~q ),
	.datac(swa_tdl_0_0),
	.datad(swa_tdl_1_0),
	.cin(gnd),
	.combout(\Mux1~1_combout ),
	.cout());
defparam \Mux1~1 .lut_mask = 16'hEFFE;
defparam \Mux1~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux5~2 (
	.dataa(\sw_1_arr[0][1]~q ),
	.datab(\sw_3_arr[0][1]~q ),
	.datac(gnd),
	.datad(swa_tdl_1_0),
	.cin(gnd),
	.combout(\Mux5~2_combout ),
	.cout());
defparam \Mux5~2 .lut_mask = 16'hAACC;
defparam \Mux5~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux3~2 (
	.dataa(\sw_1_arr[0][3]~q ),
	.datab(\sw_3_arr[0][3]~q ),
	.datac(gnd),
	.datad(swa_tdl_1_0),
	.cin(gnd),
	.combout(\Mux3~2_combout ),
	.cout());
defparam \Mux3~2 .lut_mask = 16'hAACC;
defparam \Mux3~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux1~2 (
	.dataa(\sw_1_arr[0][5]~q ),
	.datab(\sw_3_arr[0][5]~q ),
	.datac(gnd),
	.datad(swa_tdl_1_0),
	.cin(gnd),
	.combout(\Mux1~2_combout ),
	.cout());
defparam \Mux1~2 .lut_mask = 16'hAACC;
defparam \Mux1~2 .sum_lutc_input = "datac";

endmodule

module fft_asj_fft_cxb_addr_fft_120_2 (
	global_clock_enable,
	ram_in_reg_0_0,
	ram_in_reg_1_0,
	ram_in_reg_2_0,
	ram_in_reg_3_0,
	ram_in_reg_4_0,
	ram_in_reg_5_0,
	ram_in_reg_0_1,
	ram_in_reg_1_1,
	ram_in_reg_2_1,
	ram_in_reg_3_1,
	ram_in_reg_4_1,
	ram_in_reg_5_1,
	ram_in_reg_1_2,
	ram_in_reg_3_2,
	ram_in_reg_5_2,
	ram_in_reg_1_3,
	ram_in_reg_3_3,
	ram_in_reg_5_3,
	rd_addr_d_0,
	rd_addr_c_0,
	sw_0,
	rd_addr_b_1,
	rd_addr_d_1,
	sw_1,
	rd_addr_d_2,
	rd_addr_c_2,
	rd_addr_b_3,
	rd_addr_d_3,
	rd_addr_d_4,
	rd_addr_c_4,
	rd_addr_b_5,
	rd_addr_d_5,
	clk)/* synthesis synthesis_greybox=1 */;
input 	global_clock_enable;
output 	ram_in_reg_0_0;
output 	ram_in_reg_1_0;
output 	ram_in_reg_2_0;
output 	ram_in_reg_3_0;
output 	ram_in_reg_4_0;
output 	ram_in_reg_5_0;
output 	ram_in_reg_0_1;
output 	ram_in_reg_1_1;
output 	ram_in_reg_2_1;
output 	ram_in_reg_3_1;
output 	ram_in_reg_4_1;
output 	ram_in_reg_5_1;
output 	ram_in_reg_1_2;
output 	ram_in_reg_3_2;
output 	ram_in_reg_5_2;
output 	ram_in_reg_1_3;
output 	ram_in_reg_3_3;
output 	ram_in_reg_5_3;
input 	rd_addr_d_0;
input 	rd_addr_c_0;
input 	sw_0;
input 	rd_addr_b_1;
input 	rd_addr_d_1;
input 	sw_1;
input 	rd_addr_d_2;
input 	rd_addr_c_2;
input 	rd_addr_b_3;
input 	rd_addr_d_3;
input 	rd_addr_d_4;
input 	rd_addr_c_4;
input 	rd_addr_b_5;
input 	rd_addr_d_5;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Mux6~0_combout ;
wire \Mux5~0_combout ;
wire \Mux4~0_combout ;
wire \Mux3~0_combout ;
wire \Mux2~0_combout ;
wire \Mux1~0_combout ;
wire \Mux13~0_combout ;
wire \Mux5~1_combout ;
wire \Mux11~0_combout ;
wire \Mux3~1_combout ;
wire \Mux9~0_combout ;
wire \Mux1~1_combout ;
wire \Mux19~0_combout ;
wire \Mux17~0_combout ;
wire \Mux15~0_combout ;
wire \Mux5~2_combout ;
wire \Mux3~2_combout ;
wire \Mux1~2_combout ;


dffeas \ram_in_reg[0][0] (
	.clk(clk),
	.d(\Mux6~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_0_0),
	.prn(vcc));
defparam \ram_in_reg[0][0] .is_wysiwyg = "true";
defparam \ram_in_reg[0][0] .power_up = "low";

dffeas \ram_in_reg[0][1] (
	.clk(clk),
	.d(\Mux5~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_1_0),
	.prn(vcc));
defparam \ram_in_reg[0][1] .is_wysiwyg = "true";
defparam \ram_in_reg[0][1] .power_up = "low";

dffeas \ram_in_reg[0][2] (
	.clk(clk),
	.d(\Mux4~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_2_0),
	.prn(vcc));
defparam \ram_in_reg[0][2] .is_wysiwyg = "true";
defparam \ram_in_reg[0][2] .power_up = "low";

dffeas \ram_in_reg[0][3] (
	.clk(clk),
	.d(\Mux3~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_3_0),
	.prn(vcc));
defparam \ram_in_reg[0][3] .is_wysiwyg = "true";
defparam \ram_in_reg[0][3] .power_up = "low";

dffeas \ram_in_reg[0][4] (
	.clk(clk),
	.d(\Mux2~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_4_0),
	.prn(vcc));
defparam \ram_in_reg[0][4] .is_wysiwyg = "true";
defparam \ram_in_reg[0][4] .power_up = "low";

dffeas \ram_in_reg[0][5] (
	.clk(clk),
	.d(\Mux1~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_5_0),
	.prn(vcc));
defparam \ram_in_reg[0][5] .is_wysiwyg = "true";
defparam \ram_in_reg[0][5] .power_up = "low";

dffeas \ram_in_reg[1][0] (
	.clk(clk),
	.d(\Mux13~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_0_1),
	.prn(vcc));
defparam \ram_in_reg[1][0] .is_wysiwyg = "true";
defparam \ram_in_reg[1][0] .power_up = "low";

dffeas \ram_in_reg[1][1] (
	.clk(clk),
	.d(\Mux5~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_1_1),
	.prn(vcc));
defparam \ram_in_reg[1][1] .is_wysiwyg = "true";
defparam \ram_in_reg[1][1] .power_up = "low";

dffeas \ram_in_reg[1][2] (
	.clk(clk),
	.d(\Mux11~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_2_1),
	.prn(vcc));
defparam \ram_in_reg[1][2] .is_wysiwyg = "true";
defparam \ram_in_reg[1][2] .power_up = "low";

dffeas \ram_in_reg[1][3] (
	.clk(clk),
	.d(\Mux3~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_3_1),
	.prn(vcc));
defparam \ram_in_reg[1][3] .is_wysiwyg = "true";
defparam \ram_in_reg[1][3] .power_up = "low";

dffeas \ram_in_reg[1][4] (
	.clk(clk),
	.d(\Mux9~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_4_1),
	.prn(vcc));
defparam \ram_in_reg[1][4] .is_wysiwyg = "true";
defparam \ram_in_reg[1][4] .power_up = "low";

dffeas \ram_in_reg[1][5] (
	.clk(clk),
	.d(\Mux1~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_5_1),
	.prn(vcc));
defparam \ram_in_reg[1][5] .is_wysiwyg = "true";
defparam \ram_in_reg[1][5] .power_up = "low";

dffeas \ram_in_reg[2][1] (
	.clk(clk),
	.d(\Mux19~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_1_2),
	.prn(vcc));
defparam \ram_in_reg[2][1] .is_wysiwyg = "true";
defparam \ram_in_reg[2][1] .power_up = "low";

dffeas \ram_in_reg[2][3] (
	.clk(clk),
	.d(\Mux17~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_3_2),
	.prn(vcc));
defparam \ram_in_reg[2][3] .is_wysiwyg = "true";
defparam \ram_in_reg[2][3] .power_up = "low";

dffeas \ram_in_reg[2][5] (
	.clk(clk),
	.d(\Mux15~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_5_2),
	.prn(vcc));
defparam \ram_in_reg[2][5] .is_wysiwyg = "true";
defparam \ram_in_reg[2][5] .power_up = "low";

dffeas \ram_in_reg[3][1] (
	.clk(clk),
	.d(\Mux5~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_1_3),
	.prn(vcc));
defparam \ram_in_reg[3][1] .is_wysiwyg = "true";
defparam \ram_in_reg[3][1] .power_up = "low";

dffeas \ram_in_reg[3][3] (
	.clk(clk),
	.d(\Mux3~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_3_3),
	.prn(vcc));
defparam \ram_in_reg[3][3] .is_wysiwyg = "true";
defparam \ram_in_reg[3][3] .power_up = "low";

dffeas \ram_in_reg[3][5] (
	.clk(clk),
	.d(\Mux1~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_5_3),
	.prn(vcc));
defparam \ram_in_reg[3][5] .is_wysiwyg = "true";
defparam \ram_in_reg[3][5] .power_up = "low";

cycloneiii_lcell_comb \Mux6~0 (
	.dataa(rd_addr_d_0),
	.datab(rd_addr_c_0),
	.datac(gnd),
	.datad(sw_0),
	.cin(gnd),
	.combout(\Mux6~0_combout ),
	.cout());
defparam \Mux6~0 .lut_mask = 16'hAACC;
defparam \Mux6~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux5~0 (
	.dataa(rd_addr_b_1),
	.datab(rd_addr_d_1),
	.datac(sw_0),
	.datad(sw_1),
	.cin(gnd),
	.combout(\Mux5~0_combout ),
	.cout());
defparam \Mux5~0 .lut_mask = 16'hEFFE;
defparam \Mux5~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux4~0 (
	.dataa(rd_addr_d_2),
	.datab(rd_addr_c_2),
	.datac(gnd),
	.datad(sw_0),
	.cin(gnd),
	.combout(\Mux4~0_combout ),
	.cout());
defparam \Mux4~0 .lut_mask = 16'hAACC;
defparam \Mux4~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux3~0 (
	.dataa(rd_addr_b_3),
	.datab(rd_addr_d_3),
	.datac(sw_0),
	.datad(sw_1),
	.cin(gnd),
	.combout(\Mux3~0_combout ),
	.cout());
defparam \Mux3~0 .lut_mask = 16'hEFFE;
defparam \Mux3~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux2~0 (
	.dataa(rd_addr_d_4),
	.datab(rd_addr_c_4),
	.datac(gnd),
	.datad(sw_0),
	.cin(gnd),
	.combout(\Mux2~0_combout ),
	.cout());
defparam \Mux2~0 .lut_mask = 16'hAACC;
defparam \Mux2~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux1~0 (
	.dataa(rd_addr_b_5),
	.datab(rd_addr_d_5),
	.datac(sw_0),
	.datad(sw_1),
	.cin(gnd),
	.combout(\Mux1~0_combout ),
	.cout());
defparam \Mux1~0 .lut_mask = 16'hEFFE;
defparam \Mux1~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux13~0 (
	.dataa(rd_addr_c_0),
	.datab(rd_addr_d_0),
	.datac(gnd),
	.datad(sw_0),
	.cin(gnd),
	.combout(\Mux13~0_combout ),
	.cout());
defparam \Mux13~0 .lut_mask = 16'hAACC;
defparam \Mux13~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux5~1 (
	.dataa(rd_addr_d_1),
	.datab(rd_addr_b_1),
	.datac(gnd),
	.datad(sw_1),
	.cin(gnd),
	.combout(\Mux5~1_combout ),
	.cout());
defparam \Mux5~1 .lut_mask = 16'hAACC;
defparam \Mux5~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux11~0 (
	.dataa(rd_addr_c_2),
	.datab(rd_addr_d_2),
	.datac(gnd),
	.datad(sw_0),
	.cin(gnd),
	.combout(\Mux11~0_combout ),
	.cout());
defparam \Mux11~0 .lut_mask = 16'hAACC;
defparam \Mux11~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux3~1 (
	.dataa(rd_addr_d_3),
	.datab(rd_addr_b_3),
	.datac(gnd),
	.datad(sw_1),
	.cin(gnd),
	.combout(\Mux3~1_combout ),
	.cout());
defparam \Mux3~1 .lut_mask = 16'hAACC;
defparam \Mux3~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux9~0 (
	.dataa(rd_addr_c_4),
	.datab(rd_addr_d_4),
	.datac(gnd),
	.datad(sw_0),
	.cin(gnd),
	.combout(\Mux9~0_combout ),
	.cout());
defparam \Mux9~0 .lut_mask = 16'hAACC;
defparam \Mux9~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux1~1 (
	.dataa(rd_addr_d_5),
	.datab(rd_addr_b_5),
	.datac(gnd),
	.datad(sw_1),
	.cin(gnd),
	.combout(\Mux1~1_combout ),
	.cout());
defparam \Mux1~1 .lut_mask = 16'hAACC;
defparam \Mux1~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux19~0 (
	.dataa(rd_addr_d_1),
	.datab(rd_addr_b_1),
	.datac(sw_0),
	.datad(sw_1),
	.cin(gnd),
	.combout(\Mux19~0_combout ),
	.cout());
defparam \Mux19~0 .lut_mask = 16'hEFFE;
defparam \Mux19~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux17~0 (
	.dataa(rd_addr_d_3),
	.datab(rd_addr_b_3),
	.datac(sw_0),
	.datad(sw_1),
	.cin(gnd),
	.combout(\Mux17~0_combout ),
	.cout());
defparam \Mux17~0 .lut_mask = 16'hEFFE;
defparam \Mux17~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux15~0 (
	.dataa(rd_addr_d_5),
	.datab(rd_addr_b_5),
	.datac(sw_0),
	.datad(sw_1),
	.cin(gnd),
	.combout(\Mux15~0_combout ),
	.cout());
defparam \Mux15~0 .lut_mask = 16'hEFFE;
defparam \Mux15~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux5~2 (
	.dataa(rd_addr_b_1),
	.datab(rd_addr_d_1),
	.datac(gnd),
	.datad(sw_1),
	.cin(gnd),
	.combout(\Mux5~2_combout ),
	.cout());
defparam \Mux5~2 .lut_mask = 16'hAACC;
defparam \Mux5~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux3~2 (
	.dataa(rd_addr_b_3),
	.datab(rd_addr_d_3),
	.datac(gnd),
	.datad(sw_1),
	.cin(gnd),
	.combout(\Mux3~2_combout ),
	.cout());
defparam \Mux3~2 .lut_mask = 16'hAACC;
defparam \Mux3~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux1~2 (
	.dataa(rd_addr_b_5),
	.datab(rd_addr_d_5),
	.datac(gnd),
	.datad(sw_1),
	.cin(gnd),
	.combout(\Mux1~2_combout ),
	.cout());
defparam \Mux1~2 .lut_mask = 16'hAACC;
defparam \Mux1~2 .sum_lutc_input = "datac";

endmodule

module fft_asj_fft_cxb_data_fft_120 (
	ram_in_reg_1_6,
	ram_in_reg_1_5,
	ram_in_reg_1_4,
	ram_in_reg_1_7,
	ram_in_reg_0_6,
	ram_in_reg_0_5,
	ram_in_reg_0_4,
	ram_in_reg_0_7,
	ram_in_reg_7_6,
	ram_in_reg_7_5,
	ram_in_reg_7_4,
	ram_in_reg_7_7,
	ram_in_reg_6_6,
	ram_in_reg_6_5,
	ram_in_reg_6_4,
	ram_in_reg_6_7,
	ram_in_reg_5_6,
	ram_in_reg_5_5,
	ram_in_reg_5_4,
	ram_in_reg_5_7,
	ram_in_reg_4_6,
	ram_in_reg_4_5,
	ram_in_reg_4_4,
	ram_in_reg_4_7,
	ram_in_reg_3_6,
	ram_in_reg_3_5,
	ram_in_reg_3_4,
	ram_in_reg_3_7,
	ram_in_reg_2_6,
	ram_in_reg_2_5,
	ram_in_reg_2_4,
	ram_in_reg_2_7,
	ram_in_reg_1_2,
	ram_in_reg_1_1,
	ram_in_reg_1_0,
	ram_in_reg_1_3,
	ram_in_reg_0_2,
	ram_in_reg_0_1,
	ram_in_reg_0_0,
	ram_in_reg_0_3,
	ram_in_reg_7_2,
	ram_in_reg_7_1,
	ram_in_reg_7_0,
	ram_in_reg_7_3,
	ram_in_reg_6_2,
	ram_in_reg_6_1,
	ram_in_reg_6_0,
	ram_in_reg_6_3,
	ram_in_reg_5_2,
	ram_in_reg_5_1,
	ram_in_reg_5_0,
	ram_in_reg_5_3,
	ram_in_reg_4_2,
	ram_in_reg_4_1,
	ram_in_reg_4_0,
	ram_in_reg_4_3,
	ram_in_reg_3_2,
	ram_in_reg_3_1,
	ram_in_reg_3_0,
	ram_in_reg_3_3,
	ram_in_reg_2_2,
	ram_in_reg_2_1,
	ram_in_reg_2_0,
	ram_in_reg_2_3,
	r_array_out_3_0,
	i_array_out_3_0,
	r_array_out_3_1,
	i_array_out_3_1,
	r_array_out_3_2,
	i_array_out_3_2,
	r_array_out_3_3,
	i_array_out_3_3,
	r_array_out_4_0,
	i_array_out_4_0,
	r_array_out_4_1,
	i_array_out_4_1,
	r_array_out_4_2,
	i_array_out_4_2,
	r_array_out_4_3,
	i_array_out_4_3,
	r_array_out_5_0,
	i_array_out_5_0,
	r_array_out_5_1,
	i_array_out_5_1,
	r_array_out_5_2,
	i_array_out_5_2,
	r_array_out_5_3,
	i_array_out_5_3,
	i_array_out_2_2,
	i_array_out_2_1,
	i_array_out_2_0,
	i_array_out_2_3,
	r_array_out_2_2,
	r_array_out_2_1,
	r_array_out_2_0,
	r_array_out_2_3,
	global_clock_enable,
	r_array_out_7_0,
	i_array_out_7_0,
	r_array_out_7_1,
	i_array_out_7_1,
	r_array_out_7_2,
	i_array_out_7_2,
	r_array_out_7_3,
	i_array_out_7_3,
	r_array_out_6_0,
	i_array_out_6_0,
	r_array_out_6_1,
	i_array_out_6_1,
	r_array_out_6_2,
	i_array_out_6_2,
	r_array_out_6_3,
	i_array_out_6_3,
	i_array_out_1_2,
	i_array_out_1_1,
	swa_tdl_0_0,
	i_array_out_1_0,
	i_array_out_1_3,
	swa_tdl_1_0,
	i_array_out_0_2,
	i_array_out_0_1,
	i_array_out_0_0,
	i_array_out_0_3,
	r_array_out_1_2,
	r_array_out_1_1,
	r_array_out_1_0,
	r_array_out_1_3,
	r_array_out_0_2,
	r_array_out_0_1,
	r_array_out_0_0,
	r_array_out_0_3,
	clk)/* synthesis synthesis_greybox=1 */;
output 	ram_in_reg_1_6;
output 	ram_in_reg_1_5;
output 	ram_in_reg_1_4;
output 	ram_in_reg_1_7;
output 	ram_in_reg_0_6;
output 	ram_in_reg_0_5;
output 	ram_in_reg_0_4;
output 	ram_in_reg_0_7;
output 	ram_in_reg_7_6;
output 	ram_in_reg_7_5;
output 	ram_in_reg_7_4;
output 	ram_in_reg_7_7;
output 	ram_in_reg_6_6;
output 	ram_in_reg_6_5;
output 	ram_in_reg_6_4;
output 	ram_in_reg_6_7;
output 	ram_in_reg_5_6;
output 	ram_in_reg_5_5;
output 	ram_in_reg_5_4;
output 	ram_in_reg_5_7;
output 	ram_in_reg_4_6;
output 	ram_in_reg_4_5;
output 	ram_in_reg_4_4;
output 	ram_in_reg_4_7;
output 	ram_in_reg_3_6;
output 	ram_in_reg_3_5;
output 	ram_in_reg_3_4;
output 	ram_in_reg_3_7;
output 	ram_in_reg_2_6;
output 	ram_in_reg_2_5;
output 	ram_in_reg_2_4;
output 	ram_in_reg_2_7;
output 	ram_in_reg_1_2;
output 	ram_in_reg_1_1;
output 	ram_in_reg_1_0;
output 	ram_in_reg_1_3;
output 	ram_in_reg_0_2;
output 	ram_in_reg_0_1;
output 	ram_in_reg_0_0;
output 	ram_in_reg_0_3;
output 	ram_in_reg_7_2;
output 	ram_in_reg_7_1;
output 	ram_in_reg_7_0;
output 	ram_in_reg_7_3;
output 	ram_in_reg_6_2;
output 	ram_in_reg_6_1;
output 	ram_in_reg_6_0;
output 	ram_in_reg_6_3;
output 	ram_in_reg_5_2;
output 	ram_in_reg_5_1;
output 	ram_in_reg_5_0;
output 	ram_in_reg_5_3;
output 	ram_in_reg_4_2;
output 	ram_in_reg_4_1;
output 	ram_in_reg_4_0;
output 	ram_in_reg_4_3;
output 	ram_in_reg_3_2;
output 	ram_in_reg_3_1;
output 	ram_in_reg_3_0;
output 	ram_in_reg_3_3;
output 	ram_in_reg_2_2;
output 	ram_in_reg_2_1;
output 	ram_in_reg_2_0;
output 	ram_in_reg_2_3;
input 	r_array_out_3_0;
input 	i_array_out_3_0;
input 	r_array_out_3_1;
input 	i_array_out_3_1;
input 	r_array_out_3_2;
input 	i_array_out_3_2;
input 	r_array_out_3_3;
input 	i_array_out_3_3;
input 	r_array_out_4_0;
input 	i_array_out_4_0;
input 	r_array_out_4_1;
input 	i_array_out_4_1;
input 	r_array_out_4_2;
input 	i_array_out_4_2;
input 	r_array_out_4_3;
input 	i_array_out_4_3;
input 	r_array_out_5_0;
input 	i_array_out_5_0;
input 	r_array_out_5_1;
input 	i_array_out_5_1;
input 	r_array_out_5_2;
input 	i_array_out_5_2;
input 	r_array_out_5_3;
input 	i_array_out_5_3;
input 	i_array_out_2_2;
input 	i_array_out_2_1;
input 	i_array_out_2_0;
input 	i_array_out_2_3;
input 	r_array_out_2_2;
input 	r_array_out_2_1;
input 	r_array_out_2_0;
input 	r_array_out_2_3;
input 	global_clock_enable;
input 	r_array_out_7_0;
input 	i_array_out_7_0;
input 	r_array_out_7_1;
input 	i_array_out_7_1;
input 	r_array_out_7_2;
input 	i_array_out_7_2;
input 	r_array_out_7_3;
input 	i_array_out_7_3;
input 	r_array_out_6_0;
input 	i_array_out_6_0;
input 	r_array_out_6_1;
input 	i_array_out_6_1;
input 	r_array_out_6_2;
input 	i_array_out_6_2;
input 	r_array_out_6_3;
input 	i_array_out_6_3;
input 	i_array_out_1_2;
input 	i_array_out_1_1;
input 	swa_tdl_0_0;
input 	i_array_out_1_0;
input 	i_array_out_1_3;
input 	swa_tdl_1_0;
input 	i_array_out_0_2;
input 	i_array_out_0_1;
input 	i_array_out_0_0;
input 	i_array_out_0_3;
input 	r_array_out_1_2;
input 	r_array_out_1_1;
input 	r_array_out_1_0;
input 	r_array_out_1_3;
input 	r_array_out_0_2;
input 	r_array_out_0_1;
input 	r_array_out_0_0;
input 	r_array_out_0_3;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ram_in_reg[6][1]~5_combout ;
wire \ram_in_reg[4][1]~6_combout ;
wire \ram_in_reg[5][1]~4_combout ;
wire \ram_in_reg[7][1]~7_combout ;
wire \ram_in_reg[6][0]~60_combout ;
wire \ram_in_reg[4][0]~62_combout ;
wire \ram_in_reg[5][0]~61_combout ;
wire \ram_in_reg[7][0]~63_combout ;
wire \ram_in_reg[6][7]~53_combout ;
wire \ram_in_reg[4][7]~54_combout ;
wire \ram_in_reg[5][7]~52_combout ;
wire \ram_in_reg[7][7]~55_combout ;
wire \ram_in_reg[6][6]~44_combout ;
wire \ram_in_reg[4][6]~46_combout ;
wire \ram_in_reg[5][6]~45_combout ;
wire \ram_in_reg[7][6]~47_combout ;
wire \ram_in_reg[6][5]~37_combout ;
wire \ram_in_reg[4][5]~38_combout ;
wire \ram_in_reg[5][5]~36_combout ;
wire \ram_in_reg[7][5]~39_combout ;
wire \ram_in_reg[6][4]~28_combout ;
wire \ram_in_reg[4][4]~30_combout ;
wire \ram_in_reg[5][4]~29_combout ;
wire \ram_in_reg[7][4]~31_combout ;
wire \ram_in_reg[6][3]~21_combout ;
wire \ram_in_reg[4][3]~22_combout ;
wire \ram_in_reg[5][3]~20_combout ;
wire \ram_in_reg[7][3]~23_combout ;
wire \ram_in_reg[6][2]~12_combout ;
wire \ram_in_reg[4][2]~14_combout ;
wire \ram_in_reg[5][2]~13_combout ;
wire \ram_in_reg[7][2]~15_combout ;
wire \ram_in_reg[2][1]~1_combout ;
wire \ram_in_reg[0][1]~2_combout ;
wire \ram_in_reg[1][1]~0_combout ;
wire \ram_in_reg[3][1]~3_combout ;
wire \ram_in_reg[2][0]~56_combout ;
wire \ram_in_reg[0][0]~58_combout ;
wire \ram_in_reg[1][0]~57_combout ;
wire \ram_in_reg[3][0]~59_combout ;
wire \ram_in_reg[2][7]~49_combout ;
wire \ram_in_reg[0][7]~50_combout ;
wire \ram_in_reg[1][7]~48_combout ;
wire \ram_in_reg[3][7]~51_combout ;
wire \ram_in_reg[2][6]~40_combout ;
wire \ram_in_reg[0][6]~42_combout ;
wire \ram_in_reg[1][6]~41_combout ;
wire \ram_in_reg[3][6]~43_combout ;
wire \ram_in_reg[2][5]~33_combout ;
wire \ram_in_reg[0][5]~34_combout ;
wire \ram_in_reg[1][5]~32_combout ;
wire \ram_in_reg[3][5]~35_combout ;
wire \ram_in_reg[2][4]~24_combout ;
wire \ram_in_reg[0][4]~26_combout ;
wire \ram_in_reg[1][4]~25_combout ;
wire \ram_in_reg[3][4]~27_combout ;
wire \ram_in_reg[2][3]~17_combout ;
wire \ram_in_reg[0][3]~18_combout ;
wire \ram_in_reg[1][3]~16_combout ;
wire \ram_in_reg[3][3]~19_combout ;
wire \ram_in_reg[2][2]~8_combout ;
wire \ram_in_reg[0][2]~10_combout ;
wire \ram_in_reg[1][2]~9_combout ;
wire \ram_in_reg[3][2]~11_combout ;


dffeas \ram_in_reg[6][1] (
	.clk(clk),
	.d(\ram_in_reg[6][1]~5_combout ),
	.asdata(\ram_in_reg[4][1]~6_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_1_6),
	.prn(vcc));
defparam \ram_in_reg[6][1] .is_wysiwyg = "true";
defparam \ram_in_reg[6][1] .power_up = "low";

dffeas \ram_in_reg[5][1] (
	.clk(clk),
	.d(\ram_in_reg[5][1]~4_combout ),
	.asdata(\ram_in_reg[7][1]~7_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_1_5),
	.prn(vcc));
defparam \ram_in_reg[5][1] .is_wysiwyg = "true";
defparam \ram_in_reg[5][1] .power_up = "low";

dffeas \ram_in_reg[4][1] (
	.clk(clk),
	.d(\ram_in_reg[4][1]~6_combout ),
	.asdata(\ram_in_reg[6][1]~5_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_1_4),
	.prn(vcc));
defparam \ram_in_reg[4][1] .is_wysiwyg = "true";
defparam \ram_in_reg[4][1] .power_up = "low";

dffeas \ram_in_reg[7][1] (
	.clk(clk),
	.d(\ram_in_reg[7][1]~7_combout ),
	.asdata(\ram_in_reg[5][1]~4_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_1_7),
	.prn(vcc));
defparam \ram_in_reg[7][1] .is_wysiwyg = "true";
defparam \ram_in_reg[7][1] .power_up = "low";

dffeas \ram_in_reg[6][0] (
	.clk(clk),
	.d(\ram_in_reg[6][0]~60_combout ),
	.asdata(\ram_in_reg[4][0]~62_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_0_6),
	.prn(vcc));
defparam \ram_in_reg[6][0] .is_wysiwyg = "true";
defparam \ram_in_reg[6][0] .power_up = "low";

dffeas \ram_in_reg[5][0] (
	.clk(clk),
	.d(\ram_in_reg[5][0]~61_combout ),
	.asdata(\ram_in_reg[7][0]~63_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_0_5),
	.prn(vcc));
defparam \ram_in_reg[5][0] .is_wysiwyg = "true";
defparam \ram_in_reg[5][0] .power_up = "low";

dffeas \ram_in_reg[4][0] (
	.clk(clk),
	.d(\ram_in_reg[4][0]~62_combout ),
	.asdata(\ram_in_reg[6][0]~60_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_0_4),
	.prn(vcc));
defparam \ram_in_reg[4][0] .is_wysiwyg = "true";
defparam \ram_in_reg[4][0] .power_up = "low";

dffeas \ram_in_reg[7][0] (
	.clk(clk),
	.d(\ram_in_reg[7][0]~63_combout ),
	.asdata(\ram_in_reg[5][0]~61_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_0_7),
	.prn(vcc));
defparam \ram_in_reg[7][0] .is_wysiwyg = "true";
defparam \ram_in_reg[7][0] .power_up = "low";

dffeas \ram_in_reg[6][7] (
	.clk(clk),
	.d(\ram_in_reg[6][7]~53_combout ),
	.asdata(\ram_in_reg[4][7]~54_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_7_6),
	.prn(vcc));
defparam \ram_in_reg[6][7] .is_wysiwyg = "true";
defparam \ram_in_reg[6][7] .power_up = "low";

dffeas \ram_in_reg[5][7] (
	.clk(clk),
	.d(\ram_in_reg[5][7]~52_combout ),
	.asdata(\ram_in_reg[7][7]~55_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_7_5),
	.prn(vcc));
defparam \ram_in_reg[5][7] .is_wysiwyg = "true";
defparam \ram_in_reg[5][7] .power_up = "low";

dffeas \ram_in_reg[4][7] (
	.clk(clk),
	.d(\ram_in_reg[4][7]~54_combout ),
	.asdata(\ram_in_reg[6][7]~53_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_7_4),
	.prn(vcc));
defparam \ram_in_reg[4][7] .is_wysiwyg = "true";
defparam \ram_in_reg[4][7] .power_up = "low";

dffeas \ram_in_reg[7][7] (
	.clk(clk),
	.d(\ram_in_reg[7][7]~55_combout ),
	.asdata(\ram_in_reg[5][7]~52_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_7_7),
	.prn(vcc));
defparam \ram_in_reg[7][7] .is_wysiwyg = "true";
defparam \ram_in_reg[7][7] .power_up = "low";

dffeas \ram_in_reg[6][6] (
	.clk(clk),
	.d(\ram_in_reg[6][6]~44_combout ),
	.asdata(\ram_in_reg[4][6]~46_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_6_6),
	.prn(vcc));
defparam \ram_in_reg[6][6] .is_wysiwyg = "true";
defparam \ram_in_reg[6][6] .power_up = "low";

dffeas \ram_in_reg[5][6] (
	.clk(clk),
	.d(\ram_in_reg[5][6]~45_combout ),
	.asdata(\ram_in_reg[7][6]~47_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_6_5),
	.prn(vcc));
defparam \ram_in_reg[5][6] .is_wysiwyg = "true";
defparam \ram_in_reg[5][6] .power_up = "low";

dffeas \ram_in_reg[4][6] (
	.clk(clk),
	.d(\ram_in_reg[4][6]~46_combout ),
	.asdata(\ram_in_reg[6][6]~44_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_6_4),
	.prn(vcc));
defparam \ram_in_reg[4][6] .is_wysiwyg = "true";
defparam \ram_in_reg[4][6] .power_up = "low";

dffeas \ram_in_reg[7][6] (
	.clk(clk),
	.d(\ram_in_reg[7][6]~47_combout ),
	.asdata(\ram_in_reg[5][6]~45_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_6_7),
	.prn(vcc));
defparam \ram_in_reg[7][6] .is_wysiwyg = "true";
defparam \ram_in_reg[7][6] .power_up = "low";

dffeas \ram_in_reg[6][5] (
	.clk(clk),
	.d(\ram_in_reg[6][5]~37_combout ),
	.asdata(\ram_in_reg[4][5]~38_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_5_6),
	.prn(vcc));
defparam \ram_in_reg[6][5] .is_wysiwyg = "true";
defparam \ram_in_reg[6][5] .power_up = "low";

dffeas \ram_in_reg[5][5] (
	.clk(clk),
	.d(\ram_in_reg[5][5]~36_combout ),
	.asdata(\ram_in_reg[7][5]~39_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_5_5),
	.prn(vcc));
defparam \ram_in_reg[5][5] .is_wysiwyg = "true";
defparam \ram_in_reg[5][5] .power_up = "low";

dffeas \ram_in_reg[4][5] (
	.clk(clk),
	.d(\ram_in_reg[4][5]~38_combout ),
	.asdata(\ram_in_reg[6][5]~37_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_5_4),
	.prn(vcc));
defparam \ram_in_reg[4][5] .is_wysiwyg = "true";
defparam \ram_in_reg[4][5] .power_up = "low";

dffeas \ram_in_reg[7][5] (
	.clk(clk),
	.d(\ram_in_reg[7][5]~39_combout ),
	.asdata(\ram_in_reg[5][5]~36_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_5_7),
	.prn(vcc));
defparam \ram_in_reg[7][5] .is_wysiwyg = "true";
defparam \ram_in_reg[7][5] .power_up = "low";

dffeas \ram_in_reg[6][4] (
	.clk(clk),
	.d(\ram_in_reg[6][4]~28_combout ),
	.asdata(\ram_in_reg[4][4]~30_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_4_6),
	.prn(vcc));
defparam \ram_in_reg[6][4] .is_wysiwyg = "true";
defparam \ram_in_reg[6][4] .power_up = "low";

dffeas \ram_in_reg[5][4] (
	.clk(clk),
	.d(\ram_in_reg[5][4]~29_combout ),
	.asdata(\ram_in_reg[7][4]~31_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_4_5),
	.prn(vcc));
defparam \ram_in_reg[5][4] .is_wysiwyg = "true";
defparam \ram_in_reg[5][4] .power_up = "low";

dffeas \ram_in_reg[4][4] (
	.clk(clk),
	.d(\ram_in_reg[4][4]~30_combout ),
	.asdata(\ram_in_reg[6][4]~28_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_4_4),
	.prn(vcc));
defparam \ram_in_reg[4][4] .is_wysiwyg = "true";
defparam \ram_in_reg[4][4] .power_up = "low";

dffeas \ram_in_reg[7][4] (
	.clk(clk),
	.d(\ram_in_reg[7][4]~31_combout ),
	.asdata(\ram_in_reg[5][4]~29_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_4_7),
	.prn(vcc));
defparam \ram_in_reg[7][4] .is_wysiwyg = "true";
defparam \ram_in_reg[7][4] .power_up = "low";

dffeas \ram_in_reg[6][3] (
	.clk(clk),
	.d(\ram_in_reg[6][3]~21_combout ),
	.asdata(\ram_in_reg[4][3]~22_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_3_6),
	.prn(vcc));
defparam \ram_in_reg[6][3] .is_wysiwyg = "true";
defparam \ram_in_reg[6][3] .power_up = "low";

dffeas \ram_in_reg[5][3] (
	.clk(clk),
	.d(\ram_in_reg[5][3]~20_combout ),
	.asdata(\ram_in_reg[7][3]~23_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_3_5),
	.prn(vcc));
defparam \ram_in_reg[5][3] .is_wysiwyg = "true";
defparam \ram_in_reg[5][3] .power_up = "low";

dffeas \ram_in_reg[4][3] (
	.clk(clk),
	.d(\ram_in_reg[4][3]~22_combout ),
	.asdata(\ram_in_reg[6][3]~21_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_3_4),
	.prn(vcc));
defparam \ram_in_reg[4][3] .is_wysiwyg = "true";
defparam \ram_in_reg[4][3] .power_up = "low";

dffeas \ram_in_reg[7][3] (
	.clk(clk),
	.d(\ram_in_reg[7][3]~23_combout ),
	.asdata(\ram_in_reg[5][3]~20_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_3_7),
	.prn(vcc));
defparam \ram_in_reg[7][3] .is_wysiwyg = "true";
defparam \ram_in_reg[7][3] .power_up = "low";

dffeas \ram_in_reg[6][2] (
	.clk(clk),
	.d(\ram_in_reg[6][2]~12_combout ),
	.asdata(\ram_in_reg[4][2]~14_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_2_6),
	.prn(vcc));
defparam \ram_in_reg[6][2] .is_wysiwyg = "true";
defparam \ram_in_reg[6][2] .power_up = "low";

dffeas \ram_in_reg[5][2] (
	.clk(clk),
	.d(\ram_in_reg[5][2]~13_combout ),
	.asdata(\ram_in_reg[7][2]~15_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_2_5),
	.prn(vcc));
defparam \ram_in_reg[5][2] .is_wysiwyg = "true";
defparam \ram_in_reg[5][2] .power_up = "low";

dffeas \ram_in_reg[4][2] (
	.clk(clk),
	.d(\ram_in_reg[4][2]~14_combout ),
	.asdata(\ram_in_reg[6][2]~12_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_2_4),
	.prn(vcc));
defparam \ram_in_reg[4][2] .is_wysiwyg = "true";
defparam \ram_in_reg[4][2] .power_up = "low";

dffeas \ram_in_reg[7][2] (
	.clk(clk),
	.d(\ram_in_reg[7][2]~15_combout ),
	.asdata(\ram_in_reg[5][2]~13_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_2_7),
	.prn(vcc));
defparam \ram_in_reg[7][2] .is_wysiwyg = "true";
defparam \ram_in_reg[7][2] .power_up = "low";

dffeas \ram_in_reg[2][1] (
	.clk(clk),
	.d(\ram_in_reg[2][1]~1_combout ),
	.asdata(\ram_in_reg[0][1]~2_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_1_2),
	.prn(vcc));
defparam \ram_in_reg[2][1] .is_wysiwyg = "true";
defparam \ram_in_reg[2][1] .power_up = "low";

dffeas \ram_in_reg[1][1] (
	.clk(clk),
	.d(\ram_in_reg[1][1]~0_combout ),
	.asdata(\ram_in_reg[3][1]~3_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_1_1),
	.prn(vcc));
defparam \ram_in_reg[1][1] .is_wysiwyg = "true";
defparam \ram_in_reg[1][1] .power_up = "low";

dffeas \ram_in_reg[0][1] (
	.clk(clk),
	.d(\ram_in_reg[0][1]~2_combout ),
	.asdata(\ram_in_reg[2][1]~1_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_1_0),
	.prn(vcc));
defparam \ram_in_reg[0][1] .is_wysiwyg = "true";
defparam \ram_in_reg[0][1] .power_up = "low";

dffeas \ram_in_reg[3][1] (
	.clk(clk),
	.d(\ram_in_reg[3][1]~3_combout ),
	.asdata(\ram_in_reg[1][1]~0_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_1_3),
	.prn(vcc));
defparam \ram_in_reg[3][1] .is_wysiwyg = "true";
defparam \ram_in_reg[3][1] .power_up = "low";

dffeas \ram_in_reg[2][0] (
	.clk(clk),
	.d(\ram_in_reg[2][0]~56_combout ),
	.asdata(\ram_in_reg[0][0]~58_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_0_2),
	.prn(vcc));
defparam \ram_in_reg[2][0] .is_wysiwyg = "true";
defparam \ram_in_reg[2][0] .power_up = "low";

dffeas \ram_in_reg[1][0] (
	.clk(clk),
	.d(\ram_in_reg[1][0]~57_combout ),
	.asdata(\ram_in_reg[3][0]~59_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_0_1),
	.prn(vcc));
defparam \ram_in_reg[1][0] .is_wysiwyg = "true";
defparam \ram_in_reg[1][0] .power_up = "low";

dffeas \ram_in_reg[0][0] (
	.clk(clk),
	.d(\ram_in_reg[0][0]~58_combout ),
	.asdata(\ram_in_reg[2][0]~56_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_0_0),
	.prn(vcc));
defparam \ram_in_reg[0][0] .is_wysiwyg = "true";
defparam \ram_in_reg[0][0] .power_up = "low";

dffeas \ram_in_reg[3][0] (
	.clk(clk),
	.d(\ram_in_reg[3][0]~59_combout ),
	.asdata(\ram_in_reg[1][0]~57_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_0_3),
	.prn(vcc));
defparam \ram_in_reg[3][0] .is_wysiwyg = "true";
defparam \ram_in_reg[3][0] .power_up = "low";

dffeas \ram_in_reg[2][7] (
	.clk(clk),
	.d(\ram_in_reg[2][7]~49_combout ),
	.asdata(\ram_in_reg[0][7]~50_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_7_2),
	.prn(vcc));
defparam \ram_in_reg[2][7] .is_wysiwyg = "true";
defparam \ram_in_reg[2][7] .power_up = "low";

dffeas \ram_in_reg[1][7] (
	.clk(clk),
	.d(\ram_in_reg[1][7]~48_combout ),
	.asdata(\ram_in_reg[3][7]~51_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_7_1),
	.prn(vcc));
defparam \ram_in_reg[1][7] .is_wysiwyg = "true";
defparam \ram_in_reg[1][7] .power_up = "low";

dffeas \ram_in_reg[0][7] (
	.clk(clk),
	.d(\ram_in_reg[0][7]~50_combout ),
	.asdata(\ram_in_reg[2][7]~49_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_7_0),
	.prn(vcc));
defparam \ram_in_reg[0][7] .is_wysiwyg = "true";
defparam \ram_in_reg[0][7] .power_up = "low";

dffeas \ram_in_reg[3][7] (
	.clk(clk),
	.d(\ram_in_reg[3][7]~51_combout ),
	.asdata(\ram_in_reg[1][7]~48_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_7_3),
	.prn(vcc));
defparam \ram_in_reg[3][7] .is_wysiwyg = "true";
defparam \ram_in_reg[3][7] .power_up = "low";

dffeas \ram_in_reg[2][6] (
	.clk(clk),
	.d(\ram_in_reg[2][6]~40_combout ),
	.asdata(\ram_in_reg[0][6]~42_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_6_2),
	.prn(vcc));
defparam \ram_in_reg[2][6] .is_wysiwyg = "true";
defparam \ram_in_reg[2][6] .power_up = "low";

dffeas \ram_in_reg[1][6] (
	.clk(clk),
	.d(\ram_in_reg[1][6]~41_combout ),
	.asdata(\ram_in_reg[3][6]~43_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_6_1),
	.prn(vcc));
defparam \ram_in_reg[1][6] .is_wysiwyg = "true";
defparam \ram_in_reg[1][6] .power_up = "low";

dffeas \ram_in_reg[0][6] (
	.clk(clk),
	.d(\ram_in_reg[0][6]~42_combout ),
	.asdata(\ram_in_reg[2][6]~40_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_6_0),
	.prn(vcc));
defparam \ram_in_reg[0][6] .is_wysiwyg = "true";
defparam \ram_in_reg[0][6] .power_up = "low";

dffeas \ram_in_reg[3][6] (
	.clk(clk),
	.d(\ram_in_reg[3][6]~43_combout ),
	.asdata(\ram_in_reg[1][6]~41_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_6_3),
	.prn(vcc));
defparam \ram_in_reg[3][6] .is_wysiwyg = "true";
defparam \ram_in_reg[3][6] .power_up = "low";

dffeas \ram_in_reg[2][5] (
	.clk(clk),
	.d(\ram_in_reg[2][5]~33_combout ),
	.asdata(\ram_in_reg[0][5]~34_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_5_2),
	.prn(vcc));
defparam \ram_in_reg[2][5] .is_wysiwyg = "true";
defparam \ram_in_reg[2][5] .power_up = "low";

dffeas \ram_in_reg[1][5] (
	.clk(clk),
	.d(\ram_in_reg[1][5]~32_combout ),
	.asdata(\ram_in_reg[3][5]~35_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_5_1),
	.prn(vcc));
defparam \ram_in_reg[1][5] .is_wysiwyg = "true";
defparam \ram_in_reg[1][5] .power_up = "low";

dffeas \ram_in_reg[0][5] (
	.clk(clk),
	.d(\ram_in_reg[0][5]~34_combout ),
	.asdata(\ram_in_reg[2][5]~33_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_5_0),
	.prn(vcc));
defparam \ram_in_reg[0][5] .is_wysiwyg = "true";
defparam \ram_in_reg[0][5] .power_up = "low";

dffeas \ram_in_reg[3][5] (
	.clk(clk),
	.d(\ram_in_reg[3][5]~35_combout ),
	.asdata(\ram_in_reg[1][5]~32_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_5_3),
	.prn(vcc));
defparam \ram_in_reg[3][5] .is_wysiwyg = "true";
defparam \ram_in_reg[3][5] .power_up = "low";

dffeas \ram_in_reg[2][4] (
	.clk(clk),
	.d(\ram_in_reg[2][4]~24_combout ),
	.asdata(\ram_in_reg[0][4]~26_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_4_2),
	.prn(vcc));
defparam \ram_in_reg[2][4] .is_wysiwyg = "true";
defparam \ram_in_reg[2][4] .power_up = "low";

dffeas \ram_in_reg[1][4] (
	.clk(clk),
	.d(\ram_in_reg[1][4]~25_combout ),
	.asdata(\ram_in_reg[3][4]~27_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_4_1),
	.prn(vcc));
defparam \ram_in_reg[1][4] .is_wysiwyg = "true";
defparam \ram_in_reg[1][4] .power_up = "low";

dffeas \ram_in_reg[0][4] (
	.clk(clk),
	.d(\ram_in_reg[0][4]~26_combout ),
	.asdata(\ram_in_reg[2][4]~24_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_4_0),
	.prn(vcc));
defparam \ram_in_reg[0][4] .is_wysiwyg = "true";
defparam \ram_in_reg[0][4] .power_up = "low";

dffeas \ram_in_reg[3][4] (
	.clk(clk),
	.d(\ram_in_reg[3][4]~27_combout ),
	.asdata(\ram_in_reg[1][4]~25_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_4_3),
	.prn(vcc));
defparam \ram_in_reg[3][4] .is_wysiwyg = "true";
defparam \ram_in_reg[3][4] .power_up = "low";

dffeas \ram_in_reg[2][3] (
	.clk(clk),
	.d(\ram_in_reg[2][3]~17_combout ),
	.asdata(\ram_in_reg[0][3]~18_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_3_2),
	.prn(vcc));
defparam \ram_in_reg[2][3] .is_wysiwyg = "true";
defparam \ram_in_reg[2][3] .power_up = "low";

dffeas \ram_in_reg[1][3] (
	.clk(clk),
	.d(\ram_in_reg[1][3]~16_combout ),
	.asdata(\ram_in_reg[3][3]~19_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_3_1),
	.prn(vcc));
defparam \ram_in_reg[1][3] .is_wysiwyg = "true";
defparam \ram_in_reg[1][3] .power_up = "low";

dffeas \ram_in_reg[0][3] (
	.clk(clk),
	.d(\ram_in_reg[0][3]~18_combout ),
	.asdata(\ram_in_reg[2][3]~17_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_3_0),
	.prn(vcc));
defparam \ram_in_reg[0][3] .is_wysiwyg = "true";
defparam \ram_in_reg[0][3] .power_up = "low";

dffeas \ram_in_reg[3][3] (
	.clk(clk),
	.d(\ram_in_reg[3][3]~19_combout ),
	.asdata(\ram_in_reg[1][3]~16_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_3_3),
	.prn(vcc));
defparam \ram_in_reg[3][3] .is_wysiwyg = "true";
defparam \ram_in_reg[3][3] .power_up = "low";

dffeas \ram_in_reg[2][2] (
	.clk(clk),
	.d(\ram_in_reg[2][2]~8_combout ),
	.asdata(\ram_in_reg[0][2]~10_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_2_2),
	.prn(vcc));
defparam \ram_in_reg[2][2] .is_wysiwyg = "true";
defparam \ram_in_reg[2][2] .power_up = "low";

dffeas \ram_in_reg[1][2] (
	.clk(clk),
	.d(\ram_in_reg[1][2]~9_combout ),
	.asdata(\ram_in_reg[3][2]~11_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_2_1),
	.prn(vcc));
defparam \ram_in_reg[1][2] .is_wysiwyg = "true";
defparam \ram_in_reg[1][2] .power_up = "low";

dffeas \ram_in_reg[0][2] (
	.clk(clk),
	.d(\ram_in_reg[0][2]~10_combout ),
	.asdata(\ram_in_reg[2][2]~8_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_2_0),
	.prn(vcc));
defparam \ram_in_reg[0][2] .is_wysiwyg = "true";
defparam \ram_in_reg[0][2] .power_up = "low";

dffeas \ram_in_reg[3][2] (
	.clk(clk),
	.d(\ram_in_reg[3][2]~11_combout ),
	.asdata(\ram_in_reg[1][2]~9_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_0),
	.ena(global_clock_enable),
	.q(ram_in_reg_2_3),
	.prn(vcc));
defparam \ram_in_reg[3][2] .is_wysiwyg = "true";
defparam \ram_in_reg[3][2] .power_up = "low";

cycloneiii_lcell_comb \ram_in_reg[6][1]~5 (
	.dataa(i_array_out_1_2),
	.datab(i_array_out_1_1),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[6][1]~5_combout ),
	.cout());
defparam \ram_in_reg[6][1]~5 .lut_mask = 16'hAACC;
defparam \ram_in_reg[6][1]~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[4][1]~6 (
	.dataa(i_array_out_1_0),
	.datab(i_array_out_1_3),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[4][1]~6_combout ),
	.cout());
defparam \ram_in_reg[4][1]~6 .lut_mask = 16'hAACC;
defparam \ram_in_reg[4][1]~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[5][1]~4 (
	.dataa(i_array_out_1_1),
	.datab(i_array_out_1_0),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[5][1]~4_combout ),
	.cout());
defparam \ram_in_reg[5][1]~4 .lut_mask = 16'hAACC;
defparam \ram_in_reg[5][1]~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[7][1]~7 (
	.dataa(i_array_out_1_3),
	.datab(i_array_out_1_2),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[7][1]~7_combout ),
	.cout());
defparam \ram_in_reg[7][1]~7 .lut_mask = 16'hAACC;
defparam \ram_in_reg[7][1]~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[6][0]~60 (
	.dataa(i_array_out_0_2),
	.datab(i_array_out_0_1),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[6][0]~60_combout ),
	.cout());
defparam \ram_in_reg[6][0]~60 .lut_mask = 16'hAACC;
defparam \ram_in_reg[6][0]~60 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[4][0]~62 (
	.dataa(i_array_out_0_0),
	.datab(i_array_out_0_3),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[4][0]~62_combout ),
	.cout());
defparam \ram_in_reg[4][0]~62 .lut_mask = 16'hAACC;
defparam \ram_in_reg[4][0]~62 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[5][0]~61 (
	.dataa(i_array_out_0_1),
	.datab(i_array_out_0_0),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[5][0]~61_combout ),
	.cout());
defparam \ram_in_reg[5][0]~61 .lut_mask = 16'hAACC;
defparam \ram_in_reg[5][0]~61 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[7][0]~63 (
	.dataa(i_array_out_0_3),
	.datab(i_array_out_0_2),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[7][0]~63_combout ),
	.cout());
defparam \ram_in_reg[7][0]~63 .lut_mask = 16'hAACC;
defparam \ram_in_reg[7][0]~63 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[6][7]~53 (
	.dataa(i_array_out_7_2),
	.datab(i_array_out_7_1),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[6][7]~53_combout ),
	.cout());
defparam \ram_in_reg[6][7]~53 .lut_mask = 16'hAACC;
defparam \ram_in_reg[6][7]~53 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[4][7]~54 (
	.dataa(i_array_out_7_0),
	.datab(i_array_out_7_3),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[4][7]~54_combout ),
	.cout());
defparam \ram_in_reg[4][7]~54 .lut_mask = 16'hAACC;
defparam \ram_in_reg[4][7]~54 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[5][7]~52 (
	.dataa(i_array_out_7_1),
	.datab(i_array_out_7_0),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[5][7]~52_combout ),
	.cout());
defparam \ram_in_reg[5][7]~52 .lut_mask = 16'hAACC;
defparam \ram_in_reg[5][7]~52 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[7][7]~55 (
	.dataa(i_array_out_7_3),
	.datab(i_array_out_7_2),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[7][7]~55_combout ),
	.cout());
defparam \ram_in_reg[7][7]~55 .lut_mask = 16'hAACC;
defparam \ram_in_reg[7][7]~55 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[6][6]~44 (
	.dataa(i_array_out_6_2),
	.datab(i_array_out_6_1),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[6][6]~44_combout ),
	.cout());
defparam \ram_in_reg[6][6]~44 .lut_mask = 16'hAACC;
defparam \ram_in_reg[6][6]~44 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[4][6]~46 (
	.dataa(i_array_out_6_0),
	.datab(i_array_out_6_3),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[4][6]~46_combout ),
	.cout());
defparam \ram_in_reg[4][6]~46 .lut_mask = 16'hAACC;
defparam \ram_in_reg[4][6]~46 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[5][6]~45 (
	.dataa(i_array_out_6_1),
	.datab(i_array_out_6_0),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[5][6]~45_combout ),
	.cout());
defparam \ram_in_reg[5][6]~45 .lut_mask = 16'hAACC;
defparam \ram_in_reg[5][6]~45 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[7][6]~47 (
	.dataa(i_array_out_6_3),
	.datab(i_array_out_6_2),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[7][6]~47_combout ),
	.cout());
defparam \ram_in_reg[7][6]~47 .lut_mask = 16'hAACC;
defparam \ram_in_reg[7][6]~47 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[6][5]~37 (
	.dataa(i_array_out_5_2),
	.datab(i_array_out_5_1),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[6][5]~37_combout ),
	.cout());
defparam \ram_in_reg[6][5]~37 .lut_mask = 16'hAACC;
defparam \ram_in_reg[6][5]~37 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[4][5]~38 (
	.dataa(i_array_out_5_0),
	.datab(i_array_out_5_3),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[4][5]~38_combout ),
	.cout());
defparam \ram_in_reg[4][5]~38 .lut_mask = 16'hAACC;
defparam \ram_in_reg[4][5]~38 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[5][5]~36 (
	.dataa(i_array_out_5_1),
	.datab(i_array_out_5_0),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[5][5]~36_combout ),
	.cout());
defparam \ram_in_reg[5][5]~36 .lut_mask = 16'hAACC;
defparam \ram_in_reg[5][5]~36 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[7][5]~39 (
	.dataa(i_array_out_5_3),
	.datab(i_array_out_5_2),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[7][5]~39_combout ),
	.cout());
defparam \ram_in_reg[7][5]~39 .lut_mask = 16'hAACC;
defparam \ram_in_reg[7][5]~39 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[6][4]~28 (
	.dataa(i_array_out_4_2),
	.datab(i_array_out_4_1),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[6][4]~28_combout ),
	.cout());
defparam \ram_in_reg[6][4]~28 .lut_mask = 16'hAACC;
defparam \ram_in_reg[6][4]~28 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[4][4]~30 (
	.dataa(i_array_out_4_0),
	.datab(i_array_out_4_3),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[4][4]~30_combout ),
	.cout());
defparam \ram_in_reg[4][4]~30 .lut_mask = 16'hAACC;
defparam \ram_in_reg[4][4]~30 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[5][4]~29 (
	.dataa(i_array_out_4_1),
	.datab(i_array_out_4_0),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[5][4]~29_combout ),
	.cout());
defparam \ram_in_reg[5][4]~29 .lut_mask = 16'hAACC;
defparam \ram_in_reg[5][4]~29 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[7][4]~31 (
	.dataa(i_array_out_4_3),
	.datab(i_array_out_4_2),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[7][4]~31_combout ),
	.cout());
defparam \ram_in_reg[7][4]~31 .lut_mask = 16'hAACC;
defparam \ram_in_reg[7][4]~31 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[6][3]~21 (
	.dataa(i_array_out_3_2),
	.datab(i_array_out_3_1),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[6][3]~21_combout ),
	.cout());
defparam \ram_in_reg[6][3]~21 .lut_mask = 16'hAACC;
defparam \ram_in_reg[6][3]~21 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[4][3]~22 (
	.dataa(i_array_out_3_0),
	.datab(i_array_out_3_3),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[4][3]~22_combout ),
	.cout());
defparam \ram_in_reg[4][3]~22 .lut_mask = 16'hAACC;
defparam \ram_in_reg[4][3]~22 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[5][3]~20 (
	.dataa(i_array_out_3_1),
	.datab(i_array_out_3_0),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[5][3]~20_combout ),
	.cout());
defparam \ram_in_reg[5][3]~20 .lut_mask = 16'hAACC;
defparam \ram_in_reg[5][3]~20 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[7][3]~23 (
	.dataa(i_array_out_3_3),
	.datab(i_array_out_3_2),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[7][3]~23_combout ),
	.cout());
defparam \ram_in_reg[7][3]~23 .lut_mask = 16'hAACC;
defparam \ram_in_reg[7][3]~23 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[6][2]~12 (
	.dataa(i_array_out_2_2),
	.datab(i_array_out_2_1),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[6][2]~12_combout ),
	.cout());
defparam \ram_in_reg[6][2]~12 .lut_mask = 16'hAACC;
defparam \ram_in_reg[6][2]~12 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[4][2]~14 (
	.dataa(i_array_out_2_0),
	.datab(i_array_out_2_3),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[4][2]~14_combout ),
	.cout());
defparam \ram_in_reg[4][2]~14 .lut_mask = 16'hAACC;
defparam \ram_in_reg[4][2]~14 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[5][2]~13 (
	.dataa(i_array_out_2_1),
	.datab(i_array_out_2_0),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[5][2]~13_combout ),
	.cout());
defparam \ram_in_reg[5][2]~13 .lut_mask = 16'hAACC;
defparam \ram_in_reg[5][2]~13 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[7][2]~15 (
	.dataa(i_array_out_2_3),
	.datab(i_array_out_2_2),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[7][2]~15_combout ),
	.cout());
defparam \ram_in_reg[7][2]~15 .lut_mask = 16'hAACC;
defparam \ram_in_reg[7][2]~15 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[2][1]~1 (
	.dataa(r_array_out_1_2),
	.datab(r_array_out_1_1),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[2][1]~1_combout ),
	.cout());
defparam \ram_in_reg[2][1]~1 .lut_mask = 16'hAACC;
defparam \ram_in_reg[2][1]~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[0][1]~2 (
	.dataa(r_array_out_1_0),
	.datab(r_array_out_1_3),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[0][1]~2_combout ),
	.cout());
defparam \ram_in_reg[0][1]~2 .lut_mask = 16'hAACC;
defparam \ram_in_reg[0][1]~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[1][1]~0 (
	.dataa(r_array_out_1_1),
	.datab(r_array_out_1_0),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[1][1]~0_combout ),
	.cout());
defparam \ram_in_reg[1][1]~0 .lut_mask = 16'hAACC;
defparam \ram_in_reg[1][1]~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[3][1]~3 (
	.dataa(r_array_out_1_3),
	.datab(r_array_out_1_2),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[3][1]~3_combout ),
	.cout());
defparam \ram_in_reg[3][1]~3 .lut_mask = 16'hAACC;
defparam \ram_in_reg[3][1]~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[2][0]~56 (
	.dataa(r_array_out_0_2),
	.datab(r_array_out_0_1),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[2][0]~56_combout ),
	.cout());
defparam \ram_in_reg[2][0]~56 .lut_mask = 16'hAACC;
defparam \ram_in_reg[2][0]~56 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[0][0]~58 (
	.dataa(r_array_out_0_0),
	.datab(r_array_out_0_3),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[0][0]~58_combout ),
	.cout());
defparam \ram_in_reg[0][0]~58 .lut_mask = 16'hAACC;
defparam \ram_in_reg[0][0]~58 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[1][0]~57 (
	.dataa(r_array_out_0_1),
	.datab(r_array_out_0_0),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[1][0]~57_combout ),
	.cout());
defparam \ram_in_reg[1][0]~57 .lut_mask = 16'hAACC;
defparam \ram_in_reg[1][0]~57 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[3][0]~59 (
	.dataa(r_array_out_0_3),
	.datab(r_array_out_0_2),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[3][0]~59_combout ),
	.cout());
defparam \ram_in_reg[3][0]~59 .lut_mask = 16'hAACC;
defparam \ram_in_reg[3][0]~59 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[2][7]~49 (
	.dataa(r_array_out_7_2),
	.datab(r_array_out_7_1),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[2][7]~49_combout ),
	.cout());
defparam \ram_in_reg[2][7]~49 .lut_mask = 16'hAACC;
defparam \ram_in_reg[2][7]~49 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[0][7]~50 (
	.dataa(r_array_out_7_0),
	.datab(r_array_out_7_3),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[0][7]~50_combout ),
	.cout());
defparam \ram_in_reg[0][7]~50 .lut_mask = 16'hAACC;
defparam \ram_in_reg[0][7]~50 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[1][7]~48 (
	.dataa(r_array_out_7_1),
	.datab(r_array_out_7_0),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[1][7]~48_combout ),
	.cout());
defparam \ram_in_reg[1][7]~48 .lut_mask = 16'hAACC;
defparam \ram_in_reg[1][7]~48 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[3][7]~51 (
	.dataa(r_array_out_7_3),
	.datab(r_array_out_7_2),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[3][7]~51_combout ),
	.cout());
defparam \ram_in_reg[3][7]~51 .lut_mask = 16'hAACC;
defparam \ram_in_reg[3][7]~51 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[2][6]~40 (
	.dataa(r_array_out_6_2),
	.datab(r_array_out_6_1),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[2][6]~40_combout ),
	.cout());
defparam \ram_in_reg[2][6]~40 .lut_mask = 16'hAACC;
defparam \ram_in_reg[2][6]~40 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[0][6]~42 (
	.dataa(r_array_out_6_0),
	.datab(r_array_out_6_3),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[0][6]~42_combout ),
	.cout());
defparam \ram_in_reg[0][6]~42 .lut_mask = 16'hAACC;
defparam \ram_in_reg[0][6]~42 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[1][6]~41 (
	.dataa(r_array_out_6_1),
	.datab(r_array_out_6_0),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[1][6]~41_combout ),
	.cout());
defparam \ram_in_reg[1][6]~41 .lut_mask = 16'hAACC;
defparam \ram_in_reg[1][6]~41 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[3][6]~43 (
	.dataa(r_array_out_6_3),
	.datab(r_array_out_6_2),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[3][6]~43_combout ),
	.cout());
defparam \ram_in_reg[3][6]~43 .lut_mask = 16'hAACC;
defparam \ram_in_reg[3][6]~43 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[2][5]~33 (
	.dataa(r_array_out_5_2),
	.datab(r_array_out_5_1),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[2][5]~33_combout ),
	.cout());
defparam \ram_in_reg[2][5]~33 .lut_mask = 16'hAACC;
defparam \ram_in_reg[2][5]~33 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[0][5]~34 (
	.dataa(r_array_out_5_0),
	.datab(r_array_out_5_3),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[0][5]~34_combout ),
	.cout());
defparam \ram_in_reg[0][5]~34 .lut_mask = 16'hAACC;
defparam \ram_in_reg[0][5]~34 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[1][5]~32 (
	.dataa(r_array_out_5_1),
	.datab(r_array_out_5_0),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[1][5]~32_combout ),
	.cout());
defparam \ram_in_reg[1][5]~32 .lut_mask = 16'hAACC;
defparam \ram_in_reg[1][5]~32 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[3][5]~35 (
	.dataa(r_array_out_5_3),
	.datab(r_array_out_5_2),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[3][5]~35_combout ),
	.cout());
defparam \ram_in_reg[3][5]~35 .lut_mask = 16'hAACC;
defparam \ram_in_reg[3][5]~35 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[2][4]~24 (
	.dataa(r_array_out_4_2),
	.datab(r_array_out_4_1),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[2][4]~24_combout ),
	.cout());
defparam \ram_in_reg[2][4]~24 .lut_mask = 16'hAACC;
defparam \ram_in_reg[2][4]~24 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[0][4]~26 (
	.dataa(r_array_out_4_0),
	.datab(r_array_out_4_3),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[0][4]~26_combout ),
	.cout());
defparam \ram_in_reg[0][4]~26 .lut_mask = 16'hAACC;
defparam \ram_in_reg[0][4]~26 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[1][4]~25 (
	.dataa(r_array_out_4_1),
	.datab(r_array_out_4_0),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[1][4]~25_combout ),
	.cout());
defparam \ram_in_reg[1][4]~25 .lut_mask = 16'hAACC;
defparam \ram_in_reg[1][4]~25 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[3][4]~27 (
	.dataa(r_array_out_4_3),
	.datab(r_array_out_4_2),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[3][4]~27_combout ),
	.cout());
defparam \ram_in_reg[3][4]~27 .lut_mask = 16'hAACC;
defparam \ram_in_reg[3][4]~27 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[2][3]~17 (
	.dataa(r_array_out_3_2),
	.datab(r_array_out_3_1),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[2][3]~17_combout ),
	.cout());
defparam \ram_in_reg[2][3]~17 .lut_mask = 16'hAACC;
defparam \ram_in_reg[2][3]~17 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[0][3]~18 (
	.dataa(r_array_out_3_0),
	.datab(r_array_out_3_3),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[0][3]~18_combout ),
	.cout());
defparam \ram_in_reg[0][3]~18 .lut_mask = 16'hAACC;
defparam \ram_in_reg[0][3]~18 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[1][3]~16 (
	.dataa(r_array_out_3_1),
	.datab(r_array_out_3_0),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[1][3]~16_combout ),
	.cout());
defparam \ram_in_reg[1][3]~16 .lut_mask = 16'hAACC;
defparam \ram_in_reg[1][3]~16 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[3][3]~19 (
	.dataa(r_array_out_3_3),
	.datab(r_array_out_3_2),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[3][3]~19_combout ),
	.cout());
defparam \ram_in_reg[3][3]~19 .lut_mask = 16'hAACC;
defparam \ram_in_reg[3][3]~19 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[2][2]~8 (
	.dataa(r_array_out_2_2),
	.datab(r_array_out_2_1),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[2][2]~8_combout ),
	.cout());
defparam \ram_in_reg[2][2]~8 .lut_mask = 16'hAACC;
defparam \ram_in_reg[2][2]~8 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[0][2]~10 (
	.dataa(r_array_out_2_0),
	.datab(r_array_out_2_3),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[0][2]~10_combout ),
	.cout());
defparam \ram_in_reg[0][2]~10 .lut_mask = 16'hAACC;
defparam \ram_in_reg[0][2]~10 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[1][2]~9 (
	.dataa(r_array_out_2_1),
	.datab(r_array_out_2_0),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[1][2]~9_combout ),
	.cout());
defparam \ram_in_reg[1][2]~9 .lut_mask = 16'hAACC;
defparam \ram_in_reg[1][2]~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[3][2]~11 (
	.dataa(r_array_out_2_3),
	.datab(r_array_out_2_2),
	.datac(gnd),
	.datad(swa_tdl_0_0),
	.cin(gnd),
	.combout(\ram_in_reg[3][2]~11_combout ),
	.cout());
defparam \ram_in_reg[3][2]~11 .lut_mask = 16'hAACC;
defparam \ram_in_reg[3][2]~11 .sum_lutc_input = "datac";

endmodule

module fft_asj_fft_cxb_data_r_fft_120 (
	ram_in_reg_2_0,
	ram_in_reg_6_0,
	ram_in_reg_4_0,
	ram_in_reg_3_0,
	ram_in_reg_5_0,
	ram_in_reg_2_2,
	ram_in_reg_6_2,
	ram_in_reg_4_2,
	ram_in_reg_3_2,
	ram_in_reg_5_2,
	ram_in_reg_1_0,
	ram_in_reg_1_2,
	ram_in_reg_0_0,
	ram_in_reg_0_2,
	ram_in_reg_2_1,
	ram_in_reg_6_1,
	ram_in_reg_4_1,
	ram_in_reg_3_1,
	ram_in_reg_5_1,
	ram_in_reg_2_3,
	ram_in_reg_6_3,
	ram_in_reg_4_3,
	ram_in_reg_3_3,
	ram_in_reg_5_3,
	ram_in_reg_1_1,
	ram_in_reg_1_3,
	ram_in_reg_0_1,
	ram_in_reg_0_3,
	ram_in_reg_7_0,
	ram_in_reg_7_2,
	ram_in_reg_7_1,
	ram_in_reg_7_3,
	ram_in_reg_7_4,
	ram_in_reg_3_4,
	ram_in_reg_5_4,
	ram_in_reg_4_4,
	ram_in_reg_6_4,
	ram_in_reg_7_6,
	ram_in_reg_3_6,
	ram_in_reg_5_6,
	ram_in_reg_4_6,
	ram_in_reg_6_6,
	ram_in_reg_2_4,
	ram_in_reg_2_6,
	ram_in_reg_1_4,
	ram_in_reg_1_6,
	ram_in_reg_0_4,
	ram_in_reg_0_6,
	ram_in_reg_7_5,
	ram_in_reg_3_5,
	ram_in_reg_5_5,
	ram_in_reg_4_5,
	ram_in_reg_6_5,
	ram_in_reg_3_7,
	ram_in_reg_7_7,
	ram_in_reg_5_7,
	ram_in_reg_4_7,
	ram_in_reg_6_7,
	ram_in_reg_2_5,
	ram_in_reg_2_7,
	ram_in_reg_1_5,
	ram_in_reg_1_7,
	ram_in_reg_0_5,
	ram_in_reg_0_7,
	global_clock_enable,
	ram_data_out0_10,
	ram_data_out1_10,
	sw_r_tdl_0_4,
	ram_data_out2_10,
	ram_data_out3_10,
	sw_r_tdl_1_4,
	ram_data_out0_14,
	ram_data_out1_14,
	ram_data_out2_14,
	ram_data_out3_14,
	ram_data_out0_12,
	ram_data_out1_12,
	ram_data_out2_12,
	ram_data_out3_12,
	ram_data_out0_11,
	ram_data_out1_11,
	ram_data_out2_11,
	ram_data_out3_11,
	ram_data_out0_13,
	ram_data_out1_13,
	ram_data_out2_13,
	ram_data_out3_13,
	ram_data_out0_9,
	ram_data_out1_9,
	ram_data_out2_9,
	ram_data_out3_9,
	ram_data_out0_8,
	ram_data_out1_8,
	ram_data_out2_8,
	ram_data_out3_8,
	ram_data_out0_15,
	ram_data_out1_15,
	ram_data_out2_15,
	ram_data_out3_15,
	ram_data_out0_7,
	ram_data_out1_7,
	ram_data_out2_7,
	ram_data_out3_7,
	ram_data_out0_3,
	ram_data_out1_3,
	ram_data_out2_3,
	ram_data_out3_3,
	ram_data_out0_5,
	ram_data_out1_5,
	ram_data_out2_5,
	ram_data_out3_5,
	ram_data_out0_4,
	ram_data_out1_4,
	ram_data_out2_4,
	ram_data_out3_4,
	ram_data_out0_6,
	ram_data_out1_6,
	ram_data_out2_6,
	ram_data_out3_6,
	ram_data_out0_2,
	ram_data_out1_2,
	ram_data_out2_2,
	ram_data_out3_2,
	ram_data_out0_1,
	ram_data_out1_1,
	ram_data_out2_1,
	ram_data_out3_1,
	ram_data_out0_0,
	ram_data_out1_0,
	ram_data_out2_0,
	ram_data_out3_0,
	clk)/* synthesis synthesis_greybox=1 */;
output 	ram_in_reg_2_0;
output 	ram_in_reg_6_0;
output 	ram_in_reg_4_0;
output 	ram_in_reg_3_0;
output 	ram_in_reg_5_0;
output 	ram_in_reg_2_2;
output 	ram_in_reg_6_2;
output 	ram_in_reg_4_2;
output 	ram_in_reg_3_2;
output 	ram_in_reg_5_2;
output 	ram_in_reg_1_0;
output 	ram_in_reg_1_2;
output 	ram_in_reg_0_0;
output 	ram_in_reg_0_2;
output 	ram_in_reg_2_1;
output 	ram_in_reg_6_1;
output 	ram_in_reg_4_1;
output 	ram_in_reg_3_1;
output 	ram_in_reg_5_1;
output 	ram_in_reg_2_3;
output 	ram_in_reg_6_3;
output 	ram_in_reg_4_3;
output 	ram_in_reg_3_3;
output 	ram_in_reg_5_3;
output 	ram_in_reg_1_1;
output 	ram_in_reg_1_3;
output 	ram_in_reg_0_1;
output 	ram_in_reg_0_3;
output 	ram_in_reg_7_0;
output 	ram_in_reg_7_2;
output 	ram_in_reg_7_1;
output 	ram_in_reg_7_3;
output 	ram_in_reg_7_4;
output 	ram_in_reg_3_4;
output 	ram_in_reg_5_4;
output 	ram_in_reg_4_4;
output 	ram_in_reg_6_4;
output 	ram_in_reg_7_6;
output 	ram_in_reg_3_6;
output 	ram_in_reg_5_6;
output 	ram_in_reg_4_6;
output 	ram_in_reg_6_6;
output 	ram_in_reg_2_4;
output 	ram_in_reg_2_6;
output 	ram_in_reg_1_4;
output 	ram_in_reg_1_6;
output 	ram_in_reg_0_4;
output 	ram_in_reg_0_6;
output 	ram_in_reg_7_5;
output 	ram_in_reg_3_5;
output 	ram_in_reg_5_5;
output 	ram_in_reg_4_5;
output 	ram_in_reg_6_5;
output 	ram_in_reg_3_7;
output 	ram_in_reg_7_7;
output 	ram_in_reg_5_7;
output 	ram_in_reg_4_7;
output 	ram_in_reg_6_7;
output 	ram_in_reg_2_5;
output 	ram_in_reg_2_7;
output 	ram_in_reg_1_5;
output 	ram_in_reg_1_7;
output 	ram_in_reg_0_5;
output 	ram_in_reg_0_7;
input 	global_clock_enable;
input 	ram_data_out0_10;
input 	ram_data_out1_10;
input 	sw_r_tdl_0_4;
input 	ram_data_out2_10;
input 	ram_data_out3_10;
input 	sw_r_tdl_1_4;
input 	ram_data_out0_14;
input 	ram_data_out1_14;
input 	ram_data_out2_14;
input 	ram_data_out3_14;
input 	ram_data_out0_12;
input 	ram_data_out1_12;
input 	ram_data_out2_12;
input 	ram_data_out3_12;
input 	ram_data_out0_11;
input 	ram_data_out1_11;
input 	ram_data_out2_11;
input 	ram_data_out3_11;
input 	ram_data_out0_13;
input 	ram_data_out1_13;
input 	ram_data_out2_13;
input 	ram_data_out3_13;
input 	ram_data_out0_9;
input 	ram_data_out1_9;
input 	ram_data_out2_9;
input 	ram_data_out3_9;
input 	ram_data_out0_8;
input 	ram_data_out1_8;
input 	ram_data_out2_8;
input 	ram_data_out3_8;
input 	ram_data_out0_15;
input 	ram_data_out1_15;
input 	ram_data_out2_15;
input 	ram_data_out3_15;
input 	ram_data_out0_7;
input 	ram_data_out1_7;
input 	ram_data_out2_7;
input 	ram_data_out3_7;
input 	ram_data_out0_3;
input 	ram_data_out1_3;
input 	ram_data_out2_3;
input 	ram_data_out3_3;
input 	ram_data_out0_5;
input 	ram_data_out1_5;
input 	ram_data_out2_5;
input 	ram_data_out3_5;
input 	ram_data_out0_4;
input 	ram_data_out1_4;
input 	ram_data_out2_4;
input 	ram_data_out3_4;
input 	ram_data_out0_6;
input 	ram_data_out1_6;
input 	ram_data_out2_6;
input 	ram_data_out3_6;
input 	ram_data_out0_2;
input 	ram_data_out1_2;
input 	ram_data_out2_2;
input 	ram_data_out3_2;
input 	ram_data_out0_1;
input 	ram_data_out1_1;
input 	ram_data_out2_1;
input 	ram_data_out3_1;
input 	ram_data_out0_0;
input 	ram_data_out1_0;
input 	ram_data_out2_0;
input 	ram_data_out3_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ram_in_reg[0][2]~0_combout ;
wire \ram_in_reg[2][2]~5_combout ;
wire \ram_in_reg[0][6]~1_combout ;
wire \ram_in_reg[2][6]~6_combout ;
wire \ram_in_reg[0][4]~2_combout ;
wire \ram_in_reg[2][4]~7_combout ;
wire \ram_in_reg[0][3]~3_combout ;
wire \ram_in_reg[2][3]~8_combout ;
wire \ram_in_reg[0][5]~4_combout ;
wire \ram_in_reg[2][5]~9_combout ;
wire \ram_in_reg[0][1]~57_combout ;
wire \ram_in_reg[2][1]~59_combout ;
wire \ram_in_reg[0][0]~56_combout ;
wire \ram_in_reg[2][0]~58_combout ;
wire \ram_in_reg[1][2]~10_combout ;
wire \ram_in_reg[3][2]~15_combout ;
wire \ram_in_reg[1][6]~11_combout ;
wire \ram_in_reg[3][6]~16_combout ;
wire \ram_in_reg[1][4]~12_combout ;
wire \ram_in_reg[3][4]~17_combout ;
wire \ram_in_reg[1][3]~13_combout ;
wire \ram_in_reg[3][3]~18_combout ;
wire \ram_in_reg[1][5]~14_combout ;
wire \ram_in_reg[3][5]~19_combout ;
wire \ram_in_reg[1][1]~53_combout ;
wire \ram_in_reg[3][1]~55_combout ;
wire \ram_in_reg[1][0]~52_combout ;
wire \ram_in_reg[3][0]~54_combout ;
wire \ram_in_reg[0][7]~20_combout ;
wire \ram_in_reg[2][7]~21_combout ;
wire \ram_in_reg[1][7]~22_combout ;
wire \ram_in_reg[3][7]~23_combout ;
wire \ram_in_reg[4][7]~24_combout ;
wire \ram_in_reg[6][7]~29_combout ;
wire \ram_in_reg[4][3]~25_combout ;
wire \ram_in_reg[6][3]~30_combout ;
wire \ram_in_reg[4][5]~26_combout ;
wire \ram_in_reg[6][5]~31_combout ;
wire \ram_in_reg[4][4]~27_combout ;
wire \ram_in_reg[6][4]~32_combout ;
wire \ram_in_reg[4][6]~28_combout ;
wire \ram_in_reg[6][6]~33_combout ;
wire \ram_in_reg[4][2]~44_combout ;
wire \ram_in_reg[6][2]~45_combout ;
wire \ram_in_reg[4][1]~49_combout ;
wire \ram_in_reg[6][1]~51_combout ;
wire \ram_in_reg[4][0]~48_combout ;
wire \ram_in_reg[6][0]~50_combout ;
wire \ram_in_reg[5][7]~34_combout ;
wire \ram_in_reg[7][7]~40_combout ;
wire \ram_in_reg[5][3]~35_combout ;
wire \ram_in_reg[7][3]~39_combout ;
wire \ram_in_reg[5][5]~36_combout ;
wire \ram_in_reg[7][5]~41_combout ;
wire \ram_in_reg[5][4]~37_combout ;
wire \ram_in_reg[7][4]~42_combout ;
wire \ram_in_reg[5][6]~38_combout ;
wire \ram_in_reg[7][6]~43_combout ;
wire \ram_in_reg[5][2]~46_combout ;
wire \ram_in_reg[7][2]~47_combout ;
wire \ram_in_reg[5][1]~61_combout ;
wire \ram_in_reg[7][1]~63_combout ;
wire \ram_in_reg[5][0]~60_combout ;
wire \ram_in_reg[7][0]~62_combout ;


dffeas \ram_in_reg[0][2] (
	.clk(clk),
	.d(\ram_in_reg[0][2]~0_combout ),
	.asdata(\ram_in_reg[2][2]~5_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_2_0),
	.prn(vcc));
defparam \ram_in_reg[0][2] .is_wysiwyg = "true";
defparam \ram_in_reg[0][2] .power_up = "low";

dffeas \ram_in_reg[0][6] (
	.clk(clk),
	.d(\ram_in_reg[0][6]~1_combout ),
	.asdata(\ram_in_reg[2][6]~6_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_6_0),
	.prn(vcc));
defparam \ram_in_reg[0][6] .is_wysiwyg = "true";
defparam \ram_in_reg[0][6] .power_up = "low";

dffeas \ram_in_reg[0][4] (
	.clk(clk),
	.d(\ram_in_reg[0][4]~2_combout ),
	.asdata(\ram_in_reg[2][4]~7_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_4_0),
	.prn(vcc));
defparam \ram_in_reg[0][4] .is_wysiwyg = "true";
defparam \ram_in_reg[0][4] .power_up = "low";

dffeas \ram_in_reg[0][3] (
	.clk(clk),
	.d(\ram_in_reg[0][3]~3_combout ),
	.asdata(\ram_in_reg[2][3]~8_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_3_0),
	.prn(vcc));
defparam \ram_in_reg[0][3] .is_wysiwyg = "true";
defparam \ram_in_reg[0][3] .power_up = "low";

dffeas \ram_in_reg[0][5] (
	.clk(clk),
	.d(\ram_in_reg[0][5]~4_combout ),
	.asdata(\ram_in_reg[2][5]~9_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_5_0),
	.prn(vcc));
defparam \ram_in_reg[0][5] .is_wysiwyg = "true";
defparam \ram_in_reg[0][5] .power_up = "low";

dffeas \ram_in_reg[2][2] (
	.clk(clk),
	.d(\ram_in_reg[2][2]~5_combout ),
	.asdata(\ram_in_reg[0][2]~0_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_2_2),
	.prn(vcc));
defparam \ram_in_reg[2][2] .is_wysiwyg = "true";
defparam \ram_in_reg[2][2] .power_up = "low";

dffeas \ram_in_reg[2][6] (
	.clk(clk),
	.d(\ram_in_reg[2][6]~6_combout ),
	.asdata(\ram_in_reg[0][6]~1_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_6_2),
	.prn(vcc));
defparam \ram_in_reg[2][6] .is_wysiwyg = "true";
defparam \ram_in_reg[2][6] .power_up = "low";

dffeas \ram_in_reg[2][4] (
	.clk(clk),
	.d(\ram_in_reg[2][4]~7_combout ),
	.asdata(\ram_in_reg[0][4]~2_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_4_2),
	.prn(vcc));
defparam \ram_in_reg[2][4] .is_wysiwyg = "true";
defparam \ram_in_reg[2][4] .power_up = "low";

dffeas \ram_in_reg[2][3] (
	.clk(clk),
	.d(\ram_in_reg[2][3]~8_combout ),
	.asdata(\ram_in_reg[0][3]~3_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_3_2),
	.prn(vcc));
defparam \ram_in_reg[2][3] .is_wysiwyg = "true";
defparam \ram_in_reg[2][3] .power_up = "low";

dffeas \ram_in_reg[2][5] (
	.clk(clk),
	.d(\ram_in_reg[2][5]~9_combout ),
	.asdata(\ram_in_reg[0][5]~4_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_5_2),
	.prn(vcc));
defparam \ram_in_reg[2][5] .is_wysiwyg = "true";
defparam \ram_in_reg[2][5] .power_up = "low";

dffeas \ram_in_reg[0][1] (
	.clk(clk),
	.d(\ram_in_reg[0][1]~57_combout ),
	.asdata(\ram_in_reg[2][1]~59_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_1_0),
	.prn(vcc));
defparam \ram_in_reg[0][1] .is_wysiwyg = "true";
defparam \ram_in_reg[0][1] .power_up = "low";

dffeas \ram_in_reg[2][1] (
	.clk(clk),
	.d(\ram_in_reg[2][1]~59_combout ),
	.asdata(\ram_in_reg[0][1]~57_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_1_2),
	.prn(vcc));
defparam \ram_in_reg[2][1] .is_wysiwyg = "true";
defparam \ram_in_reg[2][1] .power_up = "low";

dffeas \ram_in_reg[0][0] (
	.clk(clk),
	.d(\ram_in_reg[0][0]~56_combout ),
	.asdata(\ram_in_reg[2][0]~58_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_0_0),
	.prn(vcc));
defparam \ram_in_reg[0][0] .is_wysiwyg = "true";
defparam \ram_in_reg[0][0] .power_up = "low";

dffeas \ram_in_reg[2][0] (
	.clk(clk),
	.d(\ram_in_reg[2][0]~58_combout ),
	.asdata(\ram_in_reg[0][0]~56_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_0_2),
	.prn(vcc));
defparam \ram_in_reg[2][0] .is_wysiwyg = "true";
defparam \ram_in_reg[2][0] .power_up = "low";

dffeas \ram_in_reg[1][2] (
	.clk(clk),
	.d(\ram_in_reg[1][2]~10_combout ),
	.asdata(\ram_in_reg[3][2]~15_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_2_1),
	.prn(vcc));
defparam \ram_in_reg[1][2] .is_wysiwyg = "true";
defparam \ram_in_reg[1][2] .power_up = "low";

dffeas \ram_in_reg[1][6] (
	.clk(clk),
	.d(\ram_in_reg[1][6]~11_combout ),
	.asdata(\ram_in_reg[3][6]~16_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_6_1),
	.prn(vcc));
defparam \ram_in_reg[1][6] .is_wysiwyg = "true";
defparam \ram_in_reg[1][6] .power_up = "low";

dffeas \ram_in_reg[1][4] (
	.clk(clk),
	.d(\ram_in_reg[1][4]~12_combout ),
	.asdata(\ram_in_reg[3][4]~17_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_4_1),
	.prn(vcc));
defparam \ram_in_reg[1][4] .is_wysiwyg = "true";
defparam \ram_in_reg[1][4] .power_up = "low";

dffeas \ram_in_reg[1][3] (
	.clk(clk),
	.d(\ram_in_reg[1][3]~13_combout ),
	.asdata(\ram_in_reg[3][3]~18_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_3_1),
	.prn(vcc));
defparam \ram_in_reg[1][3] .is_wysiwyg = "true";
defparam \ram_in_reg[1][3] .power_up = "low";

dffeas \ram_in_reg[1][5] (
	.clk(clk),
	.d(\ram_in_reg[1][5]~14_combout ),
	.asdata(\ram_in_reg[3][5]~19_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_5_1),
	.prn(vcc));
defparam \ram_in_reg[1][5] .is_wysiwyg = "true";
defparam \ram_in_reg[1][5] .power_up = "low";

dffeas \ram_in_reg[3][2] (
	.clk(clk),
	.d(\ram_in_reg[3][2]~15_combout ),
	.asdata(\ram_in_reg[1][2]~10_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_2_3),
	.prn(vcc));
defparam \ram_in_reg[3][2] .is_wysiwyg = "true";
defparam \ram_in_reg[3][2] .power_up = "low";

dffeas \ram_in_reg[3][6] (
	.clk(clk),
	.d(\ram_in_reg[3][6]~16_combout ),
	.asdata(\ram_in_reg[1][6]~11_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_6_3),
	.prn(vcc));
defparam \ram_in_reg[3][6] .is_wysiwyg = "true";
defparam \ram_in_reg[3][6] .power_up = "low";

dffeas \ram_in_reg[3][4] (
	.clk(clk),
	.d(\ram_in_reg[3][4]~17_combout ),
	.asdata(\ram_in_reg[1][4]~12_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_4_3),
	.prn(vcc));
defparam \ram_in_reg[3][4] .is_wysiwyg = "true";
defparam \ram_in_reg[3][4] .power_up = "low";

dffeas \ram_in_reg[3][3] (
	.clk(clk),
	.d(\ram_in_reg[3][3]~18_combout ),
	.asdata(\ram_in_reg[1][3]~13_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_3_3),
	.prn(vcc));
defparam \ram_in_reg[3][3] .is_wysiwyg = "true";
defparam \ram_in_reg[3][3] .power_up = "low";

dffeas \ram_in_reg[3][5] (
	.clk(clk),
	.d(\ram_in_reg[3][5]~19_combout ),
	.asdata(\ram_in_reg[1][5]~14_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_5_3),
	.prn(vcc));
defparam \ram_in_reg[3][5] .is_wysiwyg = "true";
defparam \ram_in_reg[3][5] .power_up = "low";

dffeas \ram_in_reg[1][1] (
	.clk(clk),
	.d(\ram_in_reg[1][1]~53_combout ),
	.asdata(\ram_in_reg[3][1]~55_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_1_1),
	.prn(vcc));
defparam \ram_in_reg[1][1] .is_wysiwyg = "true";
defparam \ram_in_reg[1][1] .power_up = "low";

dffeas \ram_in_reg[3][1] (
	.clk(clk),
	.d(\ram_in_reg[3][1]~55_combout ),
	.asdata(\ram_in_reg[1][1]~53_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_1_3),
	.prn(vcc));
defparam \ram_in_reg[3][1] .is_wysiwyg = "true";
defparam \ram_in_reg[3][1] .power_up = "low";

dffeas \ram_in_reg[1][0] (
	.clk(clk),
	.d(\ram_in_reg[1][0]~52_combout ),
	.asdata(\ram_in_reg[3][0]~54_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_0_1),
	.prn(vcc));
defparam \ram_in_reg[1][0] .is_wysiwyg = "true";
defparam \ram_in_reg[1][0] .power_up = "low";

dffeas \ram_in_reg[3][0] (
	.clk(clk),
	.d(\ram_in_reg[3][0]~54_combout ),
	.asdata(\ram_in_reg[1][0]~52_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_0_3),
	.prn(vcc));
defparam \ram_in_reg[3][0] .is_wysiwyg = "true";
defparam \ram_in_reg[3][0] .power_up = "low";

dffeas \ram_in_reg[0][7] (
	.clk(clk),
	.d(\ram_in_reg[0][7]~20_combout ),
	.asdata(\ram_in_reg[2][7]~21_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_7_0),
	.prn(vcc));
defparam \ram_in_reg[0][7] .is_wysiwyg = "true";
defparam \ram_in_reg[0][7] .power_up = "low";

dffeas \ram_in_reg[2][7] (
	.clk(clk),
	.d(\ram_in_reg[2][7]~21_combout ),
	.asdata(\ram_in_reg[0][7]~20_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_7_2),
	.prn(vcc));
defparam \ram_in_reg[2][7] .is_wysiwyg = "true";
defparam \ram_in_reg[2][7] .power_up = "low";

dffeas \ram_in_reg[1][7] (
	.clk(clk),
	.d(\ram_in_reg[1][7]~22_combout ),
	.asdata(\ram_in_reg[3][7]~23_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_7_1),
	.prn(vcc));
defparam \ram_in_reg[1][7] .is_wysiwyg = "true";
defparam \ram_in_reg[1][7] .power_up = "low";

dffeas \ram_in_reg[3][7] (
	.clk(clk),
	.d(\ram_in_reg[3][7]~23_combout ),
	.asdata(\ram_in_reg[1][7]~22_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_7_3),
	.prn(vcc));
defparam \ram_in_reg[3][7] .is_wysiwyg = "true";
defparam \ram_in_reg[3][7] .power_up = "low";

dffeas \ram_in_reg[4][7] (
	.clk(clk),
	.d(\ram_in_reg[4][7]~24_combout ),
	.asdata(\ram_in_reg[6][7]~29_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_7_4),
	.prn(vcc));
defparam \ram_in_reg[4][7] .is_wysiwyg = "true";
defparam \ram_in_reg[4][7] .power_up = "low";

dffeas \ram_in_reg[4][3] (
	.clk(clk),
	.d(\ram_in_reg[4][3]~25_combout ),
	.asdata(\ram_in_reg[6][3]~30_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_3_4),
	.prn(vcc));
defparam \ram_in_reg[4][3] .is_wysiwyg = "true";
defparam \ram_in_reg[4][3] .power_up = "low";

dffeas \ram_in_reg[4][5] (
	.clk(clk),
	.d(\ram_in_reg[4][5]~26_combout ),
	.asdata(\ram_in_reg[6][5]~31_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_5_4),
	.prn(vcc));
defparam \ram_in_reg[4][5] .is_wysiwyg = "true";
defparam \ram_in_reg[4][5] .power_up = "low";

dffeas \ram_in_reg[4][4] (
	.clk(clk),
	.d(\ram_in_reg[4][4]~27_combout ),
	.asdata(\ram_in_reg[6][4]~32_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_4_4),
	.prn(vcc));
defparam \ram_in_reg[4][4] .is_wysiwyg = "true";
defparam \ram_in_reg[4][4] .power_up = "low";

dffeas \ram_in_reg[4][6] (
	.clk(clk),
	.d(\ram_in_reg[4][6]~28_combout ),
	.asdata(\ram_in_reg[6][6]~33_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_6_4),
	.prn(vcc));
defparam \ram_in_reg[4][6] .is_wysiwyg = "true";
defparam \ram_in_reg[4][6] .power_up = "low";

dffeas \ram_in_reg[6][7] (
	.clk(clk),
	.d(\ram_in_reg[6][7]~29_combout ),
	.asdata(\ram_in_reg[4][7]~24_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_7_6),
	.prn(vcc));
defparam \ram_in_reg[6][7] .is_wysiwyg = "true";
defparam \ram_in_reg[6][7] .power_up = "low";

dffeas \ram_in_reg[6][3] (
	.clk(clk),
	.d(\ram_in_reg[6][3]~30_combout ),
	.asdata(\ram_in_reg[4][3]~25_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_3_6),
	.prn(vcc));
defparam \ram_in_reg[6][3] .is_wysiwyg = "true";
defparam \ram_in_reg[6][3] .power_up = "low";

dffeas \ram_in_reg[6][5] (
	.clk(clk),
	.d(\ram_in_reg[6][5]~31_combout ),
	.asdata(\ram_in_reg[4][5]~26_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_5_6),
	.prn(vcc));
defparam \ram_in_reg[6][5] .is_wysiwyg = "true";
defparam \ram_in_reg[6][5] .power_up = "low";

dffeas \ram_in_reg[6][4] (
	.clk(clk),
	.d(\ram_in_reg[6][4]~32_combout ),
	.asdata(\ram_in_reg[4][4]~27_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_4_6),
	.prn(vcc));
defparam \ram_in_reg[6][4] .is_wysiwyg = "true";
defparam \ram_in_reg[6][4] .power_up = "low";

dffeas \ram_in_reg[6][6] (
	.clk(clk),
	.d(\ram_in_reg[6][6]~33_combout ),
	.asdata(\ram_in_reg[4][6]~28_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_6_6),
	.prn(vcc));
defparam \ram_in_reg[6][6] .is_wysiwyg = "true";
defparam \ram_in_reg[6][6] .power_up = "low";

dffeas \ram_in_reg[4][2] (
	.clk(clk),
	.d(\ram_in_reg[4][2]~44_combout ),
	.asdata(\ram_in_reg[6][2]~45_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_2_4),
	.prn(vcc));
defparam \ram_in_reg[4][2] .is_wysiwyg = "true";
defparam \ram_in_reg[4][2] .power_up = "low";

dffeas \ram_in_reg[6][2] (
	.clk(clk),
	.d(\ram_in_reg[6][2]~45_combout ),
	.asdata(\ram_in_reg[4][2]~44_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_2_6),
	.prn(vcc));
defparam \ram_in_reg[6][2] .is_wysiwyg = "true";
defparam \ram_in_reg[6][2] .power_up = "low";

dffeas \ram_in_reg[4][1] (
	.clk(clk),
	.d(\ram_in_reg[4][1]~49_combout ),
	.asdata(\ram_in_reg[6][1]~51_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_1_4),
	.prn(vcc));
defparam \ram_in_reg[4][1] .is_wysiwyg = "true";
defparam \ram_in_reg[4][1] .power_up = "low";

dffeas \ram_in_reg[6][1] (
	.clk(clk),
	.d(\ram_in_reg[6][1]~51_combout ),
	.asdata(\ram_in_reg[4][1]~49_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_1_6),
	.prn(vcc));
defparam \ram_in_reg[6][1] .is_wysiwyg = "true";
defparam \ram_in_reg[6][1] .power_up = "low";

dffeas \ram_in_reg[4][0] (
	.clk(clk),
	.d(\ram_in_reg[4][0]~48_combout ),
	.asdata(\ram_in_reg[6][0]~50_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_0_4),
	.prn(vcc));
defparam \ram_in_reg[4][0] .is_wysiwyg = "true";
defparam \ram_in_reg[4][0] .power_up = "low";

dffeas \ram_in_reg[6][0] (
	.clk(clk),
	.d(\ram_in_reg[6][0]~50_combout ),
	.asdata(\ram_in_reg[4][0]~48_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_0_6),
	.prn(vcc));
defparam \ram_in_reg[6][0] .is_wysiwyg = "true";
defparam \ram_in_reg[6][0] .power_up = "low";

dffeas \ram_in_reg[5][7] (
	.clk(clk),
	.d(\ram_in_reg[5][7]~34_combout ),
	.asdata(\ram_in_reg[7][7]~40_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_7_5),
	.prn(vcc));
defparam \ram_in_reg[5][7] .is_wysiwyg = "true";
defparam \ram_in_reg[5][7] .power_up = "low";

dffeas \ram_in_reg[5][3] (
	.clk(clk),
	.d(\ram_in_reg[5][3]~35_combout ),
	.asdata(\ram_in_reg[7][3]~39_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_3_5),
	.prn(vcc));
defparam \ram_in_reg[5][3] .is_wysiwyg = "true";
defparam \ram_in_reg[5][3] .power_up = "low";

dffeas \ram_in_reg[5][5] (
	.clk(clk),
	.d(\ram_in_reg[5][5]~36_combout ),
	.asdata(\ram_in_reg[7][5]~41_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_5_5),
	.prn(vcc));
defparam \ram_in_reg[5][5] .is_wysiwyg = "true";
defparam \ram_in_reg[5][5] .power_up = "low";

dffeas \ram_in_reg[5][4] (
	.clk(clk),
	.d(\ram_in_reg[5][4]~37_combout ),
	.asdata(\ram_in_reg[7][4]~42_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_4_5),
	.prn(vcc));
defparam \ram_in_reg[5][4] .is_wysiwyg = "true";
defparam \ram_in_reg[5][4] .power_up = "low";

dffeas \ram_in_reg[5][6] (
	.clk(clk),
	.d(\ram_in_reg[5][6]~38_combout ),
	.asdata(\ram_in_reg[7][6]~43_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_6_5),
	.prn(vcc));
defparam \ram_in_reg[5][6] .is_wysiwyg = "true";
defparam \ram_in_reg[5][6] .power_up = "low";

dffeas \ram_in_reg[7][3] (
	.clk(clk),
	.d(\ram_in_reg[7][3]~39_combout ),
	.asdata(\ram_in_reg[5][3]~35_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_3_7),
	.prn(vcc));
defparam \ram_in_reg[7][3] .is_wysiwyg = "true";
defparam \ram_in_reg[7][3] .power_up = "low";

dffeas \ram_in_reg[7][7] (
	.clk(clk),
	.d(\ram_in_reg[7][7]~40_combout ),
	.asdata(\ram_in_reg[5][7]~34_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_7_7),
	.prn(vcc));
defparam \ram_in_reg[7][7] .is_wysiwyg = "true";
defparam \ram_in_reg[7][7] .power_up = "low";

dffeas \ram_in_reg[7][5] (
	.clk(clk),
	.d(\ram_in_reg[7][5]~41_combout ),
	.asdata(\ram_in_reg[5][5]~36_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_5_7),
	.prn(vcc));
defparam \ram_in_reg[7][5] .is_wysiwyg = "true";
defparam \ram_in_reg[7][5] .power_up = "low";

dffeas \ram_in_reg[7][4] (
	.clk(clk),
	.d(\ram_in_reg[7][4]~42_combout ),
	.asdata(\ram_in_reg[5][4]~37_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_4_7),
	.prn(vcc));
defparam \ram_in_reg[7][4] .is_wysiwyg = "true";
defparam \ram_in_reg[7][4] .power_up = "low";

dffeas \ram_in_reg[7][6] (
	.clk(clk),
	.d(\ram_in_reg[7][6]~43_combout ),
	.asdata(\ram_in_reg[5][6]~38_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_6_7),
	.prn(vcc));
defparam \ram_in_reg[7][6] .is_wysiwyg = "true";
defparam \ram_in_reg[7][6] .power_up = "low";

dffeas \ram_in_reg[5][2] (
	.clk(clk),
	.d(\ram_in_reg[5][2]~46_combout ),
	.asdata(\ram_in_reg[7][2]~47_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_2_5),
	.prn(vcc));
defparam \ram_in_reg[5][2] .is_wysiwyg = "true";
defparam \ram_in_reg[5][2] .power_up = "low";

dffeas \ram_in_reg[7][2] (
	.clk(clk),
	.d(\ram_in_reg[7][2]~47_combout ),
	.asdata(\ram_in_reg[5][2]~46_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_2_7),
	.prn(vcc));
defparam \ram_in_reg[7][2] .is_wysiwyg = "true";
defparam \ram_in_reg[7][2] .power_up = "low";

dffeas \ram_in_reg[5][1] (
	.clk(clk),
	.d(\ram_in_reg[5][1]~61_combout ),
	.asdata(\ram_in_reg[7][1]~63_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_1_5),
	.prn(vcc));
defparam \ram_in_reg[5][1] .is_wysiwyg = "true";
defparam \ram_in_reg[5][1] .power_up = "low";

dffeas \ram_in_reg[7][1] (
	.clk(clk),
	.d(\ram_in_reg[7][1]~63_combout ),
	.asdata(\ram_in_reg[5][1]~61_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_1_7),
	.prn(vcc));
defparam \ram_in_reg[7][1] .is_wysiwyg = "true";
defparam \ram_in_reg[7][1] .power_up = "low";

dffeas \ram_in_reg[5][0] (
	.clk(clk),
	.d(\ram_in_reg[5][0]~60_combout ),
	.asdata(\ram_in_reg[7][0]~62_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_0_5),
	.prn(vcc));
defparam \ram_in_reg[5][0] .is_wysiwyg = "true";
defparam \ram_in_reg[5][0] .power_up = "low";

dffeas \ram_in_reg[7][0] (
	.clk(clk),
	.d(\ram_in_reg[7][0]~62_combout ),
	.asdata(\ram_in_reg[5][0]~60_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_0_7),
	.prn(vcc));
defparam \ram_in_reg[7][0] .is_wysiwyg = "true";
defparam \ram_in_reg[7][0] .power_up = "low";

cycloneiii_lcell_comb \ram_in_reg[0][2]~0 (
	.dataa(ram_data_out0_10),
	.datab(ram_data_out1_10),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[0][2]~0_combout ),
	.cout());
defparam \ram_in_reg[0][2]~0 .lut_mask = 16'hAACC;
defparam \ram_in_reg[0][2]~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[2][2]~5 (
	.dataa(ram_data_out2_10),
	.datab(ram_data_out3_10),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[2][2]~5_combout ),
	.cout());
defparam \ram_in_reg[2][2]~5 .lut_mask = 16'hAACC;
defparam \ram_in_reg[2][2]~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[0][6]~1 (
	.dataa(ram_data_out0_14),
	.datab(ram_data_out1_14),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[0][6]~1_combout ),
	.cout());
defparam \ram_in_reg[0][6]~1 .lut_mask = 16'hAACC;
defparam \ram_in_reg[0][6]~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[2][6]~6 (
	.dataa(ram_data_out2_14),
	.datab(ram_data_out3_14),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[2][6]~6_combout ),
	.cout());
defparam \ram_in_reg[2][6]~6 .lut_mask = 16'hAACC;
defparam \ram_in_reg[2][6]~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[0][4]~2 (
	.dataa(ram_data_out0_12),
	.datab(ram_data_out1_12),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[0][4]~2_combout ),
	.cout());
defparam \ram_in_reg[0][4]~2 .lut_mask = 16'hAACC;
defparam \ram_in_reg[0][4]~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[2][4]~7 (
	.dataa(ram_data_out2_12),
	.datab(ram_data_out3_12),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[2][4]~7_combout ),
	.cout());
defparam \ram_in_reg[2][4]~7 .lut_mask = 16'hAACC;
defparam \ram_in_reg[2][4]~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[0][3]~3 (
	.dataa(ram_data_out0_11),
	.datab(ram_data_out1_11),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[0][3]~3_combout ),
	.cout());
defparam \ram_in_reg[0][3]~3 .lut_mask = 16'hAACC;
defparam \ram_in_reg[0][3]~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[2][3]~8 (
	.dataa(ram_data_out2_11),
	.datab(ram_data_out3_11),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[2][3]~8_combout ),
	.cout());
defparam \ram_in_reg[2][3]~8 .lut_mask = 16'hAACC;
defparam \ram_in_reg[2][3]~8 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[0][5]~4 (
	.dataa(ram_data_out0_13),
	.datab(ram_data_out1_13),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[0][5]~4_combout ),
	.cout());
defparam \ram_in_reg[0][5]~4 .lut_mask = 16'hAACC;
defparam \ram_in_reg[0][5]~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[2][5]~9 (
	.dataa(ram_data_out2_13),
	.datab(ram_data_out3_13),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[2][5]~9_combout ),
	.cout());
defparam \ram_in_reg[2][5]~9 .lut_mask = 16'hAACC;
defparam \ram_in_reg[2][5]~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[0][1]~57 (
	.dataa(ram_data_out0_9),
	.datab(ram_data_out1_9),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[0][1]~57_combout ),
	.cout());
defparam \ram_in_reg[0][1]~57 .lut_mask = 16'hAACC;
defparam \ram_in_reg[0][1]~57 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[2][1]~59 (
	.dataa(ram_data_out2_9),
	.datab(ram_data_out3_9),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[2][1]~59_combout ),
	.cout());
defparam \ram_in_reg[2][1]~59 .lut_mask = 16'hAACC;
defparam \ram_in_reg[2][1]~59 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[0][0]~56 (
	.dataa(ram_data_out0_8),
	.datab(ram_data_out1_8),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[0][0]~56_combout ),
	.cout());
defparam \ram_in_reg[0][0]~56 .lut_mask = 16'hAACC;
defparam \ram_in_reg[0][0]~56 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[2][0]~58 (
	.dataa(ram_data_out2_8),
	.datab(ram_data_out3_8),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[2][0]~58_combout ),
	.cout());
defparam \ram_in_reg[2][0]~58 .lut_mask = 16'hAACC;
defparam \ram_in_reg[2][0]~58 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[1][2]~10 (
	.dataa(ram_data_out1_10),
	.datab(ram_data_out2_10),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[1][2]~10_combout ),
	.cout());
defparam \ram_in_reg[1][2]~10 .lut_mask = 16'hAACC;
defparam \ram_in_reg[1][2]~10 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[3][2]~15 (
	.dataa(ram_data_out3_10),
	.datab(ram_data_out0_10),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[3][2]~15_combout ),
	.cout());
defparam \ram_in_reg[3][2]~15 .lut_mask = 16'hAACC;
defparam \ram_in_reg[3][2]~15 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[1][6]~11 (
	.dataa(ram_data_out1_14),
	.datab(ram_data_out2_14),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[1][6]~11_combout ),
	.cout());
defparam \ram_in_reg[1][6]~11 .lut_mask = 16'hAACC;
defparam \ram_in_reg[1][6]~11 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[3][6]~16 (
	.dataa(ram_data_out3_14),
	.datab(ram_data_out0_14),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[3][6]~16_combout ),
	.cout());
defparam \ram_in_reg[3][6]~16 .lut_mask = 16'hAACC;
defparam \ram_in_reg[3][6]~16 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[1][4]~12 (
	.dataa(ram_data_out1_12),
	.datab(ram_data_out2_12),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[1][4]~12_combout ),
	.cout());
defparam \ram_in_reg[1][4]~12 .lut_mask = 16'hAACC;
defparam \ram_in_reg[1][4]~12 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[3][4]~17 (
	.dataa(ram_data_out3_12),
	.datab(ram_data_out0_12),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[3][4]~17_combout ),
	.cout());
defparam \ram_in_reg[3][4]~17 .lut_mask = 16'hAACC;
defparam \ram_in_reg[3][4]~17 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[1][3]~13 (
	.dataa(ram_data_out1_11),
	.datab(ram_data_out2_11),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[1][3]~13_combout ),
	.cout());
defparam \ram_in_reg[1][3]~13 .lut_mask = 16'hAACC;
defparam \ram_in_reg[1][3]~13 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[3][3]~18 (
	.dataa(ram_data_out3_11),
	.datab(ram_data_out0_11),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[3][3]~18_combout ),
	.cout());
defparam \ram_in_reg[3][3]~18 .lut_mask = 16'hAACC;
defparam \ram_in_reg[3][3]~18 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[1][5]~14 (
	.dataa(ram_data_out1_13),
	.datab(ram_data_out2_13),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[1][5]~14_combout ),
	.cout());
defparam \ram_in_reg[1][5]~14 .lut_mask = 16'hAACC;
defparam \ram_in_reg[1][5]~14 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[3][5]~19 (
	.dataa(ram_data_out3_13),
	.datab(ram_data_out0_13),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[3][5]~19_combout ),
	.cout());
defparam \ram_in_reg[3][5]~19 .lut_mask = 16'hAACC;
defparam \ram_in_reg[3][5]~19 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[1][1]~53 (
	.dataa(ram_data_out1_9),
	.datab(ram_data_out2_9),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[1][1]~53_combout ),
	.cout());
defparam \ram_in_reg[1][1]~53 .lut_mask = 16'hAACC;
defparam \ram_in_reg[1][1]~53 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[3][1]~55 (
	.dataa(ram_data_out3_9),
	.datab(ram_data_out0_9),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[3][1]~55_combout ),
	.cout());
defparam \ram_in_reg[3][1]~55 .lut_mask = 16'hAACC;
defparam \ram_in_reg[3][1]~55 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[1][0]~52 (
	.dataa(ram_data_out1_8),
	.datab(ram_data_out2_8),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[1][0]~52_combout ),
	.cout());
defparam \ram_in_reg[1][0]~52 .lut_mask = 16'hAACC;
defparam \ram_in_reg[1][0]~52 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[3][0]~54 (
	.dataa(ram_data_out3_8),
	.datab(ram_data_out0_8),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[3][0]~54_combout ),
	.cout());
defparam \ram_in_reg[3][0]~54 .lut_mask = 16'hAACC;
defparam \ram_in_reg[3][0]~54 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[0][7]~20 (
	.dataa(ram_data_out0_15),
	.datab(ram_data_out1_15),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[0][7]~20_combout ),
	.cout());
defparam \ram_in_reg[0][7]~20 .lut_mask = 16'hAACC;
defparam \ram_in_reg[0][7]~20 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[2][7]~21 (
	.dataa(ram_data_out2_15),
	.datab(ram_data_out3_15),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[2][7]~21_combout ),
	.cout());
defparam \ram_in_reg[2][7]~21 .lut_mask = 16'hAACC;
defparam \ram_in_reg[2][7]~21 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[1][7]~22 (
	.dataa(ram_data_out1_15),
	.datab(ram_data_out2_15),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[1][7]~22_combout ),
	.cout());
defparam \ram_in_reg[1][7]~22 .lut_mask = 16'hAACC;
defparam \ram_in_reg[1][7]~22 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[3][7]~23 (
	.dataa(ram_data_out3_15),
	.datab(ram_data_out0_15),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[3][7]~23_combout ),
	.cout());
defparam \ram_in_reg[3][7]~23 .lut_mask = 16'hAACC;
defparam \ram_in_reg[3][7]~23 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[4][7]~24 (
	.dataa(ram_data_out0_7),
	.datab(ram_data_out1_7),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[4][7]~24_combout ),
	.cout());
defparam \ram_in_reg[4][7]~24 .lut_mask = 16'hAACC;
defparam \ram_in_reg[4][7]~24 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[6][7]~29 (
	.dataa(ram_data_out2_7),
	.datab(ram_data_out3_7),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[6][7]~29_combout ),
	.cout());
defparam \ram_in_reg[6][7]~29 .lut_mask = 16'hAACC;
defparam \ram_in_reg[6][7]~29 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[4][3]~25 (
	.dataa(ram_data_out0_3),
	.datab(ram_data_out1_3),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[4][3]~25_combout ),
	.cout());
defparam \ram_in_reg[4][3]~25 .lut_mask = 16'hAACC;
defparam \ram_in_reg[4][3]~25 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[6][3]~30 (
	.dataa(ram_data_out2_3),
	.datab(ram_data_out3_3),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[6][3]~30_combout ),
	.cout());
defparam \ram_in_reg[6][3]~30 .lut_mask = 16'hAACC;
defparam \ram_in_reg[6][3]~30 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[4][5]~26 (
	.dataa(ram_data_out0_5),
	.datab(ram_data_out1_5),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[4][5]~26_combout ),
	.cout());
defparam \ram_in_reg[4][5]~26 .lut_mask = 16'hAACC;
defparam \ram_in_reg[4][5]~26 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[6][5]~31 (
	.dataa(ram_data_out2_5),
	.datab(ram_data_out3_5),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[6][5]~31_combout ),
	.cout());
defparam \ram_in_reg[6][5]~31 .lut_mask = 16'hAACC;
defparam \ram_in_reg[6][5]~31 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[4][4]~27 (
	.dataa(ram_data_out0_4),
	.datab(ram_data_out1_4),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[4][4]~27_combout ),
	.cout());
defparam \ram_in_reg[4][4]~27 .lut_mask = 16'hAACC;
defparam \ram_in_reg[4][4]~27 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[6][4]~32 (
	.dataa(ram_data_out2_4),
	.datab(ram_data_out3_4),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[6][4]~32_combout ),
	.cout());
defparam \ram_in_reg[6][4]~32 .lut_mask = 16'hAACC;
defparam \ram_in_reg[6][4]~32 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[4][6]~28 (
	.dataa(ram_data_out0_6),
	.datab(ram_data_out1_6),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[4][6]~28_combout ),
	.cout());
defparam \ram_in_reg[4][6]~28 .lut_mask = 16'hAACC;
defparam \ram_in_reg[4][6]~28 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[6][6]~33 (
	.dataa(ram_data_out2_6),
	.datab(ram_data_out3_6),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[6][6]~33_combout ),
	.cout());
defparam \ram_in_reg[6][6]~33 .lut_mask = 16'hAACC;
defparam \ram_in_reg[6][6]~33 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[4][2]~44 (
	.dataa(ram_data_out0_2),
	.datab(ram_data_out1_2),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[4][2]~44_combout ),
	.cout());
defparam \ram_in_reg[4][2]~44 .lut_mask = 16'hAACC;
defparam \ram_in_reg[4][2]~44 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[6][2]~45 (
	.dataa(ram_data_out2_2),
	.datab(ram_data_out3_2),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[6][2]~45_combout ),
	.cout());
defparam \ram_in_reg[6][2]~45 .lut_mask = 16'hAACC;
defparam \ram_in_reg[6][2]~45 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[4][1]~49 (
	.dataa(ram_data_out0_1),
	.datab(ram_data_out1_1),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[4][1]~49_combout ),
	.cout());
defparam \ram_in_reg[4][1]~49 .lut_mask = 16'hAACC;
defparam \ram_in_reg[4][1]~49 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[6][1]~51 (
	.dataa(ram_data_out2_1),
	.datab(ram_data_out3_1),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[6][1]~51_combout ),
	.cout());
defparam \ram_in_reg[6][1]~51 .lut_mask = 16'hAACC;
defparam \ram_in_reg[6][1]~51 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[4][0]~48 (
	.dataa(ram_data_out0_0),
	.datab(ram_data_out1_0),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[4][0]~48_combout ),
	.cout());
defparam \ram_in_reg[4][0]~48 .lut_mask = 16'hAACC;
defparam \ram_in_reg[4][0]~48 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[6][0]~50 (
	.dataa(ram_data_out2_0),
	.datab(ram_data_out3_0),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[6][0]~50_combout ),
	.cout());
defparam \ram_in_reg[6][0]~50 .lut_mask = 16'hAACC;
defparam \ram_in_reg[6][0]~50 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[5][7]~34 (
	.dataa(ram_data_out1_7),
	.datab(ram_data_out2_7),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[5][7]~34_combout ),
	.cout());
defparam \ram_in_reg[5][7]~34 .lut_mask = 16'hAACC;
defparam \ram_in_reg[5][7]~34 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[7][7]~40 (
	.dataa(ram_data_out3_7),
	.datab(ram_data_out0_7),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[7][7]~40_combout ),
	.cout());
defparam \ram_in_reg[7][7]~40 .lut_mask = 16'hAACC;
defparam \ram_in_reg[7][7]~40 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[5][3]~35 (
	.dataa(ram_data_out1_3),
	.datab(ram_data_out2_3),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[5][3]~35_combout ),
	.cout());
defparam \ram_in_reg[5][3]~35 .lut_mask = 16'hAACC;
defparam \ram_in_reg[5][3]~35 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[7][3]~39 (
	.dataa(ram_data_out3_3),
	.datab(ram_data_out0_3),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[7][3]~39_combout ),
	.cout());
defparam \ram_in_reg[7][3]~39 .lut_mask = 16'hAACC;
defparam \ram_in_reg[7][3]~39 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[5][5]~36 (
	.dataa(ram_data_out1_5),
	.datab(ram_data_out2_5),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[5][5]~36_combout ),
	.cout());
defparam \ram_in_reg[5][5]~36 .lut_mask = 16'hAACC;
defparam \ram_in_reg[5][5]~36 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[7][5]~41 (
	.dataa(ram_data_out3_5),
	.datab(ram_data_out0_5),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[7][5]~41_combout ),
	.cout());
defparam \ram_in_reg[7][5]~41 .lut_mask = 16'hAACC;
defparam \ram_in_reg[7][5]~41 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[5][4]~37 (
	.dataa(ram_data_out1_4),
	.datab(ram_data_out2_4),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[5][4]~37_combout ),
	.cout());
defparam \ram_in_reg[5][4]~37 .lut_mask = 16'hAACC;
defparam \ram_in_reg[5][4]~37 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[7][4]~42 (
	.dataa(ram_data_out3_4),
	.datab(ram_data_out0_4),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[7][4]~42_combout ),
	.cout());
defparam \ram_in_reg[7][4]~42 .lut_mask = 16'hAACC;
defparam \ram_in_reg[7][4]~42 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[5][6]~38 (
	.dataa(ram_data_out1_6),
	.datab(ram_data_out2_6),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[5][6]~38_combout ),
	.cout());
defparam \ram_in_reg[5][6]~38 .lut_mask = 16'hAACC;
defparam \ram_in_reg[5][6]~38 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[7][6]~43 (
	.dataa(ram_data_out3_6),
	.datab(ram_data_out0_6),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[7][6]~43_combout ),
	.cout());
defparam \ram_in_reg[7][6]~43 .lut_mask = 16'hAACC;
defparam \ram_in_reg[7][6]~43 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[5][2]~46 (
	.dataa(ram_data_out1_2),
	.datab(ram_data_out2_2),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[5][2]~46_combout ),
	.cout());
defparam \ram_in_reg[5][2]~46 .lut_mask = 16'hAACC;
defparam \ram_in_reg[5][2]~46 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[7][2]~47 (
	.dataa(ram_data_out3_2),
	.datab(ram_data_out0_2),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[7][2]~47_combout ),
	.cout());
defparam \ram_in_reg[7][2]~47 .lut_mask = 16'hAACC;
defparam \ram_in_reg[7][2]~47 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[5][1]~61 (
	.dataa(ram_data_out1_1),
	.datab(ram_data_out2_1),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[5][1]~61_combout ),
	.cout());
defparam \ram_in_reg[5][1]~61 .lut_mask = 16'hAACC;
defparam \ram_in_reg[5][1]~61 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[7][1]~63 (
	.dataa(ram_data_out3_1),
	.datab(ram_data_out0_1),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[7][1]~63_combout ),
	.cout());
defparam \ram_in_reg[7][1]~63 .lut_mask = 16'hAACC;
defparam \ram_in_reg[7][1]~63 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[5][0]~60 (
	.dataa(ram_data_out1_0),
	.datab(ram_data_out2_0),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[5][0]~60_combout ),
	.cout());
defparam \ram_in_reg[5][0]~60 .lut_mask = 16'hAACC;
defparam \ram_in_reg[5][0]~60 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ram_in_reg[7][0]~62 (
	.dataa(ram_data_out3_0),
	.datab(ram_data_out0_0),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[7][0]~62_combout ),
	.cout());
defparam \ram_in_reg[7][0]~62 .lut_mask = 16'hAACC;
defparam \ram_in_reg[7][0]~62 .sum_lutc_input = "datac";

endmodule

module fft_asj_fft_dataadgen_fft_120 (
	global_clock_enable,
	rd_addr_d_0,
	rd_addr_c_0,
	rd_addr_d_1,
	rd_addr_b_1,
	rd_addr_d_2,
	rd_addr_c_2,
	rd_addr_d_3,
	rd_addr_b_3,
	rd_addr_d_4,
	rd_addr_c_4,
	rd_addr_d_5,
	rd_addr_b_5,
	rd_addr_d_6,
	tdl_arr_4_20,
	tdl_arr_6_20,
	tdl_arr_0_20,
	tdl_arr_2_20,
	tdl_arr_0_1,
	tdl_arr_2_1,
	tdl_arr_1_1,
	tdl_arr_1_20,
	tdl_arr_3_20,
	tdl_arr_5_20,
	clk)/* synthesis synthesis_greybox=1 */;
input 	global_clock_enable;
output 	rd_addr_d_0;
output 	rd_addr_c_0;
output 	rd_addr_d_1;
output 	rd_addr_b_1;
output 	rd_addr_d_2;
output 	rd_addr_c_2;
output 	rd_addr_d_3;
output 	rd_addr_b_3;
output 	rd_addr_d_4;
output 	rd_addr_c_4;
output 	rd_addr_d_5;
output 	rd_addr_b_5;
output 	rd_addr_d_6;
input 	tdl_arr_4_20;
input 	tdl_arr_6_20;
input 	tdl_arr_0_20;
input 	tdl_arr_2_20;
input 	tdl_arr_0_1;
input 	tdl_arr_2_1;
input 	tdl_arr_1_1;
input 	tdl_arr_1_20;
input 	tdl_arr_3_20;
input 	tdl_arr_5_20;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Mux7~0_combout ;
wire \Mux7~1_combout ;
wire \Mux10~0_combout ;
wire \Mux7~2_combout ;
wire \Mux13~0_combout ;
wire \Mux6~0_combout ;
wire \Mux5~0_combout ;
wire \Mux9~0_combout ;
wire \Mux5~1_combout ;
wire \Mux12~0_combout ;
wire \Mux4~0_combout ;
wire \Mux8~0_combout ;
wire \Mux3~0_combout ;
wire \Mux11~0_combout ;
wire \Mux2~0_combout ;


dffeas \rd_addr_d[0] (
	.clk(clk),
	.d(\Mux10~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_d_0),
	.prn(vcc));
defparam \rd_addr_d[0] .is_wysiwyg = "true";
defparam \rd_addr_d[0] .power_up = "low";

dffeas \rd_addr_c[0] (
	.clk(clk),
	.d(\Mux7~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_c_0),
	.prn(vcc));
defparam \rd_addr_c[0] .is_wysiwyg = "true";
defparam \rd_addr_c[0] .power_up = "low";

dffeas \rd_addr_d[1] (
	.clk(clk),
	.d(\Mux13~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_d_1),
	.prn(vcc));
defparam \rd_addr_d[1] .is_wysiwyg = "true";
defparam \rd_addr_d[1] .power_up = "low";

dffeas \rd_addr_b[1] (
	.clk(clk),
	.d(\Mux6~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_b_1),
	.prn(vcc));
defparam \rd_addr_b[1] .is_wysiwyg = "true";
defparam \rd_addr_b[1] .power_up = "low";

dffeas \rd_addr_d[2] (
	.clk(clk),
	.d(\Mux9~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_d_2),
	.prn(vcc));
defparam \rd_addr_d[2] .is_wysiwyg = "true";
defparam \rd_addr_d[2] .power_up = "low";

dffeas \rd_addr_c[2] (
	.clk(clk),
	.d(\Mux5~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_c_2),
	.prn(vcc));
defparam \rd_addr_c[2] .is_wysiwyg = "true";
defparam \rd_addr_c[2] .power_up = "low";

dffeas \rd_addr_d[3] (
	.clk(clk),
	.d(\Mux12~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_d_3),
	.prn(vcc));
defparam \rd_addr_d[3] .is_wysiwyg = "true";
defparam \rd_addr_d[3] .power_up = "low";

dffeas \rd_addr_b[3] (
	.clk(clk),
	.d(\Mux4~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_b_3),
	.prn(vcc));
defparam \rd_addr_b[3] .is_wysiwyg = "true";
defparam \rd_addr_b[3] .power_up = "low";

dffeas \rd_addr_d[4] (
	.clk(clk),
	.d(\Mux8~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_d_4),
	.prn(vcc));
defparam \rd_addr_d[4] .is_wysiwyg = "true";
defparam \rd_addr_d[4] .power_up = "low";

dffeas \rd_addr_c[4] (
	.clk(clk),
	.d(\Mux3~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_c_4),
	.prn(vcc));
defparam \rd_addr_c[4] .is_wysiwyg = "true";
defparam \rd_addr_c[4] .power_up = "low";

dffeas \rd_addr_d[5] (
	.clk(clk),
	.d(\Mux11~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_d_5),
	.prn(vcc));
defparam \rd_addr_d[5] .is_wysiwyg = "true";
defparam \rd_addr_d[5] .power_up = "low";

dffeas \rd_addr_b[5] (
	.clk(clk),
	.d(\Mux2~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_b_5),
	.prn(vcc));
defparam \rd_addr_b[5] .is_wysiwyg = "true";
defparam \rd_addr_b[5] .power_up = "low";

dffeas \rd_addr_d[6] (
	.clk(clk),
	.d(tdl_arr_6_20),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_d_6),
	.prn(vcc));
defparam \rd_addr_d[6] .is_wysiwyg = "true";
defparam \rd_addr_d[6] .power_up = "low";

cycloneiii_lcell_comb \Mux7~0 (
	.dataa(gnd),
	.datab(tdl_arr_1_1),
	.datac(tdl_arr_0_1),
	.datad(tdl_arr_2_1),
	.cin(gnd),
	.combout(\Mux7~0_combout ),
	.cout());
defparam \Mux7~0 .lut_mask = 16'h3FCF;
defparam \Mux7~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux7~1 (
	.dataa(tdl_arr_0_1),
	.datab(tdl_arr_2_1),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux7~1_combout ),
	.cout());
defparam \Mux7~1 .lut_mask = 16'hEEEE;
defparam \Mux7~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux10~0 (
	.dataa(tdl_arr_2_20),
	.datab(tdl_arr_0_20),
	.datac(\Mux7~0_combout ),
	.datad(\Mux7~1_combout ),
	.cin(gnd),
	.combout(\Mux10~0_combout ),
	.cout());
defparam \Mux10~0 .lut_mask = 16'hACFF;
defparam \Mux10~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux7~2 (
	.dataa(tdl_arr_2_20),
	.datab(\Mux7~1_combout ),
	.datac(tdl_arr_0_20),
	.datad(\Mux7~0_combout ),
	.cin(gnd),
	.combout(\Mux7~2_combout ),
	.cout());
defparam \Mux7~2 .lut_mask = 16'hFAFC;
defparam \Mux7~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux13~0 (
	.dataa(tdl_arr_3_20),
	.datab(tdl_arr_1_20),
	.datac(\Mux7~0_combout ),
	.datad(\Mux7~1_combout ),
	.cin(gnd),
	.combout(\Mux13~0_combout ),
	.cout());
defparam \Mux13~0 .lut_mask = 16'hACFF;
defparam \Mux13~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux6~0 (
	.dataa(tdl_arr_3_20),
	.datab(\Mux7~1_combout ),
	.datac(tdl_arr_1_20),
	.datad(\Mux7~0_combout ),
	.cin(gnd),
	.combout(\Mux6~0_combout ),
	.cout());
defparam \Mux6~0 .lut_mask = 16'hFAFC;
defparam \Mux6~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux5~0 (
	.dataa(tdl_arr_2_1),
	.datab(gnd),
	.datac(tdl_arr_0_1),
	.datad(tdl_arr_1_1),
	.cin(gnd),
	.combout(\Mux5~0_combout ),
	.cout());
defparam \Mux5~0 .lut_mask = 16'hA55A;
defparam \Mux5~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux9~0 (
	.dataa(tdl_arr_2_20),
	.datab(tdl_arr_4_20),
	.datac(tdl_arr_2_1),
	.datad(\Mux5~0_combout ),
	.cin(gnd),
	.combout(\Mux9~0_combout ),
	.cout());
defparam \Mux9~0 .lut_mask = 16'hAFCF;
defparam \Mux9~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux5~1 (
	.dataa(tdl_arr_2_20),
	.datab(tdl_arr_4_20),
	.datac(tdl_arr_2_1),
	.datad(\Mux5~0_combout ),
	.cin(gnd),
	.combout(\Mux5~1_combout ),
	.cout());
defparam \Mux5~1 .lut_mask = 16'hFAFC;
defparam \Mux5~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux12~0 (
	.dataa(tdl_arr_3_20),
	.datab(tdl_arr_5_20),
	.datac(tdl_arr_2_1),
	.datad(\Mux5~0_combout ),
	.cin(gnd),
	.combout(\Mux12~0_combout ),
	.cout());
defparam \Mux12~0 .lut_mask = 16'hAFCF;
defparam \Mux12~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux4~0 (
	.dataa(tdl_arr_3_20),
	.datab(tdl_arr_2_1),
	.datac(tdl_arr_5_20),
	.datad(\Mux5~0_combout ),
	.cin(gnd),
	.combout(\Mux4~0_combout ),
	.cout());
defparam \Mux4~0 .lut_mask = 16'hFAFC;
defparam \Mux4~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux8~0 (
	.dataa(tdl_arr_4_20),
	.datab(tdl_arr_2_1),
	.datac(tdl_arr_0_1),
	.datad(tdl_arr_1_1),
	.cin(gnd),
	.combout(\Mux8~0_combout ),
	.cout());
defparam \Mux8~0 .lut_mask = 16'hEFFF;
defparam \Mux8~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux3~0 (
	.dataa(tdl_arr_4_20),
	.datab(tdl_arr_0_1),
	.datac(tdl_arr_1_1),
	.datad(tdl_arr_2_1),
	.cin(gnd),
	.combout(\Mux3~0_combout ),
	.cout());
defparam \Mux3~0 .lut_mask = 16'hFEFF;
defparam \Mux3~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux11~0 (
	.dataa(tdl_arr_5_20),
	.datab(tdl_arr_2_1),
	.datac(tdl_arr_0_1),
	.datad(tdl_arr_1_1),
	.cin(gnd),
	.combout(\Mux11~0_combout ),
	.cout());
defparam \Mux11~0 .lut_mask = 16'hEFFF;
defparam \Mux11~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux2~0 (
	.dataa(tdl_arr_5_20),
	.datab(tdl_arr_0_1),
	.datac(tdl_arr_1_1),
	.datad(tdl_arr_2_1),
	.cin(gnd),
	.combout(\Mux2~0_combout ),
	.cout());
defparam \Mux2~0 .lut_mask = 16'hFEFF;
defparam \Mux2~0 .sum_lutc_input = "datac";

endmodule

module fft_asj_fft_dataadgen_fft_120_1 (
	global_clock_enable,
	p_2,
	p_0,
	p_1,
	Equal0,
	rd_addr_d_0,
	rd_addr_c_0,
	sw_0,
	rd_addr_b_1,
	rd_addr_d_1,
	sw_1,
	rd_addr_d_2,
	rd_addr_c_2,
	rd_addr_b_3,
	rd_addr_d_3,
	rd_addr_d_4,
	rd_addr_c_4,
	rd_addr_b_5,
	rd_addr_d_5,
	k_count_0,
	k_count_2,
	Mux7,
	Mux1,
	k_count_4,
	Mux11,
	k_count_1,
	k_count_3,
	k_count_5,
	k_count_6,
	clk)/* synthesis synthesis_greybox=1 */;
input 	global_clock_enable;
input 	p_2;
input 	p_0;
input 	p_1;
input 	Equal0;
output 	rd_addr_d_0;
output 	rd_addr_c_0;
output 	sw_0;
output 	rd_addr_b_1;
output 	rd_addr_d_1;
output 	sw_1;
output 	rd_addr_d_2;
output 	rd_addr_c_2;
output 	rd_addr_b_3;
output 	rd_addr_d_3;
output 	rd_addr_d_4;
output 	rd_addr_c_4;
output 	rd_addr_b_5;
output 	rd_addr_d_5;
input 	k_count_0;
input 	k_count_2;
output 	Mux7;
output 	Mux1;
input 	k_count_4;
output 	Mux11;
input 	k_count_1;
input 	k_count_3;
input 	k_count_5;
input 	k_count_6;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Mux7~0_combout ;
wire \Mux10~0_combout ;
wire \Mux7~2_combout ;
wire \Mux1~2_combout ;
wire \Mux1~3_combout ;
wire \Mux1~4_combout ;
wire \Mux1~5_combout ;
wire \Mux6~0_combout ;
wire \Mux6~1_combout ;
wire \Mux13~0_combout ;
wire \Mux0~0_combout ;
wire \Mux0~1_combout ;
wire \Mux0~2_combout ;
wire \Mux0~3_combout ;
wire \Mux0~4_combout ;
wire \Mux0~5_combout ;
wire \Mux5~0_combout ;
wire \Mux9~0_combout ;
wire \Mux5~1_combout ;
wire \Mux4~0_combout ;
wire \Mux4~1_combout ;
wire \Mux12~0_combout ;
wire \Mux8~0_combout ;
wire \Mux3~0_combout ;
wire \Mux2~0_combout ;
wire \Mux11~0_combout ;


dffeas \rd_addr_d[0] (
	.clk(clk),
	.d(\Mux10~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_d_0),
	.prn(vcc));
defparam \rd_addr_d[0] .is_wysiwyg = "true";
defparam \rd_addr_d[0] .power_up = "low";

dffeas \rd_addr_c[0] (
	.clk(clk),
	.d(\Mux7~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_c_0),
	.prn(vcc));
defparam \rd_addr_c[0] .is_wysiwyg = "true";
defparam \rd_addr_c[0] .power_up = "low";

dffeas \sw[0] (
	.clk(clk),
	.d(\Mux1~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(sw_0),
	.prn(vcc));
defparam \sw[0] .is_wysiwyg = "true";
defparam \sw[0] .power_up = "low";

dffeas \rd_addr_b[1] (
	.clk(clk),
	.d(\Mux6~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_b_1),
	.prn(vcc));
defparam \rd_addr_b[1] .is_wysiwyg = "true";
defparam \rd_addr_b[1] .power_up = "low";

dffeas \rd_addr_d[1] (
	.clk(clk),
	.d(\Mux13~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_d_1),
	.prn(vcc));
defparam \rd_addr_d[1] .is_wysiwyg = "true";
defparam \rd_addr_d[1] .power_up = "low";

dffeas \sw[1] (
	.clk(clk),
	.d(\Mux0~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(sw_1),
	.prn(vcc));
defparam \sw[1] .is_wysiwyg = "true";
defparam \sw[1] .power_up = "low";

dffeas \rd_addr_d[2] (
	.clk(clk),
	.d(\Mux9~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_d_2),
	.prn(vcc));
defparam \rd_addr_d[2] .is_wysiwyg = "true";
defparam \rd_addr_d[2] .power_up = "low";

dffeas \rd_addr_c[2] (
	.clk(clk),
	.d(\Mux5~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_c_2),
	.prn(vcc));
defparam \rd_addr_c[2] .is_wysiwyg = "true";
defparam \rd_addr_c[2] .power_up = "low";

dffeas \rd_addr_b[3] (
	.clk(clk),
	.d(\Mux4~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_b_3),
	.prn(vcc));
defparam \rd_addr_b[3] .is_wysiwyg = "true";
defparam \rd_addr_b[3] .power_up = "low";

dffeas \rd_addr_d[3] (
	.clk(clk),
	.d(\Mux12~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_d_3),
	.prn(vcc));
defparam \rd_addr_d[3] .is_wysiwyg = "true";
defparam \rd_addr_d[3] .power_up = "low";

dffeas \rd_addr_d[4] (
	.clk(clk),
	.d(\Mux8~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_d_4),
	.prn(vcc));
defparam \rd_addr_d[4] .is_wysiwyg = "true";
defparam \rd_addr_d[4] .power_up = "low";

dffeas \rd_addr_c[4] (
	.clk(clk),
	.d(\Mux3~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_c_4),
	.prn(vcc));
defparam \rd_addr_c[4] .is_wysiwyg = "true";
defparam \rd_addr_c[4] .power_up = "low";

dffeas \rd_addr_b[5] (
	.clk(clk),
	.d(\Mux2~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_b_5),
	.prn(vcc));
defparam \rd_addr_b[5] .is_wysiwyg = "true";
defparam \rd_addr_b[5] .power_up = "low";

dffeas \rd_addr_d[5] (
	.clk(clk),
	.d(\Mux11~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_d_5),
	.prn(vcc));
defparam \rd_addr_d[5] .is_wysiwyg = "true";
defparam \rd_addr_d[5] .power_up = "low";

cycloneiii_lcell_comb \Mux7~1 (
	.dataa(p_1),
	.datab(gnd),
	.datac(gnd),
	.datad(p_0),
	.cin(gnd),
	.combout(Mux7),
	.cout());
defparam \Mux7~1 .lut_mask = 16'hAAFF;
defparam \Mux7~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux1~0 (
	.dataa(k_count_0),
	.datab(gnd),
	.datac(gnd),
	.datad(p_2),
	.cin(gnd),
	.combout(Mux1),
	.cout());
defparam \Mux1~0 .lut_mask = 16'hAAFF;
defparam \Mux1~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux1~1 (
	.dataa(k_count_4),
	.datab(gnd),
	.datac(gnd),
	.datad(p_2),
	.cin(gnd),
	.combout(Mux11),
	.cout());
defparam \Mux1~1 .lut_mask = 16'hAAFF;
defparam \Mux1~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux7~0 (
	.dataa(gnd),
	.datab(p_1),
	.datac(p_0),
	.datad(p_2),
	.cin(gnd),
	.combout(\Mux7~0_combout ),
	.cout());
defparam \Mux7~0 .lut_mask = 16'h3FCF;
defparam \Mux7~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux10~0 (
	.dataa(k_count_0),
	.datab(\Mux7~0_combout ),
	.datac(k_count_2),
	.datad(Mux7),
	.cin(gnd),
	.combout(\Mux10~0_combout ),
	.cout());
defparam \Mux10~0 .lut_mask = 16'hFFB8;
defparam \Mux10~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux7~2 (
	.dataa(k_count_0),
	.datab(k_count_2),
	.datac(\Mux7~0_combout ),
	.datad(Mux7),
	.cin(gnd),
	.combout(\Mux7~2_combout ),
	.cout());
defparam \Mux7~2 .lut_mask = 16'hACFF;
defparam \Mux7~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux1~2 (
	.dataa(p_2),
	.datab(k_count_0),
	.datac(k_count_2),
	.datad(k_count_4),
	.cin(gnd),
	.combout(\Mux1~2_combout ),
	.cout());
defparam \Mux1~2 .lut_mask = 16'hEBBE;
defparam \Mux1~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux1~3 (
	.dataa(p_1),
	.datab(Mux11),
	.datac(p_0),
	.datad(\Mux1~2_combout ),
	.cin(gnd),
	.combout(\Mux1~3_combout ),
	.cout());
defparam \Mux1~3 .lut_mask = 16'hFFDE;
defparam \Mux1~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux1~4 (
	.dataa(gnd),
	.datab(k_count_0),
	.datac(k_count_2),
	.datad(p_2),
	.cin(gnd),
	.combout(\Mux1~4_combout ),
	.cout());
defparam \Mux1~4 .lut_mask = 16'h3CFF;
defparam \Mux1~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux1~5 (
	.dataa(Mux1),
	.datab(p_1),
	.datac(\Mux1~3_combout ),
	.datad(\Mux1~4_combout ),
	.cin(gnd),
	.combout(\Mux1~5_combout ),
	.cout());
defparam \Mux1~5 .lut_mask = 16'hFFBE;
defparam \Mux1~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux6~0 (
	.dataa(p_2),
	.datab(p_0),
	.datac(gnd),
	.datad(p_1),
	.cin(gnd),
	.combout(\Mux6~0_combout ),
	.cout());
defparam \Mux6~0 .lut_mask = 16'hDDEE;
defparam \Mux6~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux6~1 (
	.dataa(k_count_1),
	.datab(\Mux6~0_combout ),
	.datac(k_count_3),
	.datad(Mux7),
	.cin(gnd),
	.combout(\Mux6~1_combout ),
	.cout());
defparam \Mux6~1 .lut_mask = 16'hB8FF;
defparam \Mux6~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux13~0 (
	.dataa(k_count_1),
	.datab(Mux7),
	.datac(k_count_3),
	.datad(\Mux6~0_combout ),
	.cin(gnd),
	.combout(\Mux13~0_combout ),
	.cout());
defparam \Mux13~0 .lut_mask = 16'hFAFC;
defparam \Mux13~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux0~0 (
	.dataa(k_count_0),
	.datab(k_count_2),
	.datac(k_count_3),
	.datad(k_count_4),
	.cin(gnd),
	.combout(\Mux0~0_combout ),
	.cout());
defparam \Mux0~0 .lut_mask = 16'h6996;
defparam \Mux0~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux0~1 (
	.dataa(k_count_1),
	.datab(k_count_5),
	.datac(Equal0),
	.datad(\Mux0~0_combout ),
	.cin(gnd),
	.combout(\Mux0~1_combout ),
	.cout());
defparam \Mux0~1 .lut_mask = 16'hF9F6;
defparam \Mux0~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux0~2 (
	.dataa(p_1),
	.datab(k_count_5),
	.datac(k_count_6),
	.datad(p_2),
	.cin(gnd),
	.combout(\Mux0~2_combout ),
	.cout());
defparam \Mux0~2 .lut_mask = 16'h6996;
defparam \Mux0~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux0~3 (
	.dataa(k_count_0),
	.datab(k_count_2),
	.datac(k_count_3),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux0~3_combout ),
	.cout());
defparam \Mux0~3 .lut_mask = 16'h9696;
defparam \Mux0~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux0~4 (
	.dataa(k_count_1),
	.datab(p_0),
	.datac(\Mux0~3_combout ),
	.datad(\Mux0~2_combout ),
	.cin(gnd),
	.combout(\Mux0~4_combout ),
	.cout());
defparam \Mux0~4 .lut_mask = 16'h6996;
defparam \Mux0~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux0~5 (
	.dataa(\Mux0~1_combout ),
	.datab(p_1),
	.datac(\Mux0~2_combout ),
	.datad(\Mux0~4_combout ),
	.cin(gnd),
	.combout(\Mux0~5_combout ),
	.cout());
defparam \Mux0~5 .lut_mask = 16'hFFBE;
defparam \Mux0~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux5~0 (
	.dataa(p_2),
	.datab(gnd),
	.datac(p_0),
	.datad(p_1),
	.cin(gnd),
	.combout(\Mux5~0_combout ),
	.cout());
defparam \Mux5~0 .lut_mask = 16'hA55A;
defparam \Mux5~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux9~0 (
	.dataa(k_count_2),
	.datab(p_0),
	.datac(k_count_4),
	.datad(\Mux5~0_combout ),
	.cin(gnd),
	.combout(\Mux9~0_combout ),
	.cout());
defparam \Mux9~0 .lut_mask = 16'hFAFC;
defparam \Mux9~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux5~1 (
	.dataa(k_count_2),
	.datab(\Mux5~0_combout ),
	.datac(k_count_4),
	.datad(p_0),
	.cin(gnd),
	.combout(\Mux5~1_combout ),
	.cout());
defparam \Mux5~1 .lut_mask = 16'hB8FF;
defparam \Mux5~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux4~0 (
	.dataa(gnd),
	.datab(p_0),
	.datac(p_1),
	.datad(p_2),
	.cin(gnd),
	.combout(\Mux4~0_combout ),
	.cout());
defparam \Mux4~0 .lut_mask = 16'hC33C;
defparam \Mux4~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux4~1 (
	.dataa(k_count_3),
	.datab(k_count_5),
	.datac(\Mux4~0_combout ),
	.datad(p_1),
	.cin(gnd),
	.combout(\Mux4~1_combout ),
	.cout());
defparam \Mux4~1 .lut_mask = 16'hACFF;
defparam \Mux4~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux12~0 (
	.dataa(k_count_3),
	.datab(\Mux4~0_combout ),
	.datac(p_1),
	.datad(k_count_5),
	.cin(gnd),
	.combout(\Mux12~0_combout ),
	.cout());
defparam \Mux12~0 .lut_mask = 16'hFFB8;
defparam \Mux12~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux8~0 (
	.dataa(k_count_4),
	.datab(p_2),
	.datac(p_0),
	.datad(p_1),
	.cin(gnd),
	.combout(\Mux8~0_combout ),
	.cout());
defparam \Mux8~0 .lut_mask = 16'hEFFF;
defparam \Mux8~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux3~0 (
	.dataa(k_count_4),
	.datab(p_0),
	.datac(p_1),
	.datad(p_2),
	.cin(gnd),
	.combout(\Mux3~0_combout ),
	.cout());
defparam \Mux3~0 .lut_mask = 16'hFEFF;
defparam \Mux3~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux2~0 (
	.dataa(k_count_5),
	.datab(p_0),
	.datac(p_1),
	.datad(p_2),
	.cin(gnd),
	.combout(\Mux2~0_combout ),
	.cout());
defparam \Mux2~0 .lut_mask = 16'hFEFF;
defparam \Mux2~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux11~0 (
	.dataa(k_count_5),
	.datab(p_2),
	.datac(p_0),
	.datad(p_1),
	.cin(gnd),
	.combout(\Mux11~0_combout ),
	.cout());
defparam \Mux11~0 .lut_mask = 16'hEFFF;
defparam \Mux11~0 .sum_lutc_input = "datac";

endmodule

module fft_asj_fft_dft_bfp_fft_120 (
	r_array_out_3_0,
	i_array_out_3_0,
	r_array_out_3_1,
	i_array_out_3_1,
	r_array_out_3_2,
	i_array_out_3_2,
	r_array_out_3_3,
	i_array_out_3_3,
	r_array_out_4_0,
	i_array_out_4_0,
	r_array_out_4_1,
	i_array_out_4_1,
	r_array_out_4_2,
	i_array_out_4_2,
	r_array_out_4_3,
	i_array_out_4_3,
	r_array_out_5_0,
	i_array_out_5_0,
	r_array_out_5_1,
	i_array_out_5_1,
	r_array_out_5_2,
	i_array_out_5_2,
	r_array_out_5_3,
	i_array_out_5_3,
	i_array_out_2_2,
	i_array_out_2_1,
	i_array_out_2_0,
	i_array_out_2_3,
	r_array_out_2_2,
	r_array_out_2_1,
	r_array_out_2_0,
	r_array_out_2_3,
	ram_in_reg_2_0,
	ram_in_reg_6_0,
	ram_in_reg_4_0,
	ram_in_reg_3_0,
	ram_in_reg_5_0,
	ram_in_reg_2_2,
	ram_in_reg_6_2,
	ram_in_reg_4_2,
	ram_in_reg_3_2,
	ram_in_reg_5_2,
	ram_in_reg_1_0,
	ram_in_reg_1_2,
	ram_in_reg_0_0,
	ram_in_reg_0_2,
	ram_in_reg_2_1,
	ram_in_reg_6_1,
	ram_in_reg_4_1,
	ram_in_reg_3_1,
	ram_in_reg_5_1,
	ram_in_reg_2_3,
	ram_in_reg_6_3,
	ram_in_reg_4_3,
	ram_in_reg_3_3,
	ram_in_reg_5_3,
	ram_in_reg_1_1,
	ram_in_reg_1_3,
	ram_in_reg_0_1,
	ram_in_reg_0_3,
	ram_in_reg_7_0,
	ram_in_reg_7_2,
	ram_in_reg_7_1,
	ram_in_reg_7_3,
	ram_in_reg_7_4,
	ram_in_reg_3_4,
	ram_in_reg_5_4,
	ram_in_reg_4_4,
	ram_in_reg_6_4,
	ram_in_reg_7_6,
	ram_in_reg_3_6,
	ram_in_reg_5_6,
	ram_in_reg_4_6,
	ram_in_reg_6_6,
	ram_in_reg_2_4,
	ram_in_reg_2_6,
	ram_in_reg_1_4,
	ram_in_reg_1_6,
	ram_in_reg_0_4,
	ram_in_reg_0_6,
	ram_in_reg_7_5,
	ram_in_reg_3_5,
	ram_in_reg_5_5,
	ram_in_reg_4_5,
	ram_in_reg_6_5,
	ram_in_reg_3_7,
	ram_in_reg_7_7,
	ram_in_reg_5_7,
	ram_in_reg_4_7,
	ram_in_reg_6_7,
	ram_in_reg_2_5,
	ram_in_reg_2_7,
	ram_in_reg_1_5,
	ram_in_reg_1_7,
	ram_in_reg_0_5,
	ram_in_reg_0_7,
	global_clock_enable,
	slb_last_0,
	slb_last_1,
	slb_last_2,
	next_block,
	slb_i_0,
	slb_i_1,
	slb_i_2,
	slb_i_3,
	Mux2,
	Mux1,
	tdl_arr_4,
	tdl_arr_3,
	r_array_out_7_0,
	i_array_out_7_0,
	r_array_out_7_1,
	i_array_out_7_1,
	r_array_out_7_2,
	i_array_out_7_2,
	r_array_out_7_3,
	i_array_out_7_3,
	blk_done_vec_2,
	r_array_out_6_0,
	i_array_out_6_0,
	r_array_out_6_1,
	i_array_out_6_1,
	r_array_out_6_2,
	i_array_out_6_2,
	r_array_out_6_3,
	i_array_out_6_3,
	i_array_out_1_2,
	i_array_out_1_1,
	i_array_out_1_0,
	i_array_out_1_3,
	i_array_out_0_2,
	i_array_out_0_1,
	i_array_out_0_0,
	i_array_out_0_3,
	r_array_out_1_2,
	r_array_out_1_1,
	r_array_out_1_0,
	r_array_out_1_3,
	r_array_out_0_2,
	r_array_out_0_1,
	r_array_out_0_0,
	r_array_out_0_3,
	tdl_arr_5,
	tdl_arr_51,
	twiddle_data000,
	twiddle_data001,
	twiddle_data002,
	twiddle_data003,
	twiddle_data004,
	twiddle_data005,
	twiddle_data006,
	twiddle_data007,
	twiddle_data010,
	twiddle_data011,
	twiddle_data012,
	twiddle_data013,
	twiddle_data014,
	twiddle_data015,
	twiddle_data016,
	twiddle_data017,
	twiddle_data100,
	twiddle_data101,
	twiddle_data102,
	twiddle_data103,
	twiddle_data104,
	twiddle_data105,
	twiddle_data106,
	twiddle_data107,
	twiddle_data110,
	twiddle_data111,
	twiddle_data112,
	twiddle_data113,
	twiddle_data114,
	twiddle_data115,
	twiddle_data116,
	twiddle_data117,
	twiddle_data200,
	twiddle_data201,
	twiddle_data202,
	twiddle_data203,
	twiddle_data204,
	twiddle_data205,
	twiddle_data206,
	twiddle_data207,
	twiddle_data210,
	twiddle_data211,
	twiddle_data212,
	twiddle_data213,
	twiddle_data214,
	twiddle_data215,
	twiddle_data216,
	twiddle_data217,
	next_pass_vec_2,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	r_array_out_3_0;
output 	i_array_out_3_0;
output 	r_array_out_3_1;
output 	i_array_out_3_1;
output 	r_array_out_3_2;
output 	i_array_out_3_2;
output 	r_array_out_3_3;
output 	i_array_out_3_3;
output 	r_array_out_4_0;
output 	i_array_out_4_0;
output 	r_array_out_4_1;
output 	i_array_out_4_1;
output 	r_array_out_4_2;
output 	i_array_out_4_2;
output 	r_array_out_4_3;
output 	i_array_out_4_3;
output 	r_array_out_5_0;
output 	i_array_out_5_0;
output 	r_array_out_5_1;
output 	i_array_out_5_1;
output 	r_array_out_5_2;
output 	i_array_out_5_2;
output 	r_array_out_5_3;
output 	i_array_out_5_3;
output 	i_array_out_2_2;
output 	i_array_out_2_1;
output 	i_array_out_2_0;
output 	i_array_out_2_3;
output 	r_array_out_2_2;
output 	r_array_out_2_1;
output 	r_array_out_2_0;
output 	r_array_out_2_3;
input 	ram_in_reg_2_0;
input 	ram_in_reg_6_0;
input 	ram_in_reg_4_0;
input 	ram_in_reg_3_0;
input 	ram_in_reg_5_0;
input 	ram_in_reg_2_2;
input 	ram_in_reg_6_2;
input 	ram_in_reg_4_2;
input 	ram_in_reg_3_2;
input 	ram_in_reg_5_2;
input 	ram_in_reg_1_0;
input 	ram_in_reg_1_2;
input 	ram_in_reg_0_0;
input 	ram_in_reg_0_2;
input 	ram_in_reg_2_1;
input 	ram_in_reg_6_1;
input 	ram_in_reg_4_1;
input 	ram_in_reg_3_1;
input 	ram_in_reg_5_1;
input 	ram_in_reg_2_3;
input 	ram_in_reg_6_3;
input 	ram_in_reg_4_3;
input 	ram_in_reg_3_3;
input 	ram_in_reg_5_3;
input 	ram_in_reg_1_1;
input 	ram_in_reg_1_3;
input 	ram_in_reg_0_1;
input 	ram_in_reg_0_3;
input 	ram_in_reg_7_0;
input 	ram_in_reg_7_2;
input 	ram_in_reg_7_1;
input 	ram_in_reg_7_3;
input 	ram_in_reg_7_4;
input 	ram_in_reg_3_4;
input 	ram_in_reg_5_4;
input 	ram_in_reg_4_4;
input 	ram_in_reg_6_4;
input 	ram_in_reg_7_6;
input 	ram_in_reg_3_6;
input 	ram_in_reg_5_6;
input 	ram_in_reg_4_6;
input 	ram_in_reg_6_6;
input 	ram_in_reg_2_4;
input 	ram_in_reg_2_6;
input 	ram_in_reg_1_4;
input 	ram_in_reg_1_6;
input 	ram_in_reg_0_4;
input 	ram_in_reg_0_6;
input 	ram_in_reg_7_5;
input 	ram_in_reg_3_5;
input 	ram_in_reg_5_5;
input 	ram_in_reg_4_5;
input 	ram_in_reg_6_5;
input 	ram_in_reg_3_7;
input 	ram_in_reg_7_7;
input 	ram_in_reg_5_7;
input 	ram_in_reg_4_7;
input 	ram_in_reg_6_7;
input 	ram_in_reg_2_5;
input 	ram_in_reg_2_7;
input 	ram_in_reg_1_5;
input 	ram_in_reg_1_7;
input 	ram_in_reg_0_5;
input 	ram_in_reg_0_7;
input 	global_clock_enable;
input 	slb_last_0;
input 	slb_last_1;
input 	slb_last_2;
input 	next_block;
output 	slb_i_0;
output 	slb_i_1;
output 	slb_i_2;
output 	slb_i_3;
output 	Mux2;
output 	Mux1;
output 	tdl_arr_4;
output 	tdl_arr_3;
output 	r_array_out_7_0;
output 	i_array_out_7_0;
output 	r_array_out_7_1;
output 	i_array_out_7_1;
output 	r_array_out_7_2;
output 	i_array_out_7_2;
output 	r_array_out_7_3;
output 	i_array_out_7_3;
output 	blk_done_vec_2;
output 	r_array_out_6_0;
output 	i_array_out_6_0;
output 	r_array_out_6_1;
output 	i_array_out_6_1;
output 	r_array_out_6_2;
output 	i_array_out_6_2;
output 	r_array_out_6_3;
output 	i_array_out_6_3;
output 	i_array_out_1_2;
output 	i_array_out_1_1;
output 	i_array_out_1_0;
output 	i_array_out_1_3;
output 	i_array_out_0_2;
output 	i_array_out_0_1;
output 	i_array_out_0_0;
output 	i_array_out_0_3;
output 	r_array_out_1_2;
output 	r_array_out_1_1;
output 	r_array_out_1_0;
output 	r_array_out_1_3;
output 	r_array_out_0_2;
output 	r_array_out_0_1;
output 	r_array_out_0_0;
output 	r_array_out_0_3;
input 	tdl_arr_5;
input 	tdl_arr_51;
input 	twiddle_data000;
input 	twiddle_data001;
input 	twiddle_data002;
input 	twiddle_data003;
input 	twiddle_data004;
input 	twiddle_data005;
input 	twiddle_data006;
input 	twiddle_data007;
input 	twiddle_data010;
input 	twiddle_data011;
input 	twiddle_data012;
input 	twiddle_data013;
input 	twiddle_data014;
input 	twiddle_data015;
input 	twiddle_data016;
input 	twiddle_data017;
input 	twiddle_data100;
input 	twiddle_data101;
input 	twiddle_data102;
input 	twiddle_data103;
input 	twiddle_data104;
input 	twiddle_data105;
input 	twiddle_data106;
input 	twiddle_data107;
input 	twiddle_data110;
input 	twiddle_data111;
input 	twiddle_data112;
input 	twiddle_data113;
input 	twiddle_data114;
input 	twiddle_data115;
input 	twiddle_data116;
input 	twiddle_data117;
input 	twiddle_data200;
input 	twiddle_data201;
input 	twiddle_data202;
input 	twiddle_data203;
input 	twiddle_data204;
input 	twiddle_data205;
input 	twiddle_data206;
input 	twiddle_data207;
input 	twiddle_data210;
input 	twiddle_data211;
input 	twiddle_data212;
input 	twiddle_data213;
input 	twiddle_data214;
input 	twiddle_data215;
input 	twiddle_data216;
input 	twiddle_data217;
output 	next_pass_vec_2;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \gain_out_4pts[0]~q ;
wire \gain_out_4pts[1]~q ;
wire \gain_out_4pts[2]~q ;
wire \gain_out_4pts[3]~q ;
wire \gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ;
wire \gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ;
wire \gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ;
wire \gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ;
wire \gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ;
wire \gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ;
wire \sdft.ENABLE_DFT_O~q ;
wire \gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ;
wire \gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ;
wire \gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ;
wire \gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ;
wire \gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ;
wire \gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ;
wire \gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ;
wire \gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ;
wire \gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ;
wire \gap_reg~q ;
wire \state_cnt[2]~q ;
wire \state_cnt[3]~q ;
wire \state_cnt[4]~q ;
wire \state_cnt[5]~q ;
wire \state_cnt[0]~q ;
wire \state_cnt[1]~q ;
wire \sdft.BLOCK_DFT_I~q ;
wire \sdft.ENABLE_BFP_O~q ;
wire \state_cnt[0]~7 ;
wire \state_cnt[0]~6_combout ;
wire \state_cnt[1]~9 ;
wire \state_cnt[1]~8_combout ;
wire \state_cnt[2]~11 ;
wire \state_cnt[2]~10_combout ;
wire \state_cnt[3]~15 ;
wire \state_cnt[3]~14_combout ;
wire \state_cnt[4]~17 ;
wire \state_cnt[4]~16_combout ;
wire \state_cnt[5]~18_combout ;
wire \reg_no_twiddle[0][0][3]~q ;
wire \reg_no_twiddle[0][0][7]~q ;
wire \reg_no_twiddle[0][1][7]~q ;
wire \reg_no_twiddle[0][1][3]~q ;
wire \gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ;
wire \gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ;
wire \gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ;
wire \gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ;
wire \gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ;
wire \gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ;
wire \gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ;
wire \gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ;
wire \gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ;
wire \reg_no_twiddle[0][0][4]~q ;
wire \reg_no_twiddle[0][1][4]~q ;
wire \reg_no_twiddle[0][0][5]~q ;
wire \reg_no_twiddle[0][1][5]~q ;
wire \reg_no_twiddle[0][0][6]~q ;
wire \reg_no_twiddle[0][1][6]~q ;
wire \gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ;
wire \gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ;
wire \gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ;
wire \gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ;
wire \gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ;
wire \gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ;
wire \reg_no_twiddle[0][0][0]~2 ;
wire \reg_no_twiddle[0][0][0]~1_combout ;
wire \reg_no_twiddle[0][0][1]~2 ;
wire \reg_no_twiddle[0][0][1]~1_combout ;
wire \reg_no_twiddle[0][0][2]~2 ;
wire \reg_no_twiddle[0][0][2]~1_combout ;
wire \reg_no_twiddle[0][0][3]~2 ;
wire \reg_no_twiddle[0][0][3]~1_combout ;
wire \gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ;
wire \gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ;
wire \reg_no_twiddle[0][0][4]~2 ;
wire \reg_no_twiddle[0][0][4]~1_combout ;
wire \reg_no_twiddle[0][0][5]~2 ;
wire \reg_no_twiddle[0][0][5]~1_combout ;
wire \reg_no_twiddle[0][0][6]~2 ;
wire \reg_no_twiddle[0][0][6]~1_combout ;
wire \reg_no_twiddle[0][0][7]~1_combout ;
wire \gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ;
wire \gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ;
wire \gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ;
wire \gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ;
wire \gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ;
wire \gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ;
wire \gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ;
wire \gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ;
wire \reg_no_twiddle[0][1][0]~2 ;
wire \reg_no_twiddle[0][1][0]~1_combout ;
wire \reg_no_twiddle[0][1][1]~2 ;
wire \reg_no_twiddle[0][1][1]~1_combout ;
wire \reg_no_twiddle[0][1][2]~2 ;
wire \reg_no_twiddle[0][1][2]~1_combout ;
wire \reg_no_twiddle[0][1][3]~2 ;
wire \reg_no_twiddle[0][1][3]~1_combout ;
wire \reg_no_twiddle[0][1][4]~2 ;
wire \reg_no_twiddle[0][1][4]~1_combout ;
wire \reg_no_twiddle[0][1][5]~2 ;
wire \reg_no_twiddle[0][1][5]~1_combout ;
wire \reg_no_twiddle[0][1][6]~2 ;
wire \reg_no_twiddle[0][1][6]~1_combout ;
wire \reg_no_twiddle[0][1][7]~1_combout ;
wire \gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ;
wire \gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ;
wire \gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ;
wire \gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ;
wire \gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ;
wire \gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ;
wire \gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ;
wire \gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ;
wire \gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ;
wire \gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ;
wire \gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ;
wire \gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ;
wire \gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ;
wire \gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ;
wire \gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ;
wire \gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ;
wire \gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ;
wire \gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ;
wire \gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ;
wire \gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ;
wire \gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ;
wire \gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ;
wire \gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ;
wire \gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ;
wire \gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ;
wire \gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ;
wire \gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ;
wire \gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ;
wire \gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ;
wire \gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ;
wire \gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ;
wire \gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ;
wire \gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ;
wire \gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ;
wire \gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ;
wire \gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ;
wire \gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ;
wire \gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ;
wire \gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ;
wire \gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ;
wire \gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ;
wire \gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ;
wire \gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ;
wire \gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ;
wire \gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ;
wire \gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ;
wire \gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ;
wire \gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ;
wire \butterfly_st2[0][0][6]~q ;
wire \butterfly_st2[0][0][5]~q ;
wire \butterfly_st2[0][0][4]~q ;
wire \butterfly_st2[0][0][3]~q ;
wire \butterfly_st2[0][0][2]~q ;
wire \butterfly_st2[0][0][1]~q ;
wire \butterfly_st2[0][0][0]~q ;
wire \butterfly_st2[0][0][9]~q ;
wire \butterfly_st2[0][0][8]~q ;
wire \butterfly_st2[0][0][7]~q ;
wire \butterfly_st2[0][1][9]~q ;
wire \butterfly_st2[0][1][8]~q ;
wire \butterfly_st2[0][1][7]~q ;
wire \butterfly_st2[0][1][6]~q ;
wire \butterfly_st2[0][1][5]~q ;
wire \butterfly_st2[0][1][4]~q ;
wire \butterfly_st2[0][1][3]~q ;
wire \butterfly_st2[0][1][2]~q ;
wire \butterfly_st2[0][1][1]~q ;
wire \butterfly_st2[0][1][0]~q ;
wire \butterfly_st2[1][1][2]~q ;
wire \butterfly_st2[1][1][1]~q ;
wire \butterfly_st2[1][1][0]~q ;
wire \butterfly_st2[1][1][9]~q ;
wire \butterfly_st2[1][1][3]~q ;
wire \butterfly_st2[1][1][4]~q ;
wire \butterfly_st2[1][1][5]~q ;
wire \butterfly_st2[1][1][6]~q ;
wire \butterfly_st2[1][1][7]~q ;
wire \butterfly_st2[1][1][8]~q ;
wire \butterfly_st2[1][0][2]~q ;
wire \butterfly_st2[1][0][1]~q ;
wire \butterfly_st2[1][0][0]~q ;
wire \butterfly_st2[1][0][9]~q ;
wire \butterfly_st2[1][0][3]~q ;
wire \butterfly_st2[1][0][4]~q ;
wire \butterfly_st2[1][0][5]~q ;
wire \butterfly_st2[1][0][6]~q ;
wire \butterfly_st2[1][0][7]~q ;
wire \butterfly_st2[1][0][8]~q ;
wire \butterfly_st2[2][1][2]~q ;
wire \butterfly_st2[2][1][1]~q ;
wire \butterfly_st2[2][1][0]~q ;
wire \butterfly_st2[2][1][9]~q ;
wire \butterfly_st2[2][1][3]~q ;
wire \butterfly_st2[2][1][4]~q ;
wire \butterfly_st2[2][1][5]~q ;
wire \butterfly_st2[2][1][6]~q ;
wire \butterfly_st2[2][1][7]~q ;
wire \butterfly_st2[2][1][8]~q ;
wire \butterfly_st2[2][0][2]~q ;
wire \butterfly_st2[2][0][1]~q ;
wire \butterfly_st2[2][0][0]~q ;
wire \butterfly_st2[2][0][9]~q ;
wire \butterfly_st2[2][0][3]~q ;
wire \butterfly_st2[2][0][4]~q ;
wire \butterfly_st2[2][0][5]~q ;
wire \butterfly_st2[2][0][6]~q ;
wire \butterfly_st2[2][0][7]~q ;
wire \butterfly_st2[2][0][8]~q ;
wire \butterfly_st2[3][1][2]~q ;
wire \butterfly_st2[3][1][1]~q ;
wire \butterfly_st2[3][1][0]~q ;
wire \butterfly_st2[3][1][9]~q ;
wire \butterfly_st2[3][1][3]~q ;
wire \butterfly_st2[3][1][4]~q ;
wire \butterfly_st2[3][1][5]~q ;
wire \butterfly_st2[3][1][6]~q ;
wire \butterfly_st2[3][1][7]~q ;
wire \butterfly_st2[3][1][8]~q ;
wire \butterfly_st2[3][0][2]~q ;
wire \butterfly_st2[3][0][1]~q ;
wire \butterfly_st2[3][0][0]~q ;
wire \butterfly_st2[3][0][9]~q ;
wire \butterfly_st2[3][0][3]~q ;
wire \butterfly_st2[3][0][4]~q ;
wire \butterfly_st2[3][0][5]~q ;
wire \butterfly_st2[3][0][6]~q ;
wire \butterfly_st2[3][0][7]~q ;
wire \butterfly_st2[3][0][8]~q ;
wire \butterfly_st1[0][0][6]~q ;
wire \butterfly_st1[1][0][6]~q ;
wire \butterfly_st1[0][0][5]~q ;
wire \butterfly_st1[1][0][5]~q ;
wire \butterfly_st1[0][0][4]~q ;
wire \butterfly_st1[1][0][4]~q ;
wire \butterfly_st1[0][0][3]~q ;
wire \butterfly_st1[1][0][3]~q ;
wire \butterfly_st1[0][0][2]~q ;
wire \butterfly_st1[1][0][2]~q ;
wire \butterfly_st1[0][0][1]~q ;
wire \butterfly_st1[1][0][1]~q ;
wire \butterfly_st1[0][0][0]~q ;
wire \butterfly_st1[1][0][0]~q ;
wire \butterfly_st2[0][0][0]~2 ;
wire \butterfly_st2[0][0][0]~1_combout ;
wire \butterfly_st2[0][0][1]~2 ;
wire \butterfly_st2[0][0][1]~1_combout ;
wire \butterfly_st2[0][0][2]~2 ;
wire \butterfly_st2[0][0][2]~1_combout ;
wire \butterfly_st2[0][0][3]~2 ;
wire \butterfly_st2[0][0][3]~1_combout ;
wire \butterfly_st2[0][0][4]~2 ;
wire \butterfly_st2[0][0][4]~1_combout ;
wire \butterfly_st2[0][0][5]~2 ;
wire \butterfly_st2[0][0][5]~1_combout ;
wire \butterfly_st2[0][0][6]~2 ;
wire \butterfly_st2[0][0][6]~1_combout ;
wire \butterfly_st1[0][0][8]~q ;
wire \butterfly_st1[1][0][8]~q ;
wire \butterfly_st1[0][0][7]~q ;
wire \butterfly_st1[1][0][7]~q ;
wire \butterfly_st2[0][0][7]~2 ;
wire \butterfly_st2[0][0][7]~1_combout ;
wire \butterfly_st2[0][0][8]~2 ;
wire \butterfly_st2[0][0][8]~1_combout ;
wire \butterfly_st2[0][0][9]~1_combout ;
wire \butterfly_st1[0][1][8]~q ;
wire \butterfly_st1[1][1][8]~q ;
wire \butterfly_st1[0][1][7]~q ;
wire \butterfly_st1[1][1][7]~q ;
wire \butterfly_st1[0][1][6]~q ;
wire \butterfly_st1[1][1][6]~q ;
wire \butterfly_st1[0][1][5]~q ;
wire \butterfly_st1[1][1][5]~q ;
wire \butterfly_st1[0][1][4]~q ;
wire \butterfly_st1[1][1][4]~q ;
wire \butterfly_st1[0][1][3]~q ;
wire \butterfly_st1[1][1][3]~q ;
wire \butterfly_st1[0][1][2]~q ;
wire \butterfly_st1[1][1][2]~q ;
wire \butterfly_st1[0][1][1]~q ;
wire \butterfly_st1[1][1][1]~q ;
wire \butterfly_st1[0][1][0]~q ;
wire \butterfly_st1[1][1][0]~q ;
wire \butterfly_st2[0][1][0]~2 ;
wire \butterfly_st2[0][1][0]~1_combout ;
wire \butterfly_st2[0][1][1]~2 ;
wire \butterfly_st2[0][1][1]~1_combout ;
wire \butterfly_st2[0][1][2]~2 ;
wire \butterfly_st2[0][1][2]~1_combout ;
wire \butterfly_st2[0][1][3]~2 ;
wire \butterfly_st2[0][1][3]~1_combout ;
wire \butterfly_st2[0][1][4]~2 ;
wire \butterfly_st2[0][1][4]~1_combout ;
wire \butterfly_st2[0][1][5]~2 ;
wire \butterfly_st2[0][1][5]~1_combout ;
wire \butterfly_st2[0][1][6]~2 ;
wire \butterfly_st2[0][1][6]~1_combout ;
wire \butterfly_st2[0][1][7]~2 ;
wire \butterfly_st2[0][1][7]~1_combout ;
wire \butterfly_st2[0][1][8]~2 ;
wire \butterfly_st2[0][1][8]~1_combout ;
wire \butterfly_st2[0][1][9]~1_combout ;
wire \butterfly_st1[2][1][2]~q ;
wire \butterfly_st1[3][0][2]~q ;
wire \butterfly_st1[2][1][1]~q ;
wire \butterfly_st1[3][0][1]~q ;
wire \butterfly_st1[2][1][0]~q ;
wire \butterfly_st1[3][0][0]~q ;
wire \butterfly_st2[1][1][0]~2 ;
wire \butterfly_st2[1][1][0]~1_combout ;
wire \butterfly_st2[1][1][1]~2 ;
wire \butterfly_st2[1][1][1]~1_combout ;
wire \butterfly_st2[1][1][2]~2 ;
wire \butterfly_st2[1][1][2]~1_combout ;
wire \butterfly_st1[2][1][8]~q ;
wire \butterfly_st1[3][0][8]~q ;
wire \butterfly_st1[2][1][7]~q ;
wire \butterfly_st1[3][0][7]~q ;
wire \butterfly_st1[2][1][6]~q ;
wire \butterfly_st1[3][0][6]~q ;
wire \butterfly_st1[2][1][5]~q ;
wire \butterfly_st1[3][0][5]~q ;
wire \butterfly_st1[2][1][4]~q ;
wire \butterfly_st1[3][0][4]~q ;
wire \butterfly_st1[2][1][3]~q ;
wire \butterfly_st1[3][0][3]~q ;
wire \butterfly_st2[1][1][3]~2 ;
wire \butterfly_st2[1][1][3]~1_combout ;
wire \butterfly_st2[1][1][4]~2 ;
wire \butterfly_st2[1][1][4]~1_combout ;
wire \butterfly_st2[1][1][5]~2 ;
wire \butterfly_st2[1][1][5]~1_combout ;
wire \butterfly_st2[1][1][6]~2 ;
wire \butterfly_st2[1][1][6]~1_combout ;
wire \butterfly_st2[1][1][7]~2 ;
wire \butterfly_st2[1][1][7]~1_combout ;
wire \butterfly_st2[1][1][8]~2 ;
wire \butterfly_st2[1][1][8]~1_combout ;
wire \butterfly_st2[1][1][9]~1_combout ;
wire \butterfly_st1[2][0][2]~q ;
wire \butterfly_st1[3][1][2]~q ;
wire \butterfly_st1[2][0][1]~q ;
wire \butterfly_st1[3][1][1]~q ;
wire \butterfly_st1[2][0][0]~q ;
wire \butterfly_st1[3][1][0]~q ;
wire \butterfly_st2[1][0][0]~2 ;
wire \butterfly_st2[1][0][0]~1_combout ;
wire \butterfly_st2[1][0][1]~2 ;
wire \butterfly_st2[1][0][1]~1_combout ;
wire \butterfly_st2[1][0][2]~2 ;
wire \butterfly_st2[1][0][2]~1_combout ;
wire \butterfly_st1[2][0][8]~q ;
wire \butterfly_st1[3][1][8]~q ;
wire \butterfly_st1[2][0][7]~q ;
wire \butterfly_st1[3][1][7]~q ;
wire \butterfly_st1[2][0][6]~q ;
wire \butterfly_st1[3][1][6]~q ;
wire \butterfly_st1[2][0][5]~q ;
wire \butterfly_st1[3][1][5]~q ;
wire \butterfly_st1[2][0][4]~q ;
wire \butterfly_st1[3][1][4]~q ;
wire \butterfly_st1[2][0][3]~q ;
wire \butterfly_st1[3][1][3]~q ;
wire \butterfly_st2[1][0][3]~2 ;
wire \butterfly_st2[1][0][3]~1_combout ;
wire \butterfly_st2[1][0][4]~2 ;
wire \butterfly_st2[1][0][4]~1_combout ;
wire \butterfly_st2[1][0][5]~2 ;
wire \butterfly_st2[1][0][5]~1_combout ;
wire \butterfly_st2[1][0][6]~2 ;
wire \butterfly_st2[1][0][6]~1_combout ;
wire \butterfly_st2[1][0][7]~2 ;
wire \butterfly_st2[1][0][7]~1_combout ;
wire \butterfly_st2[1][0][8]~2 ;
wire \butterfly_st2[1][0][8]~1_combout ;
wire \butterfly_st2[1][0][9]~1_combout ;
wire \butterfly_st2[2][1][0]~2 ;
wire \butterfly_st2[2][1][0]~1_combout ;
wire \butterfly_st2[2][1][1]~2 ;
wire \butterfly_st2[2][1][1]~1_combout ;
wire \butterfly_st2[2][1][2]~2 ;
wire \butterfly_st2[2][1][2]~1_combout ;
wire \butterfly_st2[2][1][3]~2 ;
wire \butterfly_st2[2][1][3]~1_combout ;
wire \butterfly_st2[2][1][4]~2 ;
wire \butterfly_st2[2][1][4]~1_combout ;
wire \butterfly_st2[2][1][5]~2 ;
wire \butterfly_st2[2][1][5]~1_combout ;
wire \butterfly_st2[2][1][6]~2 ;
wire \butterfly_st2[2][1][6]~1_combout ;
wire \butterfly_st2[2][1][7]~2 ;
wire \butterfly_st2[2][1][7]~1_combout ;
wire \butterfly_st2[2][1][8]~2 ;
wire \butterfly_st2[2][1][8]~1_combout ;
wire \butterfly_st2[2][1][9]~1_combout ;
wire \butterfly_st2[2][0][0]~2 ;
wire \butterfly_st2[2][0][0]~1_combout ;
wire \butterfly_st2[2][0][1]~2 ;
wire \butterfly_st2[2][0][1]~1_combout ;
wire \butterfly_st2[2][0][2]~2 ;
wire \butterfly_st2[2][0][2]~1_combout ;
wire \butterfly_st2[2][0][3]~2 ;
wire \butterfly_st2[2][0][3]~1_combout ;
wire \butterfly_st2[2][0][4]~2 ;
wire \butterfly_st2[2][0][4]~1_combout ;
wire \butterfly_st2[2][0][5]~2 ;
wire \butterfly_st2[2][0][5]~1_combout ;
wire \butterfly_st2[2][0][6]~2 ;
wire \butterfly_st2[2][0][6]~1_combout ;
wire \butterfly_st2[2][0][7]~2 ;
wire \butterfly_st2[2][0][7]~1_combout ;
wire \butterfly_st2[2][0][8]~2 ;
wire \butterfly_st2[2][0][8]~1_combout ;
wire \butterfly_st2[2][0][9]~1_combout ;
wire \butterfly_st2[3][1][0]~2 ;
wire \butterfly_st2[3][1][0]~1_combout ;
wire \butterfly_st2[3][1][1]~2 ;
wire \butterfly_st2[3][1][1]~1_combout ;
wire \butterfly_st2[3][1][2]~2 ;
wire \butterfly_st2[3][1][2]~1_combout ;
wire \butterfly_st2[3][1][3]~2 ;
wire \butterfly_st2[3][1][3]~1_combout ;
wire \butterfly_st2[3][1][4]~2 ;
wire \butterfly_st2[3][1][4]~1_combout ;
wire \butterfly_st2[3][1][5]~2 ;
wire \butterfly_st2[3][1][5]~1_combout ;
wire \butterfly_st2[3][1][6]~2 ;
wire \butterfly_st2[3][1][6]~1_combout ;
wire \butterfly_st2[3][1][7]~2 ;
wire \butterfly_st2[3][1][7]~1_combout ;
wire \butterfly_st2[3][1][8]~2 ;
wire \butterfly_st2[3][1][8]~1_combout ;
wire \butterfly_st2[3][1][9]~1_combout ;
wire \butterfly_st2[3][0][0]~2 ;
wire \butterfly_st2[3][0][0]~1_combout ;
wire \butterfly_st2[3][0][1]~2 ;
wire \butterfly_st2[3][0][1]~1_combout ;
wire \butterfly_st2[3][0][2]~2 ;
wire \butterfly_st2[3][0][2]~1_combout ;
wire \butterfly_st2[3][0][3]~2 ;
wire \butterfly_st2[3][0][3]~1_combout ;
wire \butterfly_st2[3][0][4]~2 ;
wire \butterfly_st2[3][0][4]~1_combout ;
wire \butterfly_st2[3][0][5]~2 ;
wire \butterfly_st2[3][0][5]~1_combout ;
wire \butterfly_st2[3][0][6]~2 ;
wire \butterfly_st2[3][0][6]~1_combout ;
wire \butterfly_st2[3][0][7]~2 ;
wire \butterfly_st2[3][0][7]~1_combout ;
wire \butterfly_st2[3][0][8]~2 ;
wire \butterfly_st2[3][0][8]~1_combout ;
wire \butterfly_st2[3][0][9]~1_combout ;
wire \gen_cont:bfp_scale|r_array_out[0][5]~q ;
wire \gen_cont:bfp_scale|r_array_out[2][5]~q ;
wire \gen_cont:bfp_scale|r_array_out[0][4]~q ;
wire \gen_cont:bfp_scale|r_array_out[2][4]~q ;
wire \gen_cont:bfp_scale|r_array_out[0][3]~q ;
wire \gen_cont:bfp_scale|r_array_out[2][3]~q ;
wire \gen_cont:bfp_scale|r_array_out[0][2]~q ;
wire \gen_cont:bfp_scale|r_array_out[2][2]~q ;
wire \butterfly_st1[0][0][0]~2 ;
wire \butterfly_st1[0][0][0]~1_combout ;
wire \butterfly_st1[0][0][1]~2 ;
wire \butterfly_st1[0][0][1]~1_combout ;
wire \butterfly_st1[0][0][2]~2 ;
wire \butterfly_st1[0][0][2]~1_combout ;
wire \butterfly_st1[0][0][3]~2 ;
wire \butterfly_st1[0][0][3]~1_combout ;
wire \butterfly_st1[0][0][4]~2 ;
wire \butterfly_st1[0][0][4]~1_combout ;
wire \butterfly_st1[0][0][5]~2 ;
wire \butterfly_st1[0][0][5]~1_combout ;
wire \butterfly_st1[0][0][6]~2 ;
wire \butterfly_st1[0][0][6]~1_combout ;
wire \gen_cont:bfp_scale|r_array_out[1][5]~q ;
wire \gen_cont:bfp_scale|r_array_out[3][5]~q ;
wire \gen_cont:bfp_scale|r_array_out[1][4]~q ;
wire \gen_cont:bfp_scale|r_array_out[3][4]~q ;
wire \gen_cont:bfp_scale|r_array_out[1][3]~q ;
wire \gen_cont:bfp_scale|r_array_out[3][3]~q ;
wire \gen_cont:bfp_scale|r_array_out[1][2]~q ;
wire \gen_cont:bfp_scale|r_array_out[3][2]~q ;
wire \butterfly_st1[1][0][0]~2 ;
wire \butterfly_st1[1][0][0]~1_combout ;
wire \butterfly_st1[1][0][1]~2 ;
wire \butterfly_st1[1][0][1]~1_combout ;
wire \butterfly_st1[1][0][2]~2 ;
wire \butterfly_st1[1][0][2]~1_combout ;
wire \butterfly_st1[1][0][3]~2 ;
wire \butterfly_st1[1][0][3]~1_combout ;
wire \butterfly_st1[1][0][4]~2 ;
wire \butterfly_st1[1][0][4]~1_combout ;
wire \butterfly_st1[1][0][5]~2 ;
wire \butterfly_st1[1][0][5]~1_combout ;
wire \butterfly_st1[1][0][6]~2 ;
wire \butterfly_st1[1][0][6]~1_combout ;
wire \butterfly_st1[0][0][7]~2 ;
wire \butterfly_st1[0][0][7]~1_combout ;
wire \butterfly_st1[0][0][8]~1_combout ;
wire \butterfly_st1[1][0][7]~2 ;
wire \butterfly_st1[1][0][7]~1_combout ;
wire \butterfly_st1[1][0][8]~1_combout ;
wire \gen_cont:bfp_scale|i_array_out[0][5]~q ;
wire \gen_cont:bfp_scale|i_array_out[2][5]~q ;
wire \gen_cont:bfp_scale|i_array_out[0][4]~q ;
wire \gen_cont:bfp_scale|i_array_out[2][4]~q ;
wire \gen_cont:bfp_scale|i_array_out[0][3]~q ;
wire \gen_cont:bfp_scale|i_array_out[2][3]~q ;
wire \gen_cont:bfp_scale|i_array_out[0][2]~q ;
wire \gen_cont:bfp_scale|i_array_out[2][2]~q ;
wire \butterfly_st1[0][1][0]~2 ;
wire \butterfly_st1[0][1][0]~1_combout ;
wire \butterfly_st1[0][1][1]~2 ;
wire \butterfly_st1[0][1][1]~1_combout ;
wire \butterfly_st1[0][1][2]~2 ;
wire \butterfly_st1[0][1][2]~1_combout ;
wire \butterfly_st1[0][1][3]~2 ;
wire \butterfly_st1[0][1][3]~1_combout ;
wire \butterfly_st1[0][1][4]~2 ;
wire \butterfly_st1[0][1][4]~1_combout ;
wire \butterfly_st1[0][1][5]~2 ;
wire \butterfly_st1[0][1][5]~1_combout ;
wire \butterfly_st1[0][1][6]~2 ;
wire \butterfly_st1[0][1][6]~1_combout ;
wire \butterfly_st1[0][1][7]~2 ;
wire \butterfly_st1[0][1][7]~1_combout ;
wire \butterfly_st1[0][1][8]~1_combout ;
wire \gen_cont:bfp_scale|i_array_out[1][5]~q ;
wire \gen_cont:bfp_scale|i_array_out[3][5]~q ;
wire \gen_cont:bfp_scale|i_array_out[1][4]~q ;
wire \gen_cont:bfp_scale|i_array_out[3][4]~q ;
wire \gen_cont:bfp_scale|i_array_out[1][3]~q ;
wire \gen_cont:bfp_scale|i_array_out[3][3]~q ;
wire \gen_cont:bfp_scale|i_array_out[1][2]~q ;
wire \gen_cont:bfp_scale|i_array_out[3][2]~q ;
wire \butterfly_st1[1][1][0]~2 ;
wire \butterfly_st1[1][1][0]~1_combout ;
wire \butterfly_st1[1][1][1]~2 ;
wire \butterfly_st1[1][1][1]~1_combout ;
wire \butterfly_st1[1][1][2]~2 ;
wire \butterfly_st1[1][1][2]~1_combout ;
wire \butterfly_st1[1][1][3]~2 ;
wire \butterfly_st1[1][1][3]~1_combout ;
wire \butterfly_st1[1][1][4]~2 ;
wire \butterfly_st1[1][1][4]~1_combout ;
wire \butterfly_st1[1][1][5]~2 ;
wire \butterfly_st1[1][1][5]~1_combout ;
wire \butterfly_st1[1][1][6]~2 ;
wire \butterfly_st1[1][1][6]~1_combout ;
wire \butterfly_st1[1][1][7]~2 ;
wire \butterfly_st1[1][1][7]~1_combout ;
wire \butterfly_st1[1][1][8]~1_combout ;
wire \butterfly_st1[2][1][0]~2 ;
wire \butterfly_st1[2][1][0]~1_combout ;
wire \butterfly_st1[2][1][1]~2 ;
wire \butterfly_st1[2][1][1]~1_combout ;
wire \butterfly_st1[2][1][2]~2 ;
wire \butterfly_st1[2][1][2]~1_combout ;
wire \butterfly_st1[3][0][0]~2 ;
wire \butterfly_st1[3][0][0]~1_combout ;
wire \butterfly_st1[3][0][1]~2 ;
wire \butterfly_st1[3][0][1]~1_combout ;
wire \butterfly_st1[3][0][2]~2 ;
wire \butterfly_st1[3][0][2]~1_combout ;
wire \butterfly_st1[2][1][3]~2 ;
wire \butterfly_st1[2][1][3]~1_combout ;
wire \butterfly_st1[2][1][4]~2 ;
wire \butterfly_st1[2][1][4]~1_combout ;
wire \butterfly_st1[2][1][5]~2 ;
wire \butterfly_st1[2][1][5]~1_combout ;
wire \butterfly_st1[2][1][6]~2 ;
wire \butterfly_st1[2][1][6]~1_combout ;
wire \butterfly_st1[2][1][7]~2 ;
wire \butterfly_st1[2][1][7]~1_combout ;
wire \butterfly_st1[2][1][8]~1_combout ;
wire \butterfly_st1[3][0][3]~2 ;
wire \butterfly_st1[3][0][3]~1_combout ;
wire \butterfly_st1[3][0][4]~2 ;
wire \butterfly_st1[3][0][4]~1_combout ;
wire \butterfly_st1[3][0][5]~2 ;
wire \butterfly_st1[3][0][5]~1_combout ;
wire \butterfly_st1[3][0][6]~2 ;
wire \butterfly_st1[3][0][6]~1_combout ;
wire \butterfly_st1[3][0][7]~2 ;
wire \butterfly_st1[3][0][7]~1_combout ;
wire \butterfly_st1[3][0][8]~1_combout ;
wire \butterfly_st1[2][0][0]~2 ;
wire \butterfly_st1[2][0][0]~1_combout ;
wire \butterfly_st1[2][0][1]~2 ;
wire \butterfly_st1[2][0][1]~1_combout ;
wire \butterfly_st1[2][0][2]~2 ;
wire \butterfly_st1[2][0][2]~1_combout ;
wire \butterfly_st1[3][1][0]~2 ;
wire \butterfly_st1[3][1][0]~1_combout ;
wire \butterfly_st1[3][1][1]~2 ;
wire \butterfly_st1[3][1][1]~1_combout ;
wire \butterfly_st1[3][1][2]~2 ;
wire \butterfly_st1[3][1][2]~1_combout ;
wire \butterfly_st1[2][0][3]~2 ;
wire \butterfly_st1[2][0][3]~1_combout ;
wire \butterfly_st1[2][0][4]~2 ;
wire \butterfly_st1[2][0][4]~1_combout ;
wire \butterfly_st1[2][0][5]~2 ;
wire \butterfly_st1[2][0][5]~1_combout ;
wire \butterfly_st1[2][0][6]~2 ;
wire \butterfly_st1[2][0][6]~1_combout ;
wire \butterfly_st1[2][0][7]~2 ;
wire \butterfly_st1[2][0][7]~1_combout ;
wire \butterfly_st1[2][0][8]~1_combout ;
wire \butterfly_st1[3][1][3]~2 ;
wire \butterfly_st1[3][1][3]~1_combout ;
wire \butterfly_st1[3][1][4]~2 ;
wire \butterfly_st1[3][1][4]~1_combout ;
wire \butterfly_st1[3][1][5]~2 ;
wire \butterfly_st1[3][1][5]~1_combout ;
wire \butterfly_st1[3][1][6]~2 ;
wire \butterfly_st1[3][1][6]~1_combout ;
wire \butterfly_st1[3][1][7]~2 ;
wire \butterfly_st1[3][1][7]~1_combout ;
wire \butterfly_st1[3][1][8]~1_combout ;
wire \reg_no_twiddle[0][0][1]~q ;
wire \reg_no_twiddle[0][0][0]~q ;
wire \reg_no_twiddle[0][0][2]~q ;
wire \reg_no_twiddle[0][1][1]~q ;
wire \reg_no_twiddle[0][1][0]~q ;
wire \reg_no_twiddle[0][1][2]~q ;
wire \reg_no_twiddle[6][0][3]~q ;
wire \reg_no_twiddle[6][0][7]~q ;
wire \reg_no_twiddle[6][1][7]~q ;
wire \reg_no_twiddle[6][1][3]~q ;
wire \gen_da0:gen_canonic:cm1|real_out[3]~q ;
wire \gen_da0:gen_canonic:cm1|real_out[7]~q ;
wire \gen_da0:gen_canonic:cm2|real_out[3]~q ;
wire \gen_da0:gen_canonic:cm2|real_out[7]~q ;
wire \gen_da0:gen_canonic:cm3|real_out[3]~q ;
wire \gen_da0:gen_canonic:cm3|real_out[7]~q ;
wire \gen_cont:bfp_detect_1pt|gain_lut_8pts[0]~q ;
wire \Selector3~0_combout ;
wire \reg_no_twiddle[6][0][4]~q ;
wire \reg_no_twiddle[6][1][4]~q ;
wire \gen_da0:gen_canonic:cm1|real_out[4]~q ;
wire \gen_da0:gen_canonic:cm2|real_out[4]~q ;
wire \gen_da0:gen_canonic:cm3|real_out[4]~q ;
wire \gen_cont:bfp_detect_1pt|gain_lut_8pts[1]~q ;
wire \Selector2~0_combout ;
wire \reg_no_twiddle[6][0][5]~q ;
wire \reg_no_twiddle[6][1][5]~q ;
wire \gen_da0:gen_canonic:cm1|real_out[5]~q ;
wire \gen_da0:gen_canonic:cm2|real_out[5]~q ;
wire \gen_da0:gen_canonic:cm3|real_out[5]~q ;
wire \gen_cont:bfp_detect_1pt|gain_lut_8pts[2]~q ;
wire \Selector1~0_combout ;
wire \reg_no_twiddle[6][0][6]~q ;
wire \reg_no_twiddle[6][1][6]~q ;
wire \gen_da0:gen_canonic:cm1|real_out[6]~q ;
wire \gen_da0:gen_canonic:cm2|real_out[6]~q ;
wire \gen_da0:gen_canonic:cm3|real_out[6]~q ;
wire \gen_cont:bfp_detect_1pt|gain_lut_8pts[3]~q ;
wire \Selector0~0_combout ;
wire \reg_no_twiddle[5][0][3]~q ;
wire \reg_no_twiddle~0_combout ;
wire \reg_no_twiddle[5][0][7]~q ;
wire \reg_no_twiddle~1_combout ;
wire \reg_no_twiddle[5][1][7]~q ;
wire \reg_no_twiddle~2_combout ;
wire \reg_no_twiddle[5][1][3]~q ;
wire \reg_no_twiddle~3_combout ;
wire \enable_op~q ;
wire \sdft.WAIT_FOR_OUTPUT~q ;
wire \Selector14~0_combout ;
wire \gen_cont:delay_next_blk|tdl_arr[22]~q ;
wire \reg_no_twiddle[5][0][4]~q ;
wire \reg_no_twiddle~4_combout ;
wire \reg_no_twiddle[5][1][4]~q ;
wire \reg_no_twiddle~5_combout ;
wire \reg_no_twiddle[5][0][5]~q ;
wire \reg_no_twiddle~6_combout ;
wire \reg_no_twiddle[5][1][5]~q ;
wire \reg_no_twiddle~7_combout ;
wire \reg_no_twiddle[5][0][6]~q ;
wire \reg_no_twiddle~8_combout ;
wire \reg_no_twiddle[5][1][6]~q ;
wire \reg_no_twiddle~9_combout ;
wire \reg_no_twiddle[4][0][3]~q ;
wire \reg_no_twiddle~10_combout ;
wire \reg_no_twiddle[4][0][7]~q ;
wire \reg_no_twiddle~11_combout ;
wire \reg_no_twiddle[4][1][7]~q ;
wire \reg_no_twiddle~12_combout ;
wire \reg_no_twiddle[4][1][3]~q ;
wire \reg_no_twiddle~13_combout ;
wire \scale_dft_o_en~q ;
wire \do_tdl[0][0][3][3]~q ;
wire \do_tdl[0][0][3][7]~q ;
wire \do_tdl[0][0][3][4]~q ;
wire \do_tdl[0][0][3][5]~q ;
wire \do_tdl[0][0][3][6]~q ;
wire \do_tdl[0][0][3][1]~q ;
wire \do_tdl[0][0][3][0]~q ;
wire \slb_1pt[0]~combout ;
wire \do_tdl[0][0][3][2]~q ;
wire \slb_1pt[2]~0_combout ;
wire \slb_1pt[1]~combout ;
wire \do_tdl[0][1][3][3]~q ;
wire \do_tdl[0][1][3][7]~q ;
wire \do_tdl[0][1][3][4]~q ;
wire \do_tdl[0][1][3][5]~q ;
wire \do_tdl[0][1][3][6]~q ;
wire \do_tdl[0][1][3][1]~q ;
wire \do_tdl[0][1][3][0]~q ;
wire \do_tdl[0][1][3][2]~q ;
wire \do_tdl[1][0][3][3]~q ;
wire \do_tdl[1][0][3][7]~q ;
wire \do_tdl[1][0][3][4]~q ;
wire \do_tdl[1][0][3][5]~q ;
wire \do_tdl[1][0][3][6]~q ;
wire \do_tdl[1][0][3][1]~q ;
wire \do_tdl[1][0][3][0]~q ;
wire \do_tdl[1][0][3][2]~q ;
wire \do_tdl[1][1][3][3]~q ;
wire \do_tdl[1][1][3][7]~q ;
wire \do_tdl[1][1][3][4]~q ;
wire \do_tdl[1][1][3][5]~q ;
wire \do_tdl[1][1][3][6]~q ;
wire \do_tdl[1][1][3][1]~q ;
wire \do_tdl[1][1][3][0]~q ;
wire \do_tdl[1][1][3][2]~q ;
wire \do_tdl[2][0][3][3]~q ;
wire \do_tdl[2][0][3][7]~q ;
wire \do_tdl[2][0][3][4]~q ;
wire \do_tdl[2][0][3][5]~q ;
wire \do_tdl[2][0][3][6]~q ;
wire \do_tdl[2][0][3][1]~q ;
wire \do_tdl[2][0][3][0]~q ;
wire \do_tdl[2][0][3][2]~q ;
wire \do_tdl[2][1][3][3]~q ;
wire \do_tdl[2][1][3][7]~q ;
wire \do_tdl[2][1][3][4]~q ;
wire \do_tdl[2][1][3][5]~q ;
wire \do_tdl[2][1][3][6]~q ;
wire \do_tdl[2][1][3][1]~q ;
wire \do_tdl[2][1][3][0]~q ;
wire \do_tdl[2][1][3][2]~q ;
wire \do_tdl[3][0][3][3]~q ;
wire \do_tdl[3][0][3][7]~q ;
wire \do_tdl[3][0][3][4]~q ;
wire \do_tdl[3][0][3][5]~q ;
wire \do_tdl[3][0][3][6]~q ;
wire \do_tdl[3][0][3][1]~q ;
wire \do_tdl[3][0][3][0]~q ;
wire \do_tdl[3][0][3][2]~q ;
wire \do_tdl[3][1][3][3]~q ;
wire \do_tdl[3][1][3][7]~q ;
wire \do_tdl[3][1][3][4]~q ;
wire \do_tdl[3][1][3][5]~q ;
wire \do_tdl[3][1][3][6]~q ;
wire \do_tdl[3][1][3][1]~q ;
wire \do_tdl[3][1][3][0]~q ;
wire \do_tdl[3][1][3][2]~q ;
wire \gen_cont:delay_next_blk|tdl_arr[25]~q ;
wire \gap_reg~0_combout ;
wire \Equal0~0_combout ;
wire \Equal0~1_combout ;
wire \sdft~8_combout ;
wire \reg_no_twiddle[4][0][4]~q ;
wire \reg_no_twiddle~14_combout ;
wire \reg_no_twiddle[4][1][4]~q ;
wire \reg_no_twiddle~15_combout ;
wire \reg_no_twiddle[4][0][5]~q ;
wire \reg_no_twiddle~16_combout ;
wire \reg_no_twiddle[4][1][5]~q ;
wire \reg_no_twiddle~17_combout ;
wire \reg_no_twiddle[4][0][6]~q ;
wire \reg_no_twiddle~18_combout ;
wire \reg_no_twiddle[4][1][6]~q ;
wire \reg_no_twiddle~19_combout ;
wire \reg_no_twiddle[3][0][3]~q ;
wire \reg_no_twiddle~20_combout ;
wire \reg_no_twiddle[3][0][7]~q ;
wire \reg_no_twiddle~21_combout ;
wire \reg_no_twiddle[3][1][7]~q ;
wire \reg_no_twiddle~22_combout ;
wire \reg_no_twiddle[3][1][3]~q ;
wire \reg_no_twiddle~23_combout ;
wire \Selector5~0_combout ;
wire \do_tdl[0][0][2][3]~q ;
wire \do_tdl[0][0][2][7]~q ;
wire \do_tdl[0][0][2][4]~q ;
wire \do_tdl[0][0][2][5]~q ;
wire \do_tdl[0][0][2][6]~q ;
wire \do_tdl[0][0][2][1]~q ;
wire \do_tdl[0][0][2][0]~q ;
wire \do_tdl[0][0][2][2]~q ;
wire \do_tdl[0][1][2][3]~q ;
wire \do_tdl[0][1][2][7]~q ;
wire \do_tdl[0][1][2][4]~q ;
wire \do_tdl[0][1][2][5]~q ;
wire \do_tdl[0][1][2][6]~q ;
wire \do_tdl[0][1][2][1]~q ;
wire \do_tdl[0][1][2][0]~q ;
wire \do_tdl[0][1][2][2]~q ;
wire \do_tdl[1][0][2][3]~q ;
wire \do_tdl[1][0][2][7]~q ;
wire \do_tdl[1][0][2][4]~q ;
wire \do_tdl[1][0][2][5]~q ;
wire \do_tdl[1][0][2][6]~q ;
wire \do_tdl[1][0][2][1]~q ;
wire \do_tdl[1][0][2][0]~q ;
wire \do_tdl[1][0][2][2]~q ;
wire \do_tdl[1][1][2][3]~q ;
wire \do_tdl[1][1][2][7]~q ;
wire \do_tdl[1][1][2][4]~q ;
wire \do_tdl[1][1][2][5]~q ;
wire \do_tdl[1][1][2][6]~q ;
wire \do_tdl[1][1][2][1]~q ;
wire \do_tdl[1][1][2][0]~q ;
wire \do_tdl[1][1][2][2]~q ;
wire \do_tdl[2][0][2][3]~q ;
wire \do_tdl[2][0][2][7]~q ;
wire \do_tdl[2][0][2][4]~q ;
wire \do_tdl[2][0][2][5]~q ;
wire \do_tdl[2][0][2][6]~q ;
wire \do_tdl[2][0][2][1]~q ;
wire \do_tdl[2][0][2][0]~q ;
wire \do_tdl[2][0][2][2]~q ;
wire \do_tdl[2][1][2][3]~q ;
wire \do_tdl[2][1][2][7]~q ;
wire \do_tdl[2][1][2][4]~q ;
wire \do_tdl[2][1][2][5]~q ;
wire \do_tdl[2][1][2][6]~q ;
wire \do_tdl[2][1][2][1]~q ;
wire \do_tdl[2][1][2][0]~q ;
wire \do_tdl[2][1][2][2]~q ;
wire \do_tdl[3][0][2][3]~q ;
wire \do_tdl[3][0][2][7]~q ;
wire \do_tdl[3][0][2][4]~q ;
wire \do_tdl[3][0][2][5]~q ;
wire \do_tdl[3][0][2][6]~q ;
wire \do_tdl[3][0][2][1]~q ;
wire \do_tdl[3][0][2][0]~q ;
wire \do_tdl[3][0][2][2]~q ;
wire \do_tdl[3][1][2][3]~q ;
wire \do_tdl[3][1][2][7]~q ;
wire \do_tdl[3][1][2][4]~q ;
wire \do_tdl[3][1][2][5]~q ;
wire \do_tdl[3][1][2][6]~q ;
wire \do_tdl[3][1][2][1]~q ;
wire \do_tdl[3][1][2][0]~q ;
wire \do_tdl[3][1][2][2]~q ;
wire \sdft.IDLE~q ;
wire \state_cnt~12_combout ;
wire \state_cnt[0]~13_combout ;
wire \Selector13~0_combout ;
wire \reg_no_twiddle[3][0][4]~q ;
wire \reg_no_twiddle~24_combout ;
wire \reg_no_twiddle[3][1][4]~q ;
wire \reg_no_twiddle~25_combout ;
wire \reg_no_twiddle[3][0][5]~q ;
wire \reg_no_twiddle~26_combout ;
wire \reg_no_twiddle[3][1][5]~q ;
wire \reg_no_twiddle~27_combout ;
wire \reg_no_twiddle[3][0][6]~q ;
wire \reg_no_twiddle~28_combout ;
wire \reg_no_twiddle[3][1][6]~q ;
wire \reg_no_twiddle~29_combout ;
wire \reg_no_twiddle[2][0][3]~q ;
wire \reg_no_twiddle~30_combout ;
wire \reg_no_twiddle[2][0][7]~q ;
wire \reg_no_twiddle~31_combout ;
wire \reg_no_twiddle[2][1][7]~q ;
wire \reg_no_twiddle~32_combout ;
wire \reg_no_twiddle[2][1][3]~q ;
wire \reg_no_twiddle~33_combout ;
wire \Equal1~0_combout ;
wire \Selector15~0_combout ;
wire \do_tdl[0][0][1][3]~q ;
wire \do_tdl[0][0][1][7]~q ;
wire \do_tdl[0][0][1][4]~q ;
wire \do_tdl[0][0][1][5]~q ;
wire \do_tdl[0][0][1][6]~q ;
wire \do_tdl[0][0][1][1]~q ;
wire \do_tdl[0][0][1][0]~q ;
wire \do_tdl[0][0][1][2]~q ;
wire \do_tdl[0][1][1][3]~q ;
wire \do_tdl[0][1][1][7]~q ;
wire \do_tdl[0][1][1][4]~q ;
wire \do_tdl[0][1][1][5]~q ;
wire \do_tdl[0][1][1][6]~q ;
wire \do_tdl[0][1][1][1]~q ;
wire \do_tdl[0][1][1][0]~q ;
wire \do_tdl[0][1][1][2]~q ;
wire \do_tdl[1][0][1][3]~q ;
wire \do_tdl[1][0][1][7]~q ;
wire \do_tdl[1][0][1][4]~q ;
wire \do_tdl[1][0][1][5]~q ;
wire \do_tdl[1][0][1][6]~q ;
wire \do_tdl[1][0][1][1]~q ;
wire \do_tdl[1][0][1][0]~q ;
wire \do_tdl[1][0][1][2]~q ;
wire \do_tdl[1][1][1][3]~q ;
wire \do_tdl[1][1][1][7]~q ;
wire \do_tdl[1][1][1][4]~q ;
wire \do_tdl[1][1][1][5]~q ;
wire \do_tdl[1][1][1][6]~q ;
wire \do_tdl[1][1][1][1]~q ;
wire \do_tdl[1][1][1][0]~q ;
wire \do_tdl[1][1][1][2]~q ;
wire \do_tdl[2][0][1][3]~q ;
wire \do_tdl[2][0][1][7]~q ;
wire \do_tdl[2][0][1][4]~q ;
wire \do_tdl[2][0][1][5]~q ;
wire \do_tdl[2][0][1][6]~q ;
wire \do_tdl[2][0][1][1]~q ;
wire \do_tdl[2][0][1][0]~q ;
wire \do_tdl[2][0][1][2]~q ;
wire \do_tdl[2][1][1][3]~q ;
wire \do_tdl[2][1][1][7]~q ;
wire \do_tdl[2][1][1][4]~q ;
wire \do_tdl[2][1][1][5]~q ;
wire \do_tdl[2][1][1][6]~q ;
wire \do_tdl[2][1][1][1]~q ;
wire \do_tdl[2][1][1][0]~q ;
wire \do_tdl[2][1][1][2]~q ;
wire \do_tdl[3][0][1][3]~q ;
wire \do_tdl[3][0][1][7]~q ;
wire \do_tdl[3][0][1][4]~q ;
wire \do_tdl[3][0][1][5]~q ;
wire \do_tdl[3][0][1][6]~q ;
wire \do_tdl[3][0][1][1]~q ;
wire \do_tdl[3][0][1][0]~q ;
wire \do_tdl[3][0][1][2]~q ;
wire \do_tdl[3][1][1][3]~q ;
wire \do_tdl[3][1][1][7]~q ;
wire \do_tdl[3][1][1][4]~q ;
wire \do_tdl[3][1][1][5]~q ;
wire \do_tdl[3][1][1][6]~q ;
wire \do_tdl[3][1][1][1]~q ;
wire \do_tdl[3][1][1][0]~q ;
wire \do_tdl[3][1][1][2]~q ;
wire \sdft.DISABLE_DFT_O~q ;
wire \sdft.IDLE~0_combout ;
wire \reg_no_twiddle[2][0][4]~q ;
wire \reg_no_twiddle~34_combout ;
wire \reg_no_twiddle[2][1][4]~q ;
wire \reg_no_twiddle~35_combout ;
wire \reg_no_twiddle[2][0][5]~q ;
wire \reg_no_twiddle~36_combout ;
wire \reg_no_twiddle[2][1][5]~q ;
wire \reg_no_twiddle~37_combout ;
wire \reg_no_twiddle[2][0][6]~q ;
wire \reg_no_twiddle~38_combout ;
wire \reg_no_twiddle[2][1][6]~q ;
wire \reg_no_twiddle~39_combout ;
wire \reg_no_twiddle[1][0][3]~q ;
wire \reg_no_twiddle~40_combout ;
wire \reg_no_twiddle[1][0][7]~q ;
wire \reg_no_twiddle~41_combout ;
wire \reg_no_twiddle[1][1][7]~q ;
wire \reg_no_twiddle~42_combout ;
wire \reg_no_twiddle[1][1][3]~q ;
wire \reg_no_twiddle~43_combout ;
wire \do_tdl[0][0][0][3]~q ;
wire \do_tdl[0][0][0][7]~q ;
wire \do_tdl[0][0][0][4]~q ;
wire \do_tdl[0][0][0][5]~q ;
wire \do_tdl[0][0][0][6]~q ;
wire \do_tdl[0][0][0][1]~q ;
wire \do_tdl[0][0][0][0]~q ;
wire \do_tdl[0][0][0][2]~q ;
wire \do_tdl[0][1][0][3]~q ;
wire \do_tdl[0][1][0][7]~q ;
wire \do_tdl[0][1][0][4]~q ;
wire \do_tdl[0][1][0][5]~q ;
wire \do_tdl[0][1][0][6]~q ;
wire \do_tdl[0][1][0][1]~q ;
wire \do_tdl[0][1][0][0]~q ;
wire \do_tdl[0][1][0][2]~q ;
wire \do_tdl[1][0][0][3]~q ;
wire \do_tdl[1][0][0][7]~q ;
wire \do_tdl[1][0][0][4]~q ;
wire \do_tdl[1][0][0][5]~q ;
wire \do_tdl[1][0][0][6]~q ;
wire \do_tdl[1][0][0][1]~q ;
wire \do_tdl[1][0][0][0]~q ;
wire \do_tdl[1][0][0][2]~q ;
wire \do_tdl[1][1][0][3]~q ;
wire \do_tdl[1][1][0][7]~q ;
wire \do_tdl[1][1][0][4]~q ;
wire \do_tdl[1][1][0][5]~q ;
wire \do_tdl[1][1][0][6]~q ;
wire \do_tdl[1][1][0][1]~q ;
wire \do_tdl[1][1][0][0]~q ;
wire \do_tdl[1][1][0][2]~q ;
wire \do_tdl[2][0][0][3]~q ;
wire \do_tdl[2][0][0][7]~q ;
wire \do_tdl[2][0][0][4]~q ;
wire \do_tdl[2][0][0][5]~q ;
wire \do_tdl[2][0][0][6]~q ;
wire \do_tdl[2][0][0][1]~q ;
wire \do_tdl[2][0][0][0]~q ;
wire \do_tdl[2][0][0][2]~q ;
wire \do_tdl[2][1][0][3]~q ;
wire \do_tdl[2][1][0][7]~q ;
wire \do_tdl[2][1][0][4]~q ;
wire \do_tdl[2][1][0][5]~q ;
wire \do_tdl[2][1][0][6]~q ;
wire \do_tdl[2][1][0][1]~q ;
wire \do_tdl[2][1][0][0]~q ;
wire \do_tdl[2][1][0][2]~q ;
wire \do_tdl[3][0][0][3]~q ;
wire \do_tdl[3][0][0][7]~q ;
wire \do_tdl[3][0][0][4]~q ;
wire \do_tdl[3][0][0][5]~q ;
wire \do_tdl[3][0][0][6]~q ;
wire \do_tdl[3][0][0][1]~q ;
wire \do_tdl[3][0][0][0]~q ;
wire \do_tdl[3][0][0][2]~q ;
wire \do_tdl[3][1][0][3]~q ;
wire \do_tdl[3][1][0][7]~q ;
wire \do_tdl[3][1][0][4]~q ;
wire \do_tdl[3][1][0][5]~q ;
wire \do_tdl[3][1][0][6]~q ;
wire \do_tdl[3][1][0][1]~q ;
wire \do_tdl[3][1][0][0]~q ;
wire \do_tdl[3][1][0][2]~q ;
wire \sdft~9_combout ;
wire \reg_no_twiddle[1][0][4]~q ;
wire \reg_no_twiddle~44_combout ;
wire \reg_no_twiddle[1][1][4]~q ;
wire \reg_no_twiddle~45_combout ;
wire \reg_no_twiddle[1][0][5]~q ;
wire \reg_no_twiddle~46_combout ;
wire \reg_no_twiddle[1][1][5]~q ;
wire \reg_no_twiddle~47_combout ;
wire \reg_no_twiddle[1][0][6]~q ;
wire \reg_no_twiddle~48_combout ;
wire \reg_no_twiddle[1][1][6]~q ;
wire \reg_no_twiddle~49_combout ;
wire \reg_no_twiddle~50_combout ;
wire \reg_no_twiddle~51_combout ;
wire \reg_no_twiddle~52_combout ;
wire \reg_no_twiddle~53_combout ;
wire \reg_no_twiddle[6][0][1]~q ;
wire \reg_no_twiddle[6][0][0]~q ;
wire \reg_no_twiddle[6][0][2]~q ;
wire \reg_no_twiddle[6][1][1]~q ;
wire \reg_no_twiddle[6][1][0]~q ;
wire \reg_no_twiddle[6][1][2]~q ;
wire \gen_da0:gen_canonic:cm1|real_out[1]~q ;
wire \gen_da0:gen_canonic:cm1|real_out[0]~q ;
wire \gen_da0:gen_canonic:cm1|real_out[2]~q ;
wire \gen_da0:gen_canonic:cm2|real_out[1]~q ;
wire \gen_da0:gen_canonic:cm2|real_out[0]~q ;
wire \gen_da0:gen_canonic:cm2|real_out[2]~q ;
wire \gen_da0:gen_canonic:cm3|real_out[1]~q ;
wire \gen_da0:gen_canonic:cm3|real_out[0]~q ;
wire \gen_da0:gen_canonic:cm3|real_out[2]~q ;
wire \reg_no_twiddle~54_combout ;
wire \reg_no_twiddle~55_combout ;
wire \reg_no_twiddle~56_combout ;
wire \reg_no_twiddle~57_combout ;
wire \reg_no_twiddle~58_combout ;
wire \reg_no_twiddle~59_combout ;
wire \reg_no_twiddle~60_combout ;
wire \reg_no_twiddle~61_combout ;
wire \reg_no_twiddle[5][0][1]~q ;
wire \reg_no_twiddle~62_combout ;
wire \reg_no_twiddle[5][0][0]~q ;
wire \reg_no_twiddle~63_combout ;
wire \reg_no_twiddle[5][0][2]~q ;
wire \reg_no_twiddle~64_combout ;
wire \reg_no_twiddle[5][1][1]~q ;
wire \reg_no_twiddle~65_combout ;
wire \reg_no_twiddle[5][1][0]~q ;
wire \reg_no_twiddle~66_combout ;
wire \reg_no_twiddle[5][1][2]~q ;
wire \reg_no_twiddle~67_combout ;
wire \reg_no_twiddle[4][0][1]~q ;
wire \reg_no_twiddle~68_combout ;
wire \reg_no_twiddle[4][0][0]~q ;
wire \reg_no_twiddle~69_combout ;
wire \reg_no_twiddle[4][0][2]~q ;
wire \reg_no_twiddle~70_combout ;
wire \reg_no_twiddle[4][1][1]~q ;
wire \reg_no_twiddle~71_combout ;
wire \reg_no_twiddle[4][1][0]~q ;
wire \reg_no_twiddle~72_combout ;
wire \reg_no_twiddle[4][1][2]~q ;
wire \reg_no_twiddle~73_combout ;
wire \reg_no_twiddle[3][0][1]~q ;
wire \reg_no_twiddle~74_combout ;
wire \reg_no_twiddle[3][0][0]~q ;
wire \reg_no_twiddle~75_combout ;
wire \reg_no_twiddle[3][0][2]~q ;
wire \reg_no_twiddle~76_combout ;
wire \reg_no_twiddle[3][1][1]~q ;
wire \reg_no_twiddle~77_combout ;
wire \reg_no_twiddle[3][1][0]~q ;
wire \reg_no_twiddle~78_combout ;
wire \reg_no_twiddle[3][1][2]~q ;
wire \reg_no_twiddle~79_combout ;
wire \gen_cont:bfp_scale|r_array_out[0][6]~q ;
wire \gen_cont:bfp_scale|r_array_out[2][6]~q ;
wire \gen_cont:bfp_scale|r_array_out[0][1]~q ;
wire \gen_cont:bfp_scale|r_array_out[2][1]~q ;
wire \gen_cont:bfp_scale|r_array_out[0][0]~q ;
wire \gen_cont:bfp_scale|r_array_out[2][0]~q ;
wire \gen_cont:bfp_scale|r_array_out[1][6]~q ;
wire \gen_cont:bfp_scale|r_array_out[3][6]~q ;
wire \gen_cont:bfp_scale|r_array_out[1][1]~q ;
wire \gen_cont:bfp_scale|r_array_out[3][1]~q ;
wire \gen_cont:bfp_scale|r_array_out[1][0]~q ;
wire \gen_cont:bfp_scale|r_array_out[3][0]~q ;
wire \gen_cont:bfp_scale|r_array_out[0][7]~q ;
wire \gen_cont:bfp_scale|r_array_out[2][7]~q ;
wire \gen_cont:bfp_scale|r_array_out[1][7]~q ;
wire \gen_cont:bfp_scale|r_array_out[3][7]~q ;
wire \gen_cont:bfp_scale|i_array_out[0][7]~q ;
wire \gen_cont:bfp_scale|i_array_out[2][7]~q ;
wire \gen_cont:bfp_scale|i_array_out[0][6]~q ;
wire \gen_cont:bfp_scale|i_array_out[2][6]~q ;
wire \gen_cont:bfp_scale|i_array_out[0][1]~q ;
wire \gen_cont:bfp_scale|i_array_out[2][1]~q ;
wire \gen_cont:bfp_scale|i_array_out[0][0]~q ;
wire \gen_cont:bfp_scale|i_array_out[2][0]~q ;
wire \gen_cont:bfp_scale|i_array_out[1][7]~q ;
wire \gen_cont:bfp_scale|i_array_out[3][7]~q ;
wire \gen_cont:bfp_scale|i_array_out[1][6]~q ;
wire \gen_cont:bfp_scale|i_array_out[3][6]~q ;
wire \gen_cont:bfp_scale|i_array_out[1][1]~q ;
wire \gen_cont:bfp_scale|i_array_out[3][1]~q ;
wire \gen_cont:bfp_scale|i_array_out[1][0]~q ;
wire \gen_cont:bfp_scale|i_array_out[3][0]~q ;
wire \reg_no_twiddle[2][0][1]~q ;
wire \reg_no_twiddle~80_combout ;
wire \reg_no_twiddle[2][0][0]~q ;
wire \reg_no_twiddle~81_combout ;
wire \reg_no_twiddle[2][0][2]~q ;
wire \reg_no_twiddle~82_combout ;
wire \reg_no_twiddle[2][1][1]~q ;
wire \reg_no_twiddle~83_combout ;
wire \reg_no_twiddle[2][1][0]~q ;
wire \reg_no_twiddle~84_combout ;
wire \reg_no_twiddle[2][1][2]~q ;
wire \reg_no_twiddle~85_combout ;
wire \block_dft_i_en~q ;
wire \slb_nm1[1]~combout ;
wire \slb_nm1[2]~0_combout ;
wire \slb_nm1[0]~combout ;
wire \reg_no_twiddle[1][0][1]~q ;
wire \reg_no_twiddle~86_combout ;
wire \reg_no_twiddle[1][0][0]~q ;
wire \reg_no_twiddle~87_combout ;
wire \reg_no_twiddle[1][0][2]~q ;
wire \reg_no_twiddle~88_combout ;
wire \reg_no_twiddle[1][1][1]~q ;
wire \reg_no_twiddle~89_combout ;
wire \reg_no_twiddle[1][1][0]~q ;
wire \reg_no_twiddle~90_combout ;
wire \reg_no_twiddle[1][1][2]~q ;
wire \reg_no_twiddle~91_combout ;
wire \Selector4~0_combout ;
wire \reg_no_twiddle~92_combout ;
wire \reg_no_twiddle~93_combout ;
wire \reg_no_twiddle~94_combout ;
wire \reg_no_twiddle~95_combout ;
wire \reg_no_twiddle~96_combout ;
wire \reg_no_twiddle~97_combout ;
wire \blk_done_vec~2_combout ;
wire \blk_done_vec[0]~q ;
wire \blk_done_vec~1_combout ;
wire \blk_done_vec[1]~q ;
wire \blk_done_vec~0_combout ;
wire \next_pass_vec~2_combout ;
wire \next_pass_vec[0]~q ;
wire \next_pass_vec~1_combout ;
wire \next_pass_vec[1]~q ;
wire \next_pass_vec~0_combout ;


fft_asj_fft_cmult_can_fft_120_2 \gen_da0:gen_canonic:cm3 (
	.pipeline_dffe_11(\gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_15(\gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_12(\gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_13(\gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ),
	.pipeline_dffe_14(\gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_9(\gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_8(\gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_10(\gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_2(\gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_81(\gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_91(\gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_21(\gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_31(\gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_41(\gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_51(\gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_61(\gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_71(\gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_82(\gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_92(\gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.global_clock_enable(global_clock_enable),
	.real_out_3(\gen_da0:gen_canonic:cm3|real_out[3]~q ),
	.real_out_7(\gen_da0:gen_canonic:cm3|real_out[7]~q ),
	.real_out_4(\gen_da0:gen_canonic:cm3|real_out[4]~q ),
	.real_out_5(\gen_da0:gen_canonic:cm3|real_out[5]~q ),
	.real_out_6(\gen_da0:gen_canonic:cm3|real_out[6]~q ),
	.real_out_1(\gen_da0:gen_canonic:cm3|real_out[1]~q ),
	.real_out_0(\gen_da0:gen_canonic:cm3|real_out[0]~q ),
	.real_out_2(\gen_da0:gen_canonic:cm3|real_out[2]~q ),
	.twiddle_data200(twiddle_data200),
	.twiddle_data201(twiddle_data201),
	.twiddle_data202(twiddle_data202),
	.twiddle_data203(twiddle_data203),
	.twiddle_data204(twiddle_data204),
	.twiddle_data205(twiddle_data205),
	.twiddle_data206(twiddle_data206),
	.twiddle_data207(twiddle_data207),
	.twiddle_data210(twiddle_data210),
	.twiddle_data211(twiddle_data211),
	.twiddle_data212(twiddle_data212),
	.twiddle_data213(twiddle_data213),
	.twiddle_data214(twiddle_data214),
	.twiddle_data215(twiddle_data215),
	.twiddle_data216(twiddle_data216),
	.twiddle_data217(twiddle_data217),
	.clk(clk),
	.reset(reset_n));

fft_asj_fft_cmult_can_fft_120_1 \gen_da0:gen_canonic:cm2 (
	.pipeline_dffe_11(\gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_15(\gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_12(\gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_13(\gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ),
	.pipeline_dffe_14(\gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_9(\gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_8(\gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_10(\gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_2(\gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_81(\gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_91(\gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_21(\gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_31(\gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_41(\gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_51(\gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_61(\gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_71(\gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_82(\gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_92(\gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.global_clock_enable(global_clock_enable),
	.real_out_3(\gen_da0:gen_canonic:cm2|real_out[3]~q ),
	.real_out_7(\gen_da0:gen_canonic:cm2|real_out[7]~q ),
	.real_out_4(\gen_da0:gen_canonic:cm2|real_out[4]~q ),
	.real_out_5(\gen_da0:gen_canonic:cm2|real_out[5]~q ),
	.real_out_6(\gen_da0:gen_canonic:cm2|real_out[6]~q ),
	.real_out_1(\gen_da0:gen_canonic:cm2|real_out[1]~q ),
	.real_out_0(\gen_da0:gen_canonic:cm2|real_out[0]~q ),
	.real_out_2(\gen_da0:gen_canonic:cm2|real_out[2]~q ),
	.twiddle_data100(twiddle_data100),
	.twiddle_data101(twiddle_data101),
	.twiddle_data102(twiddle_data102),
	.twiddle_data103(twiddle_data103),
	.twiddle_data104(twiddle_data104),
	.twiddle_data105(twiddle_data105),
	.twiddle_data106(twiddle_data106),
	.twiddle_data107(twiddle_data107),
	.twiddle_data110(twiddle_data110),
	.twiddle_data111(twiddle_data111),
	.twiddle_data112(twiddle_data112),
	.twiddle_data113(twiddle_data113),
	.twiddle_data114(twiddle_data114),
	.twiddle_data115(twiddle_data115),
	.twiddle_data116(twiddle_data116),
	.twiddle_data117(twiddle_data117),
	.clk(clk),
	.reset(reset_n));

fft_asj_fft_cmult_can_fft_120 \gen_da0:gen_canonic:cm1 (
	.pipeline_dffe_11(\gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_15(\gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_12(\gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_13(\gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ),
	.pipeline_dffe_14(\gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_9(\gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_8(\gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_10(\gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_2(\gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_81(\gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_91(\gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_21(\gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_31(\gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_41(\gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_51(\gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_61(\gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_71(\gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_82(\gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_92(\gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.global_clock_enable(global_clock_enable),
	.real_out_3(\gen_da0:gen_canonic:cm1|real_out[3]~q ),
	.real_out_7(\gen_da0:gen_canonic:cm1|real_out[7]~q ),
	.real_out_4(\gen_da0:gen_canonic:cm1|real_out[4]~q ),
	.real_out_5(\gen_da0:gen_canonic:cm1|real_out[5]~q ),
	.real_out_6(\gen_da0:gen_canonic:cm1|real_out[6]~q ),
	.real_out_1(\gen_da0:gen_canonic:cm1|real_out[1]~q ),
	.real_out_0(\gen_da0:gen_canonic:cm1|real_out[0]~q ),
	.real_out_2(\gen_da0:gen_canonic:cm1|real_out[2]~q ),
	.twiddle_data000(twiddle_data000),
	.twiddle_data001(twiddle_data001),
	.twiddle_data002(twiddle_data002),
	.twiddle_data003(twiddle_data003),
	.twiddle_data004(twiddle_data004),
	.twiddle_data005(twiddle_data005),
	.twiddle_data006(twiddle_data006),
	.twiddle_data007(twiddle_data007),
	.twiddle_data010(twiddle_data010),
	.twiddle_data011(twiddle_data011),
	.twiddle_data012(twiddle_data012),
	.twiddle_data013(twiddle_data013),
	.twiddle_data014(twiddle_data014),
	.twiddle_data015(twiddle_data015),
	.twiddle_data016(twiddle_data016),
	.twiddle_data017(twiddle_data017),
	.clk(clk),
	.reset(reset_n));

fft_asj_fft_tdl_bit_fft_120_2 \gen_cont:delay_next_blk (
	.global_clock_enable(global_clock_enable),
	.data_in(next_block),
	.tdl_arr_4(tdl_arr_4),
	.tdl_arr_3(tdl_arr_3),
	.tdl_arr_22(\gen_cont:delay_next_blk|tdl_arr[22]~q ),
	.tdl_arr_25(\gen_cont:delay_next_blk|tdl_arr[25]~q ),
	.clk(clk));

fft_asj_fft_bfp_o_1pt_fft_120 \gen_cont:bfp_detect_1pt (
	.r_array_out_3_0(r_array_out_3_0),
	.i_array_out_3_0(i_array_out_3_0),
	.r_array_out_3_1(r_array_out_3_1),
	.i_array_out_3_1(i_array_out_3_1),
	.r_array_out_3_2(r_array_out_3_2),
	.i_array_out_3_2(i_array_out_3_2),
	.r_array_out_3_3(r_array_out_3_3),
	.i_array_out_3_3(i_array_out_3_3),
	.r_array_out_4_0(r_array_out_4_0),
	.i_array_out_4_0(i_array_out_4_0),
	.r_array_out_4_1(r_array_out_4_1),
	.i_array_out_4_1(i_array_out_4_1),
	.r_array_out_4_2(r_array_out_4_2),
	.i_array_out_4_2(i_array_out_4_2),
	.r_array_out_4_3(r_array_out_4_3),
	.i_array_out_4_3(i_array_out_4_3),
	.r_array_out_5_0(r_array_out_5_0),
	.i_array_out_5_0(i_array_out_5_0),
	.r_array_out_5_1(r_array_out_5_1),
	.i_array_out_5_1(i_array_out_5_1),
	.r_array_out_5_2(r_array_out_5_2),
	.i_array_out_5_2(i_array_out_5_2),
	.r_array_out_5_3(r_array_out_5_3),
	.i_array_out_5_3(i_array_out_5_3),
	.global_clock_enable(global_clock_enable),
	.gain_lut_8pts_0(\gen_cont:bfp_detect_1pt|gain_lut_8pts[0]~q ),
	.gain_lut_8pts_1(\gen_cont:bfp_detect_1pt|gain_lut_8pts[1]~q ),
	.gain_lut_8pts_2(\gen_cont:bfp_detect_1pt|gain_lut_8pts[2]~q ),
	.gain_lut_8pts_3(\gen_cont:bfp_detect_1pt|gain_lut_8pts[3]~q ),
	.enable_op(\enable_op~q ),
	.r_array_out_7_0(r_array_out_7_0),
	.i_array_out_7_0(i_array_out_7_0),
	.r_array_out_7_1(r_array_out_7_1),
	.i_array_out_7_1(i_array_out_7_1),
	.r_array_out_7_2(r_array_out_7_2),
	.i_array_out_7_2(i_array_out_7_2),
	.r_array_out_7_3(r_array_out_7_3),
	.i_array_out_7_3(i_array_out_7_3),
	.r_array_out_6_0(r_array_out_6_0),
	.i_array_out_6_0(i_array_out_6_0),
	.r_array_out_6_1(r_array_out_6_1),
	.i_array_out_6_1(i_array_out_6_1),
	.r_array_out_6_2(r_array_out_6_2),
	.i_array_out_6_2(i_array_out_6_2),
	.r_array_out_6_3(r_array_out_6_3),
	.i_array_out_6_3(i_array_out_6_3),
	.clk(clk),
	.reset_n(reset_n));

fft_asj_fft_bfp_o_fft_120 \gen_cont:bfp_detect (
	.gain_out_4pts_0(\gain_out_4pts[0]~q ),
	.gain_out_4pts_1(\gain_out_4pts[1]~q ),
	.gain_out_4pts_2(\gain_out_4pts[2]~q ),
	.gain_out_4pts_3(\gain_out_4pts[3]~q ),
	.pipeline_dffe_11(\gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_15(\gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_111(\gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_151(\gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_112(\gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_152(\gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_12(\gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_121(\gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_122(\gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_13(\gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ),
	.pipeline_dffe_131(\gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ),
	.pipeline_dffe_132(\gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ),
	.pipeline_dffe_14(\gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_141(\gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_142(\gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ),
	.global_clock_enable(global_clock_enable),
	.slb_i_0(slb_i_0),
	.slb_i_1(slb_i_1),
	.slb_i_2(slb_i_2),
	.slb_i_3(slb_i_3),
	.Mux2(Mux2),
	.Mux1(Mux1),
	.reg_no_twiddle603(\reg_no_twiddle[6][0][3]~q ),
	.reg_no_twiddle607(\reg_no_twiddle[6][0][7]~q ),
	.reg_no_twiddle617(\reg_no_twiddle[6][1][7]~q ),
	.reg_no_twiddle613(\reg_no_twiddle[6][1][3]~q ),
	.real_out_3(\gen_da0:gen_canonic:cm1|real_out[3]~q ),
	.real_out_7(\gen_da0:gen_canonic:cm1|real_out[7]~q ),
	.real_out_31(\gen_da0:gen_canonic:cm2|real_out[3]~q ),
	.real_out_71(\gen_da0:gen_canonic:cm2|real_out[7]~q ),
	.real_out_32(\gen_da0:gen_canonic:cm3|real_out[3]~q ),
	.real_out_72(\gen_da0:gen_canonic:cm3|real_out[7]~q ),
	.reg_no_twiddle604(\reg_no_twiddle[6][0][4]~q ),
	.reg_no_twiddle614(\reg_no_twiddle[6][1][4]~q ),
	.real_out_4(\gen_da0:gen_canonic:cm1|real_out[4]~q ),
	.real_out_41(\gen_da0:gen_canonic:cm2|real_out[4]~q ),
	.real_out_42(\gen_da0:gen_canonic:cm3|real_out[4]~q ),
	.reg_no_twiddle605(\reg_no_twiddle[6][0][5]~q ),
	.reg_no_twiddle615(\reg_no_twiddle[6][1][5]~q ),
	.real_out_5(\gen_da0:gen_canonic:cm1|real_out[5]~q ),
	.real_out_51(\gen_da0:gen_canonic:cm2|real_out[5]~q ),
	.real_out_52(\gen_da0:gen_canonic:cm3|real_out[5]~q ),
	.reg_no_twiddle606(\reg_no_twiddle[6][0][6]~q ),
	.reg_no_twiddle616(\reg_no_twiddle[6][1][6]~q ),
	.real_out_6(\gen_da0:gen_canonic:cm1|real_out[6]~q ),
	.real_out_61(\gen_da0:gen_canonic:cm2|real_out[6]~q ),
	.real_out_62(\gen_da0:gen_canonic:cm3|real_out[6]~q ),
	.blk_done_vec_2(blk_done_vec_2),
	.tdl_arr_22(\gen_cont:delay_next_blk|tdl_arr[22]~q ),
	.next_pass_vec_2(next_pass_vec_2),
	.clk(clk),
	.reset_n(reset_n));

fft_asj_fft_bfp_i_fft_120_1 \gen_cont:bfp_scale_1pt (
	.r_array_out_3_0(r_array_out_3_0),
	.i_array_out_3_0(i_array_out_3_0),
	.r_array_out_3_1(r_array_out_3_1),
	.i_array_out_3_1(i_array_out_3_1),
	.r_array_out_3_2(r_array_out_3_2),
	.i_array_out_3_2(i_array_out_3_2),
	.r_array_out_3_3(r_array_out_3_3),
	.i_array_out_3_3(i_array_out_3_3),
	.r_array_out_4_0(r_array_out_4_0),
	.i_array_out_4_0(i_array_out_4_0),
	.r_array_out_4_1(r_array_out_4_1),
	.i_array_out_4_1(i_array_out_4_1),
	.r_array_out_4_2(r_array_out_4_2),
	.i_array_out_4_2(i_array_out_4_2),
	.r_array_out_4_3(r_array_out_4_3),
	.i_array_out_4_3(i_array_out_4_3),
	.r_array_out_5_0(r_array_out_5_0),
	.i_array_out_5_0(i_array_out_5_0),
	.r_array_out_5_1(r_array_out_5_1),
	.i_array_out_5_1(i_array_out_5_1),
	.r_array_out_5_2(r_array_out_5_2),
	.i_array_out_5_2(i_array_out_5_2),
	.r_array_out_5_3(r_array_out_5_3),
	.i_array_out_5_3(i_array_out_5_3),
	.i_array_out_2_2(i_array_out_2_2),
	.i_array_out_2_1(i_array_out_2_1),
	.i_array_out_2_0(i_array_out_2_0),
	.i_array_out_2_3(i_array_out_2_3),
	.r_array_out_2_2(r_array_out_2_2),
	.r_array_out_2_1(r_array_out_2_1),
	.r_array_out_2_0(r_array_out_2_0),
	.r_array_out_2_3(r_array_out_2_3),
	.global_clock_enable(global_clock_enable),
	.slb_last_0(slb_last_0),
	.slb_last_1(slb_last_1),
	.slb_last_2(slb_last_2),
	.r_array_out_7_0(r_array_out_7_0),
	.i_array_out_7_0(i_array_out_7_0),
	.r_array_out_7_1(r_array_out_7_1),
	.i_array_out_7_1(i_array_out_7_1),
	.r_array_out_7_2(r_array_out_7_2),
	.i_array_out_7_2(i_array_out_7_2),
	.r_array_out_7_3(r_array_out_7_3),
	.i_array_out_7_3(i_array_out_7_3),
	.r_array_out_6_0(r_array_out_6_0),
	.i_array_out_6_0(i_array_out_6_0),
	.r_array_out_6_1(r_array_out_6_1),
	.i_array_out_6_1(i_array_out_6_1),
	.r_array_out_6_2(r_array_out_6_2),
	.i_array_out_6_2(i_array_out_6_2),
	.r_array_out_6_3(r_array_out_6_3),
	.i_array_out_6_3(i_array_out_6_3),
	.i_array_out_1_2(i_array_out_1_2),
	.i_array_out_1_1(i_array_out_1_1),
	.i_array_out_1_0(i_array_out_1_0),
	.i_array_out_1_3(i_array_out_1_3),
	.i_array_out_0_2(i_array_out_0_2),
	.i_array_out_0_1(i_array_out_0_1),
	.i_array_out_0_0(i_array_out_0_0),
	.i_array_out_0_3(i_array_out_0_3),
	.r_array_out_1_2(r_array_out_1_2),
	.r_array_out_1_1(r_array_out_1_1),
	.r_array_out_1_0(r_array_out_1_0),
	.r_array_out_1_3(r_array_out_1_3),
	.r_array_out_0_2(r_array_out_0_2),
	.r_array_out_0_1(r_array_out_0_1),
	.r_array_out_0_0(r_array_out_0_0),
	.r_array_out_0_3(r_array_out_0_3),
	.scale_dft_o_en(\scale_dft_o_en~q ),
	.do_tdl0033(\do_tdl[0][0][3][3]~q ),
	.do_tdl0037(\do_tdl[0][0][3][7]~q ),
	.do_tdl0034(\do_tdl[0][0][3][4]~q ),
	.do_tdl0035(\do_tdl[0][0][3][5]~q ),
	.do_tdl0036(\do_tdl[0][0][3][6]~q ),
	.do_tdl0031(\do_tdl[0][0][3][1]~q ),
	.do_tdl0030(\do_tdl[0][0][3][0]~q ),
	.slb_1pt_0(\slb_1pt[0]~combout ),
	.do_tdl0032(\do_tdl[0][0][3][2]~q ),
	.slb_1pt_2(\slb_1pt[2]~0_combout ),
	.slb_1pt_1(\slb_1pt[1]~combout ),
	.do_tdl0133(\do_tdl[0][1][3][3]~q ),
	.do_tdl0137(\do_tdl[0][1][3][7]~q ),
	.do_tdl0134(\do_tdl[0][1][3][4]~q ),
	.do_tdl0135(\do_tdl[0][1][3][5]~q ),
	.do_tdl0136(\do_tdl[0][1][3][6]~q ),
	.do_tdl0131(\do_tdl[0][1][3][1]~q ),
	.do_tdl0130(\do_tdl[0][1][3][0]~q ),
	.do_tdl0132(\do_tdl[0][1][3][2]~q ),
	.do_tdl1033(\do_tdl[1][0][3][3]~q ),
	.do_tdl1037(\do_tdl[1][0][3][7]~q ),
	.do_tdl1034(\do_tdl[1][0][3][4]~q ),
	.do_tdl1035(\do_tdl[1][0][3][5]~q ),
	.do_tdl1036(\do_tdl[1][0][3][6]~q ),
	.do_tdl1031(\do_tdl[1][0][3][1]~q ),
	.do_tdl1030(\do_tdl[1][0][3][0]~q ),
	.do_tdl1032(\do_tdl[1][0][3][2]~q ),
	.do_tdl1133(\do_tdl[1][1][3][3]~q ),
	.do_tdl1137(\do_tdl[1][1][3][7]~q ),
	.do_tdl1134(\do_tdl[1][1][3][4]~q ),
	.do_tdl1135(\do_tdl[1][1][3][5]~q ),
	.do_tdl1136(\do_tdl[1][1][3][6]~q ),
	.do_tdl1131(\do_tdl[1][1][3][1]~q ),
	.do_tdl1130(\do_tdl[1][1][3][0]~q ),
	.do_tdl1132(\do_tdl[1][1][3][2]~q ),
	.do_tdl2033(\do_tdl[2][0][3][3]~q ),
	.do_tdl2037(\do_tdl[2][0][3][7]~q ),
	.do_tdl2034(\do_tdl[2][0][3][4]~q ),
	.do_tdl2035(\do_tdl[2][0][3][5]~q ),
	.do_tdl2036(\do_tdl[2][0][3][6]~q ),
	.do_tdl2031(\do_tdl[2][0][3][1]~q ),
	.do_tdl2030(\do_tdl[2][0][3][0]~q ),
	.do_tdl2032(\do_tdl[2][0][3][2]~q ),
	.do_tdl2133(\do_tdl[2][1][3][3]~q ),
	.do_tdl2137(\do_tdl[2][1][3][7]~q ),
	.do_tdl2134(\do_tdl[2][1][3][4]~q ),
	.do_tdl2135(\do_tdl[2][1][3][5]~q ),
	.do_tdl2136(\do_tdl[2][1][3][6]~q ),
	.do_tdl2131(\do_tdl[2][1][3][1]~q ),
	.do_tdl2130(\do_tdl[2][1][3][0]~q ),
	.do_tdl2132(\do_tdl[2][1][3][2]~q ),
	.do_tdl3033(\do_tdl[3][0][3][3]~q ),
	.do_tdl3037(\do_tdl[3][0][3][7]~q ),
	.do_tdl3034(\do_tdl[3][0][3][4]~q ),
	.do_tdl3035(\do_tdl[3][0][3][5]~q ),
	.do_tdl3036(\do_tdl[3][0][3][6]~q ),
	.do_tdl3031(\do_tdl[3][0][3][1]~q ),
	.do_tdl3030(\do_tdl[3][0][3][0]~q ),
	.do_tdl3032(\do_tdl[3][0][3][2]~q ),
	.do_tdl3133(\do_tdl[3][1][3][3]~q ),
	.do_tdl3137(\do_tdl[3][1][3][7]~q ),
	.do_tdl3134(\do_tdl[3][1][3][4]~q ),
	.do_tdl3135(\do_tdl[3][1][3][5]~q ),
	.do_tdl3136(\do_tdl[3][1][3][6]~q ),
	.do_tdl3131(\do_tdl[3][1][3][1]~q ),
	.do_tdl3130(\do_tdl[3][1][3][0]~q ),
	.do_tdl3132(\do_tdl[3][1][3][2]~q ),
	.clk(clk));

fft_asj_fft_bfp_i_fft_120 \gen_cont:bfp_scale (
	.r_array_out_5_0(\gen_cont:bfp_scale|r_array_out[0][5]~q ),
	.r_array_out_5_2(\gen_cont:bfp_scale|r_array_out[2][5]~q ),
	.r_array_out_4_0(\gen_cont:bfp_scale|r_array_out[0][4]~q ),
	.r_array_out_4_2(\gen_cont:bfp_scale|r_array_out[2][4]~q ),
	.r_array_out_3_0(\gen_cont:bfp_scale|r_array_out[0][3]~q ),
	.r_array_out_3_2(\gen_cont:bfp_scale|r_array_out[2][3]~q ),
	.r_array_out_2_0(\gen_cont:bfp_scale|r_array_out[0][2]~q ),
	.r_array_out_2_2(\gen_cont:bfp_scale|r_array_out[2][2]~q ),
	.r_array_out_5_1(\gen_cont:bfp_scale|r_array_out[1][5]~q ),
	.r_array_out_5_3(\gen_cont:bfp_scale|r_array_out[3][5]~q ),
	.r_array_out_4_1(\gen_cont:bfp_scale|r_array_out[1][4]~q ),
	.r_array_out_4_3(\gen_cont:bfp_scale|r_array_out[3][4]~q ),
	.r_array_out_3_1(\gen_cont:bfp_scale|r_array_out[1][3]~q ),
	.r_array_out_3_3(\gen_cont:bfp_scale|r_array_out[3][3]~q ),
	.r_array_out_2_1(\gen_cont:bfp_scale|r_array_out[1][2]~q ),
	.r_array_out_2_3(\gen_cont:bfp_scale|r_array_out[3][2]~q ),
	.i_array_out_5_0(\gen_cont:bfp_scale|i_array_out[0][5]~q ),
	.i_array_out_5_2(\gen_cont:bfp_scale|i_array_out[2][5]~q ),
	.i_array_out_4_0(\gen_cont:bfp_scale|i_array_out[0][4]~q ),
	.i_array_out_4_2(\gen_cont:bfp_scale|i_array_out[2][4]~q ),
	.i_array_out_3_0(\gen_cont:bfp_scale|i_array_out[0][3]~q ),
	.i_array_out_3_2(\gen_cont:bfp_scale|i_array_out[2][3]~q ),
	.i_array_out_2_0(\gen_cont:bfp_scale|i_array_out[0][2]~q ),
	.i_array_out_2_2(\gen_cont:bfp_scale|i_array_out[2][2]~q ),
	.i_array_out_5_1(\gen_cont:bfp_scale|i_array_out[1][5]~q ),
	.i_array_out_5_3(\gen_cont:bfp_scale|i_array_out[3][5]~q ),
	.i_array_out_4_1(\gen_cont:bfp_scale|i_array_out[1][4]~q ),
	.i_array_out_4_3(\gen_cont:bfp_scale|i_array_out[3][4]~q ),
	.i_array_out_3_1(\gen_cont:bfp_scale|i_array_out[1][3]~q ),
	.i_array_out_3_3(\gen_cont:bfp_scale|i_array_out[3][3]~q ),
	.i_array_out_2_1(\gen_cont:bfp_scale|i_array_out[1][2]~q ),
	.i_array_out_2_3(\gen_cont:bfp_scale|i_array_out[3][2]~q ),
	.ram_in_reg_2_0(ram_in_reg_2_0),
	.ram_in_reg_6_0(ram_in_reg_6_0),
	.ram_in_reg_4_0(ram_in_reg_4_0),
	.ram_in_reg_3_0(ram_in_reg_3_0),
	.ram_in_reg_5_0(ram_in_reg_5_0),
	.ram_in_reg_2_2(ram_in_reg_2_2),
	.ram_in_reg_6_2(ram_in_reg_6_2),
	.ram_in_reg_4_2(ram_in_reg_4_2),
	.ram_in_reg_3_2(ram_in_reg_3_2),
	.ram_in_reg_5_2(ram_in_reg_5_2),
	.ram_in_reg_1_0(ram_in_reg_1_0),
	.ram_in_reg_1_2(ram_in_reg_1_2),
	.ram_in_reg_0_0(ram_in_reg_0_0),
	.ram_in_reg_0_2(ram_in_reg_0_2),
	.ram_in_reg_2_1(ram_in_reg_2_1),
	.ram_in_reg_6_1(ram_in_reg_6_1),
	.ram_in_reg_4_1(ram_in_reg_4_1),
	.ram_in_reg_3_1(ram_in_reg_3_1),
	.ram_in_reg_5_1(ram_in_reg_5_1),
	.ram_in_reg_2_3(ram_in_reg_2_3),
	.ram_in_reg_6_3(ram_in_reg_6_3),
	.ram_in_reg_4_3(ram_in_reg_4_3),
	.ram_in_reg_3_3(ram_in_reg_3_3),
	.ram_in_reg_5_3(ram_in_reg_5_3),
	.ram_in_reg_1_1(ram_in_reg_1_1),
	.ram_in_reg_1_3(ram_in_reg_1_3),
	.ram_in_reg_0_1(ram_in_reg_0_1),
	.ram_in_reg_0_3(ram_in_reg_0_3),
	.ram_in_reg_7_0(ram_in_reg_7_0),
	.ram_in_reg_7_2(ram_in_reg_7_2),
	.ram_in_reg_7_1(ram_in_reg_7_1),
	.ram_in_reg_7_3(ram_in_reg_7_3),
	.ram_in_reg_7_4(ram_in_reg_7_4),
	.ram_in_reg_3_4(ram_in_reg_3_4),
	.ram_in_reg_5_4(ram_in_reg_5_4),
	.ram_in_reg_4_4(ram_in_reg_4_4),
	.ram_in_reg_6_4(ram_in_reg_6_4),
	.ram_in_reg_7_6(ram_in_reg_7_6),
	.ram_in_reg_3_6(ram_in_reg_3_6),
	.ram_in_reg_5_6(ram_in_reg_5_6),
	.ram_in_reg_4_6(ram_in_reg_4_6),
	.ram_in_reg_6_6(ram_in_reg_6_6),
	.ram_in_reg_2_4(ram_in_reg_2_4),
	.ram_in_reg_2_6(ram_in_reg_2_6),
	.ram_in_reg_1_4(ram_in_reg_1_4),
	.ram_in_reg_1_6(ram_in_reg_1_6),
	.ram_in_reg_0_4(ram_in_reg_0_4),
	.ram_in_reg_0_6(ram_in_reg_0_6),
	.ram_in_reg_7_5(ram_in_reg_7_5),
	.ram_in_reg_3_5(ram_in_reg_3_5),
	.ram_in_reg_5_5(ram_in_reg_5_5),
	.ram_in_reg_4_5(ram_in_reg_4_5),
	.ram_in_reg_6_5(ram_in_reg_6_5),
	.ram_in_reg_3_7(ram_in_reg_3_7),
	.ram_in_reg_7_7(ram_in_reg_7_7),
	.ram_in_reg_5_7(ram_in_reg_5_7),
	.ram_in_reg_4_7(ram_in_reg_4_7),
	.ram_in_reg_6_7(ram_in_reg_6_7),
	.ram_in_reg_2_5(ram_in_reg_2_5),
	.ram_in_reg_2_7(ram_in_reg_2_7),
	.ram_in_reg_1_5(ram_in_reg_1_5),
	.ram_in_reg_1_7(ram_in_reg_1_7),
	.ram_in_reg_0_5(ram_in_reg_0_5),
	.ram_in_reg_0_7(ram_in_reg_0_7),
	.global_clock_enable(global_clock_enable),
	.slb_last_0(slb_last_0),
	.slb_last_1(slb_last_1),
	.slb_last_2(slb_last_2),
	.r_array_out_6_0(\gen_cont:bfp_scale|r_array_out[0][6]~q ),
	.r_array_out_6_2(\gen_cont:bfp_scale|r_array_out[2][6]~q ),
	.r_array_out_1_0(\gen_cont:bfp_scale|r_array_out[0][1]~q ),
	.r_array_out_1_2(\gen_cont:bfp_scale|r_array_out[2][1]~q ),
	.r_array_out_0_0(\gen_cont:bfp_scale|r_array_out[0][0]~q ),
	.r_array_out_0_2(\gen_cont:bfp_scale|r_array_out[2][0]~q ),
	.r_array_out_6_1(\gen_cont:bfp_scale|r_array_out[1][6]~q ),
	.r_array_out_6_3(\gen_cont:bfp_scale|r_array_out[3][6]~q ),
	.r_array_out_1_1(\gen_cont:bfp_scale|r_array_out[1][1]~q ),
	.r_array_out_1_3(\gen_cont:bfp_scale|r_array_out[3][1]~q ),
	.r_array_out_0_1(\gen_cont:bfp_scale|r_array_out[1][0]~q ),
	.r_array_out_0_3(\gen_cont:bfp_scale|r_array_out[3][0]~q ),
	.r_array_out_7_0(\gen_cont:bfp_scale|r_array_out[0][7]~q ),
	.r_array_out_7_2(\gen_cont:bfp_scale|r_array_out[2][7]~q ),
	.r_array_out_7_1(\gen_cont:bfp_scale|r_array_out[1][7]~q ),
	.r_array_out_7_3(\gen_cont:bfp_scale|r_array_out[3][7]~q ),
	.i_array_out_7_0(\gen_cont:bfp_scale|i_array_out[0][7]~q ),
	.i_array_out_7_2(\gen_cont:bfp_scale|i_array_out[2][7]~q ),
	.i_array_out_6_0(\gen_cont:bfp_scale|i_array_out[0][6]~q ),
	.i_array_out_6_2(\gen_cont:bfp_scale|i_array_out[2][6]~q ),
	.i_array_out_1_0(\gen_cont:bfp_scale|i_array_out[0][1]~q ),
	.i_array_out_1_2(\gen_cont:bfp_scale|i_array_out[2][1]~q ),
	.i_array_out_0_0(\gen_cont:bfp_scale|i_array_out[0][0]~q ),
	.i_array_out_0_2(\gen_cont:bfp_scale|i_array_out[2][0]~q ),
	.i_array_out_7_1(\gen_cont:bfp_scale|i_array_out[1][7]~q ),
	.i_array_out_7_3(\gen_cont:bfp_scale|i_array_out[3][7]~q ),
	.i_array_out_6_1(\gen_cont:bfp_scale|i_array_out[1][6]~q ),
	.i_array_out_6_3(\gen_cont:bfp_scale|i_array_out[3][6]~q ),
	.i_array_out_1_1(\gen_cont:bfp_scale|i_array_out[1][1]~q ),
	.i_array_out_1_3(\gen_cont:bfp_scale|i_array_out[3][1]~q ),
	.i_array_out_0_1(\gen_cont:bfp_scale|i_array_out[1][0]~q ),
	.i_array_out_0_3(\gen_cont:bfp_scale|i_array_out[3][0]~q ),
	.block_dft_i_en(\block_dft_i_en~q ),
	.slb_nm1_1(\slb_nm1[1]~combout ),
	.slb_nm1_2(\slb_nm1[2]~0_combout ),
	.slb_nm1_0(\slb_nm1[0]~combout ),
	.clk(clk));

fft_asj_fft_pround_fft_120_13 \gen_full_rnd:gen_rounding_blk:3:u1 (
	.pipeline_dffe_2(\gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.butterfly_st2312(\butterfly_st2[3][1][2]~q ),
	.butterfly_st2311(\butterfly_st2[3][1][1]~q ),
	.butterfly_st2310(\butterfly_st2[3][1][0]~q ),
	.butterfly_st2319(\butterfly_st2[3][1][9]~q ),
	.butterfly_st2313(\butterfly_st2[3][1][3]~q ),
	.butterfly_st2314(\butterfly_st2[3][1][4]~q ),
	.butterfly_st2315(\butterfly_st2[3][1][5]~q ),
	.butterfly_st2316(\butterfly_st2[3][1][6]~q ),
	.butterfly_st2317(\butterfly_st2[3][1][7]~q ),
	.butterfly_st2318(\butterfly_st2[3][1][8]~q ),
	.global_clock_enable(global_clock_enable),
	.clk(clk));

fft_asj_fft_pround_fft_120_12 \gen_full_rnd:gen_rounding_blk:3:u0 (
	.pipeline_dffe_2(\gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.butterfly_st2302(\butterfly_st2[3][0][2]~q ),
	.butterfly_st2301(\butterfly_st2[3][0][1]~q ),
	.butterfly_st2300(\butterfly_st2[3][0][0]~q ),
	.butterfly_st2309(\butterfly_st2[3][0][9]~q ),
	.butterfly_st2303(\butterfly_st2[3][0][3]~q ),
	.butterfly_st2304(\butterfly_st2[3][0][4]~q ),
	.butterfly_st2305(\butterfly_st2[3][0][5]~q ),
	.butterfly_st2306(\butterfly_st2[3][0][6]~q ),
	.butterfly_st2307(\butterfly_st2[3][0][7]~q ),
	.butterfly_st2308(\butterfly_st2[3][0][8]~q ),
	.global_clock_enable(global_clock_enable),
	.clk(clk));

fft_asj_fft_pround_fft_120_11 \gen_full_rnd:gen_rounding_blk:2:u1 (
	.pipeline_dffe_2(\gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.butterfly_st2212(\butterfly_st2[2][1][2]~q ),
	.butterfly_st2211(\butterfly_st2[2][1][1]~q ),
	.butterfly_st2210(\butterfly_st2[2][1][0]~q ),
	.butterfly_st2219(\butterfly_st2[2][1][9]~q ),
	.butterfly_st2213(\butterfly_st2[2][1][3]~q ),
	.butterfly_st2214(\butterfly_st2[2][1][4]~q ),
	.butterfly_st2215(\butterfly_st2[2][1][5]~q ),
	.butterfly_st2216(\butterfly_st2[2][1][6]~q ),
	.butterfly_st2217(\butterfly_st2[2][1][7]~q ),
	.butterfly_st2218(\butterfly_st2[2][1][8]~q ),
	.global_clock_enable(global_clock_enable),
	.clk(clk));

fft_asj_fft_pround_fft_120_10 \gen_full_rnd:gen_rounding_blk:2:u0 (
	.pipeline_dffe_2(\gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.butterfly_st2202(\butterfly_st2[2][0][2]~q ),
	.butterfly_st2201(\butterfly_st2[2][0][1]~q ),
	.butterfly_st2200(\butterfly_st2[2][0][0]~q ),
	.butterfly_st2209(\butterfly_st2[2][0][9]~q ),
	.butterfly_st2203(\butterfly_st2[2][0][3]~q ),
	.butterfly_st2204(\butterfly_st2[2][0][4]~q ),
	.butterfly_st2205(\butterfly_st2[2][0][5]~q ),
	.butterfly_st2206(\butterfly_st2[2][0][6]~q ),
	.butterfly_st2207(\butterfly_st2[2][0][7]~q ),
	.butterfly_st2208(\butterfly_st2[2][0][8]~q ),
	.global_clock_enable(global_clock_enable),
	.clk(clk));

fft_asj_fft_pround_fft_120_9 \gen_full_rnd:gen_rounding_blk:1:u1 (
	.pipeline_dffe_2(\gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.butterfly_st2112(\butterfly_st2[1][1][2]~q ),
	.butterfly_st2111(\butterfly_st2[1][1][1]~q ),
	.butterfly_st2110(\butterfly_st2[1][1][0]~q ),
	.butterfly_st2119(\butterfly_st2[1][1][9]~q ),
	.butterfly_st2113(\butterfly_st2[1][1][3]~q ),
	.butterfly_st2114(\butterfly_st2[1][1][4]~q ),
	.butterfly_st2115(\butterfly_st2[1][1][5]~q ),
	.butterfly_st2116(\butterfly_st2[1][1][6]~q ),
	.butterfly_st2117(\butterfly_st2[1][1][7]~q ),
	.butterfly_st2118(\butterfly_st2[1][1][8]~q ),
	.global_clock_enable(global_clock_enable),
	.clk(clk));

fft_asj_fft_pround_fft_120_8 \gen_full_rnd:gen_rounding_blk:1:u0 (
	.pipeline_dffe_2(\gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.butterfly_st2102(\butterfly_st2[1][0][2]~q ),
	.butterfly_st2101(\butterfly_st2[1][0][1]~q ),
	.butterfly_st2100(\butterfly_st2[1][0][0]~q ),
	.butterfly_st2109(\butterfly_st2[1][0][9]~q ),
	.butterfly_st2103(\butterfly_st2[1][0][3]~q ),
	.butterfly_st2104(\butterfly_st2[1][0][4]~q ),
	.butterfly_st2105(\butterfly_st2[1][0][5]~q ),
	.butterfly_st2106(\butterfly_st2[1][0][6]~q ),
	.butterfly_st2107(\butterfly_st2[1][0][7]~q ),
	.butterfly_st2108(\butterfly_st2[1][0][8]~q ),
	.global_clock_enable(global_clock_enable),
	.clk(clk));

fft_asj_fft_pround_fft_120_7 \gen_full_rnd:gen_rounding_blk:0:u1 (
	.pipeline_dffe_9(\gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_8(\gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_7(\gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_6(\gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_5(\gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_4(\gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_3(\gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_2(\gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.butterfly_st2019(\butterfly_st2[0][1][9]~q ),
	.butterfly_st2018(\butterfly_st2[0][1][8]~q ),
	.butterfly_st2017(\butterfly_st2[0][1][7]~q ),
	.butterfly_st2016(\butterfly_st2[0][1][6]~q ),
	.butterfly_st2015(\butterfly_st2[0][1][5]~q ),
	.butterfly_st2014(\butterfly_st2[0][1][4]~q ),
	.butterfly_st2013(\butterfly_st2[0][1][3]~q ),
	.butterfly_st2012(\butterfly_st2[0][1][2]~q ),
	.butterfly_st2011(\butterfly_st2[0][1][1]~q ),
	.butterfly_st2010(\butterfly_st2[0][1][0]~q ),
	.global_clock_enable(global_clock_enable),
	.clk(clk));

fft_asj_fft_pround_fft_120_6 \gen_full_rnd:gen_rounding_blk:0:u0 (
	.pipeline_dffe_6(\gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_5(\gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_4(\gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_3(\gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_2(\gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_9(\gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_8(\gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_7(\gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.butterfly_st2006(\butterfly_st2[0][0][6]~q ),
	.butterfly_st2005(\butterfly_st2[0][0][5]~q ),
	.butterfly_st2004(\butterfly_st2[0][0][4]~q ),
	.butterfly_st2003(\butterfly_st2[0][0][3]~q ),
	.butterfly_st2002(\butterfly_st2[0][0][2]~q ),
	.butterfly_st2001(\butterfly_st2[0][0][1]~q ),
	.butterfly_st2000(\butterfly_st2[0][0][0]~q ),
	.butterfly_st2009(\butterfly_st2[0][0][9]~q ),
	.butterfly_st2008(\butterfly_st2[0][0][8]~q ),
	.butterfly_st2007(\butterfly_st2[0][0][7]~q ),
	.global_clock_enable(global_clock_enable),
	.clk(clk));

dffeas \gain_out_4pts[0] (
	.clk(clk),
	.d(\Selector3~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\gain_out_4pts[0]~q ),
	.prn(vcc));
defparam \gain_out_4pts[0] .is_wysiwyg = "true";
defparam \gain_out_4pts[0] .power_up = "low";

dffeas \gain_out_4pts[1] (
	.clk(clk),
	.d(\Selector2~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\gain_out_4pts[1]~q ),
	.prn(vcc));
defparam \gain_out_4pts[1] .is_wysiwyg = "true";
defparam \gain_out_4pts[1] .power_up = "low";

dffeas \gain_out_4pts[2] (
	.clk(clk),
	.d(\Selector1~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\gain_out_4pts[2]~q ),
	.prn(vcc));
defparam \gain_out_4pts[2] .is_wysiwyg = "true";
defparam \gain_out_4pts[2] .power_up = "low";

dffeas \gain_out_4pts[3] (
	.clk(clk),
	.d(\Selector0~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\gain_out_4pts[3]~q ),
	.prn(vcc));
defparam \gain_out_4pts[3] .is_wysiwyg = "true";
defparam \gain_out_4pts[3] .power_up = "low";

dffeas \sdft.ENABLE_DFT_O (
	.clk(clk),
	.d(\Selector14~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sdft.ENABLE_DFT_O~q ),
	.prn(vcc));
defparam \sdft.ENABLE_DFT_O .is_wysiwyg = "true";
defparam \sdft.ENABLE_DFT_O .power_up = "low";

dffeas gap_reg(
	.clk(clk),
	.d(\gap_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\gap_reg~q ),
	.prn(vcc));
defparam gap_reg.is_wysiwyg = "true";
defparam gap_reg.power_up = "low";

dffeas \state_cnt[2] (
	.clk(clk),
	.d(\state_cnt[2]~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\state_cnt~12_combout ),
	.sload(gnd),
	.ena(\state_cnt[0]~13_combout ),
	.q(\state_cnt[2]~q ),
	.prn(vcc));
defparam \state_cnt[2] .is_wysiwyg = "true";
defparam \state_cnt[2] .power_up = "low";

dffeas \state_cnt[3] (
	.clk(clk),
	.d(\state_cnt[3]~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\state_cnt~12_combout ),
	.sload(gnd),
	.ena(\state_cnt[0]~13_combout ),
	.q(\state_cnt[3]~q ),
	.prn(vcc));
defparam \state_cnt[3] .is_wysiwyg = "true";
defparam \state_cnt[3] .power_up = "low";

dffeas \state_cnt[4] (
	.clk(clk),
	.d(\state_cnt[4]~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\state_cnt~12_combout ),
	.sload(gnd),
	.ena(\state_cnt[0]~13_combout ),
	.q(\state_cnt[4]~q ),
	.prn(vcc));
defparam \state_cnt[4] .is_wysiwyg = "true";
defparam \state_cnt[4] .power_up = "low";

dffeas \state_cnt[5] (
	.clk(clk),
	.d(\state_cnt[5]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\state_cnt~12_combout ),
	.sload(gnd),
	.ena(\state_cnt[0]~13_combout ),
	.q(\state_cnt[5]~q ),
	.prn(vcc));
defparam \state_cnt[5] .is_wysiwyg = "true";
defparam \state_cnt[5] .power_up = "low";

dffeas \state_cnt[0] (
	.clk(clk),
	.d(\state_cnt[0]~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\state_cnt~12_combout ),
	.sload(gnd),
	.ena(\state_cnt[0]~13_combout ),
	.q(\state_cnt[0]~q ),
	.prn(vcc));
defparam \state_cnt[0] .is_wysiwyg = "true";
defparam \state_cnt[0] .power_up = "low";

dffeas \state_cnt[1] (
	.clk(clk),
	.d(\state_cnt[1]~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\state_cnt~12_combout ),
	.sload(gnd),
	.ena(\state_cnt[0]~13_combout ),
	.q(\state_cnt[1]~q ),
	.prn(vcc));
defparam \state_cnt[1] .is_wysiwyg = "true";
defparam \state_cnt[1] .power_up = "low";

dffeas \sdft.BLOCK_DFT_I (
	.clk(clk),
	.d(\Selector13~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sdft.BLOCK_DFT_I~q ),
	.prn(vcc));
defparam \sdft.BLOCK_DFT_I .is_wysiwyg = "true";
defparam \sdft.BLOCK_DFT_I .power_up = "low";

dffeas \sdft.ENABLE_BFP_O (
	.clk(clk),
	.d(\Selector15~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sdft.ENABLE_BFP_O~q ),
	.prn(vcc));
defparam \sdft.ENABLE_BFP_O .is_wysiwyg = "true";
defparam \sdft.ENABLE_BFP_O .power_up = "low";

cycloneiii_lcell_comb \state_cnt[0]~6 (
	.dataa(\state_cnt[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\state_cnt[0]~6_combout ),
	.cout(\state_cnt[0]~7 ));
defparam \state_cnt[0]~6 .lut_mask = 16'h55AA;
defparam \state_cnt[0]~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \state_cnt[1]~8 (
	.dataa(\state_cnt[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\state_cnt[0]~7 ),
	.combout(\state_cnt[1]~8_combout ),
	.cout(\state_cnt[1]~9 ));
defparam \state_cnt[1]~8 .lut_mask = 16'h5A5F;
defparam \state_cnt[1]~8 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \state_cnt[2]~10 (
	.dataa(\state_cnt[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\state_cnt[1]~9 ),
	.combout(\state_cnt[2]~10_combout ),
	.cout(\state_cnt[2]~11 ));
defparam \state_cnt[2]~10 .lut_mask = 16'h5AAF;
defparam \state_cnt[2]~10 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \state_cnt[3]~14 (
	.dataa(\state_cnt[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\state_cnt[2]~11 ),
	.combout(\state_cnt[3]~14_combout ),
	.cout(\state_cnt[3]~15 ));
defparam \state_cnt[3]~14 .lut_mask = 16'h5A5F;
defparam \state_cnt[3]~14 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \state_cnt[4]~16 (
	.dataa(\state_cnt[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\state_cnt[3]~15 ),
	.combout(\state_cnt[4]~16_combout ),
	.cout(\state_cnt[4]~17 ));
defparam \state_cnt[4]~16 .lut_mask = 16'h5AAF;
defparam \state_cnt[4]~16 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \state_cnt[5]~18 (
	.dataa(\state_cnt[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\state_cnt[4]~17 ),
	.combout(\state_cnt[5]~18_combout ),
	.cout());
defparam \state_cnt[5]~18 .lut_mask = 16'h5A5A;
defparam \state_cnt[5]~18 .sum_lutc_input = "cin";

dffeas \reg_no_twiddle[0][0][3] (
	.clk(clk),
	.d(\reg_no_twiddle[0][0][3]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[0][0][3]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[0][0][3] .is_wysiwyg = "true";
defparam \reg_no_twiddle[0][0][3] .power_up = "low";

dffeas \reg_no_twiddle[0][0][7] (
	.clk(clk),
	.d(\reg_no_twiddle[0][0][7]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[0][0][7]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[0][0][7] .is_wysiwyg = "true";
defparam \reg_no_twiddle[0][0][7] .power_up = "low";

dffeas \reg_no_twiddle[0][1][7] (
	.clk(clk),
	.d(\reg_no_twiddle[0][1][7]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[0][1][7]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[0][1][7] .is_wysiwyg = "true";
defparam \reg_no_twiddle[0][1][7] .power_up = "low";

dffeas \reg_no_twiddle[0][1][3] (
	.clk(clk),
	.d(\reg_no_twiddle[0][1][3]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[0][1][3]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[0][1][3] .is_wysiwyg = "true";
defparam \reg_no_twiddle[0][1][3] .power_up = "low";

dffeas \reg_no_twiddle[0][0][4] (
	.clk(clk),
	.d(\reg_no_twiddle[0][0][4]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[0][0][4]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[0][0][4] .is_wysiwyg = "true";
defparam \reg_no_twiddle[0][0][4] .power_up = "low";

dffeas \reg_no_twiddle[0][1][4] (
	.clk(clk),
	.d(\reg_no_twiddle[0][1][4]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[0][1][4]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[0][1][4] .is_wysiwyg = "true";
defparam \reg_no_twiddle[0][1][4] .power_up = "low";

dffeas \reg_no_twiddle[0][0][5] (
	.clk(clk),
	.d(\reg_no_twiddle[0][0][5]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[0][0][5]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[0][0][5] .is_wysiwyg = "true";
defparam \reg_no_twiddle[0][0][5] .power_up = "low";

dffeas \reg_no_twiddle[0][1][5] (
	.clk(clk),
	.d(\reg_no_twiddle[0][1][5]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[0][1][5]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[0][1][5] .is_wysiwyg = "true";
defparam \reg_no_twiddle[0][1][5] .power_up = "low";

dffeas \reg_no_twiddle[0][0][6] (
	.clk(clk),
	.d(\reg_no_twiddle[0][0][6]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[0][0][6]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[0][0][6] .is_wysiwyg = "true";
defparam \reg_no_twiddle[0][0][6] .power_up = "low";

dffeas \reg_no_twiddle[0][1][6] (
	.clk(clk),
	.d(\reg_no_twiddle[0][1][6]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[0][1][6]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[0][1][6] .is_wysiwyg = "true";
defparam \reg_no_twiddle[0][1][6] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle[0][0][0]~1 (
	.dataa(\gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.datab(\reg_no_twiddle~60_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\reg_no_twiddle[0][0][0]~1_combout ),
	.cout(\reg_no_twiddle[0][0][0]~2 ));
defparam \reg_no_twiddle[0][0][0]~1 .lut_mask = 16'h66EE;
defparam \reg_no_twiddle[0][0][0]~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \reg_no_twiddle[0][0][1]~1 (
	.dataa(\gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\reg_no_twiddle[0][0][0]~2 ),
	.combout(\reg_no_twiddle[0][0][1]~1_combout ),
	.cout(\reg_no_twiddle[0][0][1]~2 ));
defparam \reg_no_twiddle[0][0][1]~1 .lut_mask = 16'h5A5F;
defparam \reg_no_twiddle[0][0][1]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \reg_no_twiddle[0][0][2]~1 (
	.dataa(\gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\reg_no_twiddle[0][0][1]~2 ),
	.combout(\reg_no_twiddle[0][0][2]~1_combout ),
	.cout(\reg_no_twiddle[0][0][2]~2 ));
defparam \reg_no_twiddle[0][0][2]~1 .lut_mask = 16'h5AAF;
defparam \reg_no_twiddle[0][0][2]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \reg_no_twiddle[0][0][3]~1 (
	.dataa(\gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\reg_no_twiddle[0][0][2]~2 ),
	.combout(\reg_no_twiddle[0][0][3]~1_combout ),
	.cout(\reg_no_twiddle[0][0][3]~2 ));
defparam \reg_no_twiddle[0][0][3]~1 .lut_mask = 16'h5A5F;
defparam \reg_no_twiddle[0][0][3]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \reg_no_twiddle[0][0][4]~1 (
	.dataa(\gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\reg_no_twiddle[0][0][3]~2 ),
	.combout(\reg_no_twiddle[0][0][4]~1_combout ),
	.cout(\reg_no_twiddle[0][0][4]~2 ));
defparam \reg_no_twiddle[0][0][4]~1 .lut_mask = 16'h5AAF;
defparam \reg_no_twiddle[0][0][4]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \reg_no_twiddle[0][0][5]~1 (
	.dataa(\gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\reg_no_twiddle[0][0][4]~2 ),
	.combout(\reg_no_twiddle[0][0][5]~1_combout ),
	.cout(\reg_no_twiddle[0][0][5]~2 ));
defparam \reg_no_twiddle[0][0][5]~1 .lut_mask = 16'h5A5F;
defparam \reg_no_twiddle[0][0][5]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \reg_no_twiddle[0][0][6]~1 (
	.dataa(\gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\reg_no_twiddle[0][0][5]~2 ),
	.combout(\reg_no_twiddle[0][0][6]~1_combout ),
	.cout(\reg_no_twiddle[0][0][6]~2 ));
defparam \reg_no_twiddle[0][0][6]~1 .lut_mask = 16'h5AAF;
defparam \reg_no_twiddle[0][0][6]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \reg_no_twiddle[0][0][7]~1 (
	.dataa(\gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\reg_no_twiddle[0][0][6]~2 ),
	.combout(\reg_no_twiddle[0][0][7]~1_combout ),
	.cout());
defparam \reg_no_twiddle[0][0][7]~1 .lut_mask = 16'h5A5A;
defparam \reg_no_twiddle[0][0][7]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \reg_no_twiddle[0][1][0]~1 (
	.dataa(\gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.datab(\reg_no_twiddle~61_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\reg_no_twiddle[0][1][0]~1_combout ),
	.cout(\reg_no_twiddle[0][1][0]~2 ));
defparam \reg_no_twiddle[0][1][0]~1 .lut_mask = 16'h66EE;
defparam \reg_no_twiddle[0][1][0]~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \reg_no_twiddle[0][1][1]~1 (
	.dataa(\gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\reg_no_twiddle[0][1][0]~2 ),
	.combout(\reg_no_twiddle[0][1][1]~1_combout ),
	.cout(\reg_no_twiddle[0][1][1]~2 ));
defparam \reg_no_twiddle[0][1][1]~1 .lut_mask = 16'h5A5F;
defparam \reg_no_twiddle[0][1][1]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \reg_no_twiddle[0][1][2]~1 (
	.dataa(\gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\reg_no_twiddle[0][1][1]~2 ),
	.combout(\reg_no_twiddle[0][1][2]~1_combout ),
	.cout(\reg_no_twiddle[0][1][2]~2 ));
defparam \reg_no_twiddle[0][1][2]~1 .lut_mask = 16'h5AAF;
defparam \reg_no_twiddle[0][1][2]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \reg_no_twiddle[0][1][3]~1 (
	.dataa(\gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\reg_no_twiddle[0][1][2]~2 ),
	.combout(\reg_no_twiddle[0][1][3]~1_combout ),
	.cout(\reg_no_twiddle[0][1][3]~2 ));
defparam \reg_no_twiddle[0][1][3]~1 .lut_mask = 16'h5A5F;
defparam \reg_no_twiddle[0][1][3]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \reg_no_twiddle[0][1][4]~1 (
	.dataa(\gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\reg_no_twiddle[0][1][3]~2 ),
	.combout(\reg_no_twiddle[0][1][4]~1_combout ),
	.cout(\reg_no_twiddle[0][1][4]~2 ));
defparam \reg_no_twiddle[0][1][4]~1 .lut_mask = 16'h5AAF;
defparam \reg_no_twiddle[0][1][4]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \reg_no_twiddle[0][1][5]~1 (
	.dataa(\gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\reg_no_twiddle[0][1][4]~2 ),
	.combout(\reg_no_twiddle[0][1][5]~1_combout ),
	.cout(\reg_no_twiddle[0][1][5]~2 ));
defparam \reg_no_twiddle[0][1][5]~1 .lut_mask = 16'h5A5F;
defparam \reg_no_twiddle[0][1][5]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \reg_no_twiddle[0][1][6]~1 (
	.dataa(\gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\reg_no_twiddle[0][1][5]~2 ),
	.combout(\reg_no_twiddle[0][1][6]~1_combout ),
	.cout(\reg_no_twiddle[0][1][6]~2 ));
defparam \reg_no_twiddle[0][1][6]~1 .lut_mask = 16'h5AAF;
defparam \reg_no_twiddle[0][1][6]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \reg_no_twiddle[0][1][7]~1 (
	.dataa(\gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\reg_no_twiddle[0][1][6]~2 ),
	.combout(\reg_no_twiddle[0][1][7]~1_combout ),
	.cout());
defparam \reg_no_twiddle[0][1][7]~1 .lut_mask = 16'h5A5A;
defparam \reg_no_twiddle[0][1][7]~1 .sum_lutc_input = "cin";

dffeas \butterfly_st2[0][0][6] (
	.clk(clk),
	.d(\butterfly_st2[0][0][6]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[0][0][6]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][0][6] .is_wysiwyg = "true";
defparam \butterfly_st2[0][0][6] .power_up = "low";

dffeas \butterfly_st2[0][0][5] (
	.clk(clk),
	.d(\butterfly_st2[0][0][5]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[0][0][5]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][0][5] .is_wysiwyg = "true";
defparam \butterfly_st2[0][0][5] .power_up = "low";

dffeas \butterfly_st2[0][0][4] (
	.clk(clk),
	.d(\butterfly_st2[0][0][4]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[0][0][4]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][0][4] .is_wysiwyg = "true";
defparam \butterfly_st2[0][0][4] .power_up = "low";

dffeas \butterfly_st2[0][0][3] (
	.clk(clk),
	.d(\butterfly_st2[0][0][3]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[0][0][3]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][0][3] .is_wysiwyg = "true";
defparam \butterfly_st2[0][0][3] .power_up = "low";

dffeas \butterfly_st2[0][0][2] (
	.clk(clk),
	.d(\butterfly_st2[0][0][2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[0][0][2]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][0][2] .is_wysiwyg = "true";
defparam \butterfly_st2[0][0][2] .power_up = "low";

dffeas \butterfly_st2[0][0][1] (
	.clk(clk),
	.d(\butterfly_st2[0][0][1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[0][0][1]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][0][1] .is_wysiwyg = "true";
defparam \butterfly_st2[0][0][1] .power_up = "low";

dffeas \butterfly_st2[0][0][0] (
	.clk(clk),
	.d(\butterfly_st2[0][0][0]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[0][0][0]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][0][0] .is_wysiwyg = "true";
defparam \butterfly_st2[0][0][0] .power_up = "low";

dffeas \butterfly_st2[0][0][9] (
	.clk(clk),
	.d(\butterfly_st2[0][0][9]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[0][0][9]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][0][9] .is_wysiwyg = "true";
defparam \butterfly_st2[0][0][9] .power_up = "low";

dffeas \butterfly_st2[0][0][8] (
	.clk(clk),
	.d(\butterfly_st2[0][0][8]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[0][0][8]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][0][8] .is_wysiwyg = "true";
defparam \butterfly_st2[0][0][8] .power_up = "low";

dffeas \butterfly_st2[0][0][7] (
	.clk(clk),
	.d(\butterfly_st2[0][0][7]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[0][0][7]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][0][7] .is_wysiwyg = "true";
defparam \butterfly_st2[0][0][7] .power_up = "low";

dffeas \butterfly_st2[0][1][9] (
	.clk(clk),
	.d(\butterfly_st2[0][1][9]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[0][1][9]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][1][9] .is_wysiwyg = "true";
defparam \butterfly_st2[0][1][9] .power_up = "low";

dffeas \butterfly_st2[0][1][8] (
	.clk(clk),
	.d(\butterfly_st2[0][1][8]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[0][1][8]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][1][8] .is_wysiwyg = "true";
defparam \butterfly_st2[0][1][8] .power_up = "low";

dffeas \butterfly_st2[0][1][7] (
	.clk(clk),
	.d(\butterfly_st2[0][1][7]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[0][1][7]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][1][7] .is_wysiwyg = "true";
defparam \butterfly_st2[0][1][7] .power_up = "low";

dffeas \butterfly_st2[0][1][6] (
	.clk(clk),
	.d(\butterfly_st2[0][1][6]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[0][1][6]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][1][6] .is_wysiwyg = "true";
defparam \butterfly_st2[0][1][6] .power_up = "low";

dffeas \butterfly_st2[0][1][5] (
	.clk(clk),
	.d(\butterfly_st2[0][1][5]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[0][1][5]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][1][5] .is_wysiwyg = "true";
defparam \butterfly_st2[0][1][5] .power_up = "low";

dffeas \butterfly_st2[0][1][4] (
	.clk(clk),
	.d(\butterfly_st2[0][1][4]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[0][1][4]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][1][4] .is_wysiwyg = "true";
defparam \butterfly_st2[0][1][4] .power_up = "low";

dffeas \butterfly_st2[0][1][3] (
	.clk(clk),
	.d(\butterfly_st2[0][1][3]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[0][1][3]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][1][3] .is_wysiwyg = "true";
defparam \butterfly_st2[0][1][3] .power_up = "low";

dffeas \butterfly_st2[0][1][2] (
	.clk(clk),
	.d(\butterfly_st2[0][1][2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[0][1][2]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][1][2] .is_wysiwyg = "true";
defparam \butterfly_st2[0][1][2] .power_up = "low";

dffeas \butterfly_st2[0][1][1] (
	.clk(clk),
	.d(\butterfly_st2[0][1][1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[0][1][1]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][1][1] .is_wysiwyg = "true";
defparam \butterfly_st2[0][1][1] .power_up = "low";

dffeas \butterfly_st2[0][1][0] (
	.clk(clk),
	.d(\butterfly_st2[0][1][0]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[0][1][0]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][1][0] .is_wysiwyg = "true";
defparam \butterfly_st2[0][1][0] .power_up = "low";

dffeas \butterfly_st2[1][1][2] (
	.clk(clk),
	.d(\butterfly_st2[1][1][2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[1][1][2]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][1][2] .is_wysiwyg = "true";
defparam \butterfly_st2[1][1][2] .power_up = "low";

dffeas \butterfly_st2[1][1][1] (
	.clk(clk),
	.d(\butterfly_st2[1][1][1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[1][1][1]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][1][1] .is_wysiwyg = "true";
defparam \butterfly_st2[1][1][1] .power_up = "low";

dffeas \butterfly_st2[1][1][0] (
	.clk(clk),
	.d(\butterfly_st2[1][1][0]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[1][1][0]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][1][0] .is_wysiwyg = "true";
defparam \butterfly_st2[1][1][0] .power_up = "low";

dffeas \butterfly_st2[1][1][9] (
	.clk(clk),
	.d(\butterfly_st2[1][1][9]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[1][1][9]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][1][9] .is_wysiwyg = "true";
defparam \butterfly_st2[1][1][9] .power_up = "low";

dffeas \butterfly_st2[1][1][3] (
	.clk(clk),
	.d(\butterfly_st2[1][1][3]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[1][1][3]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][1][3] .is_wysiwyg = "true";
defparam \butterfly_st2[1][1][3] .power_up = "low";

dffeas \butterfly_st2[1][1][4] (
	.clk(clk),
	.d(\butterfly_st2[1][1][4]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[1][1][4]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][1][4] .is_wysiwyg = "true";
defparam \butterfly_st2[1][1][4] .power_up = "low";

dffeas \butterfly_st2[1][1][5] (
	.clk(clk),
	.d(\butterfly_st2[1][1][5]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[1][1][5]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][1][5] .is_wysiwyg = "true";
defparam \butterfly_st2[1][1][5] .power_up = "low";

dffeas \butterfly_st2[1][1][6] (
	.clk(clk),
	.d(\butterfly_st2[1][1][6]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[1][1][6]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][1][6] .is_wysiwyg = "true";
defparam \butterfly_st2[1][1][6] .power_up = "low";

dffeas \butterfly_st2[1][1][7] (
	.clk(clk),
	.d(\butterfly_st2[1][1][7]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[1][1][7]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][1][7] .is_wysiwyg = "true";
defparam \butterfly_st2[1][1][7] .power_up = "low";

dffeas \butterfly_st2[1][1][8] (
	.clk(clk),
	.d(\butterfly_st2[1][1][8]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[1][1][8]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][1][8] .is_wysiwyg = "true";
defparam \butterfly_st2[1][1][8] .power_up = "low";

dffeas \butterfly_st2[1][0][2] (
	.clk(clk),
	.d(\butterfly_st2[1][0][2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[1][0][2]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][0][2] .is_wysiwyg = "true";
defparam \butterfly_st2[1][0][2] .power_up = "low";

dffeas \butterfly_st2[1][0][1] (
	.clk(clk),
	.d(\butterfly_st2[1][0][1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[1][0][1]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][0][1] .is_wysiwyg = "true";
defparam \butterfly_st2[1][0][1] .power_up = "low";

dffeas \butterfly_st2[1][0][0] (
	.clk(clk),
	.d(\butterfly_st2[1][0][0]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[1][0][0]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][0][0] .is_wysiwyg = "true";
defparam \butterfly_st2[1][0][0] .power_up = "low";

dffeas \butterfly_st2[1][0][9] (
	.clk(clk),
	.d(\butterfly_st2[1][0][9]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[1][0][9]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][0][9] .is_wysiwyg = "true";
defparam \butterfly_st2[1][0][9] .power_up = "low";

dffeas \butterfly_st2[1][0][3] (
	.clk(clk),
	.d(\butterfly_st2[1][0][3]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[1][0][3]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][0][3] .is_wysiwyg = "true";
defparam \butterfly_st2[1][0][3] .power_up = "low";

dffeas \butterfly_st2[1][0][4] (
	.clk(clk),
	.d(\butterfly_st2[1][0][4]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[1][0][4]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][0][4] .is_wysiwyg = "true";
defparam \butterfly_st2[1][0][4] .power_up = "low";

dffeas \butterfly_st2[1][0][5] (
	.clk(clk),
	.d(\butterfly_st2[1][0][5]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[1][0][5]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][0][5] .is_wysiwyg = "true";
defparam \butterfly_st2[1][0][5] .power_up = "low";

dffeas \butterfly_st2[1][0][6] (
	.clk(clk),
	.d(\butterfly_st2[1][0][6]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[1][0][6]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][0][6] .is_wysiwyg = "true";
defparam \butterfly_st2[1][0][6] .power_up = "low";

dffeas \butterfly_st2[1][0][7] (
	.clk(clk),
	.d(\butterfly_st2[1][0][7]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[1][0][7]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][0][7] .is_wysiwyg = "true";
defparam \butterfly_st2[1][0][7] .power_up = "low";

dffeas \butterfly_st2[1][0][8] (
	.clk(clk),
	.d(\butterfly_st2[1][0][8]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[1][0][8]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][0][8] .is_wysiwyg = "true";
defparam \butterfly_st2[1][0][8] .power_up = "low";

dffeas \butterfly_st2[2][1][2] (
	.clk(clk),
	.d(\butterfly_st2[2][1][2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[2][1][2]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][1][2] .is_wysiwyg = "true";
defparam \butterfly_st2[2][1][2] .power_up = "low";

dffeas \butterfly_st2[2][1][1] (
	.clk(clk),
	.d(\butterfly_st2[2][1][1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[2][1][1]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][1][1] .is_wysiwyg = "true";
defparam \butterfly_st2[2][1][1] .power_up = "low";

dffeas \butterfly_st2[2][1][0] (
	.clk(clk),
	.d(\butterfly_st2[2][1][0]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[2][1][0]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][1][0] .is_wysiwyg = "true";
defparam \butterfly_st2[2][1][0] .power_up = "low";

dffeas \butterfly_st2[2][1][9] (
	.clk(clk),
	.d(\butterfly_st2[2][1][9]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[2][1][9]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][1][9] .is_wysiwyg = "true";
defparam \butterfly_st2[2][1][9] .power_up = "low";

dffeas \butterfly_st2[2][1][3] (
	.clk(clk),
	.d(\butterfly_st2[2][1][3]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[2][1][3]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][1][3] .is_wysiwyg = "true";
defparam \butterfly_st2[2][1][3] .power_up = "low";

dffeas \butterfly_st2[2][1][4] (
	.clk(clk),
	.d(\butterfly_st2[2][1][4]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[2][1][4]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][1][4] .is_wysiwyg = "true";
defparam \butterfly_st2[2][1][4] .power_up = "low";

dffeas \butterfly_st2[2][1][5] (
	.clk(clk),
	.d(\butterfly_st2[2][1][5]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[2][1][5]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][1][5] .is_wysiwyg = "true";
defparam \butterfly_st2[2][1][5] .power_up = "low";

dffeas \butterfly_st2[2][1][6] (
	.clk(clk),
	.d(\butterfly_st2[2][1][6]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[2][1][6]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][1][6] .is_wysiwyg = "true";
defparam \butterfly_st2[2][1][6] .power_up = "low";

dffeas \butterfly_st2[2][1][7] (
	.clk(clk),
	.d(\butterfly_st2[2][1][7]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[2][1][7]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][1][7] .is_wysiwyg = "true";
defparam \butterfly_st2[2][1][7] .power_up = "low";

dffeas \butterfly_st2[2][1][8] (
	.clk(clk),
	.d(\butterfly_st2[2][1][8]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[2][1][8]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][1][8] .is_wysiwyg = "true";
defparam \butterfly_st2[2][1][8] .power_up = "low";

dffeas \butterfly_st2[2][0][2] (
	.clk(clk),
	.d(\butterfly_st2[2][0][2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[2][0][2]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][0][2] .is_wysiwyg = "true";
defparam \butterfly_st2[2][0][2] .power_up = "low";

dffeas \butterfly_st2[2][0][1] (
	.clk(clk),
	.d(\butterfly_st2[2][0][1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[2][0][1]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][0][1] .is_wysiwyg = "true";
defparam \butterfly_st2[2][0][1] .power_up = "low";

dffeas \butterfly_st2[2][0][0] (
	.clk(clk),
	.d(\butterfly_st2[2][0][0]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[2][0][0]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][0][0] .is_wysiwyg = "true";
defparam \butterfly_st2[2][0][0] .power_up = "low";

dffeas \butterfly_st2[2][0][9] (
	.clk(clk),
	.d(\butterfly_st2[2][0][9]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[2][0][9]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][0][9] .is_wysiwyg = "true";
defparam \butterfly_st2[2][0][9] .power_up = "low";

dffeas \butterfly_st2[2][0][3] (
	.clk(clk),
	.d(\butterfly_st2[2][0][3]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[2][0][3]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][0][3] .is_wysiwyg = "true";
defparam \butterfly_st2[2][0][3] .power_up = "low";

dffeas \butterfly_st2[2][0][4] (
	.clk(clk),
	.d(\butterfly_st2[2][0][4]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[2][0][4]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][0][4] .is_wysiwyg = "true";
defparam \butterfly_st2[2][0][4] .power_up = "low";

dffeas \butterfly_st2[2][0][5] (
	.clk(clk),
	.d(\butterfly_st2[2][0][5]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[2][0][5]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][0][5] .is_wysiwyg = "true";
defparam \butterfly_st2[2][0][5] .power_up = "low";

dffeas \butterfly_st2[2][0][6] (
	.clk(clk),
	.d(\butterfly_st2[2][0][6]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[2][0][6]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][0][6] .is_wysiwyg = "true";
defparam \butterfly_st2[2][0][6] .power_up = "low";

dffeas \butterfly_st2[2][0][7] (
	.clk(clk),
	.d(\butterfly_st2[2][0][7]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[2][0][7]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][0][7] .is_wysiwyg = "true";
defparam \butterfly_st2[2][0][7] .power_up = "low";

dffeas \butterfly_st2[2][0][8] (
	.clk(clk),
	.d(\butterfly_st2[2][0][8]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[2][0][8]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][0][8] .is_wysiwyg = "true";
defparam \butterfly_st2[2][0][8] .power_up = "low";

dffeas \butterfly_st2[3][1][2] (
	.clk(clk),
	.d(\butterfly_st2[3][1][2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[3][1][2]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][1][2] .is_wysiwyg = "true";
defparam \butterfly_st2[3][1][2] .power_up = "low";

dffeas \butterfly_st2[3][1][1] (
	.clk(clk),
	.d(\butterfly_st2[3][1][1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[3][1][1]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][1][1] .is_wysiwyg = "true";
defparam \butterfly_st2[3][1][1] .power_up = "low";

dffeas \butterfly_st2[3][1][0] (
	.clk(clk),
	.d(\butterfly_st2[3][1][0]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[3][1][0]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][1][0] .is_wysiwyg = "true";
defparam \butterfly_st2[3][1][0] .power_up = "low";

dffeas \butterfly_st2[3][1][9] (
	.clk(clk),
	.d(\butterfly_st2[3][1][9]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[3][1][9]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][1][9] .is_wysiwyg = "true";
defparam \butterfly_st2[3][1][9] .power_up = "low";

dffeas \butterfly_st2[3][1][3] (
	.clk(clk),
	.d(\butterfly_st2[3][1][3]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[3][1][3]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][1][3] .is_wysiwyg = "true";
defparam \butterfly_st2[3][1][3] .power_up = "low";

dffeas \butterfly_st2[3][1][4] (
	.clk(clk),
	.d(\butterfly_st2[3][1][4]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[3][1][4]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][1][4] .is_wysiwyg = "true";
defparam \butterfly_st2[3][1][4] .power_up = "low";

dffeas \butterfly_st2[3][1][5] (
	.clk(clk),
	.d(\butterfly_st2[3][1][5]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[3][1][5]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][1][5] .is_wysiwyg = "true";
defparam \butterfly_st2[3][1][5] .power_up = "low";

dffeas \butterfly_st2[3][1][6] (
	.clk(clk),
	.d(\butterfly_st2[3][1][6]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[3][1][6]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][1][6] .is_wysiwyg = "true";
defparam \butterfly_st2[3][1][6] .power_up = "low";

dffeas \butterfly_st2[3][1][7] (
	.clk(clk),
	.d(\butterfly_st2[3][1][7]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[3][1][7]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][1][7] .is_wysiwyg = "true";
defparam \butterfly_st2[3][1][7] .power_up = "low";

dffeas \butterfly_st2[3][1][8] (
	.clk(clk),
	.d(\butterfly_st2[3][1][8]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[3][1][8]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][1][8] .is_wysiwyg = "true";
defparam \butterfly_st2[3][1][8] .power_up = "low";

dffeas \butterfly_st2[3][0][2] (
	.clk(clk),
	.d(\butterfly_st2[3][0][2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[3][0][2]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][0][2] .is_wysiwyg = "true";
defparam \butterfly_st2[3][0][2] .power_up = "low";

dffeas \butterfly_st2[3][0][1] (
	.clk(clk),
	.d(\butterfly_st2[3][0][1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[3][0][1]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][0][1] .is_wysiwyg = "true";
defparam \butterfly_st2[3][0][1] .power_up = "low";

dffeas \butterfly_st2[3][0][0] (
	.clk(clk),
	.d(\butterfly_st2[3][0][0]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[3][0][0]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][0][0] .is_wysiwyg = "true";
defparam \butterfly_st2[3][0][0] .power_up = "low";

dffeas \butterfly_st2[3][0][9] (
	.clk(clk),
	.d(\butterfly_st2[3][0][9]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[3][0][9]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][0][9] .is_wysiwyg = "true";
defparam \butterfly_st2[3][0][9] .power_up = "low";

dffeas \butterfly_st2[3][0][3] (
	.clk(clk),
	.d(\butterfly_st2[3][0][3]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[3][0][3]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][0][3] .is_wysiwyg = "true";
defparam \butterfly_st2[3][0][3] .power_up = "low";

dffeas \butterfly_st2[3][0][4] (
	.clk(clk),
	.d(\butterfly_st2[3][0][4]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[3][0][4]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][0][4] .is_wysiwyg = "true";
defparam \butterfly_st2[3][0][4] .power_up = "low";

dffeas \butterfly_st2[3][0][5] (
	.clk(clk),
	.d(\butterfly_st2[3][0][5]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[3][0][5]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][0][5] .is_wysiwyg = "true";
defparam \butterfly_st2[3][0][5] .power_up = "low";

dffeas \butterfly_st2[3][0][6] (
	.clk(clk),
	.d(\butterfly_st2[3][0][6]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[3][0][6]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][0][6] .is_wysiwyg = "true";
defparam \butterfly_st2[3][0][6] .power_up = "low";

dffeas \butterfly_st2[3][0][7] (
	.clk(clk),
	.d(\butterfly_st2[3][0][7]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[3][0][7]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][0][7] .is_wysiwyg = "true";
defparam \butterfly_st2[3][0][7] .power_up = "low";

dffeas \butterfly_st2[3][0][8] (
	.clk(clk),
	.d(\butterfly_st2[3][0][8]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[3][0][8]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][0][8] .is_wysiwyg = "true";
defparam \butterfly_st2[3][0][8] .power_up = "low";

dffeas \butterfly_st1[0][0][6] (
	.clk(clk),
	.d(\butterfly_st1[0][0][6]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[0][0][6]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][0][6] .is_wysiwyg = "true";
defparam \butterfly_st1[0][0][6] .power_up = "low";

dffeas \butterfly_st1[1][0][6] (
	.clk(clk),
	.d(\butterfly_st1[1][0][6]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[1][0][6]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][0][6] .is_wysiwyg = "true";
defparam \butterfly_st1[1][0][6] .power_up = "low";

dffeas \butterfly_st1[0][0][5] (
	.clk(clk),
	.d(\butterfly_st1[0][0][5]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[0][0][5]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][0][5] .is_wysiwyg = "true";
defparam \butterfly_st1[0][0][5] .power_up = "low";

dffeas \butterfly_st1[1][0][5] (
	.clk(clk),
	.d(\butterfly_st1[1][0][5]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[1][0][5]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][0][5] .is_wysiwyg = "true";
defparam \butterfly_st1[1][0][5] .power_up = "low";

dffeas \butterfly_st1[0][0][4] (
	.clk(clk),
	.d(\butterfly_st1[0][0][4]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[0][0][4]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][0][4] .is_wysiwyg = "true";
defparam \butterfly_st1[0][0][4] .power_up = "low";

dffeas \butterfly_st1[1][0][4] (
	.clk(clk),
	.d(\butterfly_st1[1][0][4]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[1][0][4]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][0][4] .is_wysiwyg = "true";
defparam \butterfly_st1[1][0][4] .power_up = "low";

dffeas \butterfly_st1[0][0][3] (
	.clk(clk),
	.d(\butterfly_st1[0][0][3]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[0][0][3]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][0][3] .is_wysiwyg = "true";
defparam \butterfly_st1[0][0][3] .power_up = "low";

dffeas \butterfly_st1[1][0][3] (
	.clk(clk),
	.d(\butterfly_st1[1][0][3]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[1][0][3]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][0][3] .is_wysiwyg = "true";
defparam \butterfly_st1[1][0][3] .power_up = "low";

dffeas \butterfly_st1[0][0][2] (
	.clk(clk),
	.d(\butterfly_st1[0][0][2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[0][0][2]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][0][2] .is_wysiwyg = "true";
defparam \butterfly_st1[0][0][2] .power_up = "low";

dffeas \butterfly_st1[1][0][2] (
	.clk(clk),
	.d(\butterfly_st1[1][0][2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[1][0][2]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][0][2] .is_wysiwyg = "true";
defparam \butterfly_st1[1][0][2] .power_up = "low";

dffeas \butterfly_st1[0][0][1] (
	.clk(clk),
	.d(\butterfly_st1[0][0][1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[0][0][1]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][0][1] .is_wysiwyg = "true";
defparam \butterfly_st1[0][0][1] .power_up = "low";

dffeas \butterfly_st1[1][0][1] (
	.clk(clk),
	.d(\butterfly_st1[1][0][1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[1][0][1]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][0][1] .is_wysiwyg = "true";
defparam \butterfly_st1[1][0][1] .power_up = "low";

dffeas \butterfly_st1[0][0][0] (
	.clk(clk),
	.d(\butterfly_st1[0][0][0]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[0][0][0]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][0][0] .is_wysiwyg = "true";
defparam \butterfly_st1[0][0][0] .power_up = "low";

dffeas \butterfly_st1[1][0][0] (
	.clk(clk),
	.d(\butterfly_st1[1][0][0]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[1][0][0]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][0][0] .is_wysiwyg = "true";
defparam \butterfly_st1[1][0][0] .power_up = "low";

cycloneiii_lcell_comb \butterfly_st2[0][0][0]~1 (
	.dataa(\butterfly_st1[0][0][0]~q ),
	.datab(\butterfly_st1[1][0][0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\butterfly_st2[0][0][0]~1_combout ),
	.cout(\butterfly_st2[0][0][0]~2 ));
defparam \butterfly_st2[0][0][0]~1 .lut_mask = 16'h66EE;
defparam \butterfly_st2[0][0][0]~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \butterfly_st2[0][0][1]~1 (
	.dataa(\butterfly_st1[0][0][1]~q ),
	.datab(\butterfly_st1[1][0][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[0][0][0]~2 ),
	.combout(\butterfly_st2[0][0][1]~1_combout ),
	.cout(\butterfly_st2[0][0][1]~2 ));
defparam \butterfly_st2[0][0][1]~1 .lut_mask = 16'h967F;
defparam \butterfly_st2[0][0][1]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[0][0][2]~1 (
	.dataa(\butterfly_st1[0][0][2]~q ),
	.datab(\butterfly_st1[1][0][2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[0][0][1]~2 ),
	.combout(\butterfly_st2[0][0][2]~1_combout ),
	.cout(\butterfly_st2[0][0][2]~2 ));
defparam \butterfly_st2[0][0][2]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st2[0][0][2]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[0][0][3]~1 (
	.dataa(\butterfly_st1[0][0][3]~q ),
	.datab(\butterfly_st1[1][0][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[0][0][2]~2 ),
	.combout(\butterfly_st2[0][0][3]~1_combout ),
	.cout(\butterfly_st2[0][0][3]~2 ));
defparam \butterfly_st2[0][0][3]~1 .lut_mask = 16'h967F;
defparam \butterfly_st2[0][0][3]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[0][0][4]~1 (
	.dataa(\butterfly_st1[0][0][4]~q ),
	.datab(\butterfly_st1[1][0][4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[0][0][3]~2 ),
	.combout(\butterfly_st2[0][0][4]~1_combout ),
	.cout(\butterfly_st2[0][0][4]~2 ));
defparam \butterfly_st2[0][0][4]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st2[0][0][4]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[0][0][5]~1 (
	.dataa(\butterfly_st1[0][0][5]~q ),
	.datab(\butterfly_st1[1][0][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[0][0][4]~2 ),
	.combout(\butterfly_st2[0][0][5]~1_combout ),
	.cout(\butterfly_st2[0][0][5]~2 ));
defparam \butterfly_st2[0][0][5]~1 .lut_mask = 16'h967F;
defparam \butterfly_st2[0][0][5]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[0][0][6]~1 (
	.dataa(\butterfly_st1[0][0][6]~q ),
	.datab(\butterfly_st1[1][0][6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[0][0][5]~2 ),
	.combout(\butterfly_st2[0][0][6]~1_combout ),
	.cout(\butterfly_st2[0][0][6]~2 ));
defparam \butterfly_st2[0][0][6]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st2[0][0][6]~1 .sum_lutc_input = "cin";

dffeas \butterfly_st1[0][0][8] (
	.clk(clk),
	.d(\butterfly_st1[0][0][8]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[0][0][8]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][0][8] .is_wysiwyg = "true";
defparam \butterfly_st1[0][0][8] .power_up = "low";

dffeas \butterfly_st1[1][0][8] (
	.clk(clk),
	.d(\butterfly_st1[1][0][8]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[1][0][8]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][0][8] .is_wysiwyg = "true";
defparam \butterfly_st1[1][0][8] .power_up = "low";

dffeas \butterfly_st1[0][0][7] (
	.clk(clk),
	.d(\butterfly_st1[0][0][7]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[0][0][7]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][0][7] .is_wysiwyg = "true";
defparam \butterfly_st1[0][0][7] .power_up = "low";

dffeas \butterfly_st1[1][0][7] (
	.clk(clk),
	.d(\butterfly_st1[1][0][7]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[1][0][7]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][0][7] .is_wysiwyg = "true";
defparam \butterfly_st1[1][0][7] .power_up = "low";

cycloneiii_lcell_comb \butterfly_st2[0][0][7]~1 (
	.dataa(\butterfly_st1[0][0][7]~q ),
	.datab(\butterfly_st1[1][0][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[0][0][6]~2 ),
	.combout(\butterfly_st2[0][0][7]~1_combout ),
	.cout(\butterfly_st2[0][0][7]~2 ));
defparam \butterfly_st2[0][0][7]~1 .lut_mask = 16'h967F;
defparam \butterfly_st2[0][0][7]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[0][0][8]~1 (
	.dataa(\butterfly_st1[0][0][8]~q ),
	.datab(\butterfly_st1[1][0][8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[0][0][7]~2 ),
	.combout(\butterfly_st2[0][0][8]~1_combout ),
	.cout(\butterfly_st2[0][0][8]~2 ));
defparam \butterfly_st2[0][0][8]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st2[0][0][8]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[0][0][9]~1 (
	.dataa(\butterfly_st1[0][0][8]~q ),
	.datab(\butterfly_st1[1][0][8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\butterfly_st2[0][0][8]~2 ),
	.combout(\butterfly_st2[0][0][9]~1_combout ),
	.cout());
defparam \butterfly_st2[0][0][9]~1 .lut_mask = 16'h9696;
defparam \butterfly_st2[0][0][9]~1 .sum_lutc_input = "cin";

dffeas \butterfly_st1[0][1][8] (
	.clk(clk),
	.d(\butterfly_st1[0][1][8]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[0][1][8]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][1][8] .is_wysiwyg = "true";
defparam \butterfly_st1[0][1][8] .power_up = "low";

dffeas \butterfly_st1[1][1][8] (
	.clk(clk),
	.d(\butterfly_st1[1][1][8]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[1][1][8]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][1][8] .is_wysiwyg = "true";
defparam \butterfly_st1[1][1][8] .power_up = "low";

dffeas \butterfly_st1[0][1][7] (
	.clk(clk),
	.d(\butterfly_st1[0][1][7]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[0][1][7]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][1][7] .is_wysiwyg = "true";
defparam \butterfly_st1[0][1][7] .power_up = "low";

dffeas \butterfly_st1[1][1][7] (
	.clk(clk),
	.d(\butterfly_st1[1][1][7]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[1][1][7]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][1][7] .is_wysiwyg = "true";
defparam \butterfly_st1[1][1][7] .power_up = "low";

dffeas \butterfly_st1[0][1][6] (
	.clk(clk),
	.d(\butterfly_st1[0][1][6]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[0][1][6]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][1][6] .is_wysiwyg = "true";
defparam \butterfly_st1[0][1][6] .power_up = "low";

dffeas \butterfly_st1[1][1][6] (
	.clk(clk),
	.d(\butterfly_st1[1][1][6]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[1][1][6]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][1][6] .is_wysiwyg = "true";
defparam \butterfly_st1[1][1][6] .power_up = "low";

dffeas \butterfly_st1[0][1][5] (
	.clk(clk),
	.d(\butterfly_st1[0][1][5]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[0][1][5]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][1][5] .is_wysiwyg = "true";
defparam \butterfly_st1[0][1][5] .power_up = "low";

dffeas \butterfly_st1[1][1][5] (
	.clk(clk),
	.d(\butterfly_st1[1][1][5]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[1][1][5]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][1][5] .is_wysiwyg = "true";
defparam \butterfly_st1[1][1][5] .power_up = "low";

dffeas \butterfly_st1[0][1][4] (
	.clk(clk),
	.d(\butterfly_st1[0][1][4]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[0][1][4]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][1][4] .is_wysiwyg = "true";
defparam \butterfly_st1[0][1][4] .power_up = "low";

dffeas \butterfly_st1[1][1][4] (
	.clk(clk),
	.d(\butterfly_st1[1][1][4]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[1][1][4]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][1][4] .is_wysiwyg = "true";
defparam \butterfly_st1[1][1][4] .power_up = "low";

dffeas \butterfly_st1[0][1][3] (
	.clk(clk),
	.d(\butterfly_st1[0][1][3]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[0][1][3]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][1][3] .is_wysiwyg = "true";
defparam \butterfly_st1[0][1][3] .power_up = "low";

dffeas \butterfly_st1[1][1][3] (
	.clk(clk),
	.d(\butterfly_st1[1][1][3]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[1][1][3]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][1][3] .is_wysiwyg = "true";
defparam \butterfly_st1[1][1][3] .power_up = "low";

dffeas \butterfly_st1[0][1][2] (
	.clk(clk),
	.d(\butterfly_st1[0][1][2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[0][1][2]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][1][2] .is_wysiwyg = "true";
defparam \butterfly_st1[0][1][2] .power_up = "low";

dffeas \butterfly_st1[1][1][2] (
	.clk(clk),
	.d(\butterfly_st1[1][1][2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[1][1][2]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][1][2] .is_wysiwyg = "true";
defparam \butterfly_st1[1][1][2] .power_up = "low";

dffeas \butterfly_st1[0][1][1] (
	.clk(clk),
	.d(\butterfly_st1[0][1][1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[0][1][1]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][1][1] .is_wysiwyg = "true";
defparam \butterfly_st1[0][1][1] .power_up = "low";

dffeas \butterfly_st1[1][1][1] (
	.clk(clk),
	.d(\butterfly_st1[1][1][1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[1][1][1]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][1][1] .is_wysiwyg = "true";
defparam \butterfly_st1[1][1][1] .power_up = "low";

dffeas \butterfly_st1[0][1][0] (
	.clk(clk),
	.d(\butterfly_st1[0][1][0]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[0][1][0]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][1][0] .is_wysiwyg = "true";
defparam \butterfly_st1[0][1][0] .power_up = "low";

dffeas \butterfly_st1[1][1][0] (
	.clk(clk),
	.d(\butterfly_st1[1][1][0]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[1][1][0]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][1][0] .is_wysiwyg = "true";
defparam \butterfly_st1[1][1][0] .power_up = "low";

cycloneiii_lcell_comb \butterfly_st2[0][1][0]~1 (
	.dataa(\butterfly_st1[0][1][0]~q ),
	.datab(\butterfly_st1[1][1][0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\butterfly_st2[0][1][0]~1_combout ),
	.cout(\butterfly_st2[0][1][0]~2 ));
defparam \butterfly_st2[0][1][0]~1 .lut_mask = 16'h66EE;
defparam \butterfly_st2[0][1][0]~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \butterfly_st2[0][1][1]~1 (
	.dataa(\butterfly_st1[0][1][1]~q ),
	.datab(\butterfly_st1[1][1][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[0][1][0]~2 ),
	.combout(\butterfly_st2[0][1][1]~1_combout ),
	.cout(\butterfly_st2[0][1][1]~2 ));
defparam \butterfly_st2[0][1][1]~1 .lut_mask = 16'h967F;
defparam \butterfly_st2[0][1][1]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[0][1][2]~1 (
	.dataa(\butterfly_st1[0][1][2]~q ),
	.datab(\butterfly_st1[1][1][2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[0][1][1]~2 ),
	.combout(\butterfly_st2[0][1][2]~1_combout ),
	.cout(\butterfly_st2[0][1][2]~2 ));
defparam \butterfly_st2[0][1][2]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st2[0][1][2]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[0][1][3]~1 (
	.dataa(\butterfly_st1[0][1][3]~q ),
	.datab(\butterfly_st1[1][1][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[0][1][2]~2 ),
	.combout(\butterfly_st2[0][1][3]~1_combout ),
	.cout(\butterfly_st2[0][1][3]~2 ));
defparam \butterfly_st2[0][1][3]~1 .lut_mask = 16'h967F;
defparam \butterfly_st2[0][1][3]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[0][1][4]~1 (
	.dataa(\butterfly_st1[0][1][4]~q ),
	.datab(\butterfly_st1[1][1][4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[0][1][3]~2 ),
	.combout(\butterfly_st2[0][1][4]~1_combout ),
	.cout(\butterfly_st2[0][1][4]~2 ));
defparam \butterfly_st2[0][1][4]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st2[0][1][4]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[0][1][5]~1 (
	.dataa(\butterfly_st1[0][1][5]~q ),
	.datab(\butterfly_st1[1][1][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[0][1][4]~2 ),
	.combout(\butterfly_st2[0][1][5]~1_combout ),
	.cout(\butterfly_st2[0][1][5]~2 ));
defparam \butterfly_st2[0][1][5]~1 .lut_mask = 16'h967F;
defparam \butterfly_st2[0][1][5]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[0][1][6]~1 (
	.dataa(\butterfly_st1[0][1][6]~q ),
	.datab(\butterfly_st1[1][1][6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[0][1][5]~2 ),
	.combout(\butterfly_st2[0][1][6]~1_combout ),
	.cout(\butterfly_st2[0][1][6]~2 ));
defparam \butterfly_st2[0][1][6]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st2[0][1][6]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[0][1][7]~1 (
	.dataa(\butterfly_st1[0][1][7]~q ),
	.datab(\butterfly_st1[1][1][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[0][1][6]~2 ),
	.combout(\butterfly_st2[0][1][7]~1_combout ),
	.cout(\butterfly_st2[0][1][7]~2 ));
defparam \butterfly_st2[0][1][7]~1 .lut_mask = 16'h967F;
defparam \butterfly_st2[0][1][7]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[0][1][8]~1 (
	.dataa(\butterfly_st1[0][1][8]~q ),
	.datab(\butterfly_st1[1][1][8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[0][1][7]~2 ),
	.combout(\butterfly_st2[0][1][8]~1_combout ),
	.cout(\butterfly_st2[0][1][8]~2 ));
defparam \butterfly_st2[0][1][8]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st2[0][1][8]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[0][1][9]~1 (
	.dataa(\butterfly_st1[0][1][8]~q ),
	.datab(\butterfly_st1[1][1][8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\butterfly_st2[0][1][8]~2 ),
	.combout(\butterfly_st2[0][1][9]~1_combout ),
	.cout());
defparam \butterfly_st2[0][1][9]~1 .lut_mask = 16'h9696;
defparam \butterfly_st2[0][1][9]~1 .sum_lutc_input = "cin";

dffeas \butterfly_st1[2][1][2] (
	.clk(clk),
	.d(\butterfly_st1[2][1][2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[2][1][2]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][1][2] .is_wysiwyg = "true";
defparam \butterfly_st1[2][1][2] .power_up = "low";

dffeas \butterfly_st1[3][0][2] (
	.clk(clk),
	.d(\butterfly_st1[3][0][2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[3][0][2]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][0][2] .is_wysiwyg = "true";
defparam \butterfly_st1[3][0][2] .power_up = "low";

dffeas \butterfly_st1[2][1][1] (
	.clk(clk),
	.d(\butterfly_st1[2][1][1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[2][1][1]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][1][1] .is_wysiwyg = "true";
defparam \butterfly_st1[2][1][1] .power_up = "low";

dffeas \butterfly_st1[3][0][1] (
	.clk(clk),
	.d(\butterfly_st1[3][0][1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[3][0][1]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][0][1] .is_wysiwyg = "true";
defparam \butterfly_st1[3][0][1] .power_up = "low";

dffeas \butterfly_st1[2][1][0] (
	.clk(clk),
	.d(\butterfly_st1[2][1][0]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[2][1][0]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][1][0] .is_wysiwyg = "true";
defparam \butterfly_st1[2][1][0] .power_up = "low";

dffeas \butterfly_st1[3][0][0] (
	.clk(clk),
	.d(\butterfly_st1[3][0][0]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[3][0][0]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][0][0] .is_wysiwyg = "true";
defparam \butterfly_st1[3][0][0] .power_up = "low";

cycloneiii_lcell_comb \butterfly_st2[1][1][0]~1 (
	.dataa(\butterfly_st1[2][1][0]~q ),
	.datab(\butterfly_st1[3][0][0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\butterfly_st2[1][1][0]~1_combout ),
	.cout(\butterfly_st2[1][1][0]~2 ));
defparam \butterfly_st2[1][1][0]~1 .lut_mask = 16'h66BB;
defparam \butterfly_st2[1][1][0]~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \butterfly_st2[1][1][1]~1 (
	.dataa(\butterfly_st1[2][1][1]~q ),
	.datab(\butterfly_st1[3][0][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[1][1][0]~2 ),
	.combout(\butterfly_st2[1][1][1]~1_combout ),
	.cout(\butterfly_st2[1][1][1]~2 ));
defparam \butterfly_st2[1][1][1]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st2[1][1][1]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[1][1][2]~1 (
	.dataa(\butterfly_st1[2][1][2]~q ),
	.datab(\butterfly_st1[3][0][2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[1][1][1]~2 ),
	.combout(\butterfly_st2[1][1][2]~1_combout ),
	.cout(\butterfly_st2[1][1][2]~2 ));
defparam \butterfly_st2[1][1][2]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st2[1][1][2]~1 .sum_lutc_input = "cin";

dffeas \butterfly_st1[2][1][8] (
	.clk(clk),
	.d(\butterfly_st1[2][1][8]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[2][1][8]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][1][8] .is_wysiwyg = "true";
defparam \butterfly_st1[2][1][8] .power_up = "low";

dffeas \butterfly_st1[3][0][8] (
	.clk(clk),
	.d(\butterfly_st1[3][0][8]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[3][0][8]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][0][8] .is_wysiwyg = "true";
defparam \butterfly_st1[3][0][8] .power_up = "low";

dffeas \butterfly_st1[2][1][7] (
	.clk(clk),
	.d(\butterfly_st1[2][1][7]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[2][1][7]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][1][7] .is_wysiwyg = "true";
defparam \butterfly_st1[2][1][7] .power_up = "low";

dffeas \butterfly_st1[3][0][7] (
	.clk(clk),
	.d(\butterfly_st1[3][0][7]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[3][0][7]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][0][7] .is_wysiwyg = "true";
defparam \butterfly_st1[3][0][7] .power_up = "low";

dffeas \butterfly_st1[2][1][6] (
	.clk(clk),
	.d(\butterfly_st1[2][1][6]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[2][1][6]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][1][6] .is_wysiwyg = "true";
defparam \butterfly_st1[2][1][6] .power_up = "low";

dffeas \butterfly_st1[3][0][6] (
	.clk(clk),
	.d(\butterfly_st1[3][0][6]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[3][0][6]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][0][6] .is_wysiwyg = "true";
defparam \butterfly_st1[3][0][6] .power_up = "low";

dffeas \butterfly_st1[2][1][5] (
	.clk(clk),
	.d(\butterfly_st1[2][1][5]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[2][1][5]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][1][5] .is_wysiwyg = "true";
defparam \butterfly_st1[2][1][5] .power_up = "low";

dffeas \butterfly_st1[3][0][5] (
	.clk(clk),
	.d(\butterfly_st1[3][0][5]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[3][0][5]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][0][5] .is_wysiwyg = "true";
defparam \butterfly_st1[3][0][5] .power_up = "low";

dffeas \butterfly_st1[2][1][4] (
	.clk(clk),
	.d(\butterfly_st1[2][1][4]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[2][1][4]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][1][4] .is_wysiwyg = "true";
defparam \butterfly_st1[2][1][4] .power_up = "low";

dffeas \butterfly_st1[3][0][4] (
	.clk(clk),
	.d(\butterfly_st1[3][0][4]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[3][0][4]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][0][4] .is_wysiwyg = "true";
defparam \butterfly_st1[3][0][4] .power_up = "low";

dffeas \butterfly_st1[2][1][3] (
	.clk(clk),
	.d(\butterfly_st1[2][1][3]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[2][1][3]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][1][3] .is_wysiwyg = "true";
defparam \butterfly_st1[2][1][3] .power_up = "low";

dffeas \butterfly_st1[3][0][3] (
	.clk(clk),
	.d(\butterfly_st1[3][0][3]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[3][0][3]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][0][3] .is_wysiwyg = "true";
defparam \butterfly_st1[3][0][3] .power_up = "low";

cycloneiii_lcell_comb \butterfly_st2[1][1][3]~1 (
	.dataa(\butterfly_st1[2][1][3]~q ),
	.datab(\butterfly_st1[3][0][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[1][1][2]~2 ),
	.combout(\butterfly_st2[1][1][3]~1_combout ),
	.cout(\butterfly_st2[1][1][3]~2 ));
defparam \butterfly_st2[1][1][3]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st2[1][1][3]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[1][1][4]~1 (
	.dataa(\butterfly_st1[2][1][4]~q ),
	.datab(\butterfly_st1[3][0][4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[1][1][3]~2 ),
	.combout(\butterfly_st2[1][1][4]~1_combout ),
	.cout(\butterfly_st2[1][1][4]~2 ));
defparam \butterfly_st2[1][1][4]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st2[1][1][4]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[1][1][5]~1 (
	.dataa(\butterfly_st1[2][1][5]~q ),
	.datab(\butterfly_st1[3][0][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[1][1][4]~2 ),
	.combout(\butterfly_st2[1][1][5]~1_combout ),
	.cout(\butterfly_st2[1][1][5]~2 ));
defparam \butterfly_st2[1][1][5]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st2[1][1][5]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[1][1][6]~1 (
	.dataa(\butterfly_st1[2][1][6]~q ),
	.datab(\butterfly_st1[3][0][6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[1][1][5]~2 ),
	.combout(\butterfly_st2[1][1][6]~1_combout ),
	.cout(\butterfly_st2[1][1][6]~2 ));
defparam \butterfly_st2[1][1][6]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st2[1][1][6]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[1][1][7]~1 (
	.dataa(\butterfly_st1[2][1][7]~q ),
	.datab(\butterfly_st1[3][0][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[1][1][6]~2 ),
	.combout(\butterfly_st2[1][1][7]~1_combout ),
	.cout(\butterfly_st2[1][1][7]~2 ));
defparam \butterfly_st2[1][1][7]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st2[1][1][7]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[1][1][8]~1 (
	.dataa(\butterfly_st1[2][1][8]~q ),
	.datab(\butterfly_st1[3][0][8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[1][1][7]~2 ),
	.combout(\butterfly_st2[1][1][8]~1_combout ),
	.cout(\butterfly_st2[1][1][8]~2 ));
defparam \butterfly_st2[1][1][8]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st2[1][1][8]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[1][1][9]~1 (
	.dataa(\butterfly_st1[2][1][8]~q ),
	.datab(\butterfly_st1[3][0][8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\butterfly_st2[1][1][8]~2 ),
	.combout(\butterfly_st2[1][1][9]~1_combout ),
	.cout());
defparam \butterfly_st2[1][1][9]~1 .lut_mask = 16'h9696;
defparam \butterfly_st2[1][1][9]~1 .sum_lutc_input = "cin";

dffeas \butterfly_st1[2][0][2] (
	.clk(clk),
	.d(\butterfly_st1[2][0][2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[2][0][2]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][0][2] .is_wysiwyg = "true";
defparam \butterfly_st1[2][0][2] .power_up = "low";

dffeas \butterfly_st1[3][1][2] (
	.clk(clk),
	.d(\butterfly_st1[3][1][2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[3][1][2]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][1][2] .is_wysiwyg = "true";
defparam \butterfly_st1[3][1][2] .power_up = "low";

dffeas \butterfly_st1[2][0][1] (
	.clk(clk),
	.d(\butterfly_st1[2][0][1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[2][0][1]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][0][1] .is_wysiwyg = "true";
defparam \butterfly_st1[2][0][1] .power_up = "low";

dffeas \butterfly_st1[3][1][1] (
	.clk(clk),
	.d(\butterfly_st1[3][1][1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[3][1][1]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][1][1] .is_wysiwyg = "true";
defparam \butterfly_st1[3][1][1] .power_up = "low";

dffeas \butterfly_st1[2][0][0] (
	.clk(clk),
	.d(\butterfly_st1[2][0][0]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[2][0][0]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][0][0] .is_wysiwyg = "true";
defparam \butterfly_st1[2][0][0] .power_up = "low";

dffeas \butterfly_st1[3][1][0] (
	.clk(clk),
	.d(\butterfly_st1[3][1][0]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[3][1][0]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][1][0] .is_wysiwyg = "true";
defparam \butterfly_st1[3][1][0] .power_up = "low";

cycloneiii_lcell_comb \butterfly_st2[1][0][0]~1 (
	.dataa(\butterfly_st1[2][0][0]~q ),
	.datab(\butterfly_st1[3][1][0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\butterfly_st2[1][0][0]~1_combout ),
	.cout(\butterfly_st2[1][0][0]~2 ));
defparam \butterfly_st2[1][0][0]~1 .lut_mask = 16'h66EE;
defparam \butterfly_st2[1][0][0]~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \butterfly_st2[1][0][1]~1 (
	.dataa(\butterfly_st1[2][0][1]~q ),
	.datab(\butterfly_st1[3][1][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[1][0][0]~2 ),
	.combout(\butterfly_st2[1][0][1]~1_combout ),
	.cout(\butterfly_st2[1][0][1]~2 ));
defparam \butterfly_st2[1][0][1]~1 .lut_mask = 16'h967F;
defparam \butterfly_st2[1][0][1]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[1][0][2]~1 (
	.dataa(\butterfly_st1[2][0][2]~q ),
	.datab(\butterfly_st1[3][1][2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[1][0][1]~2 ),
	.combout(\butterfly_st2[1][0][2]~1_combout ),
	.cout(\butterfly_st2[1][0][2]~2 ));
defparam \butterfly_st2[1][0][2]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st2[1][0][2]~1 .sum_lutc_input = "cin";

dffeas \butterfly_st1[2][0][8] (
	.clk(clk),
	.d(\butterfly_st1[2][0][8]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[2][0][8]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][0][8] .is_wysiwyg = "true";
defparam \butterfly_st1[2][0][8] .power_up = "low";

dffeas \butterfly_st1[3][1][8] (
	.clk(clk),
	.d(\butterfly_st1[3][1][8]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[3][1][8]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][1][8] .is_wysiwyg = "true";
defparam \butterfly_st1[3][1][8] .power_up = "low";

dffeas \butterfly_st1[2][0][7] (
	.clk(clk),
	.d(\butterfly_st1[2][0][7]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[2][0][7]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][0][7] .is_wysiwyg = "true";
defparam \butterfly_st1[2][0][7] .power_up = "low";

dffeas \butterfly_st1[3][1][7] (
	.clk(clk),
	.d(\butterfly_st1[3][1][7]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[3][1][7]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][1][7] .is_wysiwyg = "true";
defparam \butterfly_st1[3][1][7] .power_up = "low";

dffeas \butterfly_st1[2][0][6] (
	.clk(clk),
	.d(\butterfly_st1[2][0][6]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[2][0][6]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][0][6] .is_wysiwyg = "true";
defparam \butterfly_st1[2][0][6] .power_up = "low";

dffeas \butterfly_st1[3][1][6] (
	.clk(clk),
	.d(\butterfly_st1[3][1][6]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[3][1][6]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][1][6] .is_wysiwyg = "true";
defparam \butterfly_st1[3][1][6] .power_up = "low";

dffeas \butterfly_st1[2][0][5] (
	.clk(clk),
	.d(\butterfly_st1[2][0][5]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[2][0][5]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][0][5] .is_wysiwyg = "true";
defparam \butterfly_st1[2][0][5] .power_up = "low";

dffeas \butterfly_st1[3][1][5] (
	.clk(clk),
	.d(\butterfly_st1[3][1][5]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[3][1][5]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][1][5] .is_wysiwyg = "true";
defparam \butterfly_st1[3][1][5] .power_up = "low";

dffeas \butterfly_st1[2][0][4] (
	.clk(clk),
	.d(\butterfly_st1[2][0][4]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[2][0][4]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][0][4] .is_wysiwyg = "true";
defparam \butterfly_st1[2][0][4] .power_up = "low";

dffeas \butterfly_st1[3][1][4] (
	.clk(clk),
	.d(\butterfly_st1[3][1][4]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[3][1][4]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][1][4] .is_wysiwyg = "true";
defparam \butterfly_st1[3][1][4] .power_up = "low";

dffeas \butterfly_st1[2][0][3] (
	.clk(clk),
	.d(\butterfly_st1[2][0][3]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[2][0][3]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][0][3] .is_wysiwyg = "true";
defparam \butterfly_st1[2][0][3] .power_up = "low";

dffeas \butterfly_st1[3][1][3] (
	.clk(clk),
	.d(\butterfly_st1[3][1][3]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[3][1][3]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][1][3] .is_wysiwyg = "true";
defparam \butterfly_st1[3][1][3] .power_up = "low";

cycloneiii_lcell_comb \butterfly_st2[1][0][3]~1 (
	.dataa(\butterfly_st1[2][0][3]~q ),
	.datab(\butterfly_st1[3][1][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[1][0][2]~2 ),
	.combout(\butterfly_st2[1][0][3]~1_combout ),
	.cout(\butterfly_st2[1][0][3]~2 ));
defparam \butterfly_st2[1][0][3]~1 .lut_mask = 16'h967F;
defparam \butterfly_st2[1][0][3]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[1][0][4]~1 (
	.dataa(\butterfly_st1[2][0][4]~q ),
	.datab(\butterfly_st1[3][1][4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[1][0][3]~2 ),
	.combout(\butterfly_st2[1][0][4]~1_combout ),
	.cout(\butterfly_st2[1][0][4]~2 ));
defparam \butterfly_st2[1][0][4]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st2[1][0][4]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[1][0][5]~1 (
	.dataa(\butterfly_st1[2][0][5]~q ),
	.datab(\butterfly_st1[3][1][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[1][0][4]~2 ),
	.combout(\butterfly_st2[1][0][5]~1_combout ),
	.cout(\butterfly_st2[1][0][5]~2 ));
defparam \butterfly_st2[1][0][5]~1 .lut_mask = 16'h967F;
defparam \butterfly_st2[1][0][5]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[1][0][6]~1 (
	.dataa(\butterfly_st1[2][0][6]~q ),
	.datab(\butterfly_st1[3][1][6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[1][0][5]~2 ),
	.combout(\butterfly_st2[1][0][6]~1_combout ),
	.cout(\butterfly_st2[1][0][6]~2 ));
defparam \butterfly_st2[1][0][6]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st2[1][0][6]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[1][0][7]~1 (
	.dataa(\butterfly_st1[2][0][7]~q ),
	.datab(\butterfly_st1[3][1][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[1][0][6]~2 ),
	.combout(\butterfly_st2[1][0][7]~1_combout ),
	.cout(\butterfly_st2[1][0][7]~2 ));
defparam \butterfly_st2[1][0][7]~1 .lut_mask = 16'h967F;
defparam \butterfly_st2[1][0][7]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[1][0][8]~1 (
	.dataa(\butterfly_st1[2][0][8]~q ),
	.datab(\butterfly_st1[3][1][8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[1][0][7]~2 ),
	.combout(\butterfly_st2[1][0][8]~1_combout ),
	.cout(\butterfly_st2[1][0][8]~2 ));
defparam \butterfly_st2[1][0][8]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st2[1][0][8]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[1][0][9]~1 (
	.dataa(\butterfly_st1[2][0][8]~q ),
	.datab(\butterfly_st1[3][1][8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\butterfly_st2[1][0][8]~2 ),
	.combout(\butterfly_st2[1][0][9]~1_combout ),
	.cout());
defparam \butterfly_st2[1][0][9]~1 .lut_mask = 16'h9696;
defparam \butterfly_st2[1][0][9]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[2][1][0]~1 (
	.dataa(\butterfly_st1[0][1][0]~q ),
	.datab(\butterfly_st1[1][1][0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\butterfly_st2[2][1][0]~1_combout ),
	.cout(\butterfly_st2[2][1][0]~2 ));
defparam \butterfly_st2[2][1][0]~1 .lut_mask = 16'h66BB;
defparam \butterfly_st2[2][1][0]~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \butterfly_st2[2][1][1]~1 (
	.dataa(\butterfly_st1[0][1][1]~q ),
	.datab(\butterfly_st1[1][1][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[2][1][0]~2 ),
	.combout(\butterfly_st2[2][1][1]~1_combout ),
	.cout(\butterfly_st2[2][1][1]~2 ));
defparam \butterfly_st2[2][1][1]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st2[2][1][1]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[2][1][2]~1 (
	.dataa(\butterfly_st1[0][1][2]~q ),
	.datab(\butterfly_st1[1][1][2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[2][1][1]~2 ),
	.combout(\butterfly_st2[2][1][2]~1_combout ),
	.cout(\butterfly_st2[2][1][2]~2 ));
defparam \butterfly_st2[2][1][2]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st2[2][1][2]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[2][1][3]~1 (
	.dataa(\butterfly_st1[0][1][3]~q ),
	.datab(\butterfly_st1[1][1][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[2][1][2]~2 ),
	.combout(\butterfly_st2[2][1][3]~1_combout ),
	.cout(\butterfly_st2[2][1][3]~2 ));
defparam \butterfly_st2[2][1][3]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st2[2][1][3]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[2][1][4]~1 (
	.dataa(\butterfly_st1[0][1][4]~q ),
	.datab(\butterfly_st1[1][1][4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[2][1][3]~2 ),
	.combout(\butterfly_st2[2][1][4]~1_combout ),
	.cout(\butterfly_st2[2][1][4]~2 ));
defparam \butterfly_st2[2][1][4]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st2[2][1][4]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[2][1][5]~1 (
	.dataa(\butterfly_st1[0][1][5]~q ),
	.datab(\butterfly_st1[1][1][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[2][1][4]~2 ),
	.combout(\butterfly_st2[2][1][5]~1_combout ),
	.cout(\butterfly_st2[2][1][5]~2 ));
defparam \butterfly_st2[2][1][5]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st2[2][1][5]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[2][1][6]~1 (
	.dataa(\butterfly_st1[0][1][6]~q ),
	.datab(\butterfly_st1[1][1][6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[2][1][5]~2 ),
	.combout(\butterfly_st2[2][1][6]~1_combout ),
	.cout(\butterfly_st2[2][1][6]~2 ));
defparam \butterfly_st2[2][1][6]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st2[2][1][6]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[2][1][7]~1 (
	.dataa(\butterfly_st1[0][1][7]~q ),
	.datab(\butterfly_st1[1][1][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[2][1][6]~2 ),
	.combout(\butterfly_st2[2][1][7]~1_combout ),
	.cout(\butterfly_st2[2][1][7]~2 ));
defparam \butterfly_st2[2][1][7]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st2[2][1][7]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[2][1][8]~1 (
	.dataa(\butterfly_st1[0][1][8]~q ),
	.datab(\butterfly_st1[1][1][8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[2][1][7]~2 ),
	.combout(\butterfly_st2[2][1][8]~1_combout ),
	.cout(\butterfly_st2[2][1][8]~2 ));
defparam \butterfly_st2[2][1][8]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st2[2][1][8]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[2][1][9]~1 (
	.dataa(\butterfly_st1[0][1][8]~q ),
	.datab(\butterfly_st1[1][1][8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\butterfly_st2[2][1][8]~2 ),
	.combout(\butterfly_st2[2][1][9]~1_combout ),
	.cout());
defparam \butterfly_st2[2][1][9]~1 .lut_mask = 16'h9696;
defparam \butterfly_st2[2][1][9]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[2][0][0]~1 (
	.dataa(\butterfly_st1[0][0][0]~q ),
	.datab(\butterfly_st1[1][0][0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\butterfly_st2[2][0][0]~1_combout ),
	.cout(\butterfly_st2[2][0][0]~2 ));
defparam \butterfly_st2[2][0][0]~1 .lut_mask = 16'h66BB;
defparam \butterfly_st2[2][0][0]~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \butterfly_st2[2][0][1]~1 (
	.dataa(\butterfly_st1[0][0][1]~q ),
	.datab(\butterfly_st1[1][0][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[2][0][0]~2 ),
	.combout(\butterfly_st2[2][0][1]~1_combout ),
	.cout(\butterfly_st2[2][0][1]~2 ));
defparam \butterfly_st2[2][0][1]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st2[2][0][1]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[2][0][2]~1 (
	.dataa(\butterfly_st1[0][0][2]~q ),
	.datab(\butterfly_st1[1][0][2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[2][0][1]~2 ),
	.combout(\butterfly_st2[2][0][2]~1_combout ),
	.cout(\butterfly_st2[2][0][2]~2 ));
defparam \butterfly_st2[2][0][2]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st2[2][0][2]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[2][0][3]~1 (
	.dataa(\butterfly_st1[0][0][3]~q ),
	.datab(\butterfly_st1[1][0][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[2][0][2]~2 ),
	.combout(\butterfly_st2[2][0][3]~1_combout ),
	.cout(\butterfly_st2[2][0][3]~2 ));
defparam \butterfly_st2[2][0][3]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st2[2][0][3]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[2][0][4]~1 (
	.dataa(\butterfly_st1[0][0][4]~q ),
	.datab(\butterfly_st1[1][0][4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[2][0][3]~2 ),
	.combout(\butterfly_st2[2][0][4]~1_combout ),
	.cout(\butterfly_st2[2][0][4]~2 ));
defparam \butterfly_st2[2][0][4]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st2[2][0][4]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[2][0][5]~1 (
	.dataa(\butterfly_st1[0][0][5]~q ),
	.datab(\butterfly_st1[1][0][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[2][0][4]~2 ),
	.combout(\butterfly_st2[2][0][5]~1_combout ),
	.cout(\butterfly_st2[2][0][5]~2 ));
defparam \butterfly_st2[2][0][5]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st2[2][0][5]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[2][0][6]~1 (
	.dataa(\butterfly_st1[0][0][6]~q ),
	.datab(\butterfly_st1[1][0][6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[2][0][5]~2 ),
	.combout(\butterfly_st2[2][0][6]~1_combout ),
	.cout(\butterfly_st2[2][0][6]~2 ));
defparam \butterfly_st2[2][0][6]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st2[2][0][6]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[2][0][7]~1 (
	.dataa(\butterfly_st1[0][0][7]~q ),
	.datab(\butterfly_st1[1][0][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[2][0][6]~2 ),
	.combout(\butterfly_st2[2][0][7]~1_combout ),
	.cout(\butterfly_st2[2][0][7]~2 ));
defparam \butterfly_st2[2][0][7]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st2[2][0][7]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[2][0][8]~1 (
	.dataa(\butterfly_st1[0][0][8]~q ),
	.datab(\butterfly_st1[1][0][8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[2][0][7]~2 ),
	.combout(\butterfly_st2[2][0][8]~1_combout ),
	.cout(\butterfly_st2[2][0][8]~2 ));
defparam \butterfly_st2[2][0][8]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st2[2][0][8]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[2][0][9]~1 (
	.dataa(\butterfly_st1[0][0][8]~q ),
	.datab(\butterfly_st1[1][0][8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\butterfly_st2[2][0][8]~2 ),
	.combout(\butterfly_st2[2][0][9]~1_combout ),
	.cout());
defparam \butterfly_st2[2][0][9]~1 .lut_mask = 16'h9696;
defparam \butterfly_st2[2][0][9]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[3][1][0]~1 (
	.dataa(\butterfly_st1[2][1][0]~q ),
	.datab(\butterfly_st1[3][0][0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\butterfly_st2[3][1][0]~1_combout ),
	.cout(\butterfly_st2[3][1][0]~2 ));
defparam \butterfly_st2[3][1][0]~1 .lut_mask = 16'h66EE;
defparam \butterfly_st2[3][1][0]~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \butterfly_st2[3][1][1]~1 (
	.dataa(\butterfly_st1[2][1][1]~q ),
	.datab(\butterfly_st1[3][0][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[3][1][0]~2 ),
	.combout(\butterfly_st2[3][1][1]~1_combout ),
	.cout(\butterfly_st2[3][1][1]~2 ));
defparam \butterfly_st2[3][1][1]~1 .lut_mask = 16'h967F;
defparam \butterfly_st2[3][1][1]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[3][1][2]~1 (
	.dataa(\butterfly_st1[2][1][2]~q ),
	.datab(\butterfly_st1[3][0][2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[3][1][1]~2 ),
	.combout(\butterfly_st2[3][1][2]~1_combout ),
	.cout(\butterfly_st2[3][1][2]~2 ));
defparam \butterfly_st2[3][1][2]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st2[3][1][2]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[3][1][3]~1 (
	.dataa(\butterfly_st1[2][1][3]~q ),
	.datab(\butterfly_st1[3][0][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[3][1][2]~2 ),
	.combout(\butterfly_st2[3][1][3]~1_combout ),
	.cout(\butterfly_st2[3][1][3]~2 ));
defparam \butterfly_st2[3][1][3]~1 .lut_mask = 16'h967F;
defparam \butterfly_st2[3][1][3]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[3][1][4]~1 (
	.dataa(\butterfly_st1[2][1][4]~q ),
	.datab(\butterfly_st1[3][0][4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[3][1][3]~2 ),
	.combout(\butterfly_st2[3][1][4]~1_combout ),
	.cout(\butterfly_st2[3][1][4]~2 ));
defparam \butterfly_st2[3][1][4]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st2[3][1][4]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[3][1][5]~1 (
	.dataa(\butterfly_st1[2][1][5]~q ),
	.datab(\butterfly_st1[3][0][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[3][1][4]~2 ),
	.combout(\butterfly_st2[3][1][5]~1_combout ),
	.cout(\butterfly_st2[3][1][5]~2 ));
defparam \butterfly_st2[3][1][5]~1 .lut_mask = 16'h967F;
defparam \butterfly_st2[3][1][5]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[3][1][6]~1 (
	.dataa(\butterfly_st1[2][1][6]~q ),
	.datab(\butterfly_st1[3][0][6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[3][1][5]~2 ),
	.combout(\butterfly_st2[3][1][6]~1_combout ),
	.cout(\butterfly_st2[3][1][6]~2 ));
defparam \butterfly_st2[3][1][6]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st2[3][1][6]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[3][1][7]~1 (
	.dataa(\butterfly_st1[2][1][7]~q ),
	.datab(\butterfly_st1[3][0][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[3][1][6]~2 ),
	.combout(\butterfly_st2[3][1][7]~1_combout ),
	.cout(\butterfly_st2[3][1][7]~2 ));
defparam \butterfly_st2[3][1][7]~1 .lut_mask = 16'h967F;
defparam \butterfly_st2[3][1][7]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[3][1][8]~1 (
	.dataa(\butterfly_st1[2][1][8]~q ),
	.datab(\butterfly_st1[3][0][8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[3][1][7]~2 ),
	.combout(\butterfly_st2[3][1][8]~1_combout ),
	.cout(\butterfly_st2[3][1][8]~2 ));
defparam \butterfly_st2[3][1][8]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st2[3][1][8]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[3][1][9]~1 (
	.dataa(\butterfly_st1[2][1][8]~q ),
	.datab(\butterfly_st1[3][0][8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\butterfly_st2[3][1][8]~2 ),
	.combout(\butterfly_st2[3][1][9]~1_combout ),
	.cout());
defparam \butterfly_st2[3][1][9]~1 .lut_mask = 16'h9696;
defparam \butterfly_st2[3][1][9]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[3][0][0]~1 (
	.dataa(\butterfly_st1[2][0][0]~q ),
	.datab(\butterfly_st1[3][1][0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\butterfly_st2[3][0][0]~1_combout ),
	.cout(\butterfly_st2[3][0][0]~2 ));
defparam \butterfly_st2[3][0][0]~1 .lut_mask = 16'h66BB;
defparam \butterfly_st2[3][0][0]~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \butterfly_st2[3][0][1]~1 (
	.dataa(\butterfly_st1[2][0][1]~q ),
	.datab(\butterfly_st1[3][1][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[3][0][0]~2 ),
	.combout(\butterfly_st2[3][0][1]~1_combout ),
	.cout(\butterfly_st2[3][0][1]~2 ));
defparam \butterfly_st2[3][0][1]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st2[3][0][1]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[3][0][2]~1 (
	.dataa(\butterfly_st1[2][0][2]~q ),
	.datab(\butterfly_st1[3][1][2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[3][0][1]~2 ),
	.combout(\butterfly_st2[3][0][2]~1_combout ),
	.cout(\butterfly_st2[3][0][2]~2 ));
defparam \butterfly_st2[3][0][2]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st2[3][0][2]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[3][0][3]~1 (
	.dataa(\butterfly_st1[2][0][3]~q ),
	.datab(\butterfly_st1[3][1][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[3][0][2]~2 ),
	.combout(\butterfly_st2[3][0][3]~1_combout ),
	.cout(\butterfly_st2[3][0][3]~2 ));
defparam \butterfly_st2[3][0][3]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st2[3][0][3]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[3][0][4]~1 (
	.dataa(\butterfly_st1[2][0][4]~q ),
	.datab(\butterfly_st1[3][1][4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[3][0][3]~2 ),
	.combout(\butterfly_st2[3][0][4]~1_combout ),
	.cout(\butterfly_st2[3][0][4]~2 ));
defparam \butterfly_st2[3][0][4]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st2[3][0][4]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[3][0][5]~1 (
	.dataa(\butterfly_st1[2][0][5]~q ),
	.datab(\butterfly_st1[3][1][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[3][0][4]~2 ),
	.combout(\butterfly_st2[3][0][5]~1_combout ),
	.cout(\butterfly_st2[3][0][5]~2 ));
defparam \butterfly_st2[3][0][5]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st2[3][0][5]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[3][0][6]~1 (
	.dataa(\butterfly_st1[2][0][6]~q ),
	.datab(\butterfly_st1[3][1][6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[3][0][5]~2 ),
	.combout(\butterfly_st2[3][0][6]~1_combout ),
	.cout(\butterfly_st2[3][0][6]~2 ));
defparam \butterfly_st2[3][0][6]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st2[3][0][6]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[3][0][7]~1 (
	.dataa(\butterfly_st1[2][0][7]~q ),
	.datab(\butterfly_st1[3][1][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[3][0][6]~2 ),
	.combout(\butterfly_st2[3][0][7]~1_combout ),
	.cout(\butterfly_st2[3][0][7]~2 ));
defparam \butterfly_st2[3][0][7]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st2[3][0][7]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[3][0][8]~1 (
	.dataa(\butterfly_st1[2][0][8]~q ),
	.datab(\butterfly_st1[3][1][8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[3][0][7]~2 ),
	.combout(\butterfly_st2[3][0][8]~1_combout ),
	.cout(\butterfly_st2[3][0][8]~2 ));
defparam \butterfly_st2[3][0][8]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st2[3][0][8]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st2[3][0][9]~1 (
	.dataa(\butterfly_st1[2][0][8]~q ),
	.datab(\butterfly_st1[3][1][8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\butterfly_st2[3][0][8]~2 ),
	.combout(\butterfly_st2[3][0][9]~1_combout ),
	.cout());
defparam \butterfly_st2[3][0][9]~1 .lut_mask = 16'h9696;
defparam \butterfly_st2[3][0][9]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[0][0][0]~1 (
	.dataa(\gen_cont:bfp_scale|r_array_out[0][0]~q ),
	.datab(\gen_cont:bfp_scale|r_array_out[2][0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\butterfly_st1[0][0][0]~1_combout ),
	.cout(\butterfly_st1[0][0][0]~2 ));
defparam \butterfly_st1[0][0][0]~1 .lut_mask = 16'h66EE;
defparam \butterfly_st1[0][0][0]~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \butterfly_st1[0][0][1]~1 (
	.dataa(\gen_cont:bfp_scale|r_array_out[0][1]~q ),
	.datab(\gen_cont:bfp_scale|r_array_out[2][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[0][0][0]~2 ),
	.combout(\butterfly_st1[0][0][1]~1_combout ),
	.cout(\butterfly_st1[0][0][1]~2 ));
defparam \butterfly_st1[0][0][1]~1 .lut_mask = 16'h967F;
defparam \butterfly_st1[0][0][1]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[0][0][2]~1 (
	.dataa(\gen_cont:bfp_scale|r_array_out[0][2]~q ),
	.datab(\gen_cont:bfp_scale|r_array_out[2][2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[0][0][1]~2 ),
	.combout(\butterfly_st1[0][0][2]~1_combout ),
	.cout(\butterfly_st1[0][0][2]~2 ));
defparam \butterfly_st1[0][0][2]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st1[0][0][2]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[0][0][3]~1 (
	.dataa(\gen_cont:bfp_scale|r_array_out[0][3]~q ),
	.datab(\gen_cont:bfp_scale|r_array_out[2][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[0][0][2]~2 ),
	.combout(\butterfly_st1[0][0][3]~1_combout ),
	.cout(\butterfly_st1[0][0][3]~2 ));
defparam \butterfly_st1[0][0][3]~1 .lut_mask = 16'h967F;
defparam \butterfly_st1[0][0][3]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[0][0][4]~1 (
	.dataa(\gen_cont:bfp_scale|r_array_out[0][4]~q ),
	.datab(\gen_cont:bfp_scale|r_array_out[2][4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[0][0][3]~2 ),
	.combout(\butterfly_st1[0][0][4]~1_combout ),
	.cout(\butterfly_st1[0][0][4]~2 ));
defparam \butterfly_st1[0][0][4]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st1[0][0][4]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[0][0][5]~1 (
	.dataa(\gen_cont:bfp_scale|r_array_out[0][5]~q ),
	.datab(\gen_cont:bfp_scale|r_array_out[2][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[0][0][4]~2 ),
	.combout(\butterfly_st1[0][0][5]~1_combout ),
	.cout(\butterfly_st1[0][0][5]~2 ));
defparam \butterfly_st1[0][0][5]~1 .lut_mask = 16'h967F;
defparam \butterfly_st1[0][0][5]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[0][0][6]~1 (
	.dataa(\gen_cont:bfp_scale|r_array_out[0][6]~q ),
	.datab(\gen_cont:bfp_scale|r_array_out[2][6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[0][0][5]~2 ),
	.combout(\butterfly_st1[0][0][6]~1_combout ),
	.cout(\butterfly_st1[0][0][6]~2 ));
defparam \butterfly_st1[0][0][6]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st1[0][0][6]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[1][0][0]~1 (
	.dataa(\gen_cont:bfp_scale|r_array_out[1][0]~q ),
	.datab(\gen_cont:bfp_scale|r_array_out[3][0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\butterfly_st1[1][0][0]~1_combout ),
	.cout(\butterfly_st1[1][0][0]~2 ));
defparam \butterfly_st1[1][0][0]~1 .lut_mask = 16'h66EE;
defparam \butterfly_st1[1][0][0]~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \butterfly_st1[1][0][1]~1 (
	.dataa(\gen_cont:bfp_scale|r_array_out[1][1]~q ),
	.datab(\gen_cont:bfp_scale|r_array_out[3][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[1][0][0]~2 ),
	.combout(\butterfly_st1[1][0][1]~1_combout ),
	.cout(\butterfly_st1[1][0][1]~2 ));
defparam \butterfly_st1[1][0][1]~1 .lut_mask = 16'h967F;
defparam \butterfly_st1[1][0][1]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[1][0][2]~1 (
	.dataa(\gen_cont:bfp_scale|r_array_out[1][2]~q ),
	.datab(\gen_cont:bfp_scale|r_array_out[3][2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[1][0][1]~2 ),
	.combout(\butterfly_st1[1][0][2]~1_combout ),
	.cout(\butterfly_st1[1][0][2]~2 ));
defparam \butterfly_st1[1][0][2]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st1[1][0][2]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[1][0][3]~1 (
	.dataa(\gen_cont:bfp_scale|r_array_out[1][3]~q ),
	.datab(\gen_cont:bfp_scale|r_array_out[3][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[1][0][2]~2 ),
	.combout(\butterfly_st1[1][0][3]~1_combout ),
	.cout(\butterfly_st1[1][0][3]~2 ));
defparam \butterfly_st1[1][0][3]~1 .lut_mask = 16'h967F;
defparam \butterfly_st1[1][0][3]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[1][0][4]~1 (
	.dataa(\gen_cont:bfp_scale|r_array_out[1][4]~q ),
	.datab(\gen_cont:bfp_scale|r_array_out[3][4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[1][0][3]~2 ),
	.combout(\butterfly_st1[1][0][4]~1_combout ),
	.cout(\butterfly_st1[1][0][4]~2 ));
defparam \butterfly_st1[1][0][4]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st1[1][0][4]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[1][0][5]~1 (
	.dataa(\gen_cont:bfp_scale|r_array_out[1][5]~q ),
	.datab(\gen_cont:bfp_scale|r_array_out[3][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[1][0][4]~2 ),
	.combout(\butterfly_st1[1][0][5]~1_combout ),
	.cout(\butterfly_st1[1][0][5]~2 ));
defparam \butterfly_st1[1][0][5]~1 .lut_mask = 16'h967F;
defparam \butterfly_st1[1][0][5]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[1][0][6]~1 (
	.dataa(\gen_cont:bfp_scale|r_array_out[1][6]~q ),
	.datab(\gen_cont:bfp_scale|r_array_out[3][6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[1][0][5]~2 ),
	.combout(\butterfly_st1[1][0][6]~1_combout ),
	.cout(\butterfly_st1[1][0][6]~2 ));
defparam \butterfly_st1[1][0][6]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st1[1][0][6]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[0][0][7]~1 (
	.dataa(\gen_cont:bfp_scale|r_array_out[0][7]~q ),
	.datab(\gen_cont:bfp_scale|r_array_out[2][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[0][0][6]~2 ),
	.combout(\butterfly_st1[0][0][7]~1_combout ),
	.cout(\butterfly_st1[0][0][7]~2 ));
defparam \butterfly_st1[0][0][7]~1 .lut_mask = 16'h967F;
defparam \butterfly_st1[0][0][7]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[0][0][8]~1 (
	.dataa(\gen_cont:bfp_scale|r_array_out[0][7]~q ),
	.datab(\gen_cont:bfp_scale|r_array_out[2][7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\butterfly_st1[0][0][7]~2 ),
	.combout(\butterfly_st1[0][0][8]~1_combout ),
	.cout());
defparam \butterfly_st1[0][0][8]~1 .lut_mask = 16'h9696;
defparam \butterfly_st1[0][0][8]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[1][0][7]~1 (
	.dataa(\gen_cont:bfp_scale|r_array_out[1][7]~q ),
	.datab(\gen_cont:bfp_scale|r_array_out[3][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[1][0][6]~2 ),
	.combout(\butterfly_st1[1][0][7]~1_combout ),
	.cout(\butterfly_st1[1][0][7]~2 ));
defparam \butterfly_st1[1][0][7]~1 .lut_mask = 16'h967F;
defparam \butterfly_st1[1][0][7]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[1][0][8]~1 (
	.dataa(\gen_cont:bfp_scale|r_array_out[1][7]~q ),
	.datab(\gen_cont:bfp_scale|r_array_out[3][7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\butterfly_st1[1][0][7]~2 ),
	.combout(\butterfly_st1[1][0][8]~1_combout ),
	.cout());
defparam \butterfly_st1[1][0][8]~1 .lut_mask = 16'h9696;
defparam \butterfly_st1[1][0][8]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[0][1][0]~1 (
	.dataa(\gen_cont:bfp_scale|i_array_out[0][0]~q ),
	.datab(\gen_cont:bfp_scale|i_array_out[2][0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\butterfly_st1[0][1][0]~1_combout ),
	.cout(\butterfly_st1[0][1][0]~2 ));
defparam \butterfly_st1[0][1][0]~1 .lut_mask = 16'h66EE;
defparam \butterfly_st1[0][1][0]~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \butterfly_st1[0][1][1]~1 (
	.dataa(\gen_cont:bfp_scale|i_array_out[0][1]~q ),
	.datab(\gen_cont:bfp_scale|i_array_out[2][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[0][1][0]~2 ),
	.combout(\butterfly_st1[0][1][1]~1_combout ),
	.cout(\butterfly_st1[0][1][1]~2 ));
defparam \butterfly_st1[0][1][1]~1 .lut_mask = 16'h967F;
defparam \butterfly_st1[0][1][1]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[0][1][2]~1 (
	.dataa(\gen_cont:bfp_scale|i_array_out[0][2]~q ),
	.datab(\gen_cont:bfp_scale|i_array_out[2][2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[0][1][1]~2 ),
	.combout(\butterfly_st1[0][1][2]~1_combout ),
	.cout(\butterfly_st1[0][1][2]~2 ));
defparam \butterfly_st1[0][1][2]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st1[0][1][2]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[0][1][3]~1 (
	.dataa(\gen_cont:bfp_scale|i_array_out[0][3]~q ),
	.datab(\gen_cont:bfp_scale|i_array_out[2][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[0][1][2]~2 ),
	.combout(\butterfly_st1[0][1][3]~1_combout ),
	.cout(\butterfly_st1[0][1][3]~2 ));
defparam \butterfly_st1[0][1][3]~1 .lut_mask = 16'h967F;
defparam \butterfly_st1[0][1][3]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[0][1][4]~1 (
	.dataa(\gen_cont:bfp_scale|i_array_out[0][4]~q ),
	.datab(\gen_cont:bfp_scale|i_array_out[2][4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[0][1][3]~2 ),
	.combout(\butterfly_st1[0][1][4]~1_combout ),
	.cout(\butterfly_st1[0][1][4]~2 ));
defparam \butterfly_st1[0][1][4]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st1[0][1][4]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[0][1][5]~1 (
	.dataa(\gen_cont:bfp_scale|i_array_out[0][5]~q ),
	.datab(\gen_cont:bfp_scale|i_array_out[2][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[0][1][4]~2 ),
	.combout(\butterfly_st1[0][1][5]~1_combout ),
	.cout(\butterfly_st1[0][1][5]~2 ));
defparam \butterfly_st1[0][1][5]~1 .lut_mask = 16'h967F;
defparam \butterfly_st1[0][1][5]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[0][1][6]~1 (
	.dataa(\gen_cont:bfp_scale|i_array_out[0][6]~q ),
	.datab(\gen_cont:bfp_scale|i_array_out[2][6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[0][1][5]~2 ),
	.combout(\butterfly_st1[0][1][6]~1_combout ),
	.cout(\butterfly_st1[0][1][6]~2 ));
defparam \butterfly_st1[0][1][6]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st1[0][1][6]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[0][1][7]~1 (
	.dataa(\gen_cont:bfp_scale|i_array_out[0][7]~q ),
	.datab(\gen_cont:bfp_scale|i_array_out[2][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[0][1][6]~2 ),
	.combout(\butterfly_st1[0][1][7]~1_combout ),
	.cout(\butterfly_st1[0][1][7]~2 ));
defparam \butterfly_st1[0][1][7]~1 .lut_mask = 16'h967F;
defparam \butterfly_st1[0][1][7]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[0][1][8]~1 (
	.dataa(\gen_cont:bfp_scale|i_array_out[0][7]~q ),
	.datab(\gen_cont:bfp_scale|i_array_out[2][7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\butterfly_st1[0][1][7]~2 ),
	.combout(\butterfly_st1[0][1][8]~1_combout ),
	.cout());
defparam \butterfly_st1[0][1][8]~1 .lut_mask = 16'h9696;
defparam \butterfly_st1[0][1][8]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[1][1][0]~1 (
	.dataa(\gen_cont:bfp_scale|i_array_out[1][0]~q ),
	.datab(\gen_cont:bfp_scale|i_array_out[3][0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\butterfly_st1[1][1][0]~1_combout ),
	.cout(\butterfly_st1[1][1][0]~2 ));
defparam \butterfly_st1[1][1][0]~1 .lut_mask = 16'h66EE;
defparam \butterfly_st1[1][1][0]~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \butterfly_st1[1][1][1]~1 (
	.dataa(\gen_cont:bfp_scale|i_array_out[1][1]~q ),
	.datab(\gen_cont:bfp_scale|i_array_out[3][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[1][1][0]~2 ),
	.combout(\butterfly_st1[1][1][1]~1_combout ),
	.cout(\butterfly_st1[1][1][1]~2 ));
defparam \butterfly_st1[1][1][1]~1 .lut_mask = 16'h967F;
defparam \butterfly_st1[1][1][1]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[1][1][2]~1 (
	.dataa(\gen_cont:bfp_scale|i_array_out[1][2]~q ),
	.datab(\gen_cont:bfp_scale|i_array_out[3][2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[1][1][1]~2 ),
	.combout(\butterfly_st1[1][1][2]~1_combout ),
	.cout(\butterfly_st1[1][1][2]~2 ));
defparam \butterfly_st1[1][1][2]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st1[1][1][2]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[1][1][3]~1 (
	.dataa(\gen_cont:bfp_scale|i_array_out[1][3]~q ),
	.datab(\gen_cont:bfp_scale|i_array_out[3][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[1][1][2]~2 ),
	.combout(\butterfly_st1[1][1][3]~1_combout ),
	.cout(\butterfly_st1[1][1][3]~2 ));
defparam \butterfly_st1[1][1][3]~1 .lut_mask = 16'h967F;
defparam \butterfly_st1[1][1][3]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[1][1][4]~1 (
	.dataa(\gen_cont:bfp_scale|i_array_out[1][4]~q ),
	.datab(\gen_cont:bfp_scale|i_array_out[3][4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[1][1][3]~2 ),
	.combout(\butterfly_st1[1][1][4]~1_combout ),
	.cout(\butterfly_st1[1][1][4]~2 ));
defparam \butterfly_st1[1][1][4]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st1[1][1][4]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[1][1][5]~1 (
	.dataa(\gen_cont:bfp_scale|i_array_out[1][5]~q ),
	.datab(\gen_cont:bfp_scale|i_array_out[3][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[1][1][4]~2 ),
	.combout(\butterfly_st1[1][1][5]~1_combout ),
	.cout(\butterfly_st1[1][1][5]~2 ));
defparam \butterfly_st1[1][1][5]~1 .lut_mask = 16'h967F;
defparam \butterfly_st1[1][1][5]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[1][1][6]~1 (
	.dataa(\gen_cont:bfp_scale|i_array_out[1][6]~q ),
	.datab(\gen_cont:bfp_scale|i_array_out[3][6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[1][1][5]~2 ),
	.combout(\butterfly_st1[1][1][6]~1_combout ),
	.cout(\butterfly_st1[1][1][6]~2 ));
defparam \butterfly_st1[1][1][6]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st1[1][1][6]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[1][1][7]~1 (
	.dataa(\gen_cont:bfp_scale|i_array_out[1][7]~q ),
	.datab(\gen_cont:bfp_scale|i_array_out[3][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[1][1][6]~2 ),
	.combout(\butterfly_st1[1][1][7]~1_combout ),
	.cout(\butterfly_st1[1][1][7]~2 ));
defparam \butterfly_st1[1][1][7]~1 .lut_mask = 16'h967F;
defparam \butterfly_st1[1][1][7]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[1][1][8]~1 (
	.dataa(\gen_cont:bfp_scale|i_array_out[1][7]~q ),
	.datab(\gen_cont:bfp_scale|i_array_out[3][7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\butterfly_st1[1][1][7]~2 ),
	.combout(\butterfly_st1[1][1][8]~1_combout ),
	.cout());
defparam \butterfly_st1[1][1][8]~1 .lut_mask = 16'h9696;
defparam \butterfly_st1[1][1][8]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[2][1][0]~1 (
	.dataa(\gen_cont:bfp_scale|i_array_out[0][0]~q ),
	.datab(\gen_cont:bfp_scale|i_array_out[2][0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\butterfly_st1[2][1][0]~1_combout ),
	.cout(\butterfly_st1[2][1][0]~2 ));
defparam \butterfly_st1[2][1][0]~1 .lut_mask = 16'h66BB;
defparam \butterfly_st1[2][1][0]~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \butterfly_st1[2][1][1]~1 (
	.dataa(\gen_cont:bfp_scale|i_array_out[0][1]~q ),
	.datab(\gen_cont:bfp_scale|i_array_out[2][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[2][1][0]~2 ),
	.combout(\butterfly_st1[2][1][1]~1_combout ),
	.cout(\butterfly_st1[2][1][1]~2 ));
defparam \butterfly_st1[2][1][1]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st1[2][1][1]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[2][1][2]~1 (
	.dataa(\gen_cont:bfp_scale|i_array_out[0][2]~q ),
	.datab(\gen_cont:bfp_scale|i_array_out[2][2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[2][1][1]~2 ),
	.combout(\butterfly_st1[2][1][2]~1_combout ),
	.cout(\butterfly_st1[2][1][2]~2 ));
defparam \butterfly_st1[2][1][2]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st1[2][1][2]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[3][0][0]~1 (
	.dataa(\gen_cont:bfp_scale|r_array_out[1][0]~q ),
	.datab(\gen_cont:bfp_scale|r_array_out[3][0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\butterfly_st1[3][0][0]~1_combout ),
	.cout(\butterfly_st1[3][0][0]~2 ));
defparam \butterfly_st1[3][0][0]~1 .lut_mask = 16'h66BB;
defparam \butterfly_st1[3][0][0]~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \butterfly_st1[3][0][1]~1 (
	.dataa(\gen_cont:bfp_scale|r_array_out[1][1]~q ),
	.datab(\gen_cont:bfp_scale|r_array_out[3][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[3][0][0]~2 ),
	.combout(\butterfly_st1[3][0][1]~1_combout ),
	.cout(\butterfly_st1[3][0][1]~2 ));
defparam \butterfly_st1[3][0][1]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st1[3][0][1]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[3][0][2]~1 (
	.dataa(\gen_cont:bfp_scale|r_array_out[1][2]~q ),
	.datab(\gen_cont:bfp_scale|r_array_out[3][2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[3][0][1]~2 ),
	.combout(\butterfly_st1[3][0][2]~1_combout ),
	.cout(\butterfly_st1[3][0][2]~2 ));
defparam \butterfly_st1[3][0][2]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st1[3][0][2]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[2][1][3]~1 (
	.dataa(\gen_cont:bfp_scale|i_array_out[0][3]~q ),
	.datab(\gen_cont:bfp_scale|i_array_out[2][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[2][1][2]~2 ),
	.combout(\butterfly_st1[2][1][3]~1_combout ),
	.cout(\butterfly_st1[2][1][3]~2 ));
defparam \butterfly_st1[2][1][3]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st1[2][1][3]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[2][1][4]~1 (
	.dataa(\gen_cont:bfp_scale|i_array_out[0][4]~q ),
	.datab(\gen_cont:bfp_scale|i_array_out[2][4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[2][1][3]~2 ),
	.combout(\butterfly_st1[2][1][4]~1_combout ),
	.cout(\butterfly_st1[2][1][4]~2 ));
defparam \butterfly_st1[2][1][4]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st1[2][1][4]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[2][1][5]~1 (
	.dataa(\gen_cont:bfp_scale|i_array_out[0][5]~q ),
	.datab(\gen_cont:bfp_scale|i_array_out[2][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[2][1][4]~2 ),
	.combout(\butterfly_st1[2][1][5]~1_combout ),
	.cout(\butterfly_st1[2][1][5]~2 ));
defparam \butterfly_st1[2][1][5]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st1[2][1][5]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[2][1][6]~1 (
	.dataa(\gen_cont:bfp_scale|i_array_out[0][6]~q ),
	.datab(\gen_cont:bfp_scale|i_array_out[2][6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[2][1][5]~2 ),
	.combout(\butterfly_st1[2][1][6]~1_combout ),
	.cout(\butterfly_st1[2][1][6]~2 ));
defparam \butterfly_st1[2][1][6]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st1[2][1][6]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[2][1][7]~1 (
	.dataa(\gen_cont:bfp_scale|i_array_out[0][7]~q ),
	.datab(\gen_cont:bfp_scale|i_array_out[2][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[2][1][6]~2 ),
	.combout(\butterfly_st1[2][1][7]~1_combout ),
	.cout(\butterfly_st1[2][1][7]~2 ));
defparam \butterfly_st1[2][1][7]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st1[2][1][7]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[2][1][8]~1 (
	.dataa(\gen_cont:bfp_scale|i_array_out[0][7]~q ),
	.datab(\gen_cont:bfp_scale|i_array_out[2][7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\butterfly_st1[2][1][7]~2 ),
	.combout(\butterfly_st1[2][1][8]~1_combout ),
	.cout());
defparam \butterfly_st1[2][1][8]~1 .lut_mask = 16'h9696;
defparam \butterfly_st1[2][1][8]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[3][0][3]~1 (
	.dataa(\gen_cont:bfp_scale|r_array_out[1][3]~q ),
	.datab(\gen_cont:bfp_scale|r_array_out[3][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[3][0][2]~2 ),
	.combout(\butterfly_st1[3][0][3]~1_combout ),
	.cout(\butterfly_st1[3][0][3]~2 ));
defparam \butterfly_st1[3][0][3]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st1[3][0][3]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[3][0][4]~1 (
	.dataa(\gen_cont:bfp_scale|r_array_out[1][4]~q ),
	.datab(\gen_cont:bfp_scale|r_array_out[3][4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[3][0][3]~2 ),
	.combout(\butterfly_st1[3][0][4]~1_combout ),
	.cout(\butterfly_st1[3][0][4]~2 ));
defparam \butterfly_st1[3][0][4]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st1[3][0][4]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[3][0][5]~1 (
	.dataa(\gen_cont:bfp_scale|r_array_out[1][5]~q ),
	.datab(\gen_cont:bfp_scale|r_array_out[3][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[3][0][4]~2 ),
	.combout(\butterfly_st1[3][0][5]~1_combout ),
	.cout(\butterfly_st1[3][0][5]~2 ));
defparam \butterfly_st1[3][0][5]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st1[3][0][5]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[3][0][6]~1 (
	.dataa(\gen_cont:bfp_scale|r_array_out[1][6]~q ),
	.datab(\gen_cont:bfp_scale|r_array_out[3][6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[3][0][5]~2 ),
	.combout(\butterfly_st1[3][0][6]~1_combout ),
	.cout(\butterfly_st1[3][0][6]~2 ));
defparam \butterfly_st1[3][0][6]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st1[3][0][6]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[3][0][7]~1 (
	.dataa(\gen_cont:bfp_scale|r_array_out[1][7]~q ),
	.datab(\gen_cont:bfp_scale|r_array_out[3][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[3][0][6]~2 ),
	.combout(\butterfly_st1[3][0][7]~1_combout ),
	.cout(\butterfly_st1[3][0][7]~2 ));
defparam \butterfly_st1[3][0][7]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st1[3][0][7]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[3][0][8]~1 (
	.dataa(\gen_cont:bfp_scale|r_array_out[1][7]~q ),
	.datab(\gen_cont:bfp_scale|r_array_out[3][7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\butterfly_st1[3][0][7]~2 ),
	.combout(\butterfly_st1[3][0][8]~1_combout ),
	.cout());
defparam \butterfly_st1[3][0][8]~1 .lut_mask = 16'h9696;
defparam \butterfly_st1[3][0][8]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[2][0][0]~1 (
	.dataa(\gen_cont:bfp_scale|r_array_out[0][0]~q ),
	.datab(\gen_cont:bfp_scale|r_array_out[2][0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\butterfly_st1[2][0][0]~1_combout ),
	.cout(\butterfly_st1[2][0][0]~2 ));
defparam \butterfly_st1[2][0][0]~1 .lut_mask = 16'h66BB;
defparam \butterfly_st1[2][0][0]~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \butterfly_st1[2][0][1]~1 (
	.dataa(\gen_cont:bfp_scale|r_array_out[0][1]~q ),
	.datab(\gen_cont:bfp_scale|r_array_out[2][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[2][0][0]~2 ),
	.combout(\butterfly_st1[2][0][1]~1_combout ),
	.cout(\butterfly_st1[2][0][1]~2 ));
defparam \butterfly_st1[2][0][1]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st1[2][0][1]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[2][0][2]~1 (
	.dataa(\gen_cont:bfp_scale|r_array_out[0][2]~q ),
	.datab(\gen_cont:bfp_scale|r_array_out[2][2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[2][0][1]~2 ),
	.combout(\butterfly_st1[2][0][2]~1_combout ),
	.cout(\butterfly_st1[2][0][2]~2 ));
defparam \butterfly_st1[2][0][2]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st1[2][0][2]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[3][1][0]~1 (
	.dataa(\gen_cont:bfp_scale|i_array_out[1][0]~q ),
	.datab(\gen_cont:bfp_scale|i_array_out[3][0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\butterfly_st1[3][1][0]~1_combout ),
	.cout(\butterfly_st1[3][1][0]~2 ));
defparam \butterfly_st1[3][1][0]~1 .lut_mask = 16'h66BB;
defparam \butterfly_st1[3][1][0]~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \butterfly_st1[3][1][1]~1 (
	.dataa(\gen_cont:bfp_scale|i_array_out[1][1]~q ),
	.datab(\gen_cont:bfp_scale|i_array_out[3][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[3][1][0]~2 ),
	.combout(\butterfly_st1[3][1][1]~1_combout ),
	.cout(\butterfly_st1[3][1][1]~2 ));
defparam \butterfly_st1[3][1][1]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st1[3][1][1]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[3][1][2]~1 (
	.dataa(\gen_cont:bfp_scale|i_array_out[1][2]~q ),
	.datab(\gen_cont:bfp_scale|i_array_out[3][2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[3][1][1]~2 ),
	.combout(\butterfly_st1[3][1][2]~1_combout ),
	.cout(\butterfly_st1[3][1][2]~2 ));
defparam \butterfly_st1[3][1][2]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st1[3][1][2]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[2][0][3]~1 (
	.dataa(\gen_cont:bfp_scale|r_array_out[0][3]~q ),
	.datab(\gen_cont:bfp_scale|r_array_out[2][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[2][0][2]~2 ),
	.combout(\butterfly_st1[2][0][3]~1_combout ),
	.cout(\butterfly_st1[2][0][3]~2 ));
defparam \butterfly_st1[2][0][3]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st1[2][0][3]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[2][0][4]~1 (
	.dataa(\gen_cont:bfp_scale|r_array_out[0][4]~q ),
	.datab(\gen_cont:bfp_scale|r_array_out[2][4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[2][0][3]~2 ),
	.combout(\butterfly_st1[2][0][4]~1_combout ),
	.cout(\butterfly_st1[2][0][4]~2 ));
defparam \butterfly_st1[2][0][4]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st1[2][0][4]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[2][0][5]~1 (
	.dataa(\gen_cont:bfp_scale|r_array_out[0][5]~q ),
	.datab(\gen_cont:bfp_scale|r_array_out[2][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[2][0][4]~2 ),
	.combout(\butterfly_st1[2][0][5]~1_combout ),
	.cout(\butterfly_st1[2][0][5]~2 ));
defparam \butterfly_st1[2][0][5]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st1[2][0][5]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[2][0][6]~1 (
	.dataa(\gen_cont:bfp_scale|r_array_out[0][6]~q ),
	.datab(\gen_cont:bfp_scale|r_array_out[2][6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[2][0][5]~2 ),
	.combout(\butterfly_st1[2][0][6]~1_combout ),
	.cout(\butterfly_st1[2][0][6]~2 ));
defparam \butterfly_st1[2][0][6]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st1[2][0][6]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[2][0][7]~1 (
	.dataa(\gen_cont:bfp_scale|r_array_out[0][7]~q ),
	.datab(\gen_cont:bfp_scale|r_array_out[2][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[2][0][6]~2 ),
	.combout(\butterfly_st1[2][0][7]~1_combout ),
	.cout(\butterfly_st1[2][0][7]~2 ));
defparam \butterfly_st1[2][0][7]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st1[2][0][7]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[2][0][8]~1 (
	.dataa(\gen_cont:bfp_scale|r_array_out[0][7]~q ),
	.datab(\gen_cont:bfp_scale|r_array_out[2][7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\butterfly_st1[2][0][7]~2 ),
	.combout(\butterfly_st1[2][0][8]~1_combout ),
	.cout());
defparam \butterfly_st1[2][0][8]~1 .lut_mask = 16'h9696;
defparam \butterfly_st1[2][0][8]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[3][1][3]~1 (
	.dataa(\gen_cont:bfp_scale|i_array_out[1][3]~q ),
	.datab(\gen_cont:bfp_scale|i_array_out[3][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[3][1][2]~2 ),
	.combout(\butterfly_st1[3][1][3]~1_combout ),
	.cout(\butterfly_st1[3][1][3]~2 ));
defparam \butterfly_st1[3][1][3]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st1[3][1][3]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[3][1][4]~1 (
	.dataa(\gen_cont:bfp_scale|i_array_out[1][4]~q ),
	.datab(\gen_cont:bfp_scale|i_array_out[3][4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[3][1][3]~2 ),
	.combout(\butterfly_st1[3][1][4]~1_combout ),
	.cout(\butterfly_st1[3][1][4]~2 ));
defparam \butterfly_st1[3][1][4]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st1[3][1][4]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[3][1][5]~1 (
	.dataa(\gen_cont:bfp_scale|i_array_out[1][5]~q ),
	.datab(\gen_cont:bfp_scale|i_array_out[3][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[3][1][4]~2 ),
	.combout(\butterfly_st1[3][1][5]~1_combout ),
	.cout(\butterfly_st1[3][1][5]~2 ));
defparam \butterfly_st1[3][1][5]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st1[3][1][5]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[3][1][6]~1 (
	.dataa(\gen_cont:bfp_scale|i_array_out[1][6]~q ),
	.datab(\gen_cont:bfp_scale|i_array_out[3][6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[3][1][5]~2 ),
	.combout(\butterfly_st1[3][1][6]~1_combout ),
	.cout(\butterfly_st1[3][1][6]~2 ));
defparam \butterfly_st1[3][1][6]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st1[3][1][6]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[3][1][7]~1 (
	.dataa(\gen_cont:bfp_scale|i_array_out[1][7]~q ),
	.datab(\gen_cont:bfp_scale|i_array_out[3][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[3][1][6]~2 ),
	.combout(\butterfly_st1[3][1][7]~1_combout ),
	.cout(\butterfly_st1[3][1][7]~2 ));
defparam \butterfly_st1[3][1][7]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st1[3][1][7]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \butterfly_st1[3][1][8]~1 (
	.dataa(\gen_cont:bfp_scale|i_array_out[1][7]~q ),
	.datab(\gen_cont:bfp_scale|i_array_out[3][7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\butterfly_st1[3][1][7]~2 ),
	.combout(\butterfly_st1[3][1][8]~1_combout ),
	.cout());
defparam \butterfly_st1[3][1][8]~1 .lut_mask = 16'h9696;
defparam \butterfly_st1[3][1][8]~1 .sum_lutc_input = "cin";

dffeas \reg_no_twiddle[0][0][1] (
	.clk(clk),
	.d(\reg_no_twiddle[0][0][1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[0][0][1]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[0][0][1] .is_wysiwyg = "true";
defparam \reg_no_twiddle[0][0][1] .power_up = "low";

dffeas \reg_no_twiddle[0][0][0] (
	.clk(clk),
	.d(\reg_no_twiddle[0][0][0]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[0][0][0]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[0][0][0] .is_wysiwyg = "true";
defparam \reg_no_twiddle[0][0][0] .power_up = "low";

dffeas \reg_no_twiddle[0][0][2] (
	.clk(clk),
	.d(\reg_no_twiddle[0][0][2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[0][0][2]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[0][0][2] .is_wysiwyg = "true";
defparam \reg_no_twiddle[0][0][2] .power_up = "low";

dffeas \reg_no_twiddle[0][1][1] (
	.clk(clk),
	.d(\reg_no_twiddle[0][1][1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[0][1][1]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[0][1][1] .is_wysiwyg = "true";
defparam \reg_no_twiddle[0][1][1] .power_up = "low";

dffeas \reg_no_twiddle[0][1][0] (
	.clk(clk),
	.d(\reg_no_twiddle[0][1][0]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[0][1][0]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[0][1][0] .is_wysiwyg = "true";
defparam \reg_no_twiddle[0][1][0] .power_up = "low";

dffeas \reg_no_twiddle[0][1][2] (
	.clk(clk),
	.d(\reg_no_twiddle[0][1][2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[0][1][2]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[0][1][2] .is_wysiwyg = "true";
defparam \reg_no_twiddle[0][1][2] .power_up = "low";

dffeas \reg_no_twiddle[6][0][3] (
	.clk(clk),
	.d(\reg_no_twiddle~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[6][0][3]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[6][0][3] .is_wysiwyg = "true";
defparam \reg_no_twiddle[6][0][3] .power_up = "low";

dffeas \reg_no_twiddle[6][0][7] (
	.clk(clk),
	.d(\reg_no_twiddle~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[6][0][7]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[6][0][7] .is_wysiwyg = "true";
defparam \reg_no_twiddle[6][0][7] .power_up = "low";

dffeas \reg_no_twiddle[6][1][7] (
	.clk(clk),
	.d(\reg_no_twiddle~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[6][1][7]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[6][1][7] .is_wysiwyg = "true";
defparam \reg_no_twiddle[6][1][7] .power_up = "low";

dffeas \reg_no_twiddle[6][1][3] (
	.clk(clk),
	.d(\reg_no_twiddle~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[6][1][3]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[6][1][3] .is_wysiwyg = "true";
defparam \reg_no_twiddle[6][1][3] .power_up = "low";

cycloneiii_lcell_comb \Selector3~0 (
	.dataa(\gain_out_4pts[0]~q ),
	.datab(\gen_cont:bfp_detect_1pt|gain_lut_8pts[0]~q ),
	.datac(gnd),
	.datad(\sdft.ENABLE_DFT_O~q ),
	.cin(gnd),
	.combout(\Selector3~0_combout ),
	.cout());
defparam \Selector3~0 .lut_mask = 16'hEEFF;
defparam \Selector3~0 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[6][0][4] (
	.clk(clk),
	.d(\reg_no_twiddle~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[6][0][4]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[6][0][4] .is_wysiwyg = "true";
defparam \reg_no_twiddle[6][0][4] .power_up = "low";

dffeas \reg_no_twiddle[6][1][4] (
	.clk(clk),
	.d(\reg_no_twiddle~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[6][1][4]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[6][1][4] .is_wysiwyg = "true";
defparam \reg_no_twiddle[6][1][4] .power_up = "low";

cycloneiii_lcell_comb \Selector2~0 (
	.dataa(\gain_out_4pts[1]~q ),
	.datab(\gen_cont:bfp_detect_1pt|gain_lut_8pts[1]~q ),
	.datac(gnd),
	.datad(\sdft.ENABLE_DFT_O~q ),
	.cin(gnd),
	.combout(\Selector2~0_combout ),
	.cout());
defparam \Selector2~0 .lut_mask = 16'hEEFF;
defparam \Selector2~0 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[6][0][5] (
	.clk(clk),
	.d(\reg_no_twiddle~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[6][0][5]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[6][0][5] .is_wysiwyg = "true";
defparam \reg_no_twiddle[6][0][5] .power_up = "low";

dffeas \reg_no_twiddle[6][1][5] (
	.clk(clk),
	.d(\reg_no_twiddle~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[6][1][5]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[6][1][5] .is_wysiwyg = "true";
defparam \reg_no_twiddle[6][1][5] .power_up = "low";

cycloneiii_lcell_comb \Selector1~0 (
	.dataa(\gain_out_4pts[2]~q ),
	.datab(\gen_cont:bfp_detect_1pt|gain_lut_8pts[2]~q ),
	.datac(gnd),
	.datad(\sdft.ENABLE_DFT_O~q ),
	.cin(gnd),
	.combout(\Selector1~0_combout ),
	.cout());
defparam \Selector1~0 .lut_mask = 16'hEEFF;
defparam \Selector1~0 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[6][0][6] (
	.clk(clk),
	.d(\reg_no_twiddle~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[6][0][6]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[6][0][6] .is_wysiwyg = "true";
defparam \reg_no_twiddle[6][0][6] .power_up = "low";

dffeas \reg_no_twiddle[6][1][6] (
	.clk(clk),
	.d(\reg_no_twiddle~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[6][1][6]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[6][1][6] .is_wysiwyg = "true";
defparam \reg_no_twiddle[6][1][6] .power_up = "low";

cycloneiii_lcell_comb \Selector0~0 (
	.dataa(\gain_out_4pts[3]~q ),
	.datab(\gen_cont:bfp_detect_1pt|gain_lut_8pts[3]~q ),
	.datac(gnd),
	.datad(\sdft.ENABLE_DFT_O~q ),
	.cin(gnd),
	.combout(\Selector0~0_combout ),
	.cout());
defparam \Selector0~0 .lut_mask = 16'hEEFF;
defparam \Selector0~0 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[5][0][3] (
	.clk(clk),
	.d(\reg_no_twiddle~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[5][0][3]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[5][0][3] .is_wysiwyg = "true";
defparam \reg_no_twiddle[5][0][3] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~0 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[5][0][3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~0_combout ),
	.cout());
defparam \reg_no_twiddle~0 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~0 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[5][0][7] (
	.clk(clk),
	.d(\reg_no_twiddle~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[5][0][7]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[5][0][7] .is_wysiwyg = "true";
defparam \reg_no_twiddle[5][0][7] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~1 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[5][0][7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~1_combout ),
	.cout());
defparam \reg_no_twiddle~1 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~1 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[5][1][7] (
	.clk(clk),
	.d(\reg_no_twiddle~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[5][1][7]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[5][1][7] .is_wysiwyg = "true";
defparam \reg_no_twiddle[5][1][7] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~2 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[5][1][7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~2_combout ),
	.cout());
defparam \reg_no_twiddle~2 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~2 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[5][1][3] (
	.clk(clk),
	.d(\reg_no_twiddle~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[5][1][3]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[5][1][3] .is_wysiwyg = "true";
defparam \reg_no_twiddle[5][1][3] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~3 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[5][1][3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~3_combout ),
	.cout());
defparam \reg_no_twiddle~3 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~3 .sum_lutc_input = "datac";

dffeas enable_op(
	.clk(clk),
	.d(\scale_dft_o_en~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\enable_op~q ),
	.prn(vcc));
defparam enable_op.is_wysiwyg = "true";
defparam enable_op.power_up = "low";

dffeas \sdft.WAIT_FOR_OUTPUT (
	.clk(clk),
	.d(\sdft~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sdft.WAIT_FOR_OUTPUT~q ),
	.prn(vcc));
defparam \sdft.WAIT_FOR_OUTPUT .is_wysiwyg = "true";
defparam \sdft.WAIT_FOR_OUTPUT .power_up = "low";

cycloneiii_lcell_comb \Selector14~0 (
	.dataa(gnd),
	.datab(\sdft.ENABLE_DFT_O~q ),
	.datac(\gap_reg~q ),
	.datad(\sdft.WAIT_FOR_OUTPUT~q ),
	.cin(gnd),
	.combout(\Selector14~0_combout ),
	.cout());
defparam \Selector14~0 .lut_mask = 16'hFFFC;
defparam \Selector14~0 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[5][0][4] (
	.clk(clk),
	.d(\reg_no_twiddle~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[5][0][4]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[5][0][4] .is_wysiwyg = "true";
defparam \reg_no_twiddle[5][0][4] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~4 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[5][0][4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~4_combout ),
	.cout());
defparam \reg_no_twiddle~4 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~4 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[5][1][4] (
	.clk(clk),
	.d(\reg_no_twiddle~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[5][1][4]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[5][1][4] .is_wysiwyg = "true";
defparam \reg_no_twiddle[5][1][4] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~5 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[5][1][4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~5_combout ),
	.cout());
defparam \reg_no_twiddle~5 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~5 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[5][0][5] (
	.clk(clk),
	.d(\reg_no_twiddle~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[5][0][5]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[5][0][5] .is_wysiwyg = "true";
defparam \reg_no_twiddle[5][0][5] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~6 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[5][0][5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~6_combout ),
	.cout());
defparam \reg_no_twiddle~6 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~6 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[5][1][5] (
	.clk(clk),
	.d(\reg_no_twiddle~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[5][1][5]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[5][1][5] .is_wysiwyg = "true";
defparam \reg_no_twiddle[5][1][5] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~7 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[5][1][5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~7_combout ),
	.cout());
defparam \reg_no_twiddle~7 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~7 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[5][0][6] (
	.clk(clk),
	.d(\reg_no_twiddle~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[5][0][6]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[5][0][6] .is_wysiwyg = "true";
defparam \reg_no_twiddle[5][0][6] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~8 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[5][0][6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~8_combout ),
	.cout());
defparam \reg_no_twiddle~8 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~8 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[5][1][6] (
	.clk(clk),
	.d(\reg_no_twiddle~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[5][1][6]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[5][1][6] .is_wysiwyg = "true";
defparam \reg_no_twiddle[5][1][6] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~9 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[5][1][6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~9_combout ),
	.cout());
defparam \reg_no_twiddle~9 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~9 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[4][0][3] (
	.clk(clk),
	.d(\reg_no_twiddle~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[4][0][3]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[4][0][3] .is_wysiwyg = "true";
defparam \reg_no_twiddle[4][0][3] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~10 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[4][0][3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~10_combout ),
	.cout());
defparam \reg_no_twiddle~10 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~10 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[4][0][7] (
	.clk(clk),
	.d(\reg_no_twiddle~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[4][0][7]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[4][0][7] .is_wysiwyg = "true";
defparam \reg_no_twiddle[4][0][7] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~11 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[4][0][7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~11_combout ),
	.cout());
defparam \reg_no_twiddle~11 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~11 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[4][1][7] (
	.clk(clk),
	.d(\reg_no_twiddle~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[4][1][7]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[4][1][7] .is_wysiwyg = "true";
defparam \reg_no_twiddle[4][1][7] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~12 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[4][1][7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~12_combout ),
	.cout());
defparam \reg_no_twiddle~12 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~12 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[4][1][3] (
	.clk(clk),
	.d(\reg_no_twiddle~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[4][1][3]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[4][1][3] .is_wysiwyg = "true";
defparam \reg_no_twiddle[4][1][3] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~13 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[4][1][3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~13_combout ),
	.cout());
defparam \reg_no_twiddle~13 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~13 .sum_lutc_input = "datac";

dffeas scale_dft_o_en(
	.clk(clk),
	.d(\Selector5~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\scale_dft_o_en~q ),
	.prn(vcc));
defparam scale_dft_o_en.is_wysiwyg = "true";
defparam scale_dft_o_en.power_up = "low";

dffeas \do_tdl[0][0][3][3] (
	.clk(clk),
	.d(\do_tdl[0][0][2][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][0][3][3]~q ),
	.prn(vcc));
defparam \do_tdl[0][0][3][3] .is_wysiwyg = "true";
defparam \do_tdl[0][0][3][3] .power_up = "low";

dffeas \do_tdl[0][0][3][7] (
	.clk(clk),
	.d(\do_tdl[0][0][2][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][0][3][7]~q ),
	.prn(vcc));
defparam \do_tdl[0][0][3][7] .is_wysiwyg = "true";
defparam \do_tdl[0][0][3][7] .power_up = "low";

dffeas \do_tdl[0][0][3][4] (
	.clk(clk),
	.d(\do_tdl[0][0][2][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][0][3][4]~q ),
	.prn(vcc));
defparam \do_tdl[0][0][3][4] .is_wysiwyg = "true";
defparam \do_tdl[0][0][3][4] .power_up = "low";

dffeas \do_tdl[0][0][3][5] (
	.clk(clk),
	.d(\do_tdl[0][0][2][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][0][3][5]~q ),
	.prn(vcc));
defparam \do_tdl[0][0][3][5] .is_wysiwyg = "true";
defparam \do_tdl[0][0][3][5] .power_up = "low";

dffeas \do_tdl[0][0][3][6] (
	.clk(clk),
	.d(\do_tdl[0][0][2][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][0][3][6]~q ),
	.prn(vcc));
defparam \do_tdl[0][0][3][6] .is_wysiwyg = "true";
defparam \do_tdl[0][0][3][6] .power_up = "low";

dffeas \do_tdl[0][0][3][1] (
	.clk(clk),
	.d(\do_tdl[0][0][2][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][0][3][1]~q ),
	.prn(vcc));
defparam \do_tdl[0][0][3][1] .is_wysiwyg = "true";
defparam \do_tdl[0][0][3][1] .power_up = "low";

dffeas \do_tdl[0][0][3][0] (
	.clk(clk),
	.d(\do_tdl[0][0][2][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][0][3][0]~q ),
	.prn(vcc));
defparam \do_tdl[0][0][3][0] .is_wysiwyg = "true";
defparam \do_tdl[0][0][3][0] .power_up = "low";

cycloneiii_lcell_comb \slb_1pt[0] (
	.dataa(slb_last_0),
	.datab(\scale_dft_o_en~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\slb_1pt[0]~combout ),
	.cout());
defparam \slb_1pt[0] .lut_mask = 16'hEEEE;
defparam \slb_1pt[0] .sum_lutc_input = "datac";

dffeas \do_tdl[0][0][3][2] (
	.clk(clk),
	.d(\do_tdl[0][0][2][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][0][3][2]~q ),
	.prn(vcc));
defparam \do_tdl[0][0][3][2] .is_wysiwyg = "true";
defparam \do_tdl[0][0][3][2] .power_up = "low";

cycloneiii_lcell_comb \slb_1pt[2]~0 (
	.dataa(slb_last_2),
	.datab(\scale_dft_o_en~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\slb_1pt[2]~0_combout ),
	.cout());
defparam \slb_1pt[2]~0 .lut_mask = 16'hEEEE;
defparam \slb_1pt[2]~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \slb_1pt[1] (
	.dataa(gnd),
	.datab(gnd),
	.datac(slb_last_1),
	.datad(\scale_dft_o_en~q ),
	.cin(gnd),
	.combout(\slb_1pt[1]~combout ),
	.cout());
defparam \slb_1pt[1] .lut_mask = 16'h0FFF;
defparam \slb_1pt[1] .sum_lutc_input = "datac";

dffeas \do_tdl[0][1][3][3] (
	.clk(clk),
	.d(\do_tdl[0][1][2][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][1][3][3]~q ),
	.prn(vcc));
defparam \do_tdl[0][1][3][3] .is_wysiwyg = "true";
defparam \do_tdl[0][1][3][3] .power_up = "low";

dffeas \do_tdl[0][1][3][7] (
	.clk(clk),
	.d(\do_tdl[0][1][2][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][1][3][7]~q ),
	.prn(vcc));
defparam \do_tdl[0][1][3][7] .is_wysiwyg = "true";
defparam \do_tdl[0][1][3][7] .power_up = "low";

dffeas \do_tdl[0][1][3][4] (
	.clk(clk),
	.d(\do_tdl[0][1][2][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][1][3][4]~q ),
	.prn(vcc));
defparam \do_tdl[0][1][3][4] .is_wysiwyg = "true";
defparam \do_tdl[0][1][3][4] .power_up = "low";

dffeas \do_tdl[0][1][3][5] (
	.clk(clk),
	.d(\do_tdl[0][1][2][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][1][3][5]~q ),
	.prn(vcc));
defparam \do_tdl[0][1][3][5] .is_wysiwyg = "true";
defparam \do_tdl[0][1][3][5] .power_up = "low";

dffeas \do_tdl[0][1][3][6] (
	.clk(clk),
	.d(\do_tdl[0][1][2][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][1][3][6]~q ),
	.prn(vcc));
defparam \do_tdl[0][1][3][6] .is_wysiwyg = "true";
defparam \do_tdl[0][1][3][6] .power_up = "low";

dffeas \do_tdl[0][1][3][1] (
	.clk(clk),
	.d(\do_tdl[0][1][2][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][1][3][1]~q ),
	.prn(vcc));
defparam \do_tdl[0][1][3][1] .is_wysiwyg = "true";
defparam \do_tdl[0][1][3][1] .power_up = "low";

dffeas \do_tdl[0][1][3][0] (
	.clk(clk),
	.d(\do_tdl[0][1][2][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][1][3][0]~q ),
	.prn(vcc));
defparam \do_tdl[0][1][3][0] .is_wysiwyg = "true";
defparam \do_tdl[0][1][3][0] .power_up = "low";

dffeas \do_tdl[0][1][3][2] (
	.clk(clk),
	.d(\do_tdl[0][1][2][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][1][3][2]~q ),
	.prn(vcc));
defparam \do_tdl[0][1][3][2] .is_wysiwyg = "true";
defparam \do_tdl[0][1][3][2] .power_up = "low";

dffeas \do_tdl[1][0][3][3] (
	.clk(clk),
	.d(\do_tdl[1][0][2][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][0][3][3]~q ),
	.prn(vcc));
defparam \do_tdl[1][0][3][3] .is_wysiwyg = "true";
defparam \do_tdl[1][0][3][3] .power_up = "low";

dffeas \do_tdl[1][0][3][7] (
	.clk(clk),
	.d(\do_tdl[1][0][2][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][0][3][7]~q ),
	.prn(vcc));
defparam \do_tdl[1][0][3][7] .is_wysiwyg = "true";
defparam \do_tdl[1][0][3][7] .power_up = "low";

dffeas \do_tdl[1][0][3][4] (
	.clk(clk),
	.d(\do_tdl[1][0][2][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][0][3][4]~q ),
	.prn(vcc));
defparam \do_tdl[1][0][3][4] .is_wysiwyg = "true";
defparam \do_tdl[1][0][3][4] .power_up = "low";

dffeas \do_tdl[1][0][3][5] (
	.clk(clk),
	.d(\do_tdl[1][0][2][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][0][3][5]~q ),
	.prn(vcc));
defparam \do_tdl[1][0][3][5] .is_wysiwyg = "true";
defparam \do_tdl[1][0][3][5] .power_up = "low";

dffeas \do_tdl[1][0][3][6] (
	.clk(clk),
	.d(\do_tdl[1][0][2][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][0][3][6]~q ),
	.prn(vcc));
defparam \do_tdl[1][0][3][6] .is_wysiwyg = "true";
defparam \do_tdl[1][0][3][6] .power_up = "low";

dffeas \do_tdl[1][0][3][1] (
	.clk(clk),
	.d(\do_tdl[1][0][2][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][0][3][1]~q ),
	.prn(vcc));
defparam \do_tdl[1][0][3][1] .is_wysiwyg = "true";
defparam \do_tdl[1][0][3][1] .power_up = "low";

dffeas \do_tdl[1][0][3][0] (
	.clk(clk),
	.d(\do_tdl[1][0][2][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][0][3][0]~q ),
	.prn(vcc));
defparam \do_tdl[1][0][3][0] .is_wysiwyg = "true";
defparam \do_tdl[1][0][3][0] .power_up = "low";

dffeas \do_tdl[1][0][3][2] (
	.clk(clk),
	.d(\do_tdl[1][0][2][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][0][3][2]~q ),
	.prn(vcc));
defparam \do_tdl[1][0][3][2] .is_wysiwyg = "true";
defparam \do_tdl[1][0][3][2] .power_up = "low";

dffeas \do_tdl[1][1][3][3] (
	.clk(clk),
	.d(\do_tdl[1][1][2][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][1][3][3]~q ),
	.prn(vcc));
defparam \do_tdl[1][1][3][3] .is_wysiwyg = "true";
defparam \do_tdl[1][1][3][3] .power_up = "low";

dffeas \do_tdl[1][1][3][7] (
	.clk(clk),
	.d(\do_tdl[1][1][2][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][1][3][7]~q ),
	.prn(vcc));
defparam \do_tdl[1][1][3][7] .is_wysiwyg = "true";
defparam \do_tdl[1][1][3][7] .power_up = "low";

dffeas \do_tdl[1][1][3][4] (
	.clk(clk),
	.d(\do_tdl[1][1][2][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][1][3][4]~q ),
	.prn(vcc));
defparam \do_tdl[1][1][3][4] .is_wysiwyg = "true";
defparam \do_tdl[1][1][3][4] .power_up = "low";

dffeas \do_tdl[1][1][3][5] (
	.clk(clk),
	.d(\do_tdl[1][1][2][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][1][3][5]~q ),
	.prn(vcc));
defparam \do_tdl[1][1][3][5] .is_wysiwyg = "true";
defparam \do_tdl[1][1][3][5] .power_up = "low";

dffeas \do_tdl[1][1][3][6] (
	.clk(clk),
	.d(\do_tdl[1][1][2][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][1][3][6]~q ),
	.prn(vcc));
defparam \do_tdl[1][1][3][6] .is_wysiwyg = "true";
defparam \do_tdl[1][1][3][6] .power_up = "low";

dffeas \do_tdl[1][1][3][1] (
	.clk(clk),
	.d(\do_tdl[1][1][2][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][1][3][1]~q ),
	.prn(vcc));
defparam \do_tdl[1][1][3][1] .is_wysiwyg = "true";
defparam \do_tdl[1][1][3][1] .power_up = "low";

dffeas \do_tdl[1][1][3][0] (
	.clk(clk),
	.d(\do_tdl[1][1][2][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][1][3][0]~q ),
	.prn(vcc));
defparam \do_tdl[1][1][3][0] .is_wysiwyg = "true";
defparam \do_tdl[1][1][3][0] .power_up = "low";

dffeas \do_tdl[1][1][3][2] (
	.clk(clk),
	.d(\do_tdl[1][1][2][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][1][3][2]~q ),
	.prn(vcc));
defparam \do_tdl[1][1][3][2] .is_wysiwyg = "true";
defparam \do_tdl[1][1][3][2] .power_up = "low";

dffeas \do_tdl[2][0][3][3] (
	.clk(clk),
	.d(\do_tdl[2][0][2][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][0][3][3]~q ),
	.prn(vcc));
defparam \do_tdl[2][0][3][3] .is_wysiwyg = "true";
defparam \do_tdl[2][0][3][3] .power_up = "low";

dffeas \do_tdl[2][0][3][7] (
	.clk(clk),
	.d(\do_tdl[2][0][2][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][0][3][7]~q ),
	.prn(vcc));
defparam \do_tdl[2][0][3][7] .is_wysiwyg = "true";
defparam \do_tdl[2][0][3][7] .power_up = "low";

dffeas \do_tdl[2][0][3][4] (
	.clk(clk),
	.d(\do_tdl[2][0][2][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][0][3][4]~q ),
	.prn(vcc));
defparam \do_tdl[2][0][3][4] .is_wysiwyg = "true";
defparam \do_tdl[2][0][3][4] .power_up = "low";

dffeas \do_tdl[2][0][3][5] (
	.clk(clk),
	.d(\do_tdl[2][0][2][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][0][3][5]~q ),
	.prn(vcc));
defparam \do_tdl[2][0][3][5] .is_wysiwyg = "true";
defparam \do_tdl[2][0][3][5] .power_up = "low";

dffeas \do_tdl[2][0][3][6] (
	.clk(clk),
	.d(\do_tdl[2][0][2][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][0][3][6]~q ),
	.prn(vcc));
defparam \do_tdl[2][0][3][6] .is_wysiwyg = "true";
defparam \do_tdl[2][0][3][6] .power_up = "low";

dffeas \do_tdl[2][0][3][1] (
	.clk(clk),
	.d(\do_tdl[2][0][2][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][0][3][1]~q ),
	.prn(vcc));
defparam \do_tdl[2][0][3][1] .is_wysiwyg = "true";
defparam \do_tdl[2][0][3][1] .power_up = "low";

dffeas \do_tdl[2][0][3][0] (
	.clk(clk),
	.d(\do_tdl[2][0][2][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][0][3][0]~q ),
	.prn(vcc));
defparam \do_tdl[2][0][3][0] .is_wysiwyg = "true";
defparam \do_tdl[2][0][3][0] .power_up = "low";

dffeas \do_tdl[2][0][3][2] (
	.clk(clk),
	.d(\do_tdl[2][0][2][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][0][3][2]~q ),
	.prn(vcc));
defparam \do_tdl[2][0][3][2] .is_wysiwyg = "true";
defparam \do_tdl[2][0][3][2] .power_up = "low";

dffeas \do_tdl[2][1][3][3] (
	.clk(clk),
	.d(\do_tdl[2][1][2][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][1][3][3]~q ),
	.prn(vcc));
defparam \do_tdl[2][1][3][3] .is_wysiwyg = "true";
defparam \do_tdl[2][1][3][3] .power_up = "low";

dffeas \do_tdl[2][1][3][7] (
	.clk(clk),
	.d(\do_tdl[2][1][2][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][1][3][7]~q ),
	.prn(vcc));
defparam \do_tdl[2][1][3][7] .is_wysiwyg = "true";
defparam \do_tdl[2][1][3][7] .power_up = "low";

dffeas \do_tdl[2][1][3][4] (
	.clk(clk),
	.d(\do_tdl[2][1][2][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][1][3][4]~q ),
	.prn(vcc));
defparam \do_tdl[2][1][3][4] .is_wysiwyg = "true";
defparam \do_tdl[2][1][3][4] .power_up = "low";

dffeas \do_tdl[2][1][3][5] (
	.clk(clk),
	.d(\do_tdl[2][1][2][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][1][3][5]~q ),
	.prn(vcc));
defparam \do_tdl[2][1][3][5] .is_wysiwyg = "true";
defparam \do_tdl[2][1][3][5] .power_up = "low";

dffeas \do_tdl[2][1][3][6] (
	.clk(clk),
	.d(\do_tdl[2][1][2][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][1][3][6]~q ),
	.prn(vcc));
defparam \do_tdl[2][1][3][6] .is_wysiwyg = "true";
defparam \do_tdl[2][1][3][6] .power_up = "low";

dffeas \do_tdl[2][1][3][1] (
	.clk(clk),
	.d(\do_tdl[2][1][2][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][1][3][1]~q ),
	.prn(vcc));
defparam \do_tdl[2][1][3][1] .is_wysiwyg = "true";
defparam \do_tdl[2][1][3][1] .power_up = "low";

dffeas \do_tdl[2][1][3][0] (
	.clk(clk),
	.d(\do_tdl[2][1][2][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][1][3][0]~q ),
	.prn(vcc));
defparam \do_tdl[2][1][3][0] .is_wysiwyg = "true";
defparam \do_tdl[2][1][3][0] .power_up = "low";

dffeas \do_tdl[2][1][3][2] (
	.clk(clk),
	.d(\do_tdl[2][1][2][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][1][3][2]~q ),
	.prn(vcc));
defparam \do_tdl[2][1][3][2] .is_wysiwyg = "true";
defparam \do_tdl[2][1][3][2] .power_up = "low";

dffeas \do_tdl[3][0][3][3] (
	.clk(clk),
	.d(\do_tdl[3][0][2][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][0][3][3]~q ),
	.prn(vcc));
defparam \do_tdl[3][0][3][3] .is_wysiwyg = "true";
defparam \do_tdl[3][0][3][3] .power_up = "low";

dffeas \do_tdl[3][0][3][7] (
	.clk(clk),
	.d(\do_tdl[3][0][2][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][0][3][7]~q ),
	.prn(vcc));
defparam \do_tdl[3][0][3][7] .is_wysiwyg = "true";
defparam \do_tdl[3][0][3][7] .power_up = "low";

dffeas \do_tdl[3][0][3][4] (
	.clk(clk),
	.d(\do_tdl[3][0][2][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][0][3][4]~q ),
	.prn(vcc));
defparam \do_tdl[3][0][3][4] .is_wysiwyg = "true";
defparam \do_tdl[3][0][3][4] .power_up = "low";

dffeas \do_tdl[3][0][3][5] (
	.clk(clk),
	.d(\do_tdl[3][0][2][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][0][3][5]~q ),
	.prn(vcc));
defparam \do_tdl[3][0][3][5] .is_wysiwyg = "true";
defparam \do_tdl[3][0][3][5] .power_up = "low";

dffeas \do_tdl[3][0][3][6] (
	.clk(clk),
	.d(\do_tdl[3][0][2][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][0][3][6]~q ),
	.prn(vcc));
defparam \do_tdl[3][0][3][6] .is_wysiwyg = "true";
defparam \do_tdl[3][0][3][6] .power_up = "low";

dffeas \do_tdl[3][0][3][1] (
	.clk(clk),
	.d(\do_tdl[3][0][2][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][0][3][1]~q ),
	.prn(vcc));
defparam \do_tdl[3][0][3][1] .is_wysiwyg = "true";
defparam \do_tdl[3][0][3][1] .power_up = "low";

dffeas \do_tdl[3][0][3][0] (
	.clk(clk),
	.d(\do_tdl[3][0][2][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][0][3][0]~q ),
	.prn(vcc));
defparam \do_tdl[3][0][3][0] .is_wysiwyg = "true";
defparam \do_tdl[3][0][3][0] .power_up = "low";

dffeas \do_tdl[3][0][3][2] (
	.clk(clk),
	.d(\do_tdl[3][0][2][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][0][3][2]~q ),
	.prn(vcc));
defparam \do_tdl[3][0][3][2] .is_wysiwyg = "true";
defparam \do_tdl[3][0][3][2] .power_up = "low";

dffeas \do_tdl[3][1][3][3] (
	.clk(clk),
	.d(\do_tdl[3][1][2][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][1][3][3]~q ),
	.prn(vcc));
defparam \do_tdl[3][1][3][3] .is_wysiwyg = "true";
defparam \do_tdl[3][1][3][3] .power_up = "low";

dffeas \do_tdl[3][1][3][7] (
	.clk(clk),
	.d(\do_tdl[3][1][2][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][1][3][7]~q ),
	.prn(vcc));
defparam \do_tdl[3][1][3][7] .is_wysiwyg = "true";
defparam \do_tdl[3][1][3][7] .power_up = "low";

dffeas \do_tdl[3][1][3][4] (
	.clk(clk),
	.d(\do_tdl[3][1][2][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][1][3][4]~q ),
	.prn(vcc));
defparam \do_tdl[3][1][3][4] .is_wysiwyg = "true";
defparam \do_tdl[3][1][3][4] .power_up = "low";

dffeas \do_tdl[3][1][3][5] (
	.clk(clk),
	.d(\do_tdl[3][1][2][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][1][3][5]~q ),
	.prn(vcc));
defparam \do_tdl[3][1][3][5] .is_wysiwyg = "true";
defparam \do_tdl[3][1][3][5] .power_up = "low";

dffeas \do_tdl[3][1][3][6] (
	.clk(clk),
	.d(\do_tdl[3][1][2][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][1][3][6]~q ),
	.prn(vcc));
defparam \do_tdl[3][1][3][6] .is_wysiwyg = "true";
defparam \do_tdl[3][1][3][6] .power_up = "low";

dffeas \do_tdl[3][1][3][1] (
	.clk(clk),
	.d(\do_tdl[3][1][2][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][1][3][1]~q ),
	.prn(vcc));
defparam \do_tdl[3][1][3][1] .is_wysiwyg = "true";
defparam \do_tdl[3][1][3][1] .power_up = "low";

dffeas \do_tdl[3][1][3][0] (
	.clk(clk),
	.d(\do_tdl[3][1][2][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][1][3][0]~q ),
	.prn(vcc));
defparam \do_tdl[3][1][3][0] .is_wysiwyg = "true";
defparam \do_tdl[3][1][3][0] .power_up = "low";

dffeas \do_tdl[3][1][3][2] (
	.clk(clk),
	.d(\do_tdl[3][1][2][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][1][3][2]~q ),
	.prn(vcc));
defparam \do_tdl[3][1][3][2] .is_wysiwyg = "true";
defparam \do_tdl[3][1][3][2] .power_up = "low";

cycloneiii_lcell_comb \gap_reg~0 (
	.dataa(tdl_arr_5),
	.datab(\gap_reg~q ),
	.datac(gnd),
	.datad(\gen_cont:delay_next_blk|tdl_arr[25]~q ),
	.cin(gnd),
	.combout(\gap_reg~0_combout ),
	.cout());
defparam \gap_reg~0 .lut_mask = 16'hEEFF;
defparam \gap_reg~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Equal0~0 (
	.dataa(\state_cnt[2]~q ),
	.datab(\state_cnt[3]~q ),
	.datac(\state_cnt[4]~q ),
	.datad(\state_cnt[5]~q ),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
defparam \Equal0~0 .lut_mask = 16'hEFFF;
defparam \Equal0~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Equal0~1 (
	.dataa(\Equal0~0_combout ),
	.datab(\state_cnt[0]~q ),
	.datac(gnd),
	.datad(\state_cnt[1]~q ),
	.cin(gnd),
	.combout(\Equal0~1_combout ),
	.cout());
defparam \Equal0~1 .lut_mask = 16'hEEFF;
defparam \Equal0~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sdft~8 (
	.dataa(reset_n),
	.datab(\Equal0~1_combout ),
	.datac(\sdft.BLOCK_DFT_I~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\sdft~8_combout ),
	.cout());
defparam \sdft~8 .lut_mask = 16'hFEFE;
defparam \sdft~8 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[4][0][4] (
	.clk(clk),
	.d(\reg_no_twiddle~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[4][0][4]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[4][0][4] .is_wysiwyg = "true";
defparam \reg_no_twiddle[4][0][4] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~14 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[4][0][4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~14_combout ),
	.cout());
defparam \reg_no_twiddle~14 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~14 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[4][1][4] (
	.clk(clk),
	.d(\reg_no_twiddle~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[4][1][4]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[4][1][4] .is_wysiwyg = "true";
defparam \reg_no_twiddle[4][1][4] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~15 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[4][1][4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~15_combout ),
	.cout());
defparam \reg_no_twiddle~15 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~15 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[4][0][5] (
	.clk(clk),
	.d(\reg_no_twiddle~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[4][0][5]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[4][0][5] .is_wysiwyg = "true";
defparam \reg_no_twiddle[4][0][5] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~16 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[4][0][5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~16_combout ),
	.cout());
defparam \reg_no_twiddle~16 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~16 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[4][1][5] (
	.clk(clk),
	.d(\reg_no_twiddle~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[4][1][5]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[4][1][5] .is_wysiwyg = "true";
defparam \reg_no_twiddle[4][1][5] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~17 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[4][1][5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~17_combout ),
	.cout());
defparam \reg_no_twiddle~17 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~17 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[4][0][6] (
	.clk(clk),
	.d(\reg_no_twiddle~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[4][0][6]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[4][0][6] .is_wysiwyg = "true";
defparam \reg_no_twiddle[4][0][6] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~18 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[4][0][6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~18_combout ),
	.cout());
defparam \reg_no_twiddle~18 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~18 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[4][1][6] (
	.clk(clk),
	.d(\reg_no_twiddle~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[4][1][6]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[4][1][6] .is_wysiwyg = "true";
defparam \reg_no_twiddle[4][1][6] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~19 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[4][1][6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~19_combout ),
	.cout());
defparam \reg_no_twiddle~19 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~19 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[3][0][3] (
	.clk(clk),
	.d(\reg_no_twiddle~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[3][0][3]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[3][0][3] .is_wysiwyg = "true";
defparam \reg_no_twiddle[3][0][3] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~20 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[3][0][3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~20_combout ),
	.cout());
defparam \reg_no_twiddle~20 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~20 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[3][0][7] (
	.clk(clk),
	.d(\reg_no_twiddle~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[3][0][7]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[3][0][7] .is_wysiwyg = "true";
defparam \reg_no_twiddle[3][0][7] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~21 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[3][0][7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~21_combout ),
	.cout());
defparam \reg_no_twiddle~21 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~21 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[3][1][7] (
	.clk(clk),
	.d(\reg_no_twiddle~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[3][1][7]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[3][1][7] .is_wysiwyg = "true";
defparam \reg_no_twiddle[3][1][7] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~22 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[3][1][7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~22_combout ),
	.cout());
defparam \reg_no_twiddle~22 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~22 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[3][1][3] (
	.clk(clk),
	.d(\reg_no_twiddle~33_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[3][1][3]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[3][1][3] .is_wysiwyg = "true";
defparam \reg_no_twiddle[3][1][3] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~23 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[3][1][3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~23_combout ),
	.cout());
defparam \reg_no_twiddle~23 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~23 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector5~0 (
	.dataa(\sdft.ENABLE_BFP_O~q ),
	.datab(\sdft.ENABLE_DFT_O~q ),
	.datac(gnd),
	.datad(\gap_reg~q ),
	.cin(gnd),
	.combout(\Selector5~0_combout ),
	.cout());
defparam \Selector5~0 .lut_mask = 16'hEEFF;
defparam \Selector5~0 .sum_lutc_input = "datac";

dffeas \do_tdl[0][0][2][3] (
	.clk(clk),
	.d(\do_tdl[0][0][1][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][0][2][3]~q ),
	.prn(vcc));
defparam \do_tdl[0][0][2][3] .is_wysiwyg = "true";
defparam \do_tdl[0][0][2][3] .power_up = "low";

dffeas \do_tdl[0][0][2][7] (
	.clk(clk),
	.d(\do_tdl[0][0][1][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][0][2][7]~q ),
	.prn(vcc));
defparam \do_tdl[0][0][2][7] .is_wysiwyg = "true";
defparam \do_tdl[0][0][2][7] .power_up = "low";

dffeas \do_tdl[0][0][2][4] (
	.clk(clk),
	.d(\do_tdl[0][0][1][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][0][2][4]~q ),
	.prn(vcc));
defparam \do_tdl[0][0][2][4] .is_wysiwyg = "true";
defparam \do_tdl[0][0][2][4] .power_up = "low";

dffeas \do_tdl[0][0][2][5] (
	.clk(clk),
	.d(\do_tdl[0][0][1][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][0][2][5]~q ),
	.prn(vcc));
defparam \do_tdl[0][0][2][5] .is_wysiwyg = "true";
defparam \do_tdl[0][0][2][5] .power_up = "low";

dffeas \do_tdl[0][0][2][6] (
	.clk(clk),
	.d(\do_tdl[0][0][1][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][0][2][6]~q ),
	.prn(vcc));
defparam \do_tdl[0][0][2][6] .is_wysiwyg = "true";
defparam \do_tdl[0][0][2][6] .power_up = "low";

dffeas \do_tdl[0][0][2][1] (
	.clk(clk),
	.d(\do_tdl[0][0][1][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][0][2][1]~q ),
	.prn(vcc));
defparam \do_tdl[0][0][2][1] .is_wysiwyg = "true";
defparam \do_tdl[0][0][2][1] .power_up = "low";

dffeas \do_tdl[0][0][2][0] (
	.clk(clk),
	.d(\do_tdl[0][0][1][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][0][2][0]~q ),
	.prn(vcc));
defparam \do_tdl[0][0][2][0] .is_wysiwyg = "true";
defparam \do_tdl[0][0][2][0] .power_up = "low";

dffeas \do_tdl[0][0][2][2] (
	.clk(clk),
	.d(\do_tdl[0][0][1][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][0][2][2]~q ),
	.prn(vcc));
defparam \do_tdl[0][0][2][2] .is_wysiwyg = "true";
defparam \do_tdl[0][0][2][2] .power_up = "low";

dffeas \do_tdl[0][1][2][3] (
	.clk(clk),
	.d(\do_tdl[0][1][1][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][1][2][3]~q ),
	.prn(vcc));
defparam \do_tdl[0][1][2][3] .is_wysiwyg = "true";
defparam \do_tdl[0][1][2][3] .power_up = "low";

dffeas \do_tdl[0][1][2][7] (
	.clk(clk),
	.d(\do_tdl[0][1][1][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][1][2][7]~q ),
	.prn(vcc));
defparam \do_tdl[0][1][2][7] .is_wysiwyg = "true";
defparam \do_tdl[0][1][2][7] .power_up = "low";

dffeas \do_tdl[0][1][2][4] (
	.clk(clk),
	.d(\do_tdl[0][1][1][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][1][2][4]~q ),
	.prn(vcc));
defparam \do_tdl[0][1][2][4] .is_wysiwyg = "true";
defparam \do_tdl[0][1][2][4] .power_up = "low";

dffeas \do_tdl[0][1][2][5] (
	.clk(clk),
	.d(\do_tdl[0][1][1][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][1][2][5]~q ),
	.prn(vcc));
defparam \do_tdl[0][1][2][5] .is_wysiwyg = "true";
defparam \do_tdl[0][1][2][5] .power_up = "low";

dffeas \do_tdl[0][1][2][6] (
	.clk(clk),
	.d(\do_tdl[0][1][1][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][1][2][6]~q ),
	.prn(vcc));
defparam \do_tdl[0][1][2][6] .is_wysiwyg = "true";
defparam \do_tdl[0][1][2][6] .power_up = "low";

dffeas \do_tdl[0][1][2][1] (
	.clk(clk),
	.d(\do_tdl[0][1][1][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][1][2][1]~q ),
	.prn(vcc));
defparam \do_tdl[0][1][2][1] .is_wysiwyg = "true";
defparam \do_tdl[0][1][2][1] .power_up = "low";

dffeas \do_tdl[0][1][2][0] (
	.clk(clk),
	.d(\do_tdl[0][1][1][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][1][2][0]~q ),
	.prn(vcc));
defparam \do_tdl[0][1][2][0] .is_wysiwyg = "true";
defparam \do_tdl[0][1][2][0] .power_up = "low";

dffeas \do_tdl[0][1][2][2] (
	.clk(clk),
	.d(\do_tdl[0][1][1][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][1][2][2]~q ),
	.prn(vcc));
defparam \do_tdl[0][1][2][2] .is_wysiwyg = "true";
defparam \do_tdl[0][1][2][2] .power_up = "low";

dffeas \do_tdl[1][0][2][3] (
	.clk(clk),
	.d(\do_tdl[1][0][1][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][0][2][3]~q ),
	.prn(vcc));
defparam \do_tdl[1][0][2][3] .is_wysiwyg = "true";
defparam \do_tdl[1][0][2][3] .power_up = "low";

dffeas \do_tdl[1][0][2][7] (
	.clk(clk),
	.d(\do_tdl[1][0][1][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][0][2][7]~q ),
	.prn(vcc));
defparam \do_tdl[1][0][2][7] .is_wysiwyg = "true";
defparam \do_tdl[1][0][2][7] .power_up = "low";

dffeas \do_tdl[1][0][2][4] (
	.clk(clk),
	.d(\do_tdl[1][0][1][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][0][2][4]~q ),
	.prn(vcc));
defparam \do_tdl[1][0][2][4] .is_wysiwyg = "true";
defparam \do_tdl[1][0][2][4] .power_up = "low";

dffeas \do_tdl[1][0][2][5] (
	.clk(clk),
	.d(\do_tdl[1][0][1][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][0][2][5]~q ),
	.prn(vcc));
defparam \do_tdl[1][0][2][5] .is_wysiwyg = "true";
defparam \do_tdl[1][0][2][5] .power_up = "low";

dffeas \do_tdl[1][0][2][6] (
	.clk(clk),
	.d(\do_tdl[1][0][1][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][0][2][6]~q ),
	.prn(vcc));
defparam \do_tdl[1][0][2][6] .is_wysiwyg = "true";
defparam \do_tdl[1][0][2][6] .power_up = "low";

dffeas \do_tdl[1][0][2][1] (
	.clk(clk),
	.d(\do_tdl[1][0][1][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][0][2][1]~q ),
	.prn(vcc));
defparam \do_tdl[1][0][2][1] .is_wysiwyg = "true";
defparam \do_tdl[1][0][2][1] .power_up = "low";

dffeas \do_tdl[1][0][2][0] (
	.clk(clk),
	.d(\do_tdl[1][0][1][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][0][2][0]~q ),
	.prn(vcc));
defparam \do_tdl[1][0][2][0] .is_wysiwyg = "true";
defparam \do_tdl[1][0][2][0] .power_up = "low";

dffeas \do_tdl[1][0][2][2] (
	.clk(clk),
	.d(\do_tdl[1][0][1][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][0][2][2]~q ),
	.prn(vcc));
defparam \do_tdl[1][0][2][2] .is_wysiwyg = "true";
defparam \do_tdl[1][0][2][2] .power_up = "low";

dffeas \do_tdl[1][1][2][3] (
	.clk(clk),
	.d(\do_tdl[1][1][1][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][1][2][3]~q ),
	.prn(vcc));
defparam \do_tdl[1][1][2][3] .is_wysiwyg = "true";
defparam \do_tdl[1][1][2][3] .power_up = "low";

dffeas \do_tdl[1][1][2][7] (
	.clk(clk),
	.d(\do_tdl[1][1][1][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][1][2][7]~q ),
	.prn(vcc));
defparam \do_tdl[1][1][2][7] .is_wysiwyg = "true";
defparam \do_tdl[1][1][2][7] .power_up = "low";

dffeas \do_tdl[1][1][2][4] (
	.clk(clk),
	.d(\do_tdl[1][1][1][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][1][2][4]~q ),
	.prn(vcc));
defparam \do_tdl[1][1][2][4] .is_wysiwyg = "true";
defparam \do_tdl[1][1][2][4] .power_up = "low";

dffeas \do_tdl[1][1][2][5] (
	.clk(clk),
	.d(\do_tdl[1][1][1][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][1][2][5]~q ),
	.prn(vcc));
defparam \do_tdl[1][1][2][5] .is_wysiwyg = "true";
defparam \do_tdl[1][1][2][5] .power_up = "low";

dffeas \do_tdl[1][1][2][6] (
	.clk(clk),
	.d(\do_tdl[1][1][1][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][1][2][6]~q ),
	.prn(vcc));
defparam \do_tdl[1][1][2][6] .is_wysiwyg = "true";
defparam \do_tdl[1][1][2][6] .power_up = "low";

dffeas \do_tdl[1][1][2][1] (
	.clk(clk),
	.d(\do_tdl[1][1][1][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][1][2][1]~q ),
	.prn(vcc));
defparam \do_tdl[1][1][2][1] .is_wysiwyg = "true";
defparam \do_tdl[1][1][2][1] .power_up = "low";

dffeas \do_tdl[1][1][2][0] (
	.clk(clk),
	.d(\do_tdl[1][1][1][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][1][2][0]~q ),
	.prn(vcc));
defparam \do_tdl[1][1][2][0] .is_wysiwyg = "true";
defparam \do_tdl[1][1][2][0] .power_up = "low";

dffeas \do_tdl[1][1][2][2] (
	.clk(clk),
	.d(\do_tdl[1][1][1][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][1][2][2]~q ),
	.prn(vcc));
defparam \do_tdl[1][1][2][2] .is_wysiwyg = "true";
defparam \do_tdl[1][1][2][2] .power_up = "low";

dffeas \do_tdl[2][0][2][3] (
	.clk(clk),
	.d(\do_tdl[2][0][1][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][0][2][3]~q ),
	.prn(vcc));
defparam \do_tdl[2][0][2][3] .is_wysiwyg = "true";
defparam \do_tdl[2][0][2][3] .power_up = "low";

dffeas \do_tdl[2][0][2][7] (
	.clk(clk),
	.d(\do_tdl[2][0][1][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][0][2][7]~q ),
	.prn(vcc));
defparam \do_tdl[2][0][2][7] .is_wysiwyg = "true";
defparam \do_tdl[2][0][2][7] .power_up = "low";

dffeas \do_tdl[2][0][2][4] (
	.clk(clk),
	.d(\do_tdl[2][0][1][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][0][2][4]~q ),
	.prn(vcc));
defparam \do_tdl[2][0][2][4] .is_wysiwyg = "true";
defparam \do_tdl[2][0][2][4] .power_up = "low";

dffeas \do_tdl[2][0][2][5] (
	.clk(clk),
	.d(\do_tdl[2][0][1][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][0][2][5]~q ),
	.prn(vcc));
defparam \do_tdl[2][0][2][5] .is_wysiwyg = "true";
defparam \do_tdl[2][0][2][5] .power_up = "low";

dffeas \do_tdl[2][0][2][6] (
	.clk(clk),
	.d(\do_tdl[2][0][1][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][0][2][6]~q ),
	.prn(vcc));
defparam \do_tdl[2][0][2][6] .is_wysiwyg = "true";
defparam \do_tdl[2][0][2][6] .power_up = "low";

dffeas \do_tdl[2][0][2][1] (
	.clk(clk),
	.d(\do_tdl[2][0][1][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][0][2][1]~q ),
	.prn(vcc));
defparam \do_tdl[2][0][2][1] .is_wysiwyg = "true";
defparam \do_tdl[2][0][2][1] .power_up = "low";

dffeas \do_tdl[2][0][2][0] (
	.clk(clk),
	.d(\do_tdl[2][0][1][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][0][2][0]~q ),
	.prn(vcc));
defparam \do_tdl[2][0][2][0] .is_wysiwyg = "true";
defparam \do_tdl[2][0][2][0] .power_up = "low";

dffeas \do_tdl[2][0][2][2] (
	.clk(clk),
	.d(\do_tdl[2][0][1][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][0][2][2]~q ),
	.prn(vcc));
defparam \do_tdl[2][0][2][2] .is_wysiwyg = "true";
defparam \do_tdl[2][0][2][2] .power_up = "low";

dffeas \do_tdl[2][1][2][3] (
	.clk(clk),
	.d(\do_tdl[2][1][1][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][1][2][3]~q ),
	.prn(vcc));
defparam \do_tdl[2][1][2][3] .is_wysiwyg = "true";
defparam \do_tdl[2][1][2][3] .power_up = "low";

dffeas \do_tdl[2][1][2][7] (
	.clk(clk),
	.d(\do_tdl[2][1][1][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][1][2][7]~q ),
	.prn(vcc));
defparam \do_tdl[2][1][2][7] .is_wysiwyg = "true";
defparam \do_tdl[2][1][2][7] .power_up = "low";

dffeas \do_tdl[2][1][2][4] (
	.clk(clk),
	.d(\do_tdl[2][1][1][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][1][2][4]~q ),
	.prn(vcc));
defparam \do_tdl[2][1][2][4] .is_wysiwyg = "true";
defparam \do_tdl[2][1][2][4] .power_up = "low";

dffeas \do_tdl[2][1][2][5] (
	.clk(clk),
	.d(\do_tdl[2][1][1][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][1][2][5]~q ),
	.prn(vcc));
defparam \do_tdl[2][1][2][5] .is_wysiwyg = "true";
defparam \do_tdl[2][1][2][5] .power_up = "low";

dffeas \do_tdl[2][1][2][6] (
	.clk(clk),
	.d(\do_tdl[2][1][1][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][1][2][6]~q ),
	.prn(vcc));
defparam \do_tdl[2][1][2][6] .is_wysiwyg = "true";
defparam \do_tdl[2][1][2][6] .power_up = "low";

dffeas \do_tdl[2][1][2][1] (
	.clk(clk),
	.d(\do_tdl[2][1][1][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][1][2][1]~q ),
	.prn(vcc));
defparam \do_tdl[2][1][2][1] .is_wysiwyg = "true";
defparam \do_tdl[2][1][2][1] .power_up = "low";

dffeas \do_tdl[2][1][2][0] (
	.clk(clk),
	.d(\do_tdl[2][1][1][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][1][2][0]~q ),
	.prn(vcc));
defparam \do_tdl[2][1][2][0] .is_wysiwyg = "true";
defparam \do_tdl[2][1][2][0] .power_up = "low";

dffeas \do_tdl[2][1][2][2] (
	.clk(clk),
	.d(\do_tdl[2][1][1][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][1][2][2]~q ),
	.prn(vcc));
defparam \do_tdl[2][1][2][2] .is_wysiwyg = "true";
defparam \do_tdl[2][1][2][2] .power_up = "low";

dffeas \do_tdl[3][0][2][3] (
	.clk(clk),
	.d(\do_tdl[3][0][1][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][0][2][3]~q ),
	.prn(vcc));
defparam \do_tdl[3][0][2][3] .is_wysiwyg = "true";
defparam \do_tdl[3][0][2][3] .power_up = "low";

dffeas \do_tdl[3][0][2][7] (
	.clk(clk),
	.d(\do_tdl[3][0][1][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][0][2][7]~q ),
	.prn(vcc));
defparam \do_tdl[3][0][2][7] .is_wysiwyg = "true";
defparam \do_tdl[3][0][2][7] .power_up = "low";

dffeas \do_tdl[3][0][2][4] (
	.clk(clk),
	.d(\do_tdl[3][0][1][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][0][2][4]~q ),
	.prn(vcc));
defparam \do_tdl[3][0][2][4] .is_wysiwyg = "true";
defparam \do_tdl[3][0][2][4] .power_up = "low";

dffeas \do_tdl[3][0][2][5] (
	.clk(clk),
	.d(\do_tdl[3][0][1][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][0][2][5]~q ),
	.prn(vcc));
defparam \do_tdl[3][0][2][5] .is_wysiwyg = "true";
defparam \do_tdl[3][0][2][5] .power_up = "low";

dffeas \do_tdl[3][0][2][6] (
	.clk(clk),
	.d(\do_tdl[3][0][1][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][0][2][6]~q ),
	.prn(vcc));
defparam \do_tdl[3][0][2][6] .is_wysiwyg = "true";
defparam \do_tdl[3][0][2][6] .power_up = "low";

dffeas \do_tdl[3][0][2][1] (
	.clk(clk),
	.d(\do_tdl[3][0][1][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][0][2][1]~q ),
	.prn(vcc));
defparam \do_tdl[3][0][2][1] .is_wysiwyg = "true";
defparam \do_tdl[3][0][2][1] .power_up = "low";

dffeas \do_tdl[3][0][2][0] (
	.clk(clk),
	.d(\do_tdl[3][0][1][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][0][2][0]~q ),
	.prn(vcc));
defparam \do_tdl[3][0][2][0] .is_wysiwyg = "true";
defparam \do_tdl[3][0][2][0] .power_up = "low";

dffeas \do_tdl[3][0][2][2] (
	.clk(clk),
	.d(\do_tdl[3][0][1][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][0][2][2]~q ),
	.prn(vcc));
defparam \do_tdl[3][0][2][2] .is_wysiwyg = "true";
defparam \do_tdl[3][0][2][2] .power_up = "low";

dffeas \do_tdl[3][1][2][3] (
	.clk(clk),
	.d(\do_tdl[3][1][1][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][1][2][3]~q ),
	.prn(vcc));
defparam \do_tdl[3][1][2][3] .is_wysiwyg = "true";
defparam \do_tdl[3][1][2][3] .power_up = "low";

dffeas \do_tdl[3][1][2][7] (
	.clk(clk),
	.d(\do_tdl[3][1][1][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][1][2][7]~q ),
	.prn(vcc));
defparam \do_tdl[3][1][2][7] .is_wysiwyg = "true";
defparam \do_tdl[3][1][2][7] .power_up = "low";

dffeas \do_tdl[3][1][2][4] (
	.clk(clk),
	.d(\do_tdl[3][1][1][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][1][2][4]~q ),
	.prn(vcc));
defparam \do_tdl[3][1][2][4] .is_wysiwyg = "true";
defparam \do_tdl[3][1][2][4] .power_up = "low";

dffeas \do_tdl[3][1][2][5] (
	.clk(clk),
	.d(\do_tdl[3][1][1][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][1][2][5]~q ),
	.prn(vcc));
defparam \do_tdl[3][1][2][5] .is_wysiwyg = "true";
defparam \do_tdl[3][1][2][5] .power_up = "low";

dffeas \do_tdl[3][1][2][6] (
	.clk(clk),
	.d(\do_tdl[3][1][1][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][1][2][6]~q ),
	.prn(vcc));
defparam \do_tdl[3][1][2][6] .is_wysiwyg = "true";
defparam \do_tdl[3][1][2][6] .power_up = "low";

dffeas \do_tdl[3][1][2][1] (
	.clk(clk),
	.d(\do_tdl[3][1][1][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][1][2][1]~q ),
	.prn(vcc));
defparam \do_tdl[3][1][2][1] .is_wysiwyg = "true";
defparam \do_tdl[3][1][2][1] .power_up = "low";

dffeas \do_tdl[3][1][2][0] (
	.clk(clk),
	.d(\do_tdl[3][1][1][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][1][2][0]~q ),
	.prn(vcc));
defparam \do_tdl[3][1][2][0] .is_wysiwyg = "true";
defparam \do_tdl[3][1][2][0] .power_up = "low";

dffeas \do_tdl[3][1][2][2] (
	.clk(clk),
	.d(\do_tdl[3][1][1][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][1][2][2]~q ),
	.prn(vcc));
defparam \do_tdl[3][1][2][2] .is_wysiwyg = "true";
defparam \do_tdl[3][1][2][2] .power_up = "low";

dffeas \sdft.IDLE (
	.clk(clk),
	.d(\sdft.IDLE~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sdft.IDLE~q ),
	.prn(vcc));
defparam \sdft.IDLE .is_wysiwyg = "true";
defparam \sdft.IDLE .power_up = "low";

cycloneiii_lcell_comb \state_cnt~12 (
	.dataa(\sdft.WAIT_FOR_OUTPUT~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\sdft.IDLE~q ),
	.cin(gnd),
	.combout(\state_cnt~12_combout ),
	.cout());
defparam \state_cnt~12 .lut_mask = 16'hAAFF;
defparam \state_cnt~12 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \state_cnt[0]~13 (
	.dataa(global_clock_enable),
	.datab(\sdft.ENABLE_DFT_O~q ),
	.datac(\gap_reg~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\state_cnt[0]~13_combout ),
	.cout());
defparam \state_cnt[0]~13 .lut_mask = 16'hBFBF;
defparam \state_cnt[0]~13 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector13~0 (
	.dataa(\sdft.BLOCK_DFT_I~q ),
	.datab(tdl_arr_51),
	.datac(\Equal0~1_combout ),
	.datad(\sdft.IDLE~q ),
	.cin(gnd),
	.combout(\Selector13~0_combout ),
	.cout());
defparam \Selector13~0 .lut_mask = 16'hEFFF;
defparam \Selector13~0 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[3][0][4] (
	.clk(clk),
	.d(\reg_no_twiddle~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[3][0][4]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[3][0][4] .is_wysiwyg = "true";
defparam \reg_no_twiddle[3][0][4] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~24 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[3][0][4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~24_combout ),
	.cout());
defparam \reg_no_twiddle~24 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~24 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[3][1][4] (
	.clk(clk),
	.d(\reg_no_twiddle~35_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[3][1][4]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[3][1][4] .is_wysiwyg = "true";
defparam \reg_no_twiddle[3][1][4] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~25 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[3][1][4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~25_combout ),
	.cout());
defparam \reg_no_twiddle~25 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~25 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[3][0][5] (
	.clk(clk),
	.d(\reg_no_twiddle~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[3][0][5]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[3][0][5] .is_wysiwyg = "true";
defparam \reg_no_twiddle[3][0][5] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~26 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[3][0][5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~26_combout ),
	.cout());
defparam \reg_no_twiddle~26 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~26 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[3][1][5] (
	.clk(clk),
	.d(\reg_no_twiddle~37_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[3][1][5]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[3][1][5] .is_wysiwyg = "true";
defparam \reg_no_twiddle[3][1][5] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~27 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[3][1][5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~27_combout ),
	.cout());
defparam \reg_no_twiddle~27 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~27 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[3][0][6] (
	.clk(clk),
	.d(\reg_no_twiddle~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[3][0][6]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[3][0][6] .is_wysiwyg = "true";
defparam \reg_no_twiddle[3][0][6] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~28 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[3][0][6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~28_combout ),
	.cout());
defparam \reg_no_twiddle~28 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~28 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[3][1][6] (
	.clk(clk),
	.d(\reg_no_twiddle~39_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[3][1][6]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[3][1][6] .is_wysiwyg = "true";
defparam \reg_no_twiddle[3][1][6] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~29 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[3][1][6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~29_combout ),
	.cout());
defparam \reg_no_twiddle~29 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~29 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[2][0][3] (
	.clk(clk),
	.d(\reg_no_twiddle~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[2][0][3]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[2][0][3] .is_wysiwyg = "true";
defparam \reg_no_twiddle[2][0][3] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~30 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[2][0][3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~30_combout ),
	.cout());
defparam \reg_no_twiddle~30 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~30 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[2][0][7] (
	.clk(clk),
	.d(\reg_no_twiddle~41_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[2][0][7]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[2][0][7] .is_wysiwyg = "true";
defparam \reg_no_twiddle[2][0][7] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~31 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[2][0][7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~31_combout ),
	.cout());
defparam \reg_no_twiddle~31 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~31 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[2][1][7] (
	.clk(clk),
	.d(\reg_no_twiddle~42_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[2][1][7]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[2][1][7] .is_wysiwyg = "true";
defparam \reg_no_twiddle[2][1][7] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~32 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[2][1][7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~32_combout ),
	.cout());
defparam \reg_no_twiddle~32 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~32 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[2][1][3] (
	.clk(clk),
	.d(\reg_no_twiddle~43_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[2][1][3]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[2][1][3] .is_wysiwyg = "true";
defparam \reg_no_twiddle[2][1][3] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~33 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[2][1][3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~33_combout ),
	.cout());
defparam \reg_no_twiddle~33 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~33 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Equal1~0 (
	.dataa(\Equal0~0_combout ),
	.datab(\state_cnt[1]~q ),
	.datac(gnd),
	.datad(\state_cnt[0]~q ),
	.cin(gnd),
	.combout(\Equal1~0_combout ),
	.cout());
defparam \Equal1~0 .lut_mask = 16'hEEFF;
defparam \Equal1~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector15~0 (
	.dataa(\sdft.ENABLE_DFT_O~q ),
	.datab(\sdft.ENABLE_BFP_O~q ),
	.datac(\gap_reg~q ),
	.datad(\Equal1~0_combout ),
	.cin(gnd),
	.combout(\Selector15~0_combout ),
	.cout());
defparam \Selector15~0 .lut_mask = 16'hEFFF;
defparam \Selector15~0 .sum_lutc_input = "datac";

dffeas \do_tdl[0][0][1][3] (
	.clk(clk),
	.d(\do_tdl[0][0][0][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][0][1][3]~q ),
	.prn(vcc));
defparam \do_tdl[0][0][1][3] .is_wysiwyg = "true";
defparam \do_tdl[0][0][1][3] .power_up = "low";

dffeas \do_tdl[0][0][1][7] (
	.clk(clk),
	.d(\do_tdl[0][0][0][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][0][1][7]~q ),
	.prn(vcc));
defparam \do_tdl[0][0][1][7] .is_wysiwyg = "true";
defparam \do_tdl[0][0][1][7] .power_up = "low";

dffeas \do_tdl[0][0][1][4] (
	.clk(clk),
	.d(\do_tdl[0][0][0][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][0][1][4]~q ),
	.prn(vcc));
defparam \do_tdl[0][0][1][4] .is_wysiwyg = "true";
defparam \do_tdl[0][0][1][4] .power_up = "low";

dffeas \do_tdl[0][0][1][5] (
	.clk(clk),
	.d(\do_tdl[0][0][0][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][0][1][5]~q ),
	.prn(vcc));
defparam \do_tdl[0][0][1][5] .is_wysiwyg = "true";
defparam \do_tdl[0][0][1][5] .power_up = "low";

dffeas \do_tdl[0][0][1][6] (
	.clk(clk),
	.d(\do_tdl[0][0][0][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][0][1][6]~q ),
	.prn(vcc));
defparam \do_tdl[0][0][1][6] .is_wysiwyg = "true";
defparam \do_tdl[0][0][1][6] .power_up = "low";

dffeas \do_tdl[0][0][1][1] (
	.clk(clk),
	.d(\do_tdl[0][0][0][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][0][1][1]~q ),
	.prn(vcc));
defparam \do_tdl[0][0][1][1] .is_wysiwyg = "true";
defparam \do_tdl[0][0][1][1] .power_up = "low";

dffeas \do_tdl[0][0][1][0] (
	.clk(clk),
	.d(\do_tdl[0][0][0][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][0][1][0]~q ),
	.prn(vcc));
defparam \do_tdl[0][0][1][0] .is_wysiwyg = "true";
defparam \do_tdl[0][0][1][0] .power_up = "low";

dffeas \do_tdl[0][0][1][2] (
	.clk(clk),
	.d(\do_tdl[0][0][0][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][0][1][2]~q ),
	.prn(vcc));
defparam \do_tdl[0][0][1][2] .is_wysiwyg = "true";
defparam \do_tdl[0][0][1][2] .power_up = "low";

dffeas \do_tdl[0][1][1][3] (
	.clk(clk),
	.d(\do_tdl[0][1][0][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][1][1][3]~q ),
	.prn(vcc));
defparam \do_tdl[0][1][1][3] .is_wysiwyg = "true";
defparam \do_tdl[0][1][1][3] .power_up = "low";

dffeas \do_tdl[0][1][1][7] (
	.clk(clk),
	.d(\do_tdl[0][1][0][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][1][1][7]~q ),
	.prn(vcc));
defparam \do_tdl[0][1][1][7] .is_wysiwyg = "true";
defparam \do_tdl[0][1][1][7] .power_up = "low";

dffeas \do_tdl[0][1][1][4] (
	.clk(clk),
	.d(\do_tdl[0][1][0][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][1][1][4]~q ),
	.prn(vcc));
defparam \do_tdl[0][1][1][4] .is_wysiwyg = "true";
defparam \do_tdl[0][1][1][4] .power_up = "low";

dffeas \do_tdl[0][1][1][5] (
	.clk(clk),
	.d(\do_tdl[0][1][0][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][1][1][5]~q ),
	.prn(vcc));
defparam \do_tdl[0][1][1][5] .is_wysiwyg = "true";
defparam \do_tdl[0][1][1][5] .power_up = "low";

dffeas \do_tdl[0][1][1][6] (
	.clk(clk),
	.d(\do_tdl[0][1][0][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][1][1][6]~q ),
	.prn(vcc));
defparam \do_tdl[0][1][1][6] .is_wysiwyg = "true";
defparam \do_tdl[0][1][1][6] .power_up = "low";

dffeas \do_tdl[0][1][1][1] (
	.clk(clk),
	.d(\do_tdl[0][1][0][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][1][1][1]~q ),
	.prn(vcc));
defparam \do_tdl[0][1][1][1] .is_wysiwyg = "true";
defparam \do_tdl[0][1][1][1] .power_up = "low";

dffeas \do_tdl[0][1][1][0] (
	.clk(clk),
	.d(\do_tdl[0][1][0][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][1][1][0]~q ),
	.prn(vcc));
defparam \do_tdl[0][1][1][0] .is_wysiwyg = "true";
defparam \do_tdl[0][1][1][0] .power_up = "low";

dffeas \do_tdl[0][1][1][2] (
	.clk(clk),
	.d(\do_tdl[0][1][0][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][1][1][2]~q ),
	.prn(vcc));
defparam \do_tdl[0][1][1][2] .is_wysiwyg = "true";
defparam \do_tdl[0][1][1][2] .power_up = "low";

dffeas \do_tdl[1][0][1][3] (
	.clk(clk),
	.d(\do_tdl[1][0][0][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][0][1][3]~q ),
	.prn(vcc));
defparam \do_tdl[1][0][1][3] .is_wysiwyg = "true";
defparam \do_tdl[1][0][1][3] .power_up = "low";

dffeas \do_tdl[1][0][1][7] (
	.clk(clk),
	.d(\do_tdl[1][0][0][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][0][1][7]~q ),
	.prn(vcc));
defparam \do_tdl[1][0][1][7] .is_wysiwyg = "true";
defparam \do_tdl[1][0][1][7] .power_up = "low";

dffeas \do_tdl[1][0][1][4] (
	.clk(clk),
	.d(\do_tdl[1][0][0][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][0][1][4]~q ),
	.prn(vcc));
defparam \do_tdl[1][0][1][4] .is_wysiwyg = "true";
defparam \do_tdl[1][0][1][4] .power_up = "low";

dffeas \do_tdl[1][0][1][5] (
	.clk(clk),
	.d(\do_tdl[1][0][0][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][0][1][5]~q ),
	.prn(vcc));
defparam \do_tdl[1][0][1][5] .is_wysiwyg = "true";
defparam \do_tdl[1][0][1][5] .power_up = "low";

dffeas \do_tdl[1][0][1][6] (
	.clk(clk),
	.d(\do_tdl[1][0][0][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][0][1][6]~q ),
	.prn(vcc));
defparam \do_tdl[1][0][1][6] .is_wysiwyg = "true";
defparam \do_tdl[1][0][1][6] .power_up = "low";

dffeas \do_tdl[1][0][1][1] (
	.clk(clk),
	.d(\do_tdl[1][0][0][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][0][1][1]~q ),
	.prn(vcc));
defparam \do_tdl[1][0][1][1] .is_wysiwyg = "true";
defparam \do_tdl[1][0][1][1] .power_up = "low";

dffeas \do_tdl[1][0][1][0] (
	.clk(clk),
	.d(\do_tdl[1][0][0][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][0][1][0]~q ),
	.prn(vcc));
defparam \do_tdl[1][0][1][0] .is_wysiwyg = "true";
defparam \do_tdl[1][0][1][0] .power_up = "low";

dffeas \do_tdl[1][0][1][2] (
	.clk(clk),
	.d(\do_tdl[1][0][0][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][0][1][2]~q ),
	.prn(vcc));
defparam \do_tdl[1][0][1][2] .is_wysiwyg = "true";
defparam \do_tdl[1][0][1][2] .power_up = "low";

dffeas \do_tdl[1][1][1][3] (
	.clk(clk),
	.d(\do_tdl[1][1][0][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][1][1][3]~q ),
	.prn(vcc));
defparam \do_tdl[1][1][1][3] .is_wysiwyg = "true";
defparam \do_tdl[1][1][1][3] .power_up = "low";

dffeas \do_tdl[1][1][1][7] (
	.clk(clk),
	.d(\do_tdl[1][1][0][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][1][1][7]~q ),
	.prn(vcc));
defparam \do_tdl[1][1][1][7] .is_wysiwyg = "true";
defparam \do_tdl[1][1][1][7] .power_up = "low";

dffeas \do_tdl[1][1][1][4] (
	.clk(clk),
	.d(\do_tdl[1][1][0][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][1][1][4]~q ),
	.prn(vcc));
defparam \do_tdl[1][1][1][4] .is_wysiwyg = "true";
defparam \do_tdl[1][1][1][4] .power_up = "low";

dffeas \do_tdl[1][1][1][5] (
	.clk(clk),
	.d(\do_tdl[1][1][0][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][1][1][5]~q ),
	.prn(vcc));
defparam \do_tdl[1][1][1][5] .is_wysiwyg = "true";
defparam \do_tdl[1][1][1][5] .power_up = "low";

dffeas \do_tdl[1][1][1][6] (
	.clk(clk),
	.d(\do_tdl[1][1][0][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][1][1][6]~q ),
	.prn(vcc));
defparam \do_tdl[1][1][1][6] .is_wysiwyg = "true";
defparam \do_tdl[1][1][1][6] .power_up = "low";

dffeas \do_tdl[1][1][1][1] (
	.clk(clk),
	.d(\do_tdl[1][1][0][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][1][1][1]~q ),
	.prn(vcc));
defparam \do_tdl[1][1][1][1] .is_wysiwyg = "true";
defparam \do_tdl[1][1][1][1] .power_up = "low";

dffeas \do_tdl[1][1][1][0] (
	.clk(clk),
	.d(\do_tdl[1][1][0][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][1][1][0]~q ),
	.prn(vcc));
defparam \do_tdl[1][1][1][0] .is_wysiwyg = "true";
defparam \do_tdl[1][1][1][0] .power_up = "low";

dffeas \do_tdl[1][1][1][2] (
	.clk(clk),
	.d(\do_tdl[1][1][0][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][1][1][2]~q ),
	.prn(vcc));
defparam \do_tdl[1][1][1][2] .is_wysiwyg = "true";
defparam \do_tdl[1][1][1][2] .power_up = "low";

dffeas \do_tdl[2][0][1][3] (
	.clk(clk),
	.d(\do_tdl[2][0][0][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][0][1][3]~q ),
	.prn(vcc));
defparam \do_tdl[2][0][1][3] .is_wysiwyg = "true";
defparam \do_tdl[2][0][1][3] .power_up = "low";

dffeas \do_tdl[2][0][1][7] (
	.clk(clk),
	.d(\do_tdl[2][0][0][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][0][1][7]~q ),
	.prn(vcc));
defparam \do_tdl[2][0][1][7] .is_wysiwyg = "true";
defparam \do_tdl[2][0][1][7] .power_up = "low";

dffeas \do_tdl[2][0][1][4] (
	.clk(clk),
	.d(\do_tdl[2][0][0][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][0][1][4]~q ),
	.prn(vcc));
defparam \do_tdl[2][0][1][4] .is_wysiwyg = "true";
defparam \do_tdl[2][0][1][4] .power_up = "low";

dffeas \do_tdl[2][0][1][5] (
	.clk(clk),
	.d(\do_tdl[2][0][0][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][0][1][5]~q ),
	.prn(vcc));
defparam \do_tdl[2][0][1][5] .is_wysiwyg = "true";
defparam \do_tdl[2][0][1][5] .power_up = "low";

dffeas \do_tdl[2][0][1][6] (
	.clk(clk),
	.d(\do_tdl[2][0][0][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][0][1][6]~q ),
	.prn(vcc));
defparam \do_tdl[2][0][1][6] .is_wysiwyg = "true";
defparam \do_tdl[2][0][1][6] .power_up = "low";

dffeas \do_tdl[2][0][1][1] (
	.clk(clk),
	.d(\do_tdl[2][0][0][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][0][1][1]~q ),
	.prn(vcc));
defparam \do_tdl[2][0][1][1] .is_wysiwyg = "true";
defparam \do_tdl[2][0][1][1] .power_up = "low";

dffeas \do_tdl[2][0][1][0] (
	.clk(clk),
	.d(\do_tdl[2][0][0][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][0][1][0]~q ),
	.prn(vcc));
defparam \do_tdl[2][0][1][0] .is_wysiwyg = "true";
defparam \do_tdl[2][0][1][0] .power_up = "low";

dffeas \do_tdl[2][0][1][2] (
	.clk(clk),
	.d(\do_tdl[2][0][0][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][0][1][2]~q ),
	.prn(vcc));
defparam \do_tdl[2][0][1][2] .is_wysiwyg = "true";
defparam \do_tdl[2][0][1][2] .power_up = "low";

dffeas \do_tdl[2][1][1][3] (
	.clk(clk),
	.d(\do_tdl[2][1][0][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][1][1][3]~q ),
	.prn(vcc));
defparam \do_tdl[2][1][1][3] .is_wysiwyg = "true";
defparam \do_tdl[2][1][1][3] .power_up = "low";

dffeas \do_tdl[2][1][1][7] (
	.clk(clk),
	.d(\do_tdl[2][1][0][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][1][1][7]~q ),
	.prn(vcc));
defparam \do_tdl[2][1][1][7] .is_wysiwyg = "true";
defparam \do_tdl[2][1][1][7] .power_up = "low";

dffeas \do_tdl[2][1][1][4] (
	.clk(clk),
	.d(\do_tdl[2][1][0][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][1][1][4]~q ),
	.prn(vcc));
defparam \do_tdl[2][1][1][4] .is_wysiwyg = "true";
defparam \do_tdl[2][1][1][4] .power_up = "low";

dffeas \do_tdl[2][1][1][5] (
	.clk(clk),
	.d(\do_tdl[2][1][0][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][1][1][5]~q ),
	.prn(vcc));
defparam \do_tdl[2][1][1][5] .is_wysiwyg = "true";
defparam \do_tdl[2][1][1][5] .power_up = "low";

dffeas \do_tdl[2][1][1][6] (
	.clk(clk),
	.d(\do_tdl[2][1][0][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][1][1][6]~q ),
	.prn(vcc));
defparam \do_tdl[2][1][1][6] .is_wysiwyg = "true";
defparam \do_tdl[2][1][1][6] .power_up = "low";

dffeas \do_tdl[2][1][1][1] (
	.clk(clk),
	.d(\do_tdl[2][1][0][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][1][1][1]~q ),
	.prn(vcc));
defparam \do_tdl[2][1][1][1] .is_wysiwyg = "true";
defparam \do_tdl[2][1][1][1] .power_up = "low";

dffeas \do_tdl[2][1][1][0] (
	.clk(clk),
	.d(\do_tdl[2][1][0][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][1][1][0]~q ),
	.prn(vcc));
defparam \do_tdl[2][1][1][0] .is_wysiwyg = "true";
defparam \do_tdl[2][1][1][0] .power_up = "low";

dffeas \do_tdl[2][1][1][2] (
	.clk(clk),
	.d(\do_tdl[2][1][0][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][1][1][2]~q ),
	.prn(vcc));
defparam \do_tdl[2][1][1][2] .is_wysiwyg = "true";
defparam \do_tdl[2][1][1][2] .power_up = "low";

dffeas \do_tdl[3][0][1][3] (
	.clk(clk),
	.d(\do_tdl[3][0][0][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][0][1][3]~q ),
	.prn(vcc));
defparam \do_tdl[3][0][1][3] .is_wysiwyg = "true";
defparam \do_tdl[3][0][1][3] .power_up = "low";

dffeas \do_tdl[3][0][1][7] (
	.clk(clk),
	.d(\do_tdl[3][0][0][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][0][1][7]~q ),
	.prn(vcc));
defparam \do_tdl[3][0][1][7] .is_wysiwyg = "true";
defparam \do_tdl[3][0][1][7] .power_up = "low";

dffeas \do_tdl[3][0][1][4] (
	.clk(clk),
	.d(\do_tdl[3][0][0][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][0][1][4]~q ),
	.prn(vcc));
defparam \do_tdl[3][0][1][4] .is_wysiwyg = "true";
defparam \do_tdl[3][0][1][4] .power_up = "low";

dffeas \do_tdl[3][0][1][5] (
	.clk(clk),
	.d(\do_tdl[3][0][0][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][0][1][5]~q ),
	.prn(vcc));
defparam \do_tdl[3][0][1][5] .is_wysiwyg = "true";
defparam \do_tdl[3][0][1][5] .power_up = "low";

dffeas \do_tdl[3][0][1][6] (
	.clk(clk),
	.d(\do_tdl[3][0][0][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][0][1][6]~q ),
	.prn(vcc));
defparam \do_tdl[3][0][1][6] .is_wysiwyg = "true";
defparam \do_tdl[3][0][1][6] .power_up = "low";

dffeas \do_tdl[3][0][1][1] (
	.clk(clk),
	.d(\do_tdl[3][0][0][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][0][1][1]~q ),
	.prn(vcc));
defparam \do_tdl[3][0][1][1] .is_wysiwyg = "true";
defparam \do_tdl[3][0][1][1] .power_up = "low";

dffeas \do_tdl[3][0][1][0] (
	.clk(clk),
	.d(\do_tdl[3][0][0][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][0][1][0]~q ),
	.prn(vcc));
defparam \do_tdl[3][0][1][0] .is_wysiwyg = "true";
defparam \do_tdl[3][0][1][0] .power_up = "low";

dffeas \do_tdl[3][0][1][2] (
	.clk(clk),
	.d(\do_tdl[3][0][0][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][0][1][2]~q ),
	.prn(vcc));
defparam \do_tdl[3][0][1][2] .is_wysiwyg = "true";
defparam \do_tdl[3][0][1][2] .power_up = "low";

dffeas \do_tdl[3][1][1][3] (
	.clk(clk),
	.d(\do_tdl[3][1][0][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][1][1][3]~q ),
	.prn(vcc));
defparam \do_tdl[3][1][1][3] .is_wysiwyg = "true";
defparam \do_tdl[3][1][1][3] .power_up = "low";

dffeas \do_tdl[3][1][1][7] (
	.clk(clk),
	.d(\do_tdl[3][1][0][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][1][1][7]~q ),
	.prn(vcc));
defparam \do_tdl[3][1][1][7] .is_wysiwyg = "true";
defparam \do_tdl[3][1][1][7] .power_up = "low";

dffeas \do_tdl[3][1][1][4] (
	.clk(clk),
	.d(\do_tdl[3][1][0][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][1][1][4]~q ),
	.prn(vcc));
defparam \do_tdl[3][1][1][4] .is_wysiwyg = "true";
defparam \do_tdl[3][1][1][4] .power_up = "low";

dffeas \do_tdl[3][1][1][5] (
	.clk(clk),
	.d(\do_tdl[3][1][0][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][1][1][5]~q ),
	.prn(vcc));
defparam \do_tdl[3][1][1][5] .is_wysiwyg = "true";
defparam \do_tdl[3][1][1][5] .power_up = "low";

dffeas \do_tdl[3][1][1][6] (
	.clk(clk),
	.d(\do_tdl[3][1][0][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][1][1][6]~q ),
	.prn(vcc));
defparam \do_tdl[3][1][1][6] .is_wysiwyg = "true";
defparam \do_tdl[3][1][1][6] .power_up = "low";

dffeas \do_tdl[3][1][1][1] (
	.clk(clk),
	.d(\do_tdl[3][1][0][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][1][1][1]~q ),
	.prn(vcc));
defparam \do_tdl[3][1][1][1] .is_wysiwyg = "true";
defparam \do_tdl[3][1][1][1] .power_up = "low";

dffeas \do_tdl[3][1][1][0] (
	.clk(clk),
	.d(\do_tdl[3][1][0][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][1][1][0]~q ),
	.prn(vcc));
defparam \do_tdl[3][1][1][0] .is_wysiwyg = "true";
defparam \do_tdl[3][1][1][0] .power_up = "low";

dffeas \do_tdl[3][1][1][2] (
	.clk(clk),
	.d(\do_tdl[3][1][0][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][1][1][2]~q ),
	.prn(vcc));
defparam \do_tdl[3][1][1][2] .is_wysiwyg = "true";
defparam \do_tdl[3][1][1][2] .power_up = "low";

dffeas \sdft.DISABLE_DFT_O (
	.clk(clk),
	.d(\sdft~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sdft.DISABLE_DFT_O~q ),
	.prn(vcc));
defparam \sdft.DISABLE_DFT_O .is_wysiwyg = "true";
defparam \sdft.DISABLE_DFT_O .power_up = "low";

cycloneiii_lcell_comb \sdft.IDLE~0 (
	.dataa(\sdft.DISABLE_DFT_O~q ),
	.datab(\sdft.IDLE~q ),
	.datac(tdl_arr_51),
	.datad(reset_n),
	.cin(gnd),
	.combout(\sdft.IDLE~0_combout ),
	.cout());
defparam \sdft.IDLE~0 .lut_mask = 16'hFFFD;
defparam \sdft.IDLE~0 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[2][0][4] (
	.clk(clk),
	.d(\reg_no_twiddle~44_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[2][0][4]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[2][0][4] .is_wysiwyg = "true";
defparam \reg_no_twiddle[2][0][4] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~34 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[2][0][4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~34_combout ),
	.cout());
defparam \reg_no_twiddle~34 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~34 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[2][1][4] (
	.clk(clk),
	.d(\reg_no_twiddle~45_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[2][1][4]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[2][1][4] .is_wysiwyg = "true";
defparam \reg_no_twiddle[2][1][4] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~35 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[2][1][4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~35_combout ),
	.cout());
defparam \reg_no_twiddle~35 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~35 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[2][0][5] (
	.clk(clk),
	.d(\reg_no_twiddle~46_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[2][0][5]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[2][0][5] .is_wysiwyg = "true";
defparam \reg_no_twiddle[2][0][5] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~36 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[2][0][5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~36_combout ),
	.cout());
defparam \reg_no_twiddle~36 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~36 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[2][1][5] (
	.clk(clk),
	.d(\reg_no_twiddle~47_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[2][1][5]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[2][1][5] .is_wysiwyg = "true";
defparam \reg_no_twiddle[2][1][5] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~37 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[2][1][5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~37_combout ),
	.cout());
defparam \reg_no_twiddle~37 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~37 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[2][0][6] (
	.clk(clk),
	.d(\reg_no_twiddle~48_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[2][0][6]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[2][0][6] .is_wysiwyg = "true";
defparam \reg_no_twiddle[2][0][6] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~38 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[2][0][6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~38_combout ),
	.cout());
defparam \reg_no_twiddle~38 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~38 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[2][1][6] (
	.clk(clk),
	.d(\reg_no_twiddle~49_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[2][1][6]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[2][1][6] .is_wysiwyg = "true";
defparam \reg_no_twiddle[2][1][6] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~39 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[2][1][6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~39_combout ),
	.cout());
defparam \reg_no_twiddle~39 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~39 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[1][0][3] (
	.clk(clk),
	.d(\reg_no_twiddle~50_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[1][0][3]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[1][0][3] .is_wysiwyg = "true";
defparam \reg_no_twiddle[1][0][3] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~40 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[1][0][3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~40_combout ),
	.cout());
defparam \reg_no_twiddle~40 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~40 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[1][0][7] (
	.clk(clk),
	.d(\reg_no_twiddle~51_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[1][0][7]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[1][0][7] .is_wysiwyg = "true";
defparam \reg_no_twiddle[1][0][7] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~41 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[1][0][7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~41_combout ),
	.cout());
defparam \reg_no_twiddle~41 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~41 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[1][1][7] (
	.clk(clk),
	.d(\reg_no_twiddle~52_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[1][1][7]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[1][1][7] .is_wysiwyg = "true";
defparam \reg_no_twiddle[1][1][7] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~42 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[1][1][7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~42_combout ),
	.cout());
defparam \reg_no_twiddle~42 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~42 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[1][1][3] (
	.clk(clk),
	.d(\reg_no_twiddle~53_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[1][1][3]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[1][1][3] .is_wysiwyg = "true";
defparam \reg_no_twiddle[1][1][3] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~43 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[1][1][3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~43_combout ),
	.cout());
defparam \reg_no_twiddle~43 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~43 .sum_lutc_input = "datac";

dffeas \do_tdl[0][0][0][3] (
	.clk(clk),
	.d(\reg_no_twiddle[6][0][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][0][0][3]~q ),
	.prn(vcc));
defparam \do_tdl[0][0][0][3] .is_wysiwyg = "true";
defparam \do_tdl[0][0][0][3] .power_up = "low";

dffeas \do_tdl[0][0][0][7] (
	.clk(clk),
	.d(\reg_no_twiddle[6][0][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][0][0][7]~q ),
	.prn(vcc));
defparam \do_tdl[0][0][0][7] .is_wysiwyg = "true";
defparam \do_tdl[0][0][0][7] .power_up = "low";

dffeas \do_tdl[0][0][0][4] (
	.clk(clk),
	.d(\reg_no_twiddle[6][0][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][0][0][4]~q ),
	.prn(vcc));
defparam \do_tdl[0][0][0][4] .is_wysiwyg = "true";
defparam \do_tdl[0][0][0][4] .power_up = "low";

dffeas \do_tdl[0][0][0][5] (
	.clk(clk),
	.d(\reg_no_twiddle[6][0][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][0][0][5]~q ),
	.prn(vcc));
defparam \do_tdl[0][0][0][5] .is_wysiwyg = "true";
defparam \do_tdl[0][0][0][5] .power_up = "low";

dffeas \do_tdl[0][0][0][6] (
	.clk(clk),
	.d(\reg_no_twiddle[6][0][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][0][0][6]~q ),
	.prn(vcc));
defparam \do_tdl[0][0][0][6] .is_wysiwyg = "true";
defparam \do_tdl[0][0][0][6] .power_up = "low";

dffeas \do_tdl[0][0][0][1] (
	.clk(clk),
	.d(\reg_no_twiddle[6][0][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][0][0][1]~q ),
	.prn(vcc));
defparam \do_tdl[0][0][0][1] .is_wysiwyg = "true";
defparam \do_tdl[0][0][0][1] .power_up = "low";

dffeas \do_tdl[0][0][0][0] (
	.clk(clk),
	.d(\reg_no_twiddle[6][0][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][0][0][0]~q ),
	.prn(vcc));
defparam \do_tdl[0][0][0][0] .is_wysiwyg = "true";
defparam \do_tdl[0][0][0][0] .power_up = "low";

dffeas \do_tdl[0][0][0][2] (
	.clk(clk),
	.d(\reg_no_twiddle[6][0][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][0][0][2]~q ),
	.prn(vcc));
defparam \do_tdl[0][0][0][2] .is_wysiwyg = "true";
defparam \do_tdl[0][0][0][2] .power_up = "low";

dffeas \do_tdl[0][1][0][3] (
	.clk(clk),
	.d(\reg_no_twiddle[6][1][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][1][0][3]~q ),
	.prn(vcc));
defparam \do_tdl[0][1][0][3] .is_wysiwyg = "true";
defparam \do_tdl[0][1][0][3] .power_up = "low";

dffeas \do_tdl[0][1][0][7] (
	.clk(clk),
	.d(\reg_no_twiddle[6][1][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][1][0][7]~q ),
	.prn(vcc));
defparam \do_tdl[0][1][0][7] .is_wysiwyg = "true";
defparam \do_tdl[0][1][0][7] .power_up = "low";

dffeas \do_tdl[0][1][0][4] (
	.clk(clk),
	.d(\reg_no_twiddle[6][1][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][1][0][4]~q ),
	.prn(vcc));
defparam \do_tdl[0][1][0][4] .is_wysiwyg = "true";
defparam \do_tdl[0][1][0][4] .power_up = "low";

dffeas \do_tdl[0][1][0][5] (
	.clk(clk),
	.d(\reg_no_twiddle[6][1][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][1][0][5]~q ),
	.prn(vcc));
defparam \do_tdl[0][1][0][5] .is_wysiwyg = "true";
defparam \do_tdl[0][1][0][5] .power_up = "low";

dffeas \do_tdl[0][1][0][6] (
	.clk(clk),
	.d(\reg_no_twiddle[6][1][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][1][0][6]~q ),
	.prn(vcc));
defparam \do_tdl[0][1][0][6] .is_wysiwyg = "true";
defparam \do_tdl[0][1][0][6] .power_up = "low";

dffeas \do_tdl[0][1][0][1] (
	.clk(clk),
	.d(\reg_no_twiddle[6][1][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][1][0][1]~q ),
	.prn(vcc));
defparam \do_tdl[0][1][0][1] .is_wysiwyg = "true";
defparam \do_tdl[0][1][0][1] .power_up = "low";

dffeas \do_tdl[0][1][0][0] (
	.clk(clk),
	.d(\reg_no_twiddle[6][1][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][1][0][0]~q ),
	.prn(vcc));
defparam \do_tdl[0][1][0][0] .is_wysiwyg = "true";
defparam \do_tdl[0][1][0][0] .power_up = "low";

dffeas \do_tdl[0][1][0][2] (
	.clk(clk),
	.d(\reg_no_twiddle[6][1][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[0][1][0][2]~q ),
	.prn(vcc));
defparam \do_tdl[0][1][0][2] .is_wysiwyg = "true";
defparam \do_tdl[0][1][0][2] .power_up = "low";

dffeas \do_tdl[1][0][0][3] (
	.clk(clk),
	.d(\gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][0][0][3]~q ),
	.prn(vcc));
defparam \do_tdl[1][0][0][3] .is_wysiwyg = "true";
defparam \do_tdl[1][0][0][3] .power_up = "low";

dffeas \do_tdl[1][0][0][7] (
	.clk(clk),
	.d(\gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][0][0][7]~q ),
	.prn(vcc));
defparam \do_tdl[1][0][0][7] .is_wysiwyg = "true";
defparam \do_tdl[1][0][0][7] .power_up = "low";

dffeas \do_tdl[1][0][0][4] (
	.clk(clk),
	.d(\gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][0][0][4]~q ),
	.prn(vcc));
defparam \do_tdl[1][0][0][4] .is_wysiwyg = "true";
defparam \do_tdl[1][0][0][4] .power_up = "low";

dffeas \do_tdl[1][0][0][5] (
	.clk(clk),
	.d(\gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][0][0][5]~q ),
	.prn(vcc));
defparam \do_tdl[1][0][0][5] .is_wysiwyg = "true";
defparam \do_tdl[1][0][0][5] .power_up = "low";

dffeas \do_tdl[1][0][0][6] (
	.clk(clk),
	.d(\gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][0][0][6]~q ),
	.prn(vcc));
defparam \do_tdl[1][0][0][6] .is_wysiwyg = "true";
defparam \do_tdl[1][0][0][6] .power_up = "low";

dffeas \do_tdl[1][0][0][1] (
	.clk(clk),
	.d(\gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][0][0][1]~q ),
	.prn(vcc));
defparam \do_tdl[1][0][0][1] .is_wysiwyg = "true";
defparam \do_tdl[1][0][0][1] .power_up = "low";

dffeas \do_tdl[1][0][0][0] (
	.clk(clk),
	.d(\gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][0][0][0]~q ),
	.prn(vcc));
defparam \do_tdl[1][0][0][0] .is_wysiwyg = "true";
defparam \do_tdl[1][0][0][0] .power_up = "low";

dffeas \do_tdl[1][0][0][2] (
	.clk(clk),
	.d(\gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][0][0][2]~q ),
	.prn(vcc));
defparam \do_tdl[1][0][0][2] .is_wysiwyg = "true";
defparam \do_tdl[1][0][0][2] .power_up = "low";

dffeas \do_tdl[1][1][0][3] (
	.clk(clk),
	.d(\gen_da0:gen_canonic:cm1|real_out[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][1][0][3]~q ),
	.prn(vcc));
defparam \do_tdl[1][1][0][3] .is_wysiwyg = "true";
defparam \do_tdl[1][1][0][3] .power_up = "low";

dffeas \do_tdl[1][1][0][7] (
	.clk(clk),
	.d(\gen_da0:gen_canonic:cm1|real_out[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][1][0][7]~q ),
	.prn(vcc));
defparam \do_tdl[1][1][0][7] .is_wysiwyg = "true";
defparam \do_tdl[1][1][0][7] .power_up = "low";

dffeas \do_tdl[1][1][0][4] (
	.clk(clk),
	.d(\gen_da0:gen_canonic:cm1|real_out[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][1][0][4]~q ),
	.prn(vcc));
defparam \do_tdl[1][1][0][4] .is_wysiwyg = "true";
defparam \do_tdl[1][1][0][4] .power_up = "low";

dffeas \do_tdl[1][1][0][5] (
	.clk(clk),
	.d(\gen_da0:gen_canonic:cm1|real_out[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][1][0][5]~q ),
	.prn(vcc));
defparam \do_tdl[1][1][0][5] .is_wysiwyg = "true";
defparam \do_tdl[1][1][0][5] .power_up = "low";

dffeas \do_tdl[1][1][0][6] (
	.clk(clk),
	.d(\gen_da0:gen_canonic:cm1|real_out[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][1][0][6]~q ),
	.prn(vcc));
defparam \do_tdl[1][1][0][6] .is_wysiwyg = "true";
defparam \do_tdl[1][1][0][6] .power_up = "low";

dffeas \do_tdl[1][1][0][1] (
	.clk(clk),
	.d(\gen_da0:gen_canonic:cm1|real_out[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][1][0][1]~q ),
	.prn(vcc));
defparam \do_tdl[1][1][0][1] .is_wysiwyg = "true";
defparam \do_tdl[1][1][0][1] .power_up = "low";

dffeas \do_tdl[1][1][0][0] (
	.clk(clk),
	.d(\gen_da0:gen_canonic:cm1|real_out[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][1][0][0]~q ),
	.prn(vcc));
defparam \do_tdl[1][1][0][0] .is_wysiwyg = "true";
defparam \do_tdl[1][1][0][0] .power_up = "low";

dffeas \do_tdl[1][1][0][2] (
	.clk(clk),
	.d(\gen_da0:gen_canonic:cm1|real_out[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[1][1][0][2]~q ),
	.prn(vcc));
defparam \do_tdl[1][1][0][2] .is_wysiwyg = "true";
defparam \do_tdl[1][1][0][2] .power_up = "low";

dffeas \do_tdl[2][0][0][3] (
	.clk(clk),
	.d(\gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][0][0][3]~q ),
	.prn(vcc));
defparam \do_tdl[2][0][0][3] .is_wysiwyg = "true";
defparam \do_tdl[2][0][0][3] .power_up = "low";

dffeas \do_tdl[2][0][0][7] (
	.clk(clk),
	.d(\gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][0][0][7]~q ),
	.prn(vcc));
defparam \do_tdl[2][0][0][7] .is_wysiwyg = "true";
defparam \do_tdl[2][0][0][7] .power_up = "low";

dffeas \do_tdl[2][0][0][4] (
	.clk(clk),
	.d(\gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][0][0][4]~q ),
	.prn(vcc));
defparam \do_tdl[2][0][0][4] .is_wysiwyg = "true";
defparam \do_tdl[2][0][0][4] .power_up = "low";

dffeas \do_tdl[2][0][0][5] (
	.clk(clk),
	.d(\gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][0][0][5]~q ),
	.prn(vcc));
defparam \do_tdl[2][0][0][5] .is_wysiwyg = "true";
defparam \do_tdl[2][0][0][5] .power_up = "low";

dffeas \do_tdl[2][0][0][6] (
	.clk(clk),
	.d(\gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][0][0][6]~q ),
	.prn(vcc));
defparam \do_tdl[2][0][0][6] .is_wysiwyg = "true";
defparam \do_tdl[2][0][0][6] .power_up = "low";

dffeas \do_tdl[2][0][0][1] (
	.clk(clk),
	.d(\gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][0][0][1]~q ),
	.prn(vcc));
defparam \do_tdl[2][0][0][1] .is_wysiwyg = "true";
defparam \do_tdl[2][0][0][1] .power_up = "low";

dffeas \do_tdl[2][0][0][0] (
	.clk(clk),
	.d(\gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][0][0][0]~q ),
	.prn(vcc));
defparam \do_tdl[2][0][0][0] .is_wysiwyg = "true";
defparam \do_tdl[2][0][0][0] .power_up = "low";

dffeas \do_tdl[2][0][0][2] (
	.clk(clk),
	.d(\gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][0][0][2]~q ),
	.prn(vcc));
defparam \do_tdl[2][0][0][2] .is_wysiwyg = "true";
defparam \do_tdl[2][0][0][2] .power_up = "low";

dffeas \do_tdl[2][1][0][3] (
	.clk(clk),
	.d(\gen_da0:gen_canonic:cm2|real_out[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][1][0][3]~q ),
	.prn(vcc));
defparam \do_tdl[2][1][0][3] .is_wysiwyg = "true";
defparam \do_tdl[2][1][0][3] .power_up = "low";

dffeas \do_tdl[2][1][0][7] (
	.clk(clk),
	.d(\gen_da0:gen_canonic:cm2|real_out[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][1][0][7]~q ),
	.prn(vcc));
defparam \do_tdl[2][1][0][7] .is_wysiwyg = "true";
defparam \do_tdl[2][1][0][7] .power_up = "low";

dffeas \do_tdl[2][1][0][4] (
	.clk(clk),
	.d(\gen_da0:gen_canonic:cm2|real_out[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][1][0][4]~q ),
	.prn(vcc));
defparam \do_tdl[2][1][0][4] .is_wysiwyg = "true";
defparam \do_tdl[2][1][0][4] .power_up = "low";

dffeas \do_tdl[2][1][0][5] (
	.clk(clk),
	.d(\gen_da0:gen_canonic:cm2|real_out[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][1][0][5]~q ),
	.prn(vcc));
defparam \do_tdl[2][1][0][5] .is_wysiwyg = "true";
defparam \do_tdl[2][1][0][5] .power_up = "low";

dffeas \do_tdl[2][1][0][6] (
	.clk(clk),
	.d(\gen_da0:gen_canonic:cm2|real_out[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][1][0][6]~q ),
	.prn(vcc));
defparam \do_tdl[2][1][0][6] .is_wysiwyg = "true";
defparam \do_tdl[2][1][0][6] .power_up = "low";

dffeas \do_tdl[2][1][0][1] (
	.clk(clk),
	.d(\gen_da0:gen_canonic:cm2|real_out[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][1][0][1]~q ),
	.prn(vcc));
defparam \do_tdl[2][1][0][1] .is_wysiwyg = "true";
defparam \do_tdl[2][1][0][1] .power_up = "low";

dffeas \do_tdl[2][1][0][0] (
	.clk(clk),
	.d(\gen_da0:gen_canonic:cm2|real_out[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][1][0][0]~q ),
	.prn(vcc));
defparam \do_tdl[2][1][0][0] .is_wysiwyg = "true";
defparam \do_tdl[2][1][0][0] .power_up = "low";

dffeas \do_tdl[2][1][0][2] (
	.clk(clk),
	.d(\gen_da0:gen_canonic:cm2|real_out[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[2][1][0][2]~q ),
	.prn(vcc));
defparam \do_tdl[2][1][0][2] .is_wysiwyg = "true";
defparam \do_tdl[2][1][0][2] .power_up = "low";

dffeas \do_tdl[3][0][0][3] (
	.clk(clk),
	.d(\gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][0][0][3]~q ),
	.prn(vcc));
defparam \do_tdl[3][0][0][3] .is_wysiwyg = "true";
defparam \do_tdl[3][0][0][3] .power_up = "low";

dffeas \do_tdl[3][0][0][7] (
	.clk(clk),
	.d(\gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][0][0][7]~q ),
	.prn(vcc));
defparam \do_tdl[3][0][0][7] .is_wysiwyg = "true";
defparam \do_tdl[3][0][0][7] .power_up = "low";

dffeas \do_tdl[3][0][0][4] (
	.clk(clk),
	.d(\gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][0][0][4]~q ),
	.prn(vcc));
defparam \do_tdl[3][0][0][4] .is_wysiwyg = "true";
defparam \do_tdl[3][0][0][4] .power_up = "low";

dffeas \do_tdl[3][0][0][5] (
	.clk(clk),
	.d(\gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][0][0][5]~q ),
	.prn(vcc));
defparam \do_tdl[3][0][0][5] .is_wysiwyg = "true";
defparam \do_tdl[3][0][0][5] .power_up = "low";

dffeas \do_tdl[3][0][0][6] (
	.clk(clk),
	.d(\gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][0][0][6]~q ),
	.prn(vcc));
defparam \do_tdl[3][0][0][6] .is_wysiwyg = "true";
defparam \do_tdl[3][0][0][6] .power_up = "low";

dffeas \do_tdl[3][0][0][1] (
	.clk(clk),
	.d(\gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][0][0][1]~q ),
	.prn(vcc));
defparam \do_tdl[3][0][0][1] .is_wysiwyg = "true";
defparam \do_tdl[3][0][0][1] .power_up = "low";

dffeas \do_tdl[3][0][0][0] (
	.clk(clk),
	.d(\gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][0][0][0]~q ),
	.prn(vcc));
defparam \do_tdl[3][0][0][0] .is_wysiwyg = "true";
defparam \do_tdl[3][0][0][0] .power_up = "low";

dffeas \do_tdl[3][0][0][2] (
	.clk(clk),
	.d(\gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][0][0][2]~q ),
	.prn(vcc));
defparam \do_tdl[3][0][0][2] .is_wysiwyg = "true";
defparam \do_tdl[3][0][0][2] .power_up = "low";

dffeas \do_tdl[3][1][0][3] (
	.clk(clk),
	.d(\gen_da0:gen_canonic:cm3|real_out[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][1][0][3]~q ),
	.prn(vcc));
defparam \do_tdl[3][1][0][3] .is_wysiwyg = "true";
defparam \do_tdl[3][1][0][3] .power_up = "low";

dffeas \do_tdl[3][1][0][7] (
	.clk(clk),
	.d(\gen_da0:gen_canonic:cm3|real_out[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][1][0][7]~q ),
	.prn(vcc));
defparam \do_tdl[3][1][0][7] .is_wysiwyg = "true";
defparam \do_tdl[3][1][0][7] .power_up = "low";

dffeas \do_tdl[3][1][0][4] (
	.clk(clk),
	.d(\gen_da0:gen_canonic:cm3|real_out[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][1][0][4]~q ),
	.prn(vcc));
defparam \do_tdl[3][1][0][4] .is_wysiwyg = "true";
defparam \do_tdl[3][1][0][4] .power_up = "low";

dffeas \do_tdl[3][1][0][5] (
	.clk(clk),
	.d(\gen_da0:gen_canonic:cm3|real_out[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][1][0][5]~q ),
	.prn(vcc));
defparam \do_tdl[3][1][0][5] .is_wysiwyg = "true";
defparam \do_tdl[3][1][0][5] .power_up = "low";

dffeas \do_tdl[3][1][0][6] (
	.clk(clk),
	.d(\gen_da0:gen_canonic:cm3|real_out[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][1][0][6]~q ),
	.prn(vcc));
defparam \do_tdl[3][1][0][6] .is_wysiwyg = "true";
defparam \do_tdl[3][1][0][6] .power_up = "low";

dffeas \do_tdl[3][1][0][1] (
	.clk(clk),
	.d(\gen_da0:gen_canonic:cm3|real_out[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][1][0][1]~q ),
	.prn(vcc));
defparam \do_tdl[3][1][0][1] .is_wysiwyg = "true";
defparam \do_tdl[3][1][0][1] .power_up = "low";

dffeas \do_tdl[3][1][0][0] (
	.clk(clk),
	.d(\gen_da0:gen_canonic:cm3|real_out[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][1][0][0]~q ),
	.prn(vcc));
defparam \do_tdl[3][1][0][0] .is_wysiwyg = "true";
defparam \do_tdl[3][1][0][0] .power_up = "low";

dffeas \do_tdl[3][1][0][2] (
	.clk(clk),
	.d(\gen_da0:gen_canonic:cm3|real_out[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\do_tdl[3][1][0][2]~q ),
	.prn(vcc));
defparam \do_tdl[3][1][0][2] .is_wysiwyg = "true";
defparam \do_tdl[3][1][0][2] .power_up = "low";

cycloneiii_lcell_comb \sdft~9 (
	.dataa(reset_n),
	.datab(\sdft.ENABLE_BFP_O~q ),
	.datac(\Equal1~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\sdft~9_combout ),
	.cout());
defparam \sdft~9 .lut_mask = 16'hFEFE;
defparam \sdft~9 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[1][0][4] (
	.clk(clk),
	.d(\reg_no_twiddle~54_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[1][0][4]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[1][0][4] .is_wysiwyg = "true";
defparam \reg_no_twiddle[1][0][4] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~44 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[1][0][4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~44_combout ),
	.cout());
defparam \reg_no_twiddle~44 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~44 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[1][1][4] (
	.clk(clk),
	.d(\reg_no_twiddle~55_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[1][1][4]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[1][1][4] .is_wysiwyg = "true";
defparam \reg_no_twiddle[1][1][4] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~45 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[1][1][4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~45_combout ),
	.cout());
defparam \reg_no_twiddle~45 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~45 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[1][0][5] (
	.clk(clk),
	.d(\reg_no_twiddle~56_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[1][0][5]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[1][0][5] .is_wysiwyg = "true";
defparam \reg_no_twiddle[1][0][5] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~46 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[1][0][5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~46_combout ),
	.cout());
defparam \reg_no_twiddle~46 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~46 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[1][1][5] (
	.clk(clk),
	.d(\reg_no_twiddle~57_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[1][1][5]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[1][1][5] .is_wysiwyg = "true";
defparam \reg_no_twiddle[1][1][5] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~47 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[1][1][5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~47_combout ),
	.cout());
defparam \reg_no_twiddle~47 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~47 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[1][0][6] (
	.clk(clk),
	.d(\reg_no_twiddle~58_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[1][0][6]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[1][0][6] .is_wysiwyg = "true";
defparam \reg_no_twiddle[1][0][6] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~48 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[1][0][6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~48_combout ),
	.cout());
defparam \reg_no_twiddle~48 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~48 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[1][1][6] (
	.clk(clk),
	.d(\reg_no_twiddle~59_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[1][1][6]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[1][1][6] .is_wysiwyg = "true";
defparam \reg_no_twiddle[1][1][6] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~49 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[1][1][6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~49_combout ),
	.cout());
defparam \reg_no_twiddle~49 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~49 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \reg_no_twiddle~50 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[0][0][3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~50_combout ),
	.cout());
defparam \reg_no_twiddle~50 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~50 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \reg_no_twiddle~51 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[0][0][7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~51_combout ),
	.cout());
defparam \reg_no_twiddle~51 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~51 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \reg_no_twiddle~52 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[0][1][7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~52_combout ),
	.cout());
defparam \reg_no_twiddle~52 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~52 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \reg_no_twiddle~53 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[0][1][3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~53_combout ),
	.cout());
defparam \reg_no_twiddle~53 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~53 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[6][0][1] (
	.clk(clk),
	.d(\reg_no_twiddle~62_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[6][0][1]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[6][0][1] .is_wysiwyg = "true";
defparam \reg_no_twiddle[6][0][1] .power_up = "low";

dffeas \reg_no_twiddle[6][0][0] (
	.clk(clk),
	.d(\reg_no_twiddle~63_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[6][0][0]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[6][0][0] .is_wysiwyg = "true";
defparam \reg_no_twiddle[6][0][0] .power_up = "low";

dffeas \reg_no_twiddle[6][0][2] (
	.clk(clk),
	.d(\reg_no_twiddle~64_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[6][0][2]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[6][0][2] .is_wysiwyg = "true";
defparam \reg_no_twiddle[6][0][2] .power_up = "low";

dffeas \reg_no_twiddle[6][1][1] (
	.clk(clk),
	.d(\reg_no_twiddle~65_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[6][1][1]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[6][1][1] .is_wysiwyg = "true";
defparam \reg_no_twiddle[6][1][1] .power_up = "low";

dffeas \reg_no_twiddle[6][1][0] (
	.clk(clk),
	.d(\reg_no_twiddle~66_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[6][1][0]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[6][1][0] .is_wysiwyg = "true";
defparam \reg_no_twiddle[6][1][0] .power_up = "low";

dffeas \reg_no_twiddle[6][1][2] (
	.clk(clk),
	.d(\reg_no_twiddle~67_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[6][1][2]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[6][1][2] .is_wysiwyg = "true";
defparam \reg_no_twiddle[6][1][2] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~54 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[0][0][4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~54_combout ),
	.cout());
defparam \reg_no_twiddle~54 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~54 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \reg_no_twiddle~55 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[0][1][4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~55_combout ),
	.cout());
defparam \reg_no_twiddle~55 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~55 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \reg_no_twiddle~56 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[0][0][5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~56_combout ),
	.cout());
defparam \reg_no_twiddle~56 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~56 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \reg_no_twiddle~57 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[0][1][5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~57_combout ),
	.cout());
defparam \reg_no_twiddle~57 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~57 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \reg_no_twiddle~58 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[0][0][6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~58_combout ),
	.cout());
defparam \reg_no_twiddle~58 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~58 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \reg_no_twiddle~59 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[0][1][6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~59_combout ),
	.cout());
defparam \reg_no_twiddle~59 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~59 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \reg_no_twiddle~60 (
	.dataa(\gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.cin(gnd),
	.combout(\reg_no_twiddle~60_combout ),
	.cout());
defparam \reg_no_twiddle~60 .lut_mask = 16'hAAFF;
defparam \reg_no_twiddle~60 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \reg_no_twiddle~61 (
	.dataa(\gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.cin(gnd),
	.combout(\reg_no_twiddle~61_combout ),
	.cout());
defparam \reg_no_twiddle~61 .lut_mask = 16'hAAFF;
defparam \reg_no_twiddle~61 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[5][0][1] (
	.clk(clk),
	.d(\reg_no_twiddle~68_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[5][0][1]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[5][0][1] .is_wysiwyg = "true";
defparam \reg_no_twiddle[5][0][1] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~62 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[5][0][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~62_combout ),
	.cout());
defparam \reg_no_twiddle~62 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~62 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[5][0][0] (
	.clk(clk),
	.d(\reg_no_twiddle~69_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[5][0][0]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[5][0][0] .is_wysiwyg = "true";
defparam \reg_no_twiddle[5][0][0] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~63 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[5][0][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~63_combout ),
	.cout());
defparam \reg_no_twiddle~63 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~63 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[5][0][2] (
	.clk(clk),
	.d(\reg_no_twiddle~70_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[5][0][2]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[5][0][2] .is_wysiwyg = "true";
defparam \reg_no_twiddle[5][0][2] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~64 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[5][0][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~64_combout ),
	.cout());
defparam \reg_no_twiddle~64 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~64 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[5][1][1] (
	.clk(clk),
	.d(\reg_no_twiddle~71_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[5][1][1]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[5][1][1] .is_wysiwyg = "true";
defparam \reg_no_twiddle[5][1][1] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~65 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[5][1][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~65_combout ),
	.cout());
defparam \reg_no_twiddle~65 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~65 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[5][1][0] (
	.clk(clk),
	.d(\reg_no_twiddle~72_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[5][1][0]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[5][1][0] .is_wysiwyg = "true";
defparam \reg_no_twiddle[5][1][0] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~66 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[5][1][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~66_combout ),
	.cout());
defparam \reg_no_twiddle~66 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~66 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[5][1][2] (
	.clk(clk),
	.d(\reg_no_twiddle~73_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[5][1][2]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[5][1][2] .is_wysiwyg = "true";
defparam \reg_no_twiddle[5][1][2] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~67 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[5][1][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~67_combout ),
	.cout());
defparam \reg_no_twiddle~67 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~67 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[4][0][1] (
	.clk(clk),
	.d(\reg_no_twiddle~74_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[4][0][1]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[4][0][1] .is_wysiwyg = "true";
defparam \reg_no_twiddle[4][0][1] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~68 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[4][0][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~68_combout ),
	.cout());
defparam \reg_no_twiddle~68 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~68 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[4][0][0] (
	.clk(clk),
	.d(\reg_no_twiddle~75_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[4][0][0]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[4][0][0] .is_wysiwyg = "true";
defparam \reg_no_twiddle[4][0][0] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~69 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[4][0][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~69_combout ),
	.cout());
defparam \reg_no_twiddle~69 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~69 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[4][0][2] (
	.clk(clk),
	.d(\reg_no_twiddle~76_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[4][0][2]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[4][0][2] .is_wysiwyg = "true";
defparam \reg_no_twiddle[4][0][2] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~70 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[4][0][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~70_combout ),
	.cout());
defparam \reg_no_twiddle~70 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~70 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[4][1][1] (
	.clk(clk),
	.d(\reg_no_twiddle~77_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[4][1][1]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[4][1][1] .is_wysiwyg = "true";
defparam \reg_no_twiddle[4][1][1] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~71 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[4][1][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~71_combout ),
	.cout());
defparam \reg_no_twiddle~71 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~71 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[4][1][0] (
	.clk(clk),
	.d(\reg_no_twiddle~78_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[4][1][0]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[4][1][0] .is_wysiwyg = "true";
defparam \reg_no_twiddle[4][1][0] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~72 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[4][1][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~72_combout ),
	.cout());
defparam \reg_no_twiddle~72 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~72 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[4][1][2] (
	.clk(clk),
	.d(\reg_no_twiddle~79_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[4][1][2]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[4][1][2] .is_wysiwyg = "true";
defparam \reg_no_twiddle[4][1][2] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~73 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[4][1][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~73_combout ),
	.cout());
defparam \reg_no_twiddle~73 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~73 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[3][0][1] (
	.clk(clk),
	.d(\reg_no_twiddle~80_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[3][0][1]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[3][0][1] .is_wysiwyg = "true";
defparam \reg_no_twiddle[3][0][1] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~74 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[3][0][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~74_combout ),
	.cout());
defparam \reg_no_twiddle~74 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~74 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[3][0][0] (
	.clk(clk),
	.d(\reg_no_twiddle~81_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[3][0][0]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[3][0][0] .is_wysiwyg = "true";
defparam \reg_no_twiddle[3][0][0] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~75 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[3][0][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~75_combout ),
	.cout());
defparam \reg_no_twiddle~75 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~75 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[3][0][2] (
	.clk(clk),
	.d(\reg_no_twiddle~82_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[3][0][2]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[3][0][2] .is_wysiwyg = "true";
defparam \reg_no_twiddle[3][0][2] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~76 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[3][0][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~76_combout ),
	.cout());
defparam \reg_no_twiddle~76 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~76 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[3][1][1] (
	.clk(clk),
	.d(\reg_no_twiddle~83_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[3][1][1]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[3][1][1] .is_wysiwyg = "true";
defparam \reg_no_twiddle[3][1][1] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~77 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[3][1][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~77_combout ),
	.cout());
defparam \reg_no_twiddle~77 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~77 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[3][1][0] (
	.clk(clk),
	.d(\reg_no_twiddle~84_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[3][1][0]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[3][1][0] .is_wysiwyg = "true";
defparam \reg_no_twiddle[3][1][0] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~78 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[3][1][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~78_combout ),
	.cout());
defparam \reg_no_twiddle~78 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~78 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[3][1][2] (
	.clk(clk),
	.d(\reg_no_twiddle~85_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[3][1][2]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[3][1][2] .is_wysiwyg = "true";
defparam \reg_no_twiddle[3][1][2] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~79 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[3][1][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~79_combout ),
	.cout());
defparam \reg_no_twiddle~79 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~79 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[2][0][1] (
	.clk(clk),
	.d(\reg_no_twiddle~86_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[2][0][1]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[2][0][1] .is_wysiwyg = "true";
defparam \reg_no_twiddle[2][0][1] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~80 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[2][0][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~80_combout ),
	.cout());
defparam \reg_no_twiddle~80 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~80 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[2][0][0] (
	.clk(clk),
	.d(\reg_no_twiddle~87_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[2][0][0]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[2][0][0] .is_wysiwyg = "true";
defparam \reg_no_twiddle[2][0][0] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~81 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[2][0][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~81_combout ),
	.cout());
defparam \reg_no_twiddle~81 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~81 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[2][0][2] (
	.clk(clk),
	.d(\reg_no_twiddle~88_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[2][0][2]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[2][0][2] .is_wysiwyg = "true";
defparam \reg_no_twiddle[2][0][2] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~82 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[2][0][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~82_combout ),
	.cout());
defparam \reg_no_twiddle~82 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~82 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[2][1][1] (
	.clk(clk),
	.d(\reg_no_twiddle~89_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[2][1][1]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[2][1][1] .is_wysiwyg = "true";
defparam \reg_no_twiddle[2][1][1] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~83 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[2][1][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~83_combout ),
	.cout());
defparam \reg_no_twiddle~83 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~83 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[2][1][0] (
	.clk(clk),
	.d(\reg_no_twiddle~90_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[2][1][0]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[2][1][0] .is_wysiwyg = "true";
defparam \reg_no_twiddle[2][1][0] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~84 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[2][1][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~84_combout ),
	.cout());
defparam \reg_no_twiddle~84 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~84 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[2][1][2] (
	.clk(clk),
	.d(\reg_no_twiddle~91_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[2][1][2]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[2][1][2] .is_wysiwyg = "true";
defparam \reg_no_twiddle[2][1][2] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~85 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[2][1][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~85_combout ),
	.cout());
defparam \reg_no_twiddle~85 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~85 .sum_lutc_input = "datac";

dffeas block_dft_i_en(
	.clk(clk),
	.d(\Selector4~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\block_dft_i_en~q ),
	.prn(vcc));
defparam block_dft_i_en.is_wysiwyg = "true";
defparam block_dft_i_en.power_up = "low";

cycloneiii_lcell_comb \slb_nm1[1] (
	.dataa(\block_dft_i_en~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\slb_nm1[1]~combout ),
	.cout());
defparam \slb_nm1[1] .lut_mask = 16'hAAFF;
defparam \slb_nm1[1] .sum_lutc_input = "datac";

cycloneiii_lcell_comb \slb_nm1[2]~0 (
	.dataa(slb_last_2),
	.datab(gnd),
	.datac(gnd),
	.datad(\block_dft_i_en~q ),
	.cin(gnd),
	.combout(\slb_nm1[2]~0_combout ),
	.cout());
defparam \slb_nm1[2]~0 .lut_mask = 16'hAAFF;
defparam \slb_nm1[2]~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \slb_nm1[0] (
	.dataa(slb_last_0),
	.datab(gnd),
	.datac(gnd),
	.datad(\block_dft_i_en~q ),
	.cin(gnd),
	.combout(\slb_nm1[0]~combout ),
	.cout());
defparam \slb_nm1[0] .lut_mask = 16'hAAFF;
defparam \slb_nm1[0] .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[1][0][1] (
	.clk(clk),
	.d(\reg_no_twiddle~92_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[1][0][1]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[1][0][1] .is_wysiwyg = "true";
defparam \reg_no_twiddle[1][0][1] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~86 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[1][0][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~86_combout ),
	.cout());
defparam \reg_no_twiddle~86 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~86 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[1][0][0] (
	.clk(clk),
	.d(\reg_no_twiddle~93_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[1][0][0]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[1][0][0] .is_wysiwyg = "true";
defparam \reg_no_twiddle[1][0][0] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~87 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[1][0][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~87_combout ),
	.cout());
defparam \reg_no_twiddle~87 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~87 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[1][0][2] (
	.clk(clk),
	.d(\reg_no_twiddle~94_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[1][0][2]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[1][0][2] .is_wysiwyg = "true";
defparam \reg_no_twiddle[1][0][2] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~88 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[1][0][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~88_combout ),
	.cout());
defparam \reg_no_twiddle~88 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~88 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[1][1][1] (
	.clk(clk),
	.d(\reg_no_twiddle~95_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[1][1][1]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[1][1][1] .is_wysiwyg = "true";
defparam \reg_no_twiddle[1][1][1] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~89 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[1][1][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~89_combout ),
	.cout());
defparam \reg_no_twiddle~89 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~89 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[1][1][0] (
	.clk(clk),
	.d(\reg_no_twiddle~96_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[1][1][0]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[1][1][0] .is_wysiwyg = "true";
defparam \reg_no_twiddle[1][1][0] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~90 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[1][1][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~90_combout ),
	.cout());
defparam \reg_no_twiddle~90 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~90 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[1][1][2] (
	.clk(clk),
	.d(\reg_no_twiddle~97_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[1][1][2]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[1][1][2] .is_wysiwyg = "true";
defparam \reg_no_twiddle[1][1][2] .power_up = "low";

cycloneiii_lcell_comb \reg_no_twiddle~91 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[1][1][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~91_combout ),
	.cout());
defparam \reg_no_twiddle~91 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~91 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector4~0 (
	.dataa(\sdft.WAIT_FOR_OUTPUT~q ),
	.datab(\sdft.BLOCK_DFT_I~q ),
	.datac(\sdft.ENABLE_DFT_O~q ),
	.datad(\gap_reg~q ),
	.cin(gnd),
	.combout(\Selector4~0_combout ),
	.cout());
defparam \Selector4~0 .lut_mask = 16'hFFFE;
defparam \Selector4~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \reg_no_twiddle~92 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[0][0][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~92_combout ),
	.cout());
defparam \reg_no_twiddle~92 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~92 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \reg_no_twiddle~93 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[0][0][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~93_combout ),
	.cout());
defparam \reg_no_twiddle~93 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~93 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \reg_no_twiddle~94 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[0][0][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~94_combout ),
	.cout());
defparam \reg_no_twiddle~94 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~94 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \reg_no_twiddle~95 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[0][1][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~95_combout ),
	.cout());
defparam \reg_no_twiddle~95 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~95 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \reg_no_twiddle~96 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[0][1][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~96_combout ),
	.cout());
defparam \reg_no_twiddle~96 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~96 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \reg_no_twiddle~97 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[0][1][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~97_combout ),
	.cout());
defparam \reg_no_twiddle~97 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~97 .sum_lutc_input = "datac";

dffeas \blk_done_vec[2] (
	.clk(clk),
	.d(\blk_done_vec~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(blk_done_vec_2),
	.prn(vcc));
defparam \blk_done_vec[2] .is_wysiwyg = "true";
defparam \blk_done_vec[2] .power_up = "low";

dffeas \next_pass_vec[2] (
	.clk(clk),
	.d(\next_pass_vec~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(next_pass_vec_2),
	.prn(vcc));
defparam \next_pass_vec[2] .is_wysiwyg = "true";
defparam \next_pass_vec[2] .power_up = "low";

cycloneiii_lcell_comb \blk_done_vec~2 (
	.dataa(reset_n),
	.datab(tdl_arr_5),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\blk_done_vec~2_combout ),
	.cout());
defparam \blk_done_vec~2 .lut_mask = 16'hEEEE;
defparam \blk_done_vec~2 .sum_lutc_input = "datac";

dffeas \blk_done_vec[0] (
	.clk(clk),
	.d(\blk_done_vec~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\blk_done_vec[0]~q ),
	.prn(vcc));
defparam \blk_done_vec[0] .is_wysiwyg = "true";
defparam \blk_done_vec[0] .power_up = "low";

cycloneiii_lcell_comb \blk_done_vec~1 (
	.dataa(reset_n),
	.datab(\blk_done_vec[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\blk_done_vec~1_combout ),
	.cout());
defparam \blk_done_vec~1 .lut_mask = 16'hEEEE;
defparam \blk_done_vec~1 .sum_lutc_input = "datac";

dffeas \blk_done_vec[1] (
	.clk(clk),
	.d(\blk_done_vec~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\blk_done_vec[1]~q ),
	.prn(vcc));
defparam \blk_done_vec[1] .is_wysiwyg = "true";
defparam \blk_done_vec[1] .power_up = "low";

cycloneiii_lcell_comb \blk_done_vec~0 (
	.dataa(reset_n),
	.datab(\blk_done_vec[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\blk_done_vec~0_combout ),
	.cout());
defparam \blk_done_vec~0 .lut_mask = 16'hEEEE;
defparam \blk_done_vec~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \next_pass_vec~2 (
	.dataa(reset_n),
	.datab(tdl_arr_51),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\next_pass_vec~2_combout ),
	.cout());
defparam \next_pass_vec~2 .lut_mask = 16'hEEEE;
defparam \next_pass_vec~2 .sum_lutc_input = "datac";

dffeas \next_pass_vec[0] (
	.clk(clk),
	.d(\next_pass_vec~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\next_pass_vec[0]~q ),
	.prn(vcc));
defparam \next_pass_vec[0] .is_wysiwyg = "true";
defparam \next_pass_vec[0] .power_up = "low";

cycloneiii_lcell_comb \next_pass_vec~1 (
	.dataa(reset_n),
	.datab(\next_pass_vec[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\next_pass_vec~1_combout ),
	.cout());
defparam \next_pass_vec~1 .lut_mask = 16'hEEEE;
defparam \next_pass_vec~1 .sum_lutc_input = "datac";

dffeas \next_pass_vec[1] (
	.clk(clk),
	.d(\next_pass_vec~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\next_pass_vec[1]~q ),
	.prn(vcc));
defparam \next_pass_vec[1] .is_wysiwyg = "true";
defparam \next_pass_vec[1] .power_up = "low";

cycloneiii_lcell_comb \next_pass_vec~0 (
	.dataa(reset_n),
	.datab(\next_pass_vec[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\next_pass_vec~0_combout ),
	.cout());
defparam \next_pass_vec~0 .lut_mask = 16'hEEEE;
defparam \next_pass_vec~0 .sum_lutc_input = "datac";

endmodule

module fft_asj_fft_bfp_i_fft_120 (
	r_array_out_5_0,
	r_array_out_5_2,
	r_array_out_4_0,
	r_array_out_4_2,
	r_array_out_3_0,
	r_array_out_3_2,
	r_array_out_2_0,
	r_array_out_2_2,
	r_array_out_5_1,
	r_array_out_5_3,
	r_array_out_4_1,
	r_array_out_4_3,
	r_array_out_3_1,
	r_array_out_3_3,
	r_array_out_2_1,
	r_array_out_2_3,
	i_array_out_5_0,
	i_array_out_5_2,
	i_array_out_4_0,
	i_array_out_4_2,
	i_array_out_3_0,
	i_array_out_3_2,
	i_array_out_2_0,
	i_array_out_2_2,
	i_array_out_5_1,
	i_array_out_5_3,
	i_array_out_4_1,
	i_array_out_4_3,
	i_array_out_3_1,
	i_array_out_3_3,
	i_array_out_2_1,
	i_array_out_2_3,
	ram_in_reg_2_0,
	ram_in_reg_6_0,
	ram_in_reg_4_0,
	ram_in_reg_3_0,
	ram_in_reg_5_0,
	ram_in_reg_2_2,
	ram_in_reg_6_2,
	ram_in_reg_4_2,
	ram_in_reg_3_2,
	ram_in_reg_5_2,
	ram_in_reg_1_0,
	ram_in_reg_1_2,
	ram_in_reg_0_0,
	ram_in_reg_0_2,
	ram_in_reg_2_1,
	ram_in_reg_6_1,
	ram_in_reg_4_1,
	ram_in_reg_3_1,
	ram_in_reg_5_1,
	ram_in_reg_2_3,
	ram_in_reg_6_3,
	ram_in_reg_4_3,
	ram_in_reg_3_3,
	ram_in_reg_5_3,
	ram_in_reg_1_1,
	ram_in_reg_1_3,
	ram_in_reg_0_1,
	ram_in_reg_0_3,
	ram_in_reg_7_0,
	ram_in_reg_7_2,
	ram_in_reg_7_1,
	ram_in_reg_7_3,
	ram_in_reg_7_4,
	ram_in_reg_3_4,
	ram_in_reg_5_4,
	ram_in_reg_4_4,
	ram_in_reg_6_4,
	ram_in_reg_7_6,
	ram_in_reg_3_6,
	ram_in_reg_5_6,
	ram_in_reg_4_6,
	ram_in_reg_6_6,
	ram_in_reg_2_4,
	ram_in_reg_2_6,
	ram_in_reg_1_4,
	ram_in_reg_1_6,
	ram_in_reg_0_4,
	ram_in_reg_0_6,
	ram_in_reg_7_5,
	ram_in_reg_3_5,
	ram_in_reg_5_5,
	ram_in_reg_4_5,
	ram_in_reg_6_5,
	ram_in_reg_3_7,
	ram_in_reg_7_7,
	ram_in_reg_5_7,
	ram_in_reg_4_7,
	ram_in_reg_6_7,
	ram_in_reg_2_5,
	ram_in_reg_2_7,
	ram_in_reg_1_5,
	ram_in_reg_1_7,
	ram_in_reg_0_5,
	ram_in_reg_0_7,
	global_clock_enable,
	slb_last_0,
	slb_last_1,
	slb_last_2,
	r_array_out_6_0,
	r_array_out_6_2,
	r_array_out_1_0,
	r_array_out_1_2,
	r_array_out_0_0,
	r_array_out_0_2,
	r_array_out_6_1,
	r_array_out_6_3,
	r_array_out_1_1,
	r_array_out_1_3,
	r_array_out_0_1,
	r_array_out_0_3,
	r_array_out_7_0,
	r_array_out_7_2,
	r_array_out_7_1,
	r_array_out_7_3,
	i_array_out_7_0,
	i_array_out_7_2,
	i_array_out_6_0,
	i_array_out_6_2,
	i_array_out_1_0,
	i_array_out_1_2,
	i_array_out_0_0,
	i_array_out_0_2,
	i_array_out_7_1,
	i_array_out_7_3,
	i_array_out_6_1,
	i_array_out_6_3,
	i_array_out_1_1,
	i_array_out_1_3,
	i_array_out_0_1,
	i_array_out_0_3,
	block_dft_i_en,
	slb_nm1_1,
	slb_nm1_2,
	slb_nm1_0,
	clk)/* synthesis synthesis_greybox=1 */;
output 	r_array_out_5_0;
output 	r_array_out_5_2;
output 	r_array_out_4_0;
output 	r_array_out_4_2;
output 	r_array_out_3_0;
output 	r_array_out_3_2;
output 	r_array_out_2_0;
output 	r_array_out_2_2;
output 	r_array_out_5_1;
output 	r_array_out_5_3;
output 	r_array_out_4_1;
output 	r_array_out_4_3;
output 	r_array_out_3_1;
output 	r_array_out_3_3;
output 	r_array_out_2_1;
output 	r_array_out_2_3;
output 	i_array_out_5_0;
output 	i_array_out_5_2;
output 	i_array_out_4_0;
output 	i_array_out_4_2;
output 	i_array_out_3_0;
output 	i_array_out_3_2;
output 	i_array_out_2_0;
output 	i_array_out_2_2;
output 	i_array_out_5_1;
output 	i_array_out_5_3;
output 	i_array_out_4_1;
output 	i_array_out_4_3;
output 	i_array_out_3_1;
output 	i_array_out_3_3;
output 	i_array_out_2_1;
output 	i_array_out_2_3;
input 	ram_in_reg_2_0;
input 	ram_in_reg_6_0;
input 	ram_in_reg_4_0;
input 	ram_in_reg_3_0;
input 	ram_in_reg_5_0;
input 	ram_in_reg_2_2;
input 	ram_in_reg_6_2;
input 	ram_in_reg_4_2;
input 	ram_in_reg_3_2;
input 	ram_in_reg_5_2;
input 	ram_in_reg_1_0;
input 	ram_in_reg_1_2;
input 	ram_in_reg_0_0;
input 	ram_in_reg_0_2;
input 	ram_in_reg_2_1;
input 	ram_in_reg_6_1;
input 	ram_in_reg_4_1;
input 	ram_in_reg_3_1;
input 	ram_in_reg_5_1;
input 	ram_in_reg_2_3;
input 	ram_in_reg_6_3;
input 	ram_in_reg_4_3;
input 	ram_in_reg_3_3;
input 	ram_in_reg_5_3;
input 	ram_in_reg_1_1;
input 	ram_in_reg_1_3;
input 	ram_in_reg_0_1;
input 	ram_in_reg_0_3;
input 	ram_in_reg_7_0;
input 	ram_in_reg_7_2;
input 	ram_in_reg_7_1;
input 	ram_in_reg_7_3;
input 	ram_in_reg_7_4;
input 	ram_in_reg_3_4;
input 	ram_in_reg_5_4;
input 	ram_in_reg_4_4;
input 	ram_in_reg_6_4;
input 	ram_in_reg_7_6;
input 	ram_in_reg_3_6;
input 	ram_in_reg_5_6;
input 	ram_in_reg_4_6;
input 	ram_in_reg_6_6;
input 	ram_in_reg_2_4;
input 	ram_in_reg_2_6;
input 	ram_in_reg_1_4;
input 	ram_in_reg_1_6;
input 	ram_in_reg_0_4;
input 	ram_in_reg_0_6;
input 	ram_in_reg_7_5;
input 	ram_in_reg_3_5;
input 	ram_in_reg_5_5;
input 	ram_in_reg_4_5;
input 	ram_in_reg_6_5;
input 	ram_in_reg_3_7;
input 	ram_in_reg_7_7;
input 	ram_in_reg_5_7;
input 	ram_in_reg_4_7;
input 	ram_in_reg_6_7;
input 	ram_in_reg_2_5;
input 	ram_in_reg_2_7;
input 	ram_in_reg_1_5;
input 	ram_in_reg_1_7;
input 	ram_in_reg_0_5;
input 	ram_in_reg_0_7;
input 	global_clock_enable;
input 	slb_last_0;
input 	slb_last_1;
input 	slb_last_2;
output 	r_array_out_6_0;
output 	r_array_out_6_2;
output 	r_array_out_1_0;
output 	r_array_out_1_2;
output 	r_array_out_0_0;
output 	r_array_out_0_2;
output 	r_array_out_6_1;
output 	r_array_out_6_3;
output 	r_array_out_1_1;
output 	r_array_out_1_3;
output 	r_array_out_0_1;
output 	r_array_out_0_3;
output 	r_array_out_7_0;
output 	r_array_out_7_2;
output 	r_array_out_7_1;
output 	r_array_out_7_3;
output 	i_array_out_7_0;
output 	i_array_out_7_2;
output 	i_array_out_6_0;
output 	i_array_out_6_2;
output 	i_array_out_1_0;
output 	i_array_out_1_2;
output 	i_array_out_0_0;
output 	i_array_out_0_2;
output 	i_array_out_7_1;
output 	i_array_out_7_3;
output 	i_array_out_6_1;
output 	i_array_out_6_3;
output 	i_array_out_1_1;
output 	i_array_out_1_3;
output 	i_array_out_0_1;
output 	i_array_out_0_3;
input 	block_dft_i_en;
input 	slb_nm1_1;
input 	slb_nm1_2;
input 	slb_nm1_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Mux0~1_combout ;
wire \Mux0~2_combout ;
wire \r_array_out[0][5]~14_combout ;
wire \Mux16~1_combout ;
wire \Mux16~2_combout ;
wire \r_array_out[2][5]~15_combout ;
wire \r_array_out[0][2]~8_combout ;
wire \Mux0~0_combout ;
wire \r_array_out[0][4]~12_combout ;
wire \r_array_out[2][2]~9_combout ;
wire \Mux16~0_combout ;
wire \r_array_out[2][4]~13_combout ;
wire \r_array_out[0][3]~10_combout ;
wire \r_array_out[2][3]~11_combout ;
wire \Mux0~3_combout ;
wire \Mux16~3_combout ;
wire \Mux8~1_combout ;
wire \Mux8~2_combout ;
wire \r_array_out[1][5]~6_combout ;
wire \Mux24~1_combout ;
wire \Mux24~2_combout ;
wire \r_array_out[3][5]~7_combout ;
wire \r_array_out[1][2]~0_combout ;
wire \Mux8~0_combout ;
wire \r_array_out[1][4]~4_combout ;
wire \r_array_out[3][2]~1_combout ;
wire \Mux24~0_combout ;
wire \r_array_out[3][4]~5_combout ;
wire \r_array_out[1][3]~2_combout ;
wire \r_array_out[3][3]~3_combout ;
wire \Mux8~3_combout ;
wire \Mux24~3_combout ;
wire \Mux32~4_combout ;
wire \Mux32~0_combout ;
wire \i_array_out[0][5]~6_combout ;
wire \Mux48~4_combout ;
wire \Mux48~0_combout ;
wire \i_array_out[2][5]~7_combout ;
wire \i_array_out[0][2]~0_combout ;
wire \Mux32~3_combout ;
wire \i_array_out[0][4]~4_combout ;
wire \i_array_out[2][2]~1_combout ;
wire \Mux48~3_combout ;
wire \i_array_out[2][4]~5_combout ;
wire \i_array_out[0][3]~2_combout ;
wire \i_array_out[2][3]~3_combout ;
wire \Mux32~5_combout ;
wire \Mux48~5_combout ;
wire \Mux40~4_combout ;
wire \Mux40~0_combout ;
wire \i_array_out[1][5]~14_combout ;
wire \Mux56~4_combout ;
wire \Mux56~0_combout ;
wire \i_array_out[3][5]~15_combout ;
wire \i_array_out[1][2]~8_combout ;
wire \Mux40~3_combout ;
wire \i_array_out[1][4]~12_combout ;
wire \i_array_out[3][2]~9_combout ;
wire \Mux56~3_combout ;
wire \i_array_out[3][4]~13_combout ;
wire \i_array_out[1][3]~10_combout ;
wire \i_array_out[3][3]~11_combout ;
wire \Mux40~5_combout ;
wire \Mux56~5_combout ;
wire \r_array_out[2][6]~16_combout ;
wire \r_array_out[2][6]~17_combout ;
wire \Mux1~0_combout ;
wire \Mux1~1_combout ;
wire \Mux17~0_combout ;
wire \Mux17~1_combout ;
wire \Mux6~2_combout ;
wire \Mux22~2_combout ;
wire \Mux7~0_combout ;
wire \Mux7~1_combout ;
wire \Mux23~0_combout ;
wire \Mux9~0_combout ;
wire \Mux9~1_combout ;
wire \Mux25~0_combout ;
wire \Mux25~1_combout ;
wire \Mux14~2_combout ;
wire \Mux30~2_combout ;
wire \Mux15~0_combout ;
wire \Mux31~0_combout ;
wire \Mux0~4_combout ;
wire \Mux0~5_combout ;
wire \Mux16~4_combout ;
wire \Mux16~5_combout ;
wire \Mux8~4_combout ;
wire \Mux8~5_combout ;
wire \Mux24~4_combout ;
wire \Mux24~5_combout ;
wire \Mux32~1_combout ;
wire \Mux32~2_combout ;
wire \Mux48~1_combout ;
wire \Mux48~2_combout ;
wire \Mux33~0_combout ;
wire \Mux33~1_combout ;
wire \Mux49~0_combout ;
wire \Mux49~1_combout ;
wire \Mux38~2_combout ;
wire \Mux54~2_combout ;
wire \Mux39~0_combout ;
wire \Mux55~0_combout ;
wire \Mux40~1_combout ;
wire \Mux40~2_combout ;
wire \Mux56~1_combout ;
wire \Mux56~2_combout ;
wire \Mux41~0_combout ;
wire \Mux41~1_combout ;
wire \Mux57~0_combout ;
wire \Mux57~1_combout ;
wire \Mux46~2_combout ;
wire \Mux62~2_combout ;
wire \Mux47~0_combout ;
wire \Mux63~0_combout ;


dffeas \r_array_out[0][5] (
	.clk(clk),
	.d(\r_array_out[0][5]~14_combout ),
	.asdata(ram_in_reg_1_0),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_nm1_2),
	.ena(global_clock_enable),
	.q(r_array_out_5_0),
	.prn(vcc));
defparam \r_array_out[0][5] .is_wysiwyg = "true";
defparam \r_array_out[0][5] .power_up = "low";

dffeas \r_array_out[2][5] (
	.clk(clk),
	.d(\r_array_out[2][5]~15_combout ),
	.asdata(ram_in_reg_1_2),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_nm1_2),
	.ena(global_clock_enable),
	.q(r_array_out_5_2),
	.prn(vcc));
defparam \r_array_out[2][5] .is_wysiwyg = "true";
defparam \r_array_out[2][5] .power_up = "low";

dffeas \r_array_out[0][4] (
	.clk(clk),
	.d(\r_array_out[0][4]~12_combout ),
	.asdata(ram_in_reg_0_0),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_nm1_2),
	.ena(global_clock_enable),
	.q(r_array_out_4_0),
	.prn(vcc));
defparam \r_array_out[0][4] .is_wysiwyg = "true";
defparam \r_array_out[0][4] .power_up = "low";

dffeas \r_array_out[2][4] (
	.clk(clk),
	.d(\r_array_out[2][4]~13_combout ),
	.asdata(ram_in_reg_0_2),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_nm1_2),
	.ena(global_clock_enable),
	.q(r_array_out_4_2),
	.prn(vcc));
defparam \r_array_out[2][4] .is_wysiwyg = "true";
defparam \r_array_out[2][4] .power_up = "low";

dffeas \r_array_out[0][3] (
	.clk(clk),
	.d(\r_array_out[0][3]~10_combout ),
	.asdata(\Mux0~1_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_nm1_2),
	.sload(slb_nm1_1),
	.ena(global_clock_enable),
	.q(r_array_out_3_0),
	.prn(vcc));
defparam \r_array_out[0][3] .is_wysiwyg = "true";
defparam \r_array_out[0][3] .power_up = "low";

dffeas \r_array_out[2][3] (
	.clk(clk),
	.d(\r_array_out[2][3]~11_combout ),
	.asdata(\Mux16~1_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_nm1_2),
	.sload(slb_nm1_1),
	.ena(global_clock_enable),
	.q(r_array_out_3_2),
	.prn(vcc));
defparam \r_array_out[2][3] .is_wysiwyg = "true";
defparam \r_array_out[2][3] .power_up = "low";

dffeas \r_array_out[0][2] (
	.clk(clk),
	.d(\r_array_out[0][2]~8_combout ),
	.asdata(\Mux0~3_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_nm1_2),
	.sload(!slb_nm1_1),
	.ena(global_clock_enable),
	.q(r_array_out_2_0),
	.prn(vcc));
defparam \r_array_out[0][2] .is_wysiwyg = "true";
defparam \r_array_out[0][2] .power_up = "low";

dffeas \r_array_out[2][2] (
	.clk(clk),
	.d(\r_array_out[2][2]~9_combout ),
	.asdata(\Mux16~3_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_nm1_2),
	.sload(!slb_nm1_1),
	.ena(global_clock_enable),
	.q(r_array_out_2_2),
	.prn(vcc));
defparam \r_array_out[2][2] .is_wysiwyg = "true";
defparam \r_array_out[2][2] .power_up = "low";

dffeas \r_array_out[1][5] (
	.clk(clk),
	.d(\r_array_out[1][5]~6_combout ),
	.asdata(ram_in_reg_1_1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_nm1_2),
	.ena(global_clock_enable),
	.q(r_array_out_5_1),
	.prn(vcc));
defparam \r_array_out[1][5] .is_wysiwyg = "true";
defparam \r_array_out[1][5] .power_up = "low";

dffeas \r_array_out[3][5] (
	.clk(clk),
	.d(\r_array_out[3][5]~7_combout ),
	.asdata(ram_in_reg_1_3),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_nm1_2),
	.ena(global_clock_enable),
	.q(r_array_out_5_3),
	.prn(vcc));
defparam \r_array_out[3][5] .is_wysiwyg = "true";
defparam \r_array_out[3][5] .power_up = "low";

dffeas \r_array_out[1][4] (
	.clk(clk),
	.d(\r_array_out[1][4]~4_combout ),
	.asdata(ram_in_reg_0_1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_nm1_2),
	.ena(global_clock_enable),
	.q(r_array_out_4_1),
	.prn(vcc));
defparam \r_array_out[1][4] .is_wysiwyg = "true";
defparam \r_array_out[1][4] .power_up = "low";

dffeas \r_array_out[3][4] (
	.clk(clk),
	.d(\r_array_out[3][4]~5_combout ),
	.asdata(ram_in_reg_0_3),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_nm1_2),
	.ena(global_clock_enable),
	.q(r_array_out_4_3),
	.prn(vcc));
defparam \r_array_out[3][4] .is_wysiwyg = "true";
defparam \r_array_out[3][4] .power_up = "low";

dffeas \r_array_out[1][3] (
	.clk(clk),
	.d(\r_array_out[1][3]~2_combout ),
	.asdata(\Mux8~1_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_nm1_2),
	.sload(slb_nm1_1),
	.ena(global_clock_enable),
	.q(r_array_out_3_1),
	.prn(vcc));
defparam \r_array_out[1][3] .is_wysiwyg = "true";
defparam \r_array_out[1][3] .power_up = "low";

dffeas \r_array_out[3][3] (
	.clk(clk),
	.d(\r_array_out[3][3]~3_combout ),
	.asdata(\Mux24~1_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_nm1_2),
	.sload(slb_nm1_1),
	.ena(global_clock_enable),
	.q(r_array_out_3_3),
	.prn(vcc));
defparam \r_array_out[3][3] .is_wysiwyg = "true";
defparam \r_array_out[3][3] .power_up = "low";

dffeas \r_array_out[1][2] (
	.clk(clk),
	.d(\r_array_out[1][2]~0_combout ),
	.asdata(\Mux8~3_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_nm1_2),
	.sload(!slb_nm1_1),
	.ena(global_clock_enable),
	.q(r_array_out_2_1),
	.prn(vcc));
defparam \r_array_out[1][2] .is_wysiwyg = "true";
defparam \r_array_out[1][2] .power_up = "low";

dffeas \r_array_out[3][2] (
	.clk(clk),
	.d(\r_array_out[3][2]~1_combout ),
	.asdata(\Mux24~3_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_nm1_2),
	.sload(!slb_nm1_1),
	.ena(global_clock_enable),
	.q(r_array_out_2_3),
	.prn(vcc));
defparam \r_array_out[3][2] .is_wysiwyg = "true";
defparam \r_array_out[3][2] .power_up = "low";

dffeas \i_array_out[0][5] (
	.clk(clk),
	.d(\i_array_out[0][5]~6_combout ),
	.asdata(ram_in_reg_1_4),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_nm1_2),
	.ena(global_clock_enable),
	.q(i_array_out_5_0),
	.prn(vcc));
defparam \i_array_out[0][5] .is_wysiwyg = "true";
defparam \i_array_out[0][5] .power_up = "low";

dffeas \i_array_out[2][5] (
	.clk(clk),
	.d(\i_array_out[2][5]~7_combout ),
	.asdata(ram_in_reg_1_6),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_nm1_2),
	.ena(global_clock_enable),
	.q(i_array_out_5_2),
	.prn(vcc));
defparam \i_array_out[2][5] .is_wysiwyg = "true";
defparam \i_array_out[2][5] .power_up = "low";

dffeas \i_array_out[0][4] (
	.clk(clk),
	.d(\i_array_out[0][4]~4_combout ),
	.asdata(ram_in_reg_0_4),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_nm1_2),
	.ena(global_clock_enable),
	.q(i_array_out_4_0),
	.prn(vcc));
defparam \i_array_out[0][4] .is_wysiwyg = "true";
defparam \i_array_out[0][4] .power_up = "low";

dffeas \i_array_out[2][4] (
	.clk(clk),
	.d(\i_array_out[2][4]~5_combout ),
	.asdata(ram_in_reg_0_6),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_nm1_2),
	.ena(global_clock_enable),
	.q(i_array_out_4_2),
	.prn(vcc));
defparam \i_array_out[2][4] .is_wysiwyg = "true";
defparam \i_array_out[2][4] .power_up = "low";

dffeas \i_array_out[0][3] (
	.clk(clk),
	.d(\i_array_out[0][3]~2_combout ),
	.asdata(\Mux32~4_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_nm1_2),
	.sload(slb_nm1_1),
	.ena(global_clock_enable),
	.q(i_array_out_3_0),
	.prn(vcc));
defparam \i_array_out[0][3] .is_wysiwyg = "true";
defparam \i_array_out[0][3] .power_up = "low";

dffeas \i_array_out[2][3] (
	.clk(clk),
	.d(\i_array_out[2][3]~3_combout ),
	.asdata(\Mux48~4_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_nm1_2),
	.sload(slb_nm1_1),
	.ena(global_clock_enable),
	.q(i_array_out_3_2),
	.prn(vcc));
defparam \i_array_out[2][3] .is_wysiwyg = "true";
defparam \i_array_out[2][3] .power_up = "low";

dffeas \i_array_out[0][2] (
	.clk(clk),
	.d(\i_array_out[0][2]~0_combout ),
	.asdata(\Mux32~5_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_nm1_2),
	.sload(!slb_nm1_1),
	.ena(global_clock_enable),
	.q(i_array_out_2_0),
	.prn(vcc));
defparam \i_array_out[0][2] .is_wysiwyg = "true";
defparam \i_array_out[0][2] .power_up = "low";

dffeas \i_array_out[2][2] (
	.clk(clk),
	.d(\i_array_out[2][2]~1_combout ),
	.asdata(\Mux48~5_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_nm1_2),
	.sload(!slb_nm1_1),
	.ena(global_clock_enable),
	.q(i_array_out_2_2),
	.prn(vcc));
defparam \i_array_out[2][2] .is_wysiwyg = "true";
defparam \i_array_out[2][2] .power_up = "low";

dffeas \i_array_out[1][5] (
	.clk(clk),
	.d(\i_array_out[1][5]~14_combout ),
	.asdata(ram_in_reg_1_5),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_nm1_2),
	.ena(global_clock_enable),
	.q(i_array_out_5_1),
	.prn(vcc));
defparam \i_array_out[1][5] .is_wysiwyg = "true";
defparam \i_array_out[1][5] .power_up = "low";

dffeas \i_array_out[3][5] (
	.clk(clk),
	.d(\i_array_out[3][5]~15_combout ),
	.asdata(ram_in_reg_1_7),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_nm1_2),
	.ena(global_clock_enable),
	.q(i_array_out_5_3),
	.prn(vcc));
defparam \i_array_out[3][5] .is_wysiwyg = "true";
defparam \i_array_out[3][5] .power_up = "low";

dffeas \i_array_out[1][4] (
	.clk(clk),
	.d(\i_array_out[1][4]~12_combout ),
	.asdata(ram_in_reg_0_5),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_nm1_2),
	.ena(global_clock_enable),
	.q(i_array_out_4_1),
	.prn(vcc));
defparam \i_array_out[1][4] .is_wysiwyg = "true";
defparam \i_array_out[1][4] .power_up = "low";

dffeas \i_array_out[3][4] (
	.clk(clk),
	.d(\i_array_out[3][4]~13_combout ),
	.asdata(ram_in_reg_0_7),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_nm1_2),
	.ena(global_clock_enable),
	.q(i_array_out_4_3),
	.prn(vcc));
defparam \i_array_out[3][4] .is_wysiwyg = "true";
defparam \i_array_out[3][4] .power_up = "low";

dffeas \i_array_out[1][3] (
	.clk(clk),
	.d(\i_array_out[1][3]~10_combout ),
	.asdata(\Mux40~4_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_nm1_2),
	.sload(slb_nm1_1),
	.ena(global_clock_enable),
	.q(i_array_out_3_1),
	.prn(vcc));
defparam \i_array_out[1][3] .is_wysiwyg = "true";
defparam \i_array_out[1][3] .power_up = "low";

dffeas \i_array_out[3][3] (
	.clk(clk),
	.d(\i_array_out[3][3]~11_combout ),
	.asdata(\Mux56~4_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_nm1_2),
	.sload(slb_nm1_1),
	.ena(global_clock_enable),
	.q(i_array_out_3_3),
	.prn(vcc));
defparam \i_array_out[3][3] .is_wysiwyg = "true";
defparam \i_array_out[3][3] .power_up = "low";

dffeas \i_array_out[1][2] (
	.clk(clk),
	.d(\i_array_out[1][2]~8_combout ),
	.asdata(\Mux40~5_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_nm1_2),
	.sload(!slb_nm1_1),
	.ena(global_clock_enable),
	.q(i_array_out_2_1),
	.prn(vcc));
defparam \i_array_out[1][2] .is_wysiwyg = "true";
defparam \i_array_out[1][2] .power_up = "low";

dffeas \i_array_out[3][2] (
	.clk(clk),
	.d(\i_array_out[3][2]~9_combout ),
	.asdata(\Mux56~5_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_nm1_2),
	.sload(!slb_nm1_1),
	.ena(global_clock_enable),
	.q(i_array_out_2_3),
	.prn(vcc));
defparam \i_array_out[3][2] .is_wysiwyg = "true";
defparam \i_array_out[3][2] .power_up = "low";

dffeas \r_array_out[0][6] (
	.clk(clk),
	.d(\Mux1~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_6_0),
	.prn(vcc));
defparam \r_array_out[0][6] .is_wysiwyg = "true";
defparam \r_array_out[0][6] .power_up = "low";

dffeas \r_array_out[2][6] (
	.clk(clk),
	.d(\Mux17~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_6_2),
	.prn(vcc));
defparam \r_array_out[2][6] .is_wysiwyg = "true";
defparam \r_array_out[2][6] .power_up = "low";

dffeas \r_array_out[0][1] (
	.clk(clk),
	.d(\Mux6~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_1_0),
	.prn(vcc));
defparam \r_array_out[0][1] .is_wysiwyg = "true";
defparam \r_array_out[0][1] .power_up = "low";

dffeas \r_array_out[2][1] (
	.clk(clk),
	.d(\Mux22~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_1_2),
	.prn(vcc));
defparam \r_array_out[2][1] .is_wysiwyg = "true";
defparam \r_array_out[2][1] .power_up = "low";

dffeas \r_array_out[0][0] (
	.clk(clk),
	.d(\Mux7~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_0_0),
	.prn(vcc));
defparam \r_array_out[0][0] .is_wysiwyg = "true";
defparam \r_array_out[0][0] .power_up = "low";

dffeas \r_array_out[2][0] (
	.clk(clk),
	.d(\Mux23~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_0_2),
	.prn(vcc));
defparam \r_array_out[2][0] .is_wysiwyg = "true";
defparam \r_array_out[2][0] .power_up = "low";

dffeas \r_array_out[1][6] (
	.clk(clk),
	.d(\Mux9~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_6_1),
	.prn(vcc));
defparam \r_array_out[1][6] .is_wysiwyg = "true";
defparam \r_array_out[1][6] .power_up = "low";

dffeas \r_array_out[3][6] (
	.clk(clk),
	.d(\Mux25~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_6_3),
	.prn(vcc));
defparam \r_array_out[3][6] .is_wysiwyg = "true";
defparam \r_array_out[3][6] .power_up = "low";

dffeas \r_array_out[1][1] (
	.clk(clk),
	.d(\Mux14~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_1_1),
	.prn(vcc));
defparam \r_array_out[1][1] .is_wysiwyg = "true";
defparam \r_array_out[1][1] .power_up = "low";

dffeas \r_array_out[3][1] (
	.clk(clk),
	.d(\Mux30~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_1_3),
	.prn(vcc));
defparam \r_array_out[3][1] .is_wysiwyg = "true";
defparam \r_array_out[3][1] .power_up = "low";

dffeas \r_array_out[1][0] (
	.clk(clk),
	.d(\Mux15~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_0_1),
	.prn(vcc));
defparam \r_array_out[1][0] .is_wysiwyg = "true";
defparam \r_array_out[1][0] .power_up = "low";

dffeas \r_array_out[3][0] (
	.clk(clk),
	.d(\Mux31~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_0_3),
	.prn(vcc));
defparam \r_array_out[3][0] .is_wysiwyg = "true";
defparam \r_array_out[3][0] .power_up = "low";

dffeas \r_array_out[0][7] (
	.clk(clk),
	.d(\Mux0~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_7_0),
	.prn(vcc));
defparam \r_array_out[0][7] .is_wysiwyg = "true";
defparam \r_array_out[0][7] .power_up = "low";

dffeas \r_array_out[2][7] (
	.clk(clk),
	.d(\Mux16~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_7_2),
	.prn(vcc));
defparam \r_array_out[2][7] .is_wysiwyg = "true";
defparam \r_array_out[2][7] .power_up = "low";

dffeas \r_array_out[1][7] (
	.clk(clk),
	.d(\Mux8~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_7_1),
	.prn(vcc));
defparam \r_array_out[1][7] .is_wysiwyg = "true";
defparam \r_array_out[1][7] .power_up = "low";

dffeas \r_array_out[3][7] (
	.clk(clk),
	.d(\Mux24~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_7_3),
	.prn(vcc));
defparam \r_array_out[3][7] .is_wysiwyg = "true";
defparam \r_array_out[3][7] .power_up = "low";

dffeas \i_array_out[0][7] (
	.clk(clk),
	.d(\Mux32~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_7_0),
	.prn(vcc));
defparam \i_array_out[0][7] .is_wysiwyg = "true";
defparam \i_array_out[0][7] .power_up = "low";

dffeas \i_array_out[2][7] (
	.clk(clk),
	.d(\Mux48~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_7_2),
	.prn(vcc));
defparam \i_array_out[2][7] .is_wysiwyg = "true";
defparam \i_array_out[2][7] .power_up = "low";

dffeas \i_array_out[0][6] (
	.clk(clk),
	.d(\Mux33~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_6_0),
	.prn(vcc));
defparam \i_array_out[0][6] .is_wysiwyg = "true";
defparam \i_array_out[0][6] .power_up = "low";

dffeas \i_array_out[2][6] (
	.clk(clk),
	.d(\Mux49~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_6_2),
	.prn(vcc));
defparam \i_array_out[2][6] .is_wysiwyg = "true";
defparam \i_array_out[2][6] .power_up = "low";

dffeas \i_array_out[0][1] (
	.clk(clk),
	.d(\Mux38~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_1_0),
	.prn(vcc));
defparam \i_array_out[0][1] .is_wysiwyg = "true";
defparam \i_array_out[0][1] .power_up = "low";

dffeas \i_array_out[2][1] (
	.clk(clk),
	.d(\Mux54~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_1_2),
	.prn(vcc));
defparam \i_array_out[2][1] .is_wysiwyg = "true";
defparam \i_array_out[2][1] .power_up = "low";

dffeas \i_array_out[0][0] (
	.clk(clk),
	.d(\Mux39~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_0_0),
	.prn(vcc));
defparam \i_array_out[0][0] .is_wysiwyg = "true";
defparam \i_array_out[0][0] .power_up = "low";

dffeas \i_array_out[2][0] (
	.clk(clk),
	.d(\Mux55~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_0_2),
	.prn(vcc));
defparam \i_array_out[2][0] .is_wysiwyg = "true";
defparam \i_array_out[2][0] .power_up = "low";

dffeas \i_array_out[1][7] (
	.clk(clk),
	.d(\Mux40~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_7_1),
	.prn(vcc));
defparam \i_array_out[1][7] .is_wysiwyg = "true";
defparam \i_array_out[1][7] .power_up = "low";

dffeas \i_array_out[3][7] (
	.clk(clk),
	.d(\Mux56~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_7_3),
	.prn(vcc));
defparam \i_array_out[3][7] .is_wysiwyg = "true";
defparam \i_array_out[3][7] .power_up = "low";

dffeas \i_array_out[1][6] (
	.clk(clk),
	.d(\Mux41~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_6_1),
	.prn(vcc));
defparam \i_array_out[1][6] .is_wysiwyg = "true";
defparam \i_array_out[1][6] .power_up = "low";

dffeas \i_array_out[3][6] (
	.clk(clk),
	.d(\Mux57~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_6_3),
	.prn(vcc));
defparam \i_array_out[3][6] .is_wysiwyg = "true";
defparam \i_array_out[3][6] .power_up = "low";

dffeas \i_array_out[1][1] (
	.clk(clk),
	.d(\Mux46~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_1_1),
	.prn(vcc));
defparam \i_array_out[1][1] .is_wysiwyg = "true";
defparam \i_array_out[1][1] .power_up = "low";

dffeas \i_array_out[3][1] (
	.clk(clk),
	.d(\Mux62~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_1_3),
	.prn(vcc));
defparam \i_array_out[3][1] .is_wysiwyg = "true";
defparam \i_array_out[3][1] .power_up = "low";

dffeas \i_array_out[1][0] (
	.clk(clk),
	.d(\Mux47~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_0_1),
	.prn(vcc));
defparam \i_array_out[1][0] .is_wysiwyg = "true";
defparam \i_array_out[1][0] .power_up = "low";

dffeas \i_array_out[3][0] (
	.clk(clk),
	.d(\Mux63~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_0_3),
	.prn(vcc));
defparam \i_array_out[3][0] .is_wysiwyg = "true";
defparam \i_array_out[3][0] .power_up = "low";

cycloneiii_lcell_comb \Mux0~1 (
	.dataa(ram_in_reg_3_0),
	.datab(ram_in_reg_2_0),
	.datac(slb_last_0),
	.datad(block_dft_i_en),
	.cin(gnd),
	.combout(\Mux0~1_combout ),
	.cout());
defparam \Mux0~1 .lut_mask = 16'hEFFE;
defparam \Mux0~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux0~2 (
	.dataa(ram_in_reg_5_0),
	.datab(ram_in_reg_4_0),
	.datac(slb_last_0),
	.datad(block_dft_i_en),
	.cin(gnd),
	.combout(\Mux0~2_combout ),
	.cout());
defparam \Mux0~2 .lut_mask = 16'hEFFE;
defparam \Mux0~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \r_array_out[0][5]~14 (
	.dataa(\Mux0~1_combout ),
	.datab(\Mux0~2_combout ),
	.datac(gnd),
	.datad(slb_nm1_1),
	.cin(gnd),
	.combout(\r_array_out[0][5]~14_combout ),
	.cout());
defparam \r_array_out[0][5]~14 .lut_mask = 16'hAACC;
defparam \r_array_out[0][5]~14 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux16~1 (
	.dataa(ram_in_reg_3_2),
	.datab(ram_in_reg_2_2),
	.datac(slb_last_0),
	.datad(block_dft_i_en),
	.cin(gnd),
	.combout(\Mux16~1_combout ),
	.cout());
defparam \Mux16~1 .lut_mask = 16'hEFFE;
defparam \Mux16~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux16~2 (
	.dataa(ram_in_reg_5_2),
	.datab(ram_in_reg_4_2),
	.datac(slb_last_0),
	.datad(block_dft_i_en),
	.cin(gnd),
	.combout(\Mux16~2_combout ),
	.cout());
defparam \Mux16~2 .lut_mask = 16'hEFFE;
defparam \Mux16~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \r_array_out[2][5]~15 (
	.dataa(\Mux16~1_combout ),
	.datab(\Mux16~2_combout ),
	.datac(gnd),
	.datad(slb_nm1_1),
	.cin(gnd),
	.combout(\r_array_out[2][5]~15_combout ),
	.cout());
defparam \r_array_out[2][5]~15 .lut_mask = 16'hAACC;
defparam \r_array_out[2][5]~15 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \r_array_out[0][2]~8 (
	.dataa(ram_in_reg_2_0),
	.datab(ram_in_reg_1_0),
	.datac(gnd),
	.datad(slb_nm1_0),
	.cin(gnd),
	.combout(\r_array_out[0][2]~8_combout ),
	.cout());
defparam \r_array_out[0][2]~8 .lut_mask = 16'hAACC;
defparam \r_array_out[0][2]~8 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux0~0 (
	.dataa(ram_in_reg_4_0),
	.datab(ram_in_reg_3_0),
	.datac(slb_last_0),
	.datad(block_dft_i_en),
	.cin(gnd),
	.combout(\Mux0~0_combout ),
	.cout());
defparam \Mux0~0 .lut_mask = 16'hEFFE;
defparam \Mux0~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \r_array_out[0][4]~12 (
	.dataa(\r_array_out[0][2]~8_combout ),
	.datab(\Mux0~0_combout ),
	.datac(gnd),
	.datad(slb_nm1_1),
	.cin(gnd),
	.combout(\r_array_out[0][4]~12_combout ),
	.cout());
defparam \r_array_out[0][4]~12 .lut_mask = 16'hAACC;
defparam \r_array_out[0][4]~12 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \r_array_out[2][2]~9 (
	.dataa(ram_in_reg_2_2),
	.datab(ram_in_reg_1_2),
	.datac(slb_last_0),
	.datad(block_dft_i_en),
	.cin(gnd),
	.combout(\r_array_out[2][2]~9_combout ),
	.cout());
defparam \r_array_out[2][2]~9 .lut_mask = 16'hEFFE;
defparam \r_array_out[2][2]~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux16~0 (
	.dataa(ram_in_reg_4_2),
	.datab(ram_in_reg_3_2),
	.datac(slb_last_0),
	.datad(block_dft_i_en),
	.cin(gnd),
	.combout(\Mux16~0_combout ),
	.cout());
defparam \Mux16~0 .lut_mask = 16'hEFFE;
defparam \Mux16~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \r_array_out[2][4]~13 (
	.dataa(\r_array_out[2][2]~9_combout ),
	.datab(\Mux16~0_combout ),
	.datac(gnd),
	.datad(slb_nm1_1),
	.cin(gnd),
	.combout(\r_array_out[2][4]~13_combout ),
	.cout());
defparam \r_array_out[2][4]~13 .lut_mask = 16'hAACC;
defparam \r_array_out[2][4]~13 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \r_array_out[0][3]~10 (
	.dataa(ram_in_reg_1_0),
	.datab(ram_in_reg_0_0),
	.datac(gnd),
	.datad(slb_nm1_0),
	.cin(gnd),
	.combout(\r_array_out[0][3]~10_combout ),
	.cout());
defparam \r_array_out[0][3]~10 .lut_mask = 16'hAACC;
defparam \r_array_out[0][3]~10 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \r_array_out[2][3]~11 (
	.dataa(ram_in_reg_1_2),
	.datab(ram_in_reg_0_2),
	.datac(gnd),
	.datad(slb_nm1_0),
	.cin(gnd),
	.combout(\r_array_out[2][3]~11_combout ),
	.cout());
defparam \r_array_out[2][3]~11 .lut_mask = 16'hAACC;
defparam \r_array_out[2][3]~11 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux0~3 (
	.dataa(ram_in_reg_0_0),
	.datab(block_dft_i_en),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux0~3_combout ),
	.cout());
defparam \Mux0~3 .lut_mask = 16'hEEFF;
defparam \Mux0~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux16~3 (
	.dataa(ram_in_reg_0_2),
	.datab(block_dft_i_en),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux16~3_combout ),
	.cout());
defparam \Mux16~3 .lut_mask = 16'hEEFF;
defparam \Mux16~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux8~1 (
	.dataa(ram_in_reg_3_1),
	.datab(ram_in_reg_2_1),
	.datac(slb_last_0),
	.datad(block_dft_i_en),
	.cin(gnd),
	.combout(\Mux8~1_combout ),
	.cout());
defparam \Mux8~1 .lut_mask = 16'hEFFE;
defparam \Mux8~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux8~2 (
	.dataa(ram_in_reg_5_1),
	.datab(ram_in_reg_4_1),
	.datac(slb_last_0),
	.datad(block_dft_i_en),
	.cin(gnd),
	.combout(\Mux8~2_combout ),
	.cout());
defparam \Mux8~2 .lut_mask = 16'hEFFE;
defparam \Mux8~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \r_array_out[1][5]~6 (
	.dataa(\Mux8~1_combout ),
	.datab(\Mux8~2_combout ),
	.datac(gnd),
	.datad(slb_nm1_1),
	.cin(gnd),
	.combout(\r_array_out[1][5]~6_combout ),
	.cout());
defparam \r_array_out[1][5]~6 .lut_mask = 16'hAACC;
defparam \r_array_out[1][5]~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux24~1 (
	.dataa(ram_in_reg_3_3),
	.datab(ram_in_reg_2_3),
	.datac(slb_last_0),
	.datad(block_dft_i_en),
	.cin(gnd),
	.combout(\Mux24~1_combout ),
	.cout());
defparam \Mux24~1 .lut_mask = 16'hEFFE;
defparam \Mux24~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux24~2 (
	.dataa(ram_in_reg_5_3),
	.datab(ram_in_reg_4_3),
	.datac(slb_last_0),
	.datad(block_dft_i_en),
	.cin(gnd),
	.combout(\Mux24~2_combout ),
	.cout());
defparam \Mux24~2 .lut_mask = 16'hEFFE;
defparam \Mux24~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \r_array_out[3][5]~7 (
	.dataa(\Mux24~1_combout ),
	.datab(\Mux24~2_combout ),
	.datac(gnd),
	.datad(slb_nm1_1),
	.cin(gnd),
	.combout(\r_array_out[3][5]~7_combout ),
	.cout());
defparam \r_array_out[3][5]~7 .lut_mask = 16'hAACC;
defparam \r_array_out[3][5]~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \r_array_out[1][2]~0 (
	.dataa(ram_in_reg_2_1),
	.datab(ram_in_reg_1_1),
	.datac(slb_last_0),
	.datad(block_dft_i_en),
	.cin(gnd),
	.combout(\r_array_out[1][2]~0_combout ),
	.cout());
defparam \r_array_out[1][2]~0 .lut_mask = 16'hEFFE;
defparam \r_array_out[1][2]~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux8~0 (
	.dataa(ram_in_reg_4_1),
	.datab(ram_in_reg_3_1),
	.datac(slb_last_0),
	.datad(block_dft_i_en),
	.cin(gnd),
	.combout(\Mux8~0_combout ),
	.cout());
defparam \Mux8~0 .lut_mask = 16'hEFFE;
defparam \Mux8~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \r_array_out[1][4]~4 (
	.dataa(\r_array_out[1][2]~0_combout ),
	.datab(\Mux8~0_combout ),
	.datac(gnd),
	.datad(slb_nm1_1),
	.cin(gnd),
	.combout(\r_array_out[1][4]~4_combout ),
	.cout());
defparam \r_array_out[1][4]~4 .lut_mask = 16'hAACC;
defparam \r_array_out[1][4]~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \r_array_out[3][2]~1 (
	.dataa(ram_in_reg_2_3),
	.datab(ram_in_reg_1_3),
	.datac(slb_last_0),
	.datad(block_dft_i_en),
	.cin(gnd),
	.combout(\r_array_out[3][2]~1_combout ),
	.cout());
defparam \r_array_out[3][2]~1 .lut_mask = 16'hEFFE;
defparam \r_array_out[3][2]~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux24~0 (
	.dataa(ram_in_reg_4_3),
	.datab(ram_in_reg_3_3),
	.datac(slb_last_0),
	.datad(block_dft_i_en),
	.cin(gnd),
	.combout(\Mux24~0_combout ),
	.cout());
defparam \Mux24~0 .lut_mask = 16'hEFFE;
defparam \Mux24~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \r_array_out[3][4]~5 (
	.dataa(\r_array_out[3][2]~1_combout ),
	.datab(\Mux24~0_combout ),
	.datac(gnd),
	.datad(slb_nm1_1),
	.cin(gnd),
	.combout(\r_array_out[3][4]~5_combout ),
	.cout());
defparam \r_array_out[3][4]~5 .lut_mask = 16'hAACC;
defparam \r_array_out[3][4]~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \r_array_out[1][3]~2 (
	.dataa(ram_in_reg_1_1),
	.datab(ram_in_reg_0_1),
	.datac(gnd),
	.datad(slb_nm1_0),
	.cin(gnd),
	.combout(\r_array_out[1][3]~2_combout ),
	.cout());
defparam \r_array_out[1][3]~2 .lut_mask = 16'hAACC;
defparam \r_array_out[1][3]~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \r_array_out[3][3]~3 (
	.dataa(ram_in_reg_1_3),
	.datab(ram_in_reg_0_3),
	.datac(gnd),
	.datad(slb_nm1_0),
	.cin(gnd),
	.combout(\r_array_out[3][3]~3_combout ),
	.cout());
defparam \r_array_out[3][3]~3 .lut_mask = 16'hAACC;
defparam \r_array_out[3][3]~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux8~3 (
	.dataa(ram_in_reg_0_1),
	.datab(block_dft_i_en),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux8~3_combout ),
	.cout());
defparam \Mux8~3 .lut_mask = 16'hEEFF;
defparam \Mux8~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux24~3 (
	.dataa(ram_in_reg_0_3),
	.datab(block_dft_i_en),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux24~3_combout ),
	.cout());
defparam \Mux24~3 .lut_mask = 16'hEEFF;
defparam \Mux24~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux32~4 (
	.dataa(ram_in_reg_3_4),
	.datab(ram_in_reg_2_4),
	.datac(slb_last_0),
	.datad(block_dft_i_en),
	.cin(gnd),
	.combout(\Mux32~4_combout ),
	.cout());
defparam \Mux32~4 .lut_mask = 16'hEFFE;
defparam \Mux32~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux32~0 (
	.dataa(ram_in_reg_5_4),
	.datab(ram_in_reg_4_4),
	.datac(slb_last_0),
	.datad(block_dft_i_en),
	.cin(gnd),
	.combout(\Mux32~0_combout ),
	.cout());
defparam \Mux32~0 .lut_mask = 16'hEFFE;
defparam \Mux32~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \i_array_out[0][5]~6 (
	.dataa(\Mux32~4_combout ),
	.datab(\Mux32~0_combout ),
	.datac(gnd),
	.datad(slb_nm1_1),
	.cin(gnd),
	.combout(\i_array_out[0][5]~6_combout ),
	.cout());
defparam \i_array_out[0][5]~6 .lut_mask = 16'hAACC;
defparam \i_array_out[0][5]~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux48~4 (
	.dataa(ram_in_reg_3_6),
	.datab(ram_in_reg_2_6),
	.datac(slb_last_0),
	.datad(block_dft_i_en),
	.cin(gnd),
	.combout(\Mux48~4_combout ),
	.cout());
defparam \Mux48~4 .lut_mask = 16'hEFFE;
defparam \Mux48~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux48~0 (
	.dataa(ram_in_reg_5_6),
	.datab(ram_in_reg_4_6),
	.datac(slb_last_0),
	.datad(block_dft_i_en),
	.cin(gnd),
	.combout(\Mux48~0_combout ),
	.cout());
defparam \Mux48~0 .lut_mask = 16'hEFFE;
defparam \Mux48~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \i_array_out[2][5]~7 (
	.dataa(\Mux48~4_combout ),
	.datab(\Mux48~0_combout ),
	.datac(gnd),
	.datad(slb_nm1_1),
	.cin(gnd),
	.combout(\i_array_out[2][5]~7_combout ),
	.cout());
defparam \i_array_out[2][5]~7 .lut_mask = 16'hAACC;
defparam \i_array_out[2][5]~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \i_array_out[0][2]~0 (
	.dataa(ram_in_reg_2_4),
	.datab(ram_in_reg_1_4),
	.datac(slb_last_0),
	.datad(block_dft_i_en),
	.cin(gnd),
	.combout(\i_array_out[0][2]~0_combout ),
	.cout());
defparam \i_array_out[0][2]~0 .lut_mask = 16'hEFFE;
defparam \i_array_out[0][2]~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux32~3 (
	.dataa(ram_in_reg_4_4),
	.datab(ram_in_reg_3_4),
	.datac(slb_last_0),
	.datad(block_dft_i_en),
	.cin(gnd),
	.combout(\Mux32~3_combout ),
	.cout());
defparam \Mux32~3 .lut_mask = 16'hEFFE;
defparam \Mux32~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \i_array_out[0][4]~4 (
	.dataa(\i_array_out[0][2]~0_combout ),
	.datab(\Mux32~3_combout ),
	.datac(gnd),
	.datad(slb_nm1_1),
	.cin(gnd),
	.combout(\i_array_out[0][4]~4_combout ),
	.cout());
defparam \i_array_out[0][4]~4 .lut_mask = 16'hAACC;
defparam \i_array_out[0][4]~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \i_array_out[2][2]~1 (
	.dataa(ram_in_reg_2_6),
	.datab(ram_in_reg_1_6),
	.datac(slb_last_0),
	.datad(block_dft_i_en),
	.cin(gnd),
	.combout(\i_array_out[2][2]~1_combout ),
	.cout());
defparam \i_array_out[2][2]~1 .lut_mask = 16'hEFFE;
defparam \i_array_out[2][2]~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux48~3 (
	.dataa(ram_in_reg_4_6),
	.datab(ram_in_reg_3_6),
	.datac(slb_last_0),
	.datad(block_dft_i_en),
	.cin(gnd),
	.combout(\Mux48~3_combout ),
	.cout());
defparam \Mux48~3 .lut_mask = 16'hEFFE;
defparam \Mux48~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \i_array_out[2][4]~5 (
	.dataa(\i_array_out[2][2]~1_combout ),
	.datab(\Mux48~3_combout ),
	.datac(gnd),
	.datad(slb_nm1_1),
	.cin(gnd),
	.combout(\i_array_out[2][4]~5_combout ),
	.cout());
defparam \i_array_out[2][4]~5 .lut_mask = 16'hAACC;
defparam \i_array_out[2][4]~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \i_array_out[0][3]~2 (
	.dataa(ram_in_reg_1_4),
	.datab(ram_in_reg_0_4),
	.datac(gnd),
	.datad(slb_nm1_0),
	.cin(gnd),
	.combout(\i_array_out[0][3]~2_combout ),
	.cout());
defparam \i_array_out[0][3]~2 .lut_mask = 16'hAACC;
defparam \i_array_out[0][3]~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \i_array_out[2][3]~3 (
	.dataa(ram_in_reg_1_6),
	.datab(ram_in_reg_0_6),
	.datac(gnd),
	.datad(slb_nm1_0),
	.cin(gnd),
	.combout(\i_array_out[2][3]~3_combout ),
	.cout());
defparam \i_array_out[2][3]~3 .lut_mask = 16'hAACC;
defparam \i_array_out[2][3]~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux32~5 (
	.dataa(ram_in_reg_0_4),
	.datab(block_dft_i_en),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux32~5_combout ),
	.cout());
defparam \Mux32~5 .lut_mask = 16'hEEFF;
defparam \Mux32~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux48~5 (
	.dataa(ram_in_reg_0_6),
	.datab(block_dft_i_en),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux48~5_combout ),
	.cout());
defparam \Mux48~5 .lut_mask = 16'hEEFF;
defparam \Mux48~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux40~4 (
	.dataa(ram_in_reg_3_5),
	.datab(ram_in_reg_2_5),
	.datac(slb_last_0),
	.datad(block_dft_i_en),
	.cin(gnd),
	.combout(\Mux40~4_combout ),
	.cout());
defparam \Mux40~4 .lut_mask = 16'hEFFE;
defparam \Mux40~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux40~0 (
	.dataa(ram_in_reg_5_5),
	.datab(ram_in_reg_4_5),
	.datac(slb_last_0),
	.datad(block_dft_i_en),
	.cin(gnd),
	.combout(\Mux40~0_combout ),
	.cout());
defparam \Mux40~0 .lut_mask = 16'hEFFE;
defparam \Mux40~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \i_array_out[1][5]~14 (
	.dataa(\Mux40~4_combout ),
	.datab(\Mux40~0_combout ),
	.datac(gnd),
	.datad(slb_nm1_1),
	.cin(gnd),
	.combout(\i_array_out[1][5]~14_combout ),
	.cout());
defparam \i_array_out[1][5]~14 .lut_mask = 16'hAACC;
defparam \i_array_out[1][5]~14 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux56~4 (
	.dataa(ram_in_reg_3_7),
	.datab(ram_in_reg_2_7),
	.datac(slb_last_0),
	.datad(block_dft_i_en),
	.cin(gnd),
	.combout(\Mux56~4_combout ),
	.cout());
defparam \Mux56~4 .lut_mask = 16'hEFFE;
defparam \Mux56~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux56~0 (
	.dataa(ram_in_reg_5_7),
	.datab(ram_in_reg_4_7),
	.datac(slb_last_0),
	.datad(block_dft_i_en),
	.cin(gnd),
	.combout(\Mux56~0_combout ),
	.cout());
defparam \Mux56~0 .lut_mask = 16'hEFFE;
defparam \Mux56~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \i_array_out[3][5]~15 (
	.dataa(\Mux56~4_combout ),
	.datab(\Mux56~0_combout ),
	.datac(gnd),
	.datad(slb_nm1_1),
	.cin(gnd),
	.combout(\i_array_out[3][5]~15_combout ),
	.cout());
defparam \i_array_out[3][5]~15 .lut_mask = 16'hAACC;
defparam \i_array_out[3][5]~15 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \i_array_out[1][2]~8 (
	.dataa(ram_in_reg_2_5),
	.datab(ram_in_reg_1_5),
	.datac(slb_last_0),
	.datad(block_dft_i_en),
	.cin(gnd),
	.combout(\i_array_out[1][2]~8_combout ),
	.cout());
defparam \i_array_out[1][2]~8 .lut_mask = 16'hEFFE;
defparam \i_array_out[1][2]~8 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux40~3 (
	.dataa(ram_in_reg_4_5),
	.datab(ram_in_reg_3_5),
	.datac(slb_last_0),
	.datad(block_dft_i_en),
	.cin(gnd),
	.combout(\Mux40~3_combout ),
	.cout());
defparam \Mux40~3 .lut_mask = 16'hEFFE;
defparam \Mux40~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \i_array_out[1][4]~12 (
	.dataa(\i_array_out[1][2]~8_combout ),
	.datab(\Mux40~3_combout ),
	.datac(gnd),
	.datad(slb_nm1_1),
	.cin(gnd),
	.combout(\i_array_out[1][4]~12_combout ),
	.cout());
defparam \i_array_out[1][4]~12 .lut_mask = 16'hAACC;
defparam \i_array_out[1][4]~12 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \i_array_out[3][2]~9 (
	.dataa(ram_in_reg_2_7),
	.datab(ram_in_reg_1_7),
	.datac(slb_last_0),
	.datad(block_dft_i_en),
	.cin(gnd),
	.combout(\i_array_out[3][2]~9_combout ),
	.cout());
defparam \i_array_out[3][2]~9 .lut_mask = 16'hEFFE;
defparam \i_array_out[3][2]~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux56~3 (
	.dataa(ram_in_reg_4_7),
	.datab(ram_in_reg_3_7),
	.datac(slb_last_0),
	.datad(block_dft_i_en),
	.cin(gnd),
	.combout(\Mux56~3_combout ),
	.cout());
defparam \Mux56~3 .lut_mask = 16'hEFFE;
defparam \Mux56~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \i_array_out[3][4]~13 (
	.dataa(\i_array_out[3][2]~9_combout ),
	.datab(\Mux56~3_combout ),
	.datac(gnd),
	.datad(slb_nm1_1),
	.cin(gnd),
	.combout(\i_array_out[3][4]~13_combout ),
	.cout());
defparam \i_array_out[3][4]~13 .lut_mask = 16'hAACC;
defparam \i_array_out[3][4]~13 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \i_array_out[1][3]~10 (
	.dataa(ram_in_reg_1_5),
	.datab(ram_in_reg_0_5),
	.datac(gnd),
	.datad(slb_nm1_0),
	.cin(gnd),
	.combout(\i_array_out[1][3]~10_combout ),
	.cout());
defparam \i_array_out[1][3]~10 .lut_mask = 16'hAACC;
defparam \i_array_out[1][3]~10 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \i_array_out[3][3]~11 (
	.dataa(ram_in_reg_1_7),
	.datab(ram_in_reg_0_7),
	.datac(gnd),
	.datad(slb_nm1_0),
	.cin(gnd),
	.combout(\i_array_out[3][3]~11_combout ),
	.cout());
defparam \i_array_out[3][3]~11 .lut_mask = 16'hAACC;
defparam \i_array_out[3][3]~11 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux40~5 (
	.dataa(ram_in_reg_0_5),
	.datab(block_dft_i_en),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux40~5_combout ),
	.cout());
defparam \Mux40~5 .lut_mask = 16'hEEFF;
defparam \Mux40~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux56~5 (
	.dataa(ram_in_reg_0_7),
	.datab(block_dft_i_en),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux56~5_combout ),
	.cout());
defparam \Mux56~5 .lut_mask = 16'hEEFF;
defparam \Mux56~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \r_array_out[2][6]~16 (
	.dataa(slb_last_2),
	.datab(slb_last_0),
	.datac(slb_last_1),
	.datad(block_dft_i_en),
	.cin(gnd),
	.combout(\r_array_out[2][6]~16_combout ),
	.cout());
defparam \r_array_out[2][6]~16 .lut_mask = 16'hEFFF;
defparam \r_array_out[2][6]~16 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \r_array_out[2][6]~17 (
	.dataa(slb_last_1),
	.datab(slb_last_2),
	.datac(gnd),
	.datad(block_dft_i_en),
	.cin(gnd),
	.combout(\r_array_out[2][6]~17_combout ),
	.cout());
defparam \r_array_out[2][6]~17 .lut_mask = 16'hEEFF;
defparam \r_array_out[2][6]~17 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux1~0 (
	.dataa(\r_array_out[2][6]~16_combout ),
	.datab(ram_in_reg_6_0),
	.datac(\r_array_out[2][6]~17_combout ),
	.datad(\Mux0~0_combout ),
	.cin(gnd),
	.combout(\Mux1~0_combout ),
	.cout());
defparam \Mux1~0 .lut_mask = 16'hFFDE;
defparam \Mux1~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux1~1 (
	.dataa(ram_in_reg_2_0),
	.datab(\r_array_out[2][6]~16_combout ),
	.datac(\Mux1~0_combout ),
	.datad(ram_in_reg_5_0),
	.cin(gnd),
	.combout(\Mux1~1_combout ),
	.cout());
defparam \Mux1~1 .lut_mask = 16'hFFBE;
defparam \Mux1~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux17~0 (
	.dataa(\r_array_out[2][6]~16_combout ),
	.datab(ram_in_reg_6_2),
	.datac(\r_array_out[2][6]~17_combout ),
	.datad(\Mux16~0_combout ),
	.cin(gnd),
	.combout(\Mux17~0_combout ),
	.cout());
defparam \Mux17~0 .lut_mask = 16'hFFDE;
defparam \Mux17~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux17~1 (
	.dataa(ram_in_reg_2_2),
	.datab(\r_array_out[2][6]~16_combout ),
	.datac(\Mux17~0_combout ),
	.datad(ram_in_reg_5_2),
	.cin(gnd),
	.combout(\Mux17~1_combout ),
	.cout());
defparam \Mux17~1 .lut_mask = 16'hFFBE;
defparam \Mux17~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux6~2 (
	.dataa(slb_last_1),
	.datab(slb_last_2),
	.datac(block_dft_i_en),
	.datad(\r_array_out[0][3]~10_combout ),
	.cin(gnd),
	.combout(\Mux6~2_combout ),
	.cout());
defparam \Mux6~2 .lut_mask = 16'hFFF7;
defparam \Mux6~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux22~2 (
	.dataa(slb_last_1),
	.datab(slb_last_2),
	.datac(block_dft_i_en),
	.datad(\r_array_out[2][3]~11_combout ),
	.cin(gnd),
	.combout(\Mux22~2_combout ),
	.cout());
defparam \Mux22~2 .lut_mask = 16'hFFF7;
defparam \Mux22~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux7~0 (
	.dataa(slb_last_0),
	.datab(slb_last_1),
	.datac(slb_last_2),
	.datad(block_dft_i_en),
	.cin(gnd),
	.combout(\Mux7~0_combout ),
	.cout());
defparam \Mux7~0 .lut_mask = 16'hFEFF;
defparam \Mux7~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux7~1 (
	.dataa(ram_in_reg_0_0),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mux7~0_combout ),
	.cin(gnd),
	.combout(\Mux7~1_combout ),
	.cout());
defparam \Mux7~1 .lut_mask = 16'hAAFF;
defparam \Mux7~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux23~0 (
	.dataa(ram_in_reg_0_2),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mux7~0_combout ),
	.cin(gnd),
	.combout(\Mux23~0_combout ),
	.cout());
defparam \Mux23~0 .lut_mask = 16'hAAFF;
defparam \Mux23~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux9~0 (
	.dataa(\r_array_out[2][6]~16_combout ),
	.datab(ram_in_reg_6_1),
	.datac(\r_array_out[2][6]~17_combout ),
	.datad(\Mux8~0_combout ),
	.cin(gnd),
	.combout(\Mux9~0_combout ),
	.cout());
defparam \Mux9~0 .lut_mask = 16'hFFDE;
defparam \Mux9~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux9~1 (
	.dataa(ram_in_reg_2_1),
	.datab(\r_array_out[2][6]~16_combout ),
	.datac(\Mux9~0_combout ),
	.datad(ram_in_reg_5_1),
	.cin(gnd),
	.combout(\Mux9~1_combout ),
	.cout());
defparam \Mux9~1 .lut_mask = 16'hFFBE;
defparam \Mux9~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux25~0 (
	.dataa(\r_array_out[2][6]~16_combout ),
	.datab(ram_in_reg_6_3),
	.datac(\r_array_out[2][6]~17_combout ),
	.datad(\Mux24~0_combout ),
	.cin(gnd),
	.combout(\Mux25~0_combout ),
	.cout());
defparam \Mux25~0 .lut_mask = 16'hFFDE;
defparam \Mux25~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux25~1 (
	.dataa(ram_in_reg_2_3),
	.datab(\r_array_out[2][6]~16_combout ),
	.datac(\Mux25~0_combout ),
	.datad(ram_in_reg_5_3),
	.cin(gnd),
	.combout(\Mux25~1_combout ),
	.cout());
defparam \Mux25~1 .lut_mask = 16'hFFBE;
defparam \Mux25~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux14~2 (
	.dataa(slb_last_1),
	.datab(slb_last_2),
	.datac(block_dft_i_en),
	.datad(\r_array_out[1][3]~2_combout ),
	.cin(gnd),
	.combout(\Mux14~2_combout ),
	.cout());
defparam \Mux14~2 .lut_mask = 16'hFFF7;
defparam \Mux14~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux30~2 (
	.dataa(slb_last_1),
	.datab(slb_last_2),
	.datac(block_dft_i_en),
	.datad(\r_array_out[3][3]~3_combout ),
	.cin(gnd),
	.combout(\Mux30~2_combout ),
	.cout());
defparam \Mux30~2 .lut_mask = 16'hFFF7;
defparam \Mux30~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux15~0 (
	.dataa(ram_in_reg_0_1),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mux7~0_combout ),
	.cin(gnd),
	.combout(\Mux15~0_combout ),
	.cout());
defparam \Mux15~0 .lut_mask = 16'hAAFF;
defparam \Mux15~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux31~0 (
	.dataa(ram_in_reg_0_3),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mux7~0_combout ),
	.cin(gnd),
	.combout(\Mux31~0_combout ),
	.cout());
defparam \Mux31~0 .lut_mask = 16'hAAFF;
defparam \Mux31~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux0~4 (
	.dataa(\r_array_out[2][6]~16_combout ),
	.datab(ram_in_reg_7_0),
	.datac(\r_array_out[2][6]~17_combout ),
	.datad(\Mux0~2_combout ),
	.cin(gnd),
	.combout(\Mux0~4_combout ),
	.cout());
defparam \Mux0~4 .lut_mask = 16'hFFDE;
defparam \Mux0~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux0~5 (
	.dataa(ram_in_reg_3_0),
	.datab(\r_array_out[2][6]~16_combout ),
	.datac(\Mux0~4_combout ),
	.datad(ram_in_reg_6_0),
	.cin(gnd),
	.combout(\Mux0~5_combout ),
	.cout());
defparam \Mux0~5 .lut_mask = 16'hFFBE;
defparam \Mux0~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux16~4 (
	.dataa(\r_array_out[2][6]~16_combout ),
	.datab(ram_in_reg_7_2),
	.datac(\r_array_out[2][6]~17_combout ),
	.datad(\Mux16~2_combout ),
	.cin(gnd),
	.combout(\Mux16~4_combout ),
	.cout());
defparam \Mux16~4 .lut_mask = 16'hFFDE;
defparam \Mux16~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux16~5 (
	.dataa(ram_in_reg_3_2),
	.datab(\r_array_out[2][6]~16_combout ),
	.datac(\Mux16~4_combout ),
	.datad(ram_in_reg_6_2),
	.cin(gnd),
	.combout(\Mux16~5_combout ),
	.cout());
defparam \Mux16~5 .lut_mask = 16'hFFBE;
defparam \Mux16~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux8~4 (
	.dataa(\r_array_out[2][6]~16_combout ),
	.datab(ram_in_reg_7_1),
	.datac(\r_array_out[2][6]~17_combout ),
	.datad(\Mux8~2_combout ),
	.cin(gnd),
	.combout(\Mux8~4_combout ),
	.cout());
defparam \Mux8~4 .lut_mask = 16'hFFDE;
defparam \Mux8~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux8~5 (
	.dataa(ram_in_reg_3_1),
	.datab(\r_array_out[2][6]~16_combout ),
	.datac(\Mux8~4_combout ),
	.datad(ram_in_reg_6_1),
	.cin(gnd),
	.combout(\Mux8~5_combout ),
	.cout());
defparam \Mux8~5 .lut_mask = 16'hFFBE;
defparam \Mux8~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux24~4 (
	.dataa(\r_array_out[2][6]~16_combout ),
	.datab(ram_in_reg_7_3),
	.datac(\r_array_out[2][6]~17_combout ),
	.datad(\Mux24~2_combout ),
	.cin(gnd),
	.combout(\Mux24~4_combout ),
	.cout());
defparam \Mux24~4 .lut_mask = 16'hFFDE;
defparam \Mux24~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux24~5 (
	.dataa(ram_in_reg_3_3),
	.datab(\r_array_out[2][6]~16_combout ),
	.datac(\Mux24~4_combout ),
	.datad(ram_in_reg_6_3),
	.cin(gnd),
	.combout(\Mux24~5_combout ),
	.cout());
defparam \Mux24~5 .lut_mask = 16'hFFBE;
defparam \Mux24~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux32~1 (
	.dataa(\r_array_out[2][6]~17_combout ),
	.datab(ram_in_reg_3_4),
	.datac(\r_array_out[2][6]~16_combout ),
	.datad(\Mux32~0_combout ),
	.cin(gnd),
	.combout(\Mux32~1_combout ),
	.cout());
defparam \Mux32~1 .lut_mask = 16'hFFDE;
defparam \Mux32~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux32~2 (
	.dataa(ram_in_reg_7_4),
	.datab(\r_array_out[2][6]~17_combout ),
	.datac(\Mux32~1_combout ),
	.datad(ram_in_reg_6_4),
	.cin(gnd),
	.combout(\Mux32~2_combout ),
	.cout());
defparam \Mux32~2 .lut_mask = 16'hFFBE;
defparam \Mux32~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux48~1 (
	.dataa(\r_array_out[2][6]~17_combout ),
	.datab(ram_in_reg_3_6),
	.datac(\r_array_out[2][6]~16_combout ),
	.datad(\Mux48~0_combout ),
	.cin(gnd),
	.combout(\Mux48~1_combout ),
	.cout());
defparam \Mux48~1 .lut_mask = 16'hFFDE;
defparam \Mux48~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux48~2 (
	.dataa(ram_in_reg_7_6),
	.datab(\r_array_out[2][6]~17_combout ),
	.datac(\Mux48~1_combout ),
	.datad(ram_in_reg_6_6),
	.cin(gnd),
	.combout(\Mux48~2_combout ),
	.cout());
defparam \Mux48~2 .lut_mask = 16'hFFBE;
defparam \Mux48~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux33~0 (
	.dataa(\r_array_out[2][6]~16_combout ),
	.datab(ram_in_reg_6_4),
	.datac(\r_array_out[2][6]~17_combout ),
	.datad(\Mux32~3_combout ),
	.cin(gnd),
	.combout(\Mux33~0_combout ),
	.cout());
defparam \Mux33~0 .lut_mask = 16'hFFDE;
defparam \Mux33~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux33~1 (
	.dataa(ram_in_reg_2_4),
	.datab(\r_array_out[2][6]~16_combout ),
	.datac(\Mux33~0_combout ),
	.datad(ram_in_reg_5_4),
	.cin(gnd),
	.combout(\Mux33~1_combout ),
	.cout());
defparam \Mux33~1 .lut_mask = 16'hFFBE;
defparam \Mux33~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux49~0 (
	.dataa(\r_array_out[2][6]~16_combout ),
	.datab(ram_in_reg_6_6),
	.datac(\r_array_out[2][6]~17_combout ),
	.datad(\Mux48~3_combout ),
	.cin(gnd),
	.combout(\Mux49~0_combout ),
	.cout());
defparam \Mux49~0 .lut_mask = 16'hFFDE;
defparam \Mux49~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux49~1 (
	.dataa(ram_in_reg_2_6),
	.datab(\r_array_out[2][6]~16_combout ),
	.datac(\Mux49~0_combout ),
	.datad(ram_in_reg_5_6),
	.cin(gnd),
	.combout(\Mux49~1_combout ),
	.cout());
defparam \Mux49~1 .lut_mask = 16'hFFBE;
defparam \Mux49~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux38~2 (
	.dataa(slb_last_1),
	.datab(slb_last_2),
	.datac(block_dft_i_en),
	.datad(\i_array_out[0][3]~2_combout ),
	.cin(gnd),
	.combout(\Mux38~2_combout ),
	.cout());
defparam \Mux38~2 .lut_mask = 16'hFFF7;
defparam \Mux38~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux54~2 (
	.dataa(slb_last_1),
	.datab(slb_last_2),
	.datac(block_dft_i_en),
	.datad(\i_array_out[2][3]~3_combout ),
	.cin(gnd),
	.combout(\Mux54~2_combout ),
	.cout());
defparam \Mux54~2 .lut_mask = 16'hFFF7;
defparam \Mux54~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux39~0 (
	.dataa(ram_in_reg_0_4),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mux7~0_combout ),
	.cin(gnd),
	.combout(\Mux39~0_combout ),
	.cout());
defparam \Mux39~0 .lut_mask = 16'hAAFF;
defparam \Mux39~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux55~0 (
	.dataa(ram_in_reg_0_6),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mux7~0_combout ),
	.cin(gnd),
	.combout(\Mux55~0_combout ),
	.cout());
defparam \Mux55~0 .lut_mask = 16'hAAFF;
defparam \Mux55~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux40~1 (
	.dataa(\r_array_out[2][6]~17_combout ),
	.datab(ram_in_reg_3_5),
	.datac(\r_array_out[2][6]~16_combout ),
	.datad(\Mux40~0_combout ),
	.cin(gnd),
	.combout(\Mux40~1_combout ),
	.cout());
defparam \Mux40~1 .lut_mask = 16'hFFDE;
defparam \Mux40~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux40~2 (
	.dataa(ram_in_reg_7_5),
	.datab(\r_array_out[2][6]~17_combout ),
	.datac(\Mux40~1_combout ),
	.datad(ram_in_reg_6_5),
	.cin(gnd),
	.combout(\Mux40~2_combout ),
	.cout());
defparam \Mux40~2 .lut_mask = 16'hFFBE;
defparam \Mux40~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux56~1 (
	.dataa(\r_array_out[2][6]~16_combout ),
	.datab(ram_in_reg_7_7),
	.datac(\r_array_out[2][6]~17_combout ),
	.datad(\Mux56~0_combout ),
	.cin(gnd),
	.combout(\Mux56~1_combout ),
	.cout());
defparam \Mux56~1 .lut_mask = 16'hFFDE;
defparam \Mux56~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux56~2 (
	.dataa(ram_in_reg_3_7),
	.datab(\r_array_out[2][6]~16_combout ),
	.datac(\Mux56~1_combout ),
	.datad(ram_in_reg_6_7),
	.cin(gnd),
	.combout(\Mux56~2_combout ),
	.cout());
defparam \Mux56~2 .lut_mask = 16'hFFBE;
defparam \Mux56~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux41~0 (
	.dataa(\r_array_out[2][6]~16_combout ),
	.datab(ram_in_reg_6_5),
	.datac(\r_array_out[2][6]~17_combout ),
	.datad(\Mux40~3_combout ),
	.cin(gnd),
	.combout(\Mux41~0_combout ),
	.cout());
defparam \Mux41~0 .lut_mask = 16'hFFDE;
defparam \Mux41~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux41~1 (
	.dataa(ram_in_reg_2_5),
	.datab(\r_array_out[2][6]~16_combout ),
	.datac(\Mux41~0_combout ),
	.datad(ram_in_reg_5_5),
	.cin(gnd),
	.combout(\Mux41~1_combout ),
	.cout());
defparam \Mux41~1 .lut_mask = 16'hFFBE;
defparam \Mux41~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux57~0 (
	.dataa(\r_array_out[2][6]~16_combout ),
	.datab(ram_in_reg_6_7),
	.datac(\r_array_out[2][6]~17_combout ),
	.datad(\Mux56~3_combout ),
	.cin(gnd),
	.combout(\Mux57~0_combout ),
	.cout());
defparam \Mux57~0 .lut_mask = 16'hFFDE;
defparam \Mux57~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux57~1 (
	.dataa(ram_in_reg_2_7),
	.datab(\r_array_out[2][6]~16_combout ),
	.datac(\Mux57~0_combout ),
	.datad(ram_in_reg_5_7),
	.cin(gnd),
	.combout(\Mux57~1_combout ),
	.cout());
defparam \Mux57~1 .lut_mask = 16'hFFBE;
defparam \Mux57~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux46~2 (
	.dataa(slb_last_1),
	.datab(slb_last_2),
	.datac(block_dft_i_en),
	.datad(\i_array_out[1][3]~10_combout ),
	.cin(gnd),
	.combout(\Mux46~2_combout ),
	.cout());
defparam \Mux46~2 .lut_mask = 16'hFFF7;
defparam \Mux46~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux62~2 (
	.dataa(slb_last_1),
	.datab(slb_last_2),
	.datac(block_dft_i_en),
	.datad(\i_array_out[3][3]~11_combout ),
	.cin(gnd),
	.combout(\Mux62~2_combout ),
	.cout());
defparam \Mux62~2 .lut_mask = 16'hFFF7;
defparam \Mux62~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux47~0 (
	.dataa(ram_in_reg_0_5),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mux7~0_combout ),
	.cin(gnd),
	.combout(\Mux47~0_combout ),
	.cout());
defparam \Mux47~0 .lut_mask = 16'hAAFF;
defparam \Mux47~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux63~0 (
	.dataa(ram_in_reg_0_7),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mux7~0_combout ),
	.cin(gnd),
	.combout(\Mux63~0_combout ),
	.cout());
defparam \Mux63~0 .lut_mask = 16'hAAFF;
defparam \Mux63~0 .sum_lutc_input = "datac";

endmodule

module fft_asj_fft_bfp_i_fft_120_1 (
	r_array_out_3_0,
	i_array_out_3_0,
	r_array_out_3_1,
	i_array_out_3_1,
	r_array_out_3_2,
	i_array_out_3_2,
	r_array_out_3_3,
	i_array_out_3_3,
	r_array_out_4_0,
	i_array_out_4_0,
	r_array_out_4_1,
	i_array_out_4_1,
	r_array_out_4_2,
	i_array_out_4_2,
	r_array_out_4_3,
	i_array_out_4_3,
	r_array_out_5_0,
	i_array_out_5_0,
	r_array_out_5_1,
	i_array_out_5_1,
	r_array_out_5_2,
	i_array_out_5_2,
	r_array_out_5_3,
	i_array_out_5_3,
	i_array_out_2_2,
	i_array_out_2_1,
	i_array_out_2_0,
	i_array_out_2_3,
	r_array_out_2_2,
	r_array_out_2_1,
	r_array_out_2_0,
	r_array_out_2_3,
	global_clock_enable,
	slb_last_0,
	slb_last_1,
	slb_last_2,
	r_array_out_7_0,
	i_array_out_7_0,
	r_array_out_7_1,
	i_array_out_7_1,
	r_array_out_7_2,
	i_array_out_7_2,
	r_array_out_7_3,
	i_array_out_7_3,
	r_array_out_6_0,
	i_array_out_6_0,
	r_array_out_6_1,
	i_array_out_6_1,
	r_array_out_6_2,
	i_array_out_6_2,
	r_array_out_6_3,
	i_array_out_6_3,
	i_array_out_1_2,
	i_array_out_1_1,
	i_array_out_1_0,
	i_array_out_1_3,
	i_array_out_0_2,
	i_array_out_0_1,
	i_array_out_0_0,
	i_array_out_0_3,
	r_array_out_1_2,
	r_array_out_1_1,
	r_array_out_1_0,
	r_array_out_1_3,
	r_array_out_0_2,
	r_array_out_0_1,
	r_array_out_0_0,
	r_array_out_0_3,
	scale_dft_o_en,
	do_tdl0033,
	do_tdl0037,
	do_tdl0034,
	do_tdl0035,
	do_tdl0036,
	do_tdl0031,
	do_tdl0030,
	slb_1pt_0,
	do_tdl0032,
	slb_1pt_2,
	slb_1pt_1,
	do_tdl0133,
	do_tdl0137,
	do_tdl0134,
	do_tdl0135,
	do_tdl0136,
	do_tdl0131,
	do_tdl0130,
	do_tdl0132,
	do_tdl1033,
	do_tdl1037,
	do_tdl1034,
	do_tdl1035,
	do_tdl1036,
	do_tdl1031,
	do_tdl1030,
	do_tdl1032,
	do_tdl1133,
	do_tdl1137,
	do_tdl1134,
	do_tdl1135,
	do_tdl1136,
	do_tdl1131,
	do_tdl1130,
	do_tdl1132,
	do_tdl2033,
	do_tdl2037,
	do_tdl2034,
	do_tdl2035,
	do_tdl2036,
	do_tdl2031,
	do_tdl2030,
	do_tdl2032,
	do_tdl2133,
	do_tdl2137,
	do_tdl2134,
	do_tdl2135,
	do_tdl2136,
	do_tdl2131,
	do_tdl2130,
	do_tdl2132,
	do_tdl3033,
	do_tdl3037,
	do_tdl3034,
	do_tdl3035,
	do_tdl3036,
	do_tdl3031,
	do_tdl3030,
	do_tdl3032,
	do_tdl3133,
	do_tdl3137,
	do_tdl3134,
	do_tdl3135,
	do_tdl3136,
	do_tdl3131,
	do_tdl3130,
	do_tdl3132,
	clk)/* synthesis synthesis_greybox=1 */;
output 	r_array_out_3_0;
output 	i_array_out_3_0;
output 	r_array_out_3_1;
output 	i_array_out_3_1;
output 	r_array_out_3_2;
output 	i_array_out_3_2;
output 	r_array_out_3_3;
output 	i_array_out_3_3;
output 	r_array_out_4_0;
output 	i_array_out_4_0;
output 	r_array_out_4_1;
output 	i_array_out_4_1;
output 	r_array_out_4_2;
output 	i_array_out_4_2;
output 	r_array_out_4_3;
output 	i_array_out_4_3;
output 	r_array_out_5_0;
output 	i_array_out_5_0;
output 	r_array_out_5_1;
output 	i_array_out_5_1;
output 	r_array_out_5_2;
output 	i_array_out_5_2;
output 	r_array_out_5_3;
output 	i_array_out_5_3;
output 	i_array_out_2_2;
output 	i_array_out_2_1;
output 	i_array_out_2_0;
output 	i_array_out_2_3;
output 	r_array_out_2_2;
output 	r_array_out_2_1;
output 	r_array_out_2_0;
output 	r_array_out_2_3;
input 	global_clock_enable;
input 	slb_last_0;
input 	slb_last_1;
input 	slb_last_2;
output 	r_array_out_7_0;
output 	i_array_out_7_0;
output 	r_array_out_7_1;
output 	i_array_out_7_1;
output 	r_array_out_7_2;
output 	i_array_out_7_2;
output 	r_array_out_7_3;
output 	i_array_out_7_3;
output 	r_array_out_6_0;
output 	i_array_out_6_0;
output 	r_array_out_6_1;
output 	i_array_out_6_1;
output 	r_array_out_6_2;
output 	i_array_out_6_2;
output 	r_array_out_6_3;
output 	i_array_out_6_3;
output 	i_array_out_1_2;
output 	i_array_out_1_1;
output 	i_array_out_1_0;
output 	i_array_out_1_3;
output 	i_array_out_0_2;
output 	i_array_out_0_1;
output 	i_array_out_0_0;
output 	i_array_out_0_3;
output 	r_array_out_1_2;
output 	r_array_out_1_1;
output 	r_array_out_1_0;
output 	r_array_out_1_3;
output 	r_array_out_0_2;
output 	r_array_out_0_1;
output 	r_array_out_0_0;
output 	r_array_out_0_3;
input 	scale_dft_o_en;
input 	do_tdl0033;
input 	do_tdl0037;
input 	do_tdl0034;
input 	do_tdl0035;
input 	do_tdl0036;
input 	do_tdl0031;
input 	do_tdl0030;
input 	slb_1pt_0;
input 	do_tdl0032;
input 	slb_1pt_2;
input 	slb_1pt_1;
input 	do_tdl0133;
input 	do_tdl0137;
input 	do_tdl0134;
input 	do_tdl0135;
input 	do_tdl0136;
input 	do_tdl0131;
input 	do_tdl0130;
input 	do_tdl0132;
input 	do_tdl1033;
input 	do_tdl1037;
input 	do_tdl1034;
input 	do_tdl1035;
input 	do_tdl1036;
input 	do_tdl1031;
input 	do_tdl1030;
input 	do_tdl1032;
input 	do_tdl1133;
input 	do_tdl1137;
input 	do_tdl1134;
input 	do_tdl1135;
input 	do_tdl1136;
input 	do_tdl1131;
input 	do_tdl1130;
input 	do_tdl1132;
input 	do_tdl2033;
input 	do_tdl2037;
input 	do_tdl2034;
input 	do_tdl2035;
input 	do_tdl2036;
input 	do_tdl2031;
input 	do_tdl2030;
input 	do_tdl2032;
input 	do_tdl2133;
input 	do_tdl2137;
input 	do_tdl2134;
input 	do_tdl2135;
input 	do_tdl2136;
input 	do_tdl2131;
input 	do_tdl2130;
input 	do_tdl2132;
input 	do_tdl3033;
input 	do_tdl3037;
input 	do_tdl3034;
input 	do_tdl3035;
input 	do_tdl3036;
input 	do_tdl3031;
input 	do_tdl3030;
input 	do_tdl3032;
input 	do_tdl3133;
input 	do_tdl3137;
input 	do_tdl3134;
input 	do_tdl3135;
input 	do_tdl3136;
input 	do_tdl3131;
input 	do_tdl3130;
input 	do_tdl3132;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \r_array_out[0][3]~0_combout ;
wire \Mux1~1_combout ;
wire \i_array_out[0][3]~0_combout ;
wire \Mux33~1_combout ;
wire \r_array_out[1][3]~1_combout ;
wire \Mux9~1_combout ;
wire \i_array_out[1][3]~1_combout ;
wire \Mux41~1_combout ;
wire \r_array_out[2][3]~2_combout ;
wire \Mux17~1_combout ;
wire \i_array_out[2][3]~2_combout ;
wire \Mux49~1_combout ;
wire \r_array_out[3][3]~3_combout ;
wire \Mux25~1_combout ;
wire \i_array_out[3][3]~3_combout ;
wire \Mux57~1_combout ;
wire \r_array_out[0][2]~14_combout ;
wire \Mux1~2_combout ;
wire \r_array_out[0][4]~4_combout ;
wire \i_array_out[0][2]~14_combout ;
wire \Mux33~2_combout ;
wire \i_array_out[0][4]~4_combout ;
wire \r_array_out[1][2]~13_combout ;
wire \Mux9~2_combout ;
wire \r_array_out[1][4]~5_combout ;
wire \i_array_out[1][2]~13_combout ;
wire \Mux41~2_combout ;
wire \i_array_out[1][4]~5_combout ;
wire \r_array_out[2][2]~12_combout ;
wire \Mux17~2_combout ;
wire \r_array_out[2][4]~6_combout ;
wire \i_array_out[2][2]~12_combout ;
wire \Mux49~2_combout ;
wire \i_array_out[2][4]~6_combout ;
wire \r_array_out[3][2]~15_combout ;
wire \Mux25~2_combout ;
wire \r_array_out[3][4]~7_combout ;
wire \i_array_out[3][2]~15_combout ;
wire \Mux57~2_combout ;
wire \i_array_out[3][4]~7_combout ;
wire \Mux1~0_combout ;
wire \r_array_out[0][5]~8_combout ;
wire \Mux33~0_combout ;
wire \i_array_out[0][5]~8_combout ;
wire \Mux9~0_combout ;
wire \r_array_out[1][5]~9_combout ;
wire \Mux41~0_combout ;
wire \i_array_out[1][5]~9_combout ;
wire \Mux17~0_combout ;
wire \r_array_out[2][5]~10_combout ;
wire \Mux49~0_combout ;
wire \i_array_out[2][5]~10_combout ;
wire \Mux25~0_combout ;
wire \r_array_out[3][5]~11_combout ;
wire \Mux57~0_combout ;
wire \i_array_out[3][5]~11_combout ;
wire \Mux49~5_combout ;
wire \Mux41~5_combout ;
wire \Mux33~5_combout ;
wire \Mux57~5_combout ;
wire \Mux17~5_combout ;
wire \Mux9~5_combout ;
wire \Mux1~5_combout ;
wire \Mux25~5_combout ;
wire \i_array_out[0][6]~16_combout ;
wire \i_array_out[0][6]~17_combout ;
wire \Mux0~0_combout ;
wire \Mux0~1_combout ;
wire \Mux32~0_combout ;
wire \Mux32~1_combout ;
wire \Mux8~0_combout ;
wire \Mux8~1_combout ;
wire \Mux40~0_combout ;
wire \Mux40~1_combout ;
wire \Mux16~0_combout ;
wire \Mux16~1_combout ;
wire \Mux48~0_combout ;
wire \Mux48~1_combout ;
wire \Mux24~0_combout ;
wire \Mux24~1_combout ;
wire \Mux56~0_combout ;
wire \Mux56~1_combout ;
wire \Mux1~3_combout ;
wire \Mux1~4_combout ;
wire \Mux33~3_combout ;
wire \Mux33~4_combout ;
wire \Mux9~3_combout ;
wire \Mux9~4_combout ;
wire \Mux41~3_combout ;
wire \Mux41~4_combout ;
wire \Mux17~3_combout ;
wire \Mux17~4_combout ;
wire \Mux49~3_combout ;
wire \Mux49~4_combout ;
wire \Mux25~3_combout ;
wire \Mux25~4_combout ;
wire \Mux57~3_combout ;
wire \Mux57~4_combout ;
wire \Mux54~2_combout ;
wire \Mux46~2_combout ;
wire \Mux38~2_combout ;
wire \Mux62~2_combout ;
wire \Mux7~0_combout ;
wire \Mux55~0_combout ;
wire \Mux47~0_combout ;
wire \Mux39~0_combout ;
wire \Mux63~0_combout ;
wire \Mux22~2_combout ;
wire \Mux14~2_combout ;
wire \Mux6~2_combout ;
wire \Mux30~2_combout ;
wire \Mux23~0_combout ;
wire \Mux15~0_combout ;
wire \Mux7~1_combout ;
wire \Mux31~0_combout ;


dffeas \r_array_out[0][3] (
	.clk(clk),
	.d(\r_array_out[0][3]~0_combout ),
	.asdata(\Mux1~1_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_1pt_2),
	.sload(slb_1pt_1),
	.ena(global_clock_enable),
	.q(r_array_out_3_0),
	.prn(vcc));
defparam \r_array_out[0][3] .is_wysiwyg = "true";
defparam \r_array_out[0][3] .power_up = "low";

dffeas \i_array_out[0][3] (
	.clk(clk),
	.d(\i_array_out[0][3]~0_combout ),
	.asdata(\Mux33~1_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_1pt_2),
	.sload(slb_1pt_1),
	.ena(global_clock_enable),
	.q(i_array_out_3_0),
	.prn(vcc));
defparam \i_array_out[0][3] .is_wysiwyg = "true";
defparam \i_array_out[0][3] .power_up = "low";

dffeas \r_array_out[1][3] (
	.clk(clk),
	.d(\r_array_out[1][3]~1_combout ),
	.asdata(\Mux9~1_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_1pt_2),
	.sload(slb_1pt_1),
	.ena(global_clock_enable),
	.q(r_array_out_3_1),
	.prn(vcc));
defparam \r_array_out[1][3] .is_wysiwyg = "true";
defparam \r_array_out[1][3] .power_up = "low";

dffeas \i_array_out[1][3] (
	.clk(clk),
	.d(\i_array_out[1][3]~1_combout ),
	.asdata(\Mux41~1_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_1pt_2),
	.sload(slb_1pt_1),
	.ena(global_clock_enable),
	.q(i_array_out_3_1),
	.prn(vcc));
defparam \i_array_out[1][3] .is_wysiwyg = "true";
defparam \i_array_out[1][3] .power_up = "low";

dffeas \r_array_out[2][3] (
	.clk(clk),
	.d(\r_array_out[2][3]~2_combout ),
	.asdata(\Mux17~1_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_1pt_2),
	.sload(slb_1pt_1),
	.ena(global_clock_enable),
	.q(r_array_out_3_2),
	.prn(vcc));
defparam \r_array_out[2][3] .is_wysiwyg = "true";
defparam \r_array_out[2][3] .power_up = "low";

dffeas \i_array_out[2][3] (
	.clk(clk),
	.d(\i_array_out[2][3]~2_combout ),
	.asdata(\Mux49~1_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_1pt_2),
	.sload(slb_1pt_1),
	.ena(global_clock_enable),
	.q(i_array_out_3_2),
	.prn(vcc));
defparam \i_array_out[2][3] .is_wysiwyg = "true";
defparam \i_array_out[2][3] .power_up = "low";

dffeas \r_array_out[3][3] (
	.clk(clk),
	.d(\r_array_out[3][3]~3_combout ),
	.asdata(\Mux25~1_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_1pt_2),
	.sload(slb_1pt_1),
	.ena(global_clock_enable),
	.q(r_array_out_3_3),
	.prn(vcc));
defparam \r_array_out[3][3] .is_wysiwyg = "true";
defparam \r_array_out[3][3] .power_up = "low";

dffeas \i_array_out[3][3] (
	.clk(clk),
	.d(\i_array_out[3][3]~3_combout ),
	.asdata(\Mux57~1_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_1pt_2),
	.sload(slb_1pt_1),
	.ena(global_clock_enable),
	.q(i_array_out_3_3),
	.prn(vcc));
defparam \i_array_out[3][3] .is_wysiwyg = "true";
defparam \i_array_out[3][3] .power_up = "low";

dffeas \r_array_out[0][4] (
	.clk(clk),
	.d(\r_array_out[0][4]~4_combout ),
	.asdata(do_tdl0030),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_1pt_2),
	.ena(global_clock_enable),
	.q(r_array_out_4_0),
	.prn(vcc));
defparam \r_array_out[0][4] .is_wysiwyg = "true";
defparam \r_array_out[0][4] .power_up = "low";

dffeas \i_array_out[0][4] (
	.clk(clk),
	.d(\i_array_out[0][4]~4_combout ),
	.asdata(do_tdl0130),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_1pt_2),
	.ena(global_clock_enable),
	.q(i_array_out_4_0),
	.prn(vcc));
defparam \i_array_out[0][4] .is_wysiwyg = "true";
defparam \i_array_out[0][4] .power_up = "low";

dffeas \r_array_out[1][4] (
	.clk(clk),
	.d(\r_array_out[1][4]~5_combout ),
	.asdata(do_tdl1030),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_1pt_2),
	.ena(global_clock_enable),
	.q(r_array_out_4_1),
	.prn(vcc));
defparam \r_array_out[1][4] .is_wysiwyg = "true";
defparam \r_array_out[1][4] .power_up = "low";

dffeas \i_array_out[1][4] (
	.clk(clk),
	.d(\i_array_out[1][4]~5_combout ),
	.asdata(do_tdl1130),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_1pt_2),
	.ena(global_clock_enable),
	.q(i_array_out_4_1),
	.prn(vcc));
defparam \i_array_out[1][4] .is_wysiwyg = "true";
defparam \i_array_out[1][4] .power_up = "low";

dffeas \r_array_out[2][4] (
	.clk(clk),
	.d(\r_array_out[2][4]~6_combout ),
	.asdata(do_tdl2030),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_1pt_2),
	.ena(global_clock_enable),
	.q(r_array_out_4_2),
	.prn(vcc));
defparam \r_array_out[2][4] .is_wysiwyg = "true";
defparam \r_array_out[2][4] .power_up = "low";

dffeas \i_array_out[2][4] (
	.clk(clk),
	.d(\i_array_out[2][4]~6_combout ),
	.asdata(do_tdl2130),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_1pt_2),
	.ena(global_clock_enable),
	.q(i_array_out_4_2),
	.prn(vcc));
defparam \i_array_out[2][4] .is_wysiwyg = "true";
defparam \i_array_out[2][4] .power_up = "low";

dffeas \r_array_out[3][4] (
	.clk(clk),
	.d(\r_array_out[3][4]~7_combout ),
	.asdata(do_tdl3030),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_1pt_2),
	.ena(global_clock_enable),
	.q(r_array_out_4_3),
	.prn(vcc));
defparam \r_array_out[3][4] .is_wysiwyg = "true";
defparam \r_array_out[3][4] .power_up = "low";

dffeas \i_array_out[3][4] (
	.clk(clk),
	.d(\i_array_out[3][4]~7_combout ),
	.asdata(do_tdl3130),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_1pt_2),
	.ena(global_clock_enable),
	.q(i_array_out_4_3),
	.prn(vcc));
defparam \i_array_out[3][4] .is_wysiwyg = "true";
defparam \i_array_out[3][4] .power_up = "low";

dffeas \r_array_out[0][5] (
	.clk(clk),
	.d(\r_array_out[0][5]~8_combout ),
	.asdata(do_tdl0031),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_1pt_2),
	.ena(global_clock_enable),
	.q(r_array_out_5_0),
	.prn(vcc));
defparam \r_array_out[0][5] .is_wysiwyg = "true";
defparam \r_array_out[0][5] .power_up = "low";

dffeas \i_array_out[0][5] (
	.clk(clk),
	.d(\i_array_out[0][5]~8_combout ),
	.asdata(do_tdl0131),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_1pt_2),
	.ena(global_clock_enable),
	.q(i_array_out_5_0),
	.prn(vcc));
defparam \i_array_out[0][5] .is_wysiwyg = "true";
defparam \i_array_out[0][5] .power_up = "low";

dffeas \r_array_out[1][5] (
	.clk(clk),
	.d(\r_array_out[1][5]~9_combout ),
	.asdata(do_tdl1031),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_1pt_2),
	.ena(global_clock_enable),
	.q(r_array_out_5_1),
	.prn(vcc));
defparam \r_array_out[1][5] .is_wysiwyg = "true";
defparam \r_array_out[1][5] .power_up = "low";

dffeas \i_array_out[1][5] (
	.clk(clk),
	.d(\i_array_out[1][5]~9_combout ),
	.asdata(do_tdl1131),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_1pt_2),
	.ena(global_clock_enable),
	.q(i_array_out_5_1),
	.prn(vcc));
defparam \i_array_out[1][5] .is_wysiwyg = "true";
defparam \i_array_out[1][5] .power_up = "low";

dffeas \r_array_out[2][5] (
	.clk(clk),
	.d(\r_array_out[2][5]~10_combout ),
	.asdata(do_tdl2031),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_1pt_2),
	.ena(global_clock_enable),
	.q(r_array_out_5_2),
	.prn(vcc));
defparam \r_array_out[2][5] .is_wysiwyg = "true";
defparam \r_array_out[2][5] .power_up = "low";

dffeas \i_array_out[2][5] (
	.clk(clk),
	.d(\i_array_out[2][5]~10_combout ),
	.asdata(do_tdl2131),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_1pt_2),
	.ena(global_clock_enable),
	.q(i_array_out_5_2),
	.prn(vcc));
defparam \i_array_out[2][5] .is_wysiwyg = "true";
defparam \i_array_out[2][5] .power_up = "low";

dffeas \r_array_out[3][5] (
	.clk(clk),
	.d(\r_array_out[3][5]~11_combout ),
	.asdata(do_tdl3031),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_1pt_2),
	.ena(global_clock_enable),
	.q(r_array_out_5_3),
	.prn(vcc));
defparam \r_array_out[3][5] .is_wysiwyg = "true";
defparam \r_array_out[3][5] .power_up = "low";

dffeas \i_array_out[3][5] (
	.clk(clk),
	.d(\i_array_out[3][5]~11_combout ),
	.asdata(do_tdl3131),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_1pt_2),
	.ena(global_clock_enable),
	.q(i_array_out_5_3),
	.prn(vcc));
defparam \i_array_out[3][5] .is_wysiwyg = "true";
defparam \i_array_out[3][5] .power_up = "low";

dffeas \i_array_out[2][2] (
	.clk(clk),
	.d(\i_array_out[2][2]~12_combout ),
	.asdata(\Mux49~5_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_1pt_2),
	.sload(!slb_1pt_1),
	.ena(global_clock_enable),
	.q(i_array_out_2_2),
	.prn(vcc));
defparam \i_array_out[2][2] .is_wysiwyg = "true";
defparam \i_array_out[2][2] .power_up = "low";

dffeas \i_array_out[1][2] (
	.clk(clk),
	.d(\i_array_out[1][2]~13_combout ),
	.asdata(\Mux41~5_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_1pt_2),
	.sload(!slb_1pt_1),
	.ena(global_clock_enable),
	.q(i_array_out_2_1),
	.prn(vcc));
defparam \i_array_out[1][2] .is_wysiwyg = "true";
defparam \i_array_out[1][2] .power_up = "low";

dffeas \i_array_out[0][2] (
	.clk(clk),
	.d(\i_array_out[0][2]~14_combout ),
	.asdata(\Mux33~5_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_1pt_2),
	.sload(!slb_1pt_1),
	.ena(global_clock_enable),
	.q(i_array_out_2_0),
	.prn(vcc));
defparam \i_array_out[0][2] .is_wysiwyg = "true";
defparam \i_array_out[0][2] .power_up = "low";

dffeas \i_array_out[3][2] (
	.clk(clk),
	.d(\i_array_out[3][2]~15_combout ),
	.asdata(\Mux57~5_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_1pt_2),
	.sload(!slb_1pt_1),
	.ena(global_clock_enable),
	.q(i_array_out_2_3),
	.prn(vcc));
defparam \i_array_out[3][2] .is_wysiwyg = "true";
defparam \i_array_out[3][2] .power_up = "low";

dffeas \r_array_out[2][2] (
	.clk(clk),
	.d(\r_array_out[2][2]~12_combout ),
	.asdata(\Mux17~5_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_1pt_2),
	.sload(!slb_1pt_1),
	.ena(global_clock_enable),
	.q(r_array_out_2_2),
	.prn(vcc));
defparam \r_array_out[2][2] .is_wysiwyg = "true";
defparam \r_array_out[2][2] .power_up = "low";

dffeas \r_array_out[1][2] (
	.clk(clk),
	.d(\r_array_out[1][2]~13_combout ),
	.asdata(\Mux9~5_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_1pt_2),
	.sload(!slb_1pt_1),
	.ena(global_clock_enable),
	.q(r_array_out_2_1),
	.prn(vcc));
defparam \r_array_out[1][2] .is_wysiwyg = "true";
defparam \r_array_out[1][2] .power_up = "low";

dffeas \r_array_out[0][2] (
	.clk(clk),
	.d(\r_array_out[0][2]~14_combout ),
	.asdata(\Mux1~5_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_1pt_2),
	.sload(!slb_1pt_1),
	.ena(global_clock_enable),
	.q(r_array_out_2_0),
	.prn(vcc));
defparam \r_array_out[0][2] .is_wysiwyg = "true";
defparam \r_array_out[0][2] .power_up = "low";

dffeas \r_array_out[3][2] (
	.clk(clk),
	.d(\r_array_out[3][2]~15_combout ),
	.asdata(\Mux25~5_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_1pt_2),
	.sload(!slb_1pt_1),
	.ena(global_clock_enable),
	.q(r_array_out_2_3),
	.prn(vcc));
defparam \r_array_out[3][2] .is_wysiwyg = "true";
defparam \r_array_out[3][2] .power_up = "low";

dffeas \r_array_out[0][7] (
	.clk(clk),
	.d(\Mux0~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_7_0),
	.prn(vcc));
defparam \r_array_out[0][7] .is_wysiwyg = "true";
defparam \r_array_out[0][7] .power_up = "low";

dffeas \i_array_out[0][7] (
	.clk(clk),
	.d(\Mux32~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_7_0),
	.prn(vcc));
defparam \i_array_out[0][7] .is_wysiwyg = "true";
defparam \i_array_out[0][7] .power_up = "low";

dffeas \r_array_out[1][7] (
	.clk(clk),
	.d(\Mux8~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_7_1),
	.prn(vcc));
defparam \r_array_out[1][7] .is_wysiwyg = "true";
defparam \r_array_out[1][7] .power_up = "low";

dffeas \i_array_out[1][7] (
	.clk(clk),
	.d(\Mux40~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_7_1),
	.prn(vcc));
defparam \i_array_out[1][7] .is_wysiwyg = "true";
defparam \i_array_out[1][7] .power_up = "low";

dffeas \r_array_out[2][7] (
	.clk(clk),
	.d(\Mux16~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_7_2),
	.prn(vcc));
defparam \r_array_out[2][7] .is_wysiwyg = "true";
defparam \r_array_out[2][7] .power_up = "low";

dffeas \i_array_out[2][7] (
	.clk(clk),
	.d(\Mux48~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_7_2),
	.prn(vcc));
defparam \i_array_out[2][7] .is_wysiwyg = "true";
defparam \i_array_out[2][7] .power_up = "low";

dffeas \r_array_out[3][7] (
	.clk(clk),
	.d(\Mux24~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_7_3),
	.prn(vcc));
defparam \r_array_out[3][7] .is_wysiwyg = "true";
defparam \r_array_out[3][7] .power_up = "low";

dffeas \i_array_out[3][7] (
	.clk(clk),
	.d(\Mux56~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_7_3),
	.prn(vcc));
defparam \i_array_out[3][7] .is_wysiwyg = "true";
defparam \i_array_out[3][7] .power_up = "low";

dffeas \r_array_out[0][6] (
	.clk(clk),
	.d(\Mux1~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_6_0),
	.prn(vcc));
defparam \r_array_out[0][6] .is_wysiwyg = "true";
defparam \r_array_out[0][6] .power_up = "low";

dffeas \i_array_out[0][6] (
	.clk(clk),
	.d(\Mux33~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_6_0),
	.prn(vcc));
defparam \i_array_out[0][6] .is_wysiwyg = "true";
defparam \i_array_out[0][6] .power_up = "low";

dffeas \r_array_out[1][6] (
	.clk(clk),
	.d(\Mux9~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_6_1),
	.prn(vcc));
defparam \r_array_out[1][6] .is_wysiwyg = "true";
defparam \r_array_out[1][6] .power_up = "low";

dffeas \i_array_out[1][6] (
	.clk(clk),
	.d(\Mux41~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_6_1),
	.prn(vcc));
defparam \i_array_out[1][6] .is_wysiwyg = "true";
defparam \i_array_out[1][6] .power_up = "low";

dffeas \r_array_out[2][6] (
	.clk(clk),
	.d(\Mux17~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_6_2),
	.prn(vcc));
defparam \r_array_out[2][6] .is_wysiwyg = "true";
defparam \r_array_out[2][6] .power_up = "low";

dffeas \i_array_out[2][6] (
	.clk(clk),
	.d(\Mux49~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_6_2),
	.prn(vcc));
defparam \i_array_out[2][6] .is_wysiwyg = "true";
defparam \i_array_out[2][6] .power_up = "low";

dffeas \r_array_out[3][6] (
	.clk(clk),
	.d(\Mux25~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_6_3),
	.prn(vcc));
defparam \r_array_out[3][6] .is_wysiwyg = "true";
defparam \r_array_out[3][6] .power_up = "low";

dffeas \i_array_out[3][6] (
	.clk(clk),
	.d(\Mux57~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_6_3),
	.prn(vcc));
defparam \i_array_out[3][6] .is_wysiwyg = "true";
defparam \i_array_out[3][6] .power_up = "low";

dffeas \i_array_out[2][1] (
	.clk(clk),
	.d(\Mux54~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_1_2),
	.prn(vcc));
defparam \i_array_out[2][1] .is_wysiwyg = "true";
defparam \i_array_out[2][1] .power_up = "low";

dffeas \i_array_out[1][1] (
	.clk(clk),
	.d(\Mux46~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_1_1),
	.prn(vcc));
defparam \i_array_out[1][1] .is_wysiwyg = "true";
defparam \i_array_out[1][1] .power_up = "low";

dffeas \i_array_out[0][1] (
	.clk(clk),
	.d(\Mux38~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_1_0),
	.prn(vcc));
defparam \i_array_out[0][1] .is_wysiwyg = "true";
defparam \i_array_out[0][1] .power_up = "low";

dffeas \i_array_out[3][1] (
	.clk(clk),
	.d(\Mux62~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_1_3),
	.prn(vcc));
defparam \i_array_out[3][1] .is_wysiwyg = "true";
defparam \i_array_out[3][1] .power_up = "low";

dffeas \i_array_out[2][0] (
	.clk(clk),
	.d(\Mux55~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_0_2),
	.prn(vcc));
defparam \i_array_out[2][0] .is_wysiwyg = "true";
defparam \i_array_out[2][0] .power_up = "low";

dffeas \i_array_out[1][0] (
	.clk(clk),
	.d(\Mux47~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_0_1),
	.prn(vcc));
defparam \i_array_out[1][0] .is_wysiwyg = "true";
defparam \i_array_out[1][0] .power_up = "low";

dffeas \i_array_out[0][0] (
	.clk(clk),
	.d(\Mux39~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_0_0),
	.prn(vcc));
defparam \i_array_out[0][0] .is_wysiwyg = "true";
defparam \i_array_out[0][0] .power_up = "low";

dffeas \i_array_out[3][0] (
	.clk(clk),
	.d(\Mux63~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_0_3),
	.prn(vcc));
defparam \i_array_out[3][0] .is_wysiwyg = "true";
defparam \i_array_out[3][0] .power_up = "low";

dffeas \r_array_out[2][1] (
	.clk(clk),
	.d(\Mux22~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_1_2),
	.prn(vcc));
defparam \r_array_out[2][1] .is_wysiwyg = "true";
defparam \r_array_out[2][1] .power_up = "low";

dffeas \r_array_out[1][1] (
	.clk(clk),
	.d(\Mux14~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_1_1),
	.prn(vcc));
defparam \r_array_out[1][1] .is_wysiwyg = "true";
defparam \r_array_out[1][1] .power_up = "low";

dffeas \r_array_out[0][1] (
	.clk(clk),
	.d(\Mux6~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_1_0),
	.prn(vcc));
defparam \r_array_out[0][1] .is_wysiwyg = "true";
defparam \r_array_out[0][1] .power_up = "low";

dffeas \r_array_out[3][1] (
	.clk(clk),
	.d(\Mux30~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_1_3),
	.prn(vcc));
defparam \r_array_out[3][1] .is_wysiwyg = "true";
defparam \r_array_out[3][1] .power_up = "low";

dffeas \r_array_out[2][0] (
	.clk(clk),
	.d(\Mux23~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_0_2),
	.prn(vcc));
defparam \r_array_out[2][0] .is_wysiwyg = "true";
defparam \r_array_out[2][0] .power_up = "low";

dffeas \r_array_out[1][0] (
	.clk(clk),
	.d(\Mux15~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_0_1),
	.prn(vcc));
defparam \r_array_out[1][0] .is_wysiwyg = "true";
defparam \r_array_out[1][0] .power_up = "low";

dffeas \r_array_out[0][0] (
	.clk(clk),
	.d(\Mux7~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_0_0),
	.prn(vcc));
defparam \r_array_out[0][0] .is_wysiwyg = "true";
defparam \r_array_out[0][0] .power_up = "low";

dffeas \r_array_out[3][0] (
	.clk(clk),
	.d(\Mux31~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_0_3),
	.prn(vcc));
defparam \r_array_out[3][0] .is_wysiwyg = "true";
defparam \r_array_out[3][0] .power_up = "low";

cycloneiii_lcell_comb \r_array_out[0][3]~0 (
	.dataa(do_tdl0031),
	.datab(do_tdl0030),
	.datac(gnd),
	.datad(slb_1pt_0),
	.cin(gnd),
	.combout(\r_array_out[0][3]~0_combout ),
	.cout());
defparam \r_array_out[0][3]~0 .lut_mask = 16'hAACC;
defparam \r_array_out[0][3]~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux1~1 (
	.dataa(do_tdl0032),
	.datab(do_tdl0033),
	.datac(slb_last_0),
	.datad(scale_dft_o_en),
	.cin(gnd),
	.combout(\Mux1~1_combout ),
	.cout());
defparam \Mux1~1 .lut_mask = 16'hEFFE;
defparam \Mux1~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \i_array_out[0][3]~0 (
	.dataa(do_tdl0131),
	.datab(do_tdl0130),
	.datac(gnd),
	.datad(slb_1pt_0),
	.cin(gnd),
	.combout(\i_array_out[0][3]~0_combout ),
	.cout());
defparam \i_array_out[0][3]~0 .lut_mask = 16'hAACC;
defparam \i_array_out[0][3]~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux33~1 (
	.dataa(do_tdl0132),
	.datab(do_tdl0133),
	.datac(slb_last_0),
	.datad(scale_dft_o_en),
	.cin(gnd),
	.combout(\Mux33~1_combout ),
	.cout());
defparam \Mux33~1 .lut_mask = 16'hEFFE;
defparam \Mux33~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \r_array_out[1][3]~1 (
	.dataa(do_tdl1031),
	.datab(do_tdl1030),
	.datac(gnd),
	.datad(slb_1pt_0),
	.cin(gnd),
	.combout(\r_array_out[1][3]~1_combout ),
	.cout());
defparam \r_array_out[1][3]~1 .lut_mask = 16'hAACC;
defparam \r_array_out[1][3]~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux9~1 (
	.dataa(do_tdl1032),
	.datab(do_tdl1033),
	.datac(slb_last_0),
	.datad(scale_dft_o_en),
	.cin(gnd),
	.combout(\Mux9~1_combout ),
	.cout());
defparam \Mux9~1 .lut_mask = 16'hEFFE;
defparam \Mux9~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \i_array_out[1][3]~1 (
	.dataa(do_tdl1131),
	.datab(do_tdl1130),
	.datac(gnd),
	.datad(slb_1pt_0),
	.cin(gnd),
	.combout(\i_array_out[1][3]~1_combout ),
	.cout());
defparam \i_array_out[1][3]~1 .lut_mask = 16'hAACC;
defparam \i_array_out[1][3]~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux41~1 (
	.dataa(do_tdl1132),
	.datab(do_tdl1133),
	.datac(slb_last_0),
	.datad(scale_dft_o_en),
	.cin(gnd),
	.combout(\Mux41~1_combout ),
	.cout());
defparam \Mux41~1 .lut_mask = 16'hEFFE;
defparam \Mux41~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \r_array_out[2][3]~2 (
	.dataa(do_tdl2031),
	.datab(do_tdl2030),
	.datac(gnd),
	.datad(slb_1pt_0),
	.cin(gnd),
	.combout(\r_array_out[2][3]~2_combout ),
	.cout());
defparam \r_array_out[2][3]~2 .lut_mask = 16'hAACC;
defparam \r_array_out[2][3]~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux17~1 (
	.dataa(do_tdl2032),
	.datab(do_tdl2033),
	.datac(slb_last_0),
	.datad(scale_dft_o_en),
	.cin(gnd),
	.combout(\Mux17~1_combout ),
	.cout());
defparam \Mux17~1 .lut_mask = 16'hEFFE;
defparam \Mux17~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \i_array_out[2][3]~2 (
	.dataa(do_tdl2131),
	.datab(do_tdl2130),
	.datac(gnd),
	.datad(slb_1pt_0),
	.cin(gnd),
	.combout(\i_array_out[2][3]~2_combout ),
	.cout());
defparam \i_array_out[2][3]~2 .lut_mask = 16'hAACC;
defparam \i_array_out[2][3]~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux49~1 (
	.dataa(do_tdl2132),
	.datab(do_tdl2133),
	.datac(slb_last_0),
	.datad(scale_dft_o_en),
	.cin(gnd),
	.combout(\Mux49~1_combout ),
	.cout());
defparam \Mux49~1 .lut_mask = 16'hEFFE;
defparam \Mux49~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \r_array_out[3][3]~3 (
	.dataa(do_tdl3031),
	.datab(do_tdl3030),
	.datac(gnd),
	.datad(slb_1pt_0),
	.cin(gnd),
	.combout(\r_array_out[3][3]~3_combout ),
	.cout());
defparam \r_array_out[3][3]~3 .lut_mask = 16'hAACC;
defparam \r_array_out[3][3]~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux25~1 (
	.dataa(do_tdl3032),
	.datab(do_tdl3033),
	.datac(slb_last_0),
	.datad(scale_dft_o_en),
	.cin(gnd),
	.combout(\Mux25~1_combout ),
	.cout());
defparam \Mux25~1 .lut_mask = 16'hEFFE;
defparam \Mux25~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \i_array_out[3][3]~3 (
	.dataa(do_tdl3131),
	.datab(do_tdl3130),
	.datac(gnd),
	.datad(slb_1pt_0),
	.cin(gnd),
	.combout(\i_array_out[3][3]~3_combout ),
	.cout());
defparam \i_array_out[3][3]~3 .lut_mask = 16'hAACC;
defparam \i_array_out[3][3]~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux57~1 (
	.dataa(do_tdl3132),
	.datab(do_tdl3133),
	.datac(slb_last_0),
	.datad(scale_dft_o_en),
	.cin(gnd),
	.combout(\Mux57~1_combout ),
	.cout());
defparam \Mux57~1 .lut_mask = 16'hEFFE;
defparam \Mux57~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \r_array_out[0][2]~14 (
	.dataa(do_tdl0032),
	.datab(do_tdl0031),
	.datac(slb_last_0),
	.datad(scale_dft_o_en),
	.cin(gnd),
	.combout(\r_array_out[0][2]~14_combout ),
	.cout());
defparam \r_array_out[0][2]~14 .lut_mask = 16'hEFFE;
defparam \r_array_out[0][2]~14 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux1~2 (
	.dataa(do_tdl0033),
	.datab(do_tdl0034),
	.datac(slb_last_0),
	.datad(scale_dft_o_en),
	.cin(gnd),
	.combout(\Mux1~2_combout ),
	.cout());
defparam \Mux1~2 .lut_mask = 16'hEFFE;
defparam \Mux1~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \r_array_out[0][4]~4 (
	.dataa(\r_array_out[0][2]~14_combout ),
	.datab(\Mux1~2_combout ),
	.datac(gnd),
	.datad(slb_1pt_1),
	.cin(gnd),
	.combout(\r_array_out[0][4]~4_combout ),
	.cout());
defparam \r_array_out[0][4]~4 .lut_mask = 16'hAACC;
defparam \r_array_out[0][4]~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \i_array_out[0][2]~14 (
	.dataa(do_tdl0132),
	.datab(do_tdl0131),
	.datac(gnd),
	.datad(slb_1pt_0),
	.cin(gnd),
	.combout(\i_array_out[0][2]~14_combout ),
	.cout());
defparam \i_array_out[0][2]~14 .lut_mask = 16'hAACC;
defparam \i_array_out[0][2]~14 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux33~2 (
	.dataa(do_tdl0133),
	.datab(do_tdl0134),
	.datac(slb_last_0),
	.datad(scale_dft_o_en),
	.cin(gnd),
	.combout(\Mux33~2_combout ),
	.cout());
defparam \Mux33~2 .lut_mask = 16'hEFFE;
defparam \Mux33~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \i_array_out[0][4]~4 (
	.dataa(\i_array_out[0][2]~14_combout ),
	.datab(\Mux33~2_combout ),
	.datac(gnd),
	.datad(slb_1pt_1),
	.cin(gnd),
	.combout(\i_array_out[0][4]~4_combout ),
	.cout());
defparam \i_array_out[0][4]~4 .lut_mask = 16'hAACC;
defparam \i_array_out[0][4]~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \r_array_out[1][2]~13 (
	.dataa(do_tdl1032),
	.datab(do_tdl1031),
	.datac(slb_last_0),
	.datad(scale_dft_o_en),
	.cin(gnd),
	.combout(\r_array_out[1][2]~13_combout ),
	.cout());
defparam \r_array_out[1][2]~13 .lut_mask = 16'hEFFE;
defparam \r_array_out[1][2]~13 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux9~2 (
	.dataa(do_tdl1033),
	.datab(do_tdl1034),
	.datac(slb_last_0),
	.datad(scale_dft_o_en),
	.cin(gnd),
	.combout(\Mux9~2_combout ),
	.cout());
defparam \Mux9~2 .lut_mask = 16'hEFFE;
defparam \Mux9~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \r_array_out[1][4]~5 (
	.dataa(\r_array_out[1][2]~13_combout ),
	.datab(\Mux9~2_combout ),
	.datac(gnd),
	.datad(slb_1pt_1),
	.cin(gnd),
	.combout(\r_array_out[1][4]~5_combout ),
	.cout());
defparam \r_array_out[1][4]~5 .lut_mask = 16'hAACC;
defparam \r_array_out[1][4]~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \i_array_out[1][2]~13 (
	.dataa(do_tdl1132),
	.datab(do_tdl1131),
	.datac(gnd),
	.datad(slb_1pt_0),
	.cin(gnd),
	.combout(\i_array_out[1][2]~13_combout ),
	.cout());
defparam \i_array_out[1][2]~13 .lut_mask = 16'hAACC;
defparam \i_array_out[1][2]~13 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux41~2 (
	.dataa(do_tdl1133),
	.datab(do_tdl1134),
	.datac(slb_last_0),
	.datad(scale_dft_o_en),
	.cin(gnd),
	.combout(\Mux41~2_combout ),
	.cout());
defparam \Mux41~2 .lut_mask = 16'hEFFE;
defparam \Mux41~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \i_array_out[1][4]~5 (
	.dataa(\i_array_out[1][2]~13_combout ),
	.datab(\Mux41~2_combout ),
	.datac(gnd),
	.datad(slb_1pt_1),
	.cin(gnd),
	.combout(\i_array_out[1][4]~5_combout ),
	.cout());
defparam \i_array_out[1][4]~5 .lut_mask = 16'hAACC;
defparam \i_array_out[1][4]~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \r_array_out[2][2]~12 (
	.dataa(do_tdl2032),
	.datab(do_tdl2031),
	.datac(gnd),
	.datad(slb_1pt_0),
	.cin(gnd),
	.combout(\r_array_out[2][2]~12_combout ),
	.cout());
defparam \r_array_out[2][2]~12 .lut_mask = 16'hAACC;
defparam \r_array_out[2][2]~12 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux17~2 (
	.dataa(do_tdl2033),
	.datab(do_tdl2034),
	.datac(slb_last_0),
	.datad(scale_dft_o_en),
	.cin(gnd),
	.combout(\Mux17~2_combout ),
	.cout());
defparam \Mux17~2 .lut_mask = 16'hEFFE;
defparam \Mux17~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \r_array_out[2][4]~6 (
	.dataa(\r_array_out[2][2]~12_combout ),
	.datab(\Mux17~2_combout ),
	.datac(gnd),
	.datad(slb_1pt_1),
	.cin(gnd),
	.combout(\r_array_out[2][4]~6_combout ),
	.cout());
defparam \r_array_out[2][4]~6 .lut_mask = 16'hAACC;
defparam \r_array_out[2][4]~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \i_array_out[2][2]~12 (
	.dataa(do_tdl2132),
	.datab(do_tdl2131),
	.datac(slb_last_0),
	.datad(scale_dft_o_en),
	.cin(gnd),
	.combout(\i_array_out[2][2]~12_combout ),
	.cout());
defparam \i_array_out[2][2]~12 .lut_mask = 16'hEFFE;
defparam \i_array_out[2][2]~12 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux49~2 (
	.dataa(do_tdl2133),
	.datab(do_tdl2134),
	.datac(slb_last_0),
	.datad(scale_dft_o_en),
	.cin(gnd),
	.combout(\Mux49~2_combout ),
	.cout());
defparam \Mux49~2 .lut_mask = 16'hEFFE;
defparam \Mux49~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \i_array_out[2][4]~6 (
	.dataa(\i_array_out[2][2]~12_combout ),
	.datab(\Mux49~2_combout ),
	.datac(gnd),
	.datad(slb_1pt_1),
	.cin(gnd),
	.combout(\i_array_out[2][4]~6_combout ),
	.cout());
defparam \i_array_out[2][4]~6 .lut_mask = 16'hAACC;
defparam \i_array_out[2][4]~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \r_array_out[3][2]~15 (
	.dataa(do_tdl3032),
	.datab(do_tdl3031),
	.datac(slb_last_0),
	.datad(scale_dft_o_en),
	.cin(gnd),
	.combout(\r_array_out[3][2]~15_combout ),
	.cout());
defparam \r_array_out[3][2]~15 .lut_mask = 16'hEFFE;
defparam \r_array_out[3][2]~15 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux25~2 (
	.dataa(do_tdl3033),
	.datab(do_tdl3034),
	.datac(slb_last_0),
	.datad(scale_dft_o_en),
	.cin(gnd),
	.combout(\Mux25~2_combout ),
	.cout());
defparam \Mux25~2 .lut_mask = 16'hEFFE;
defparam \Mux25~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \r_array_out[3][4]~7 (
	.dataa(\r_array_out[3][2]~15_combout ),
	.datab(\Mux25~2_combout ),
	.datac(gnd),
	.datad(slb_1pt_1),
	.cin(gnd),
	.combout(\r_array_out[3][4]~7_combout ),
	.cout());
defparam \r_array_out[3][4]~7 .lut_mask = 16'hAACC;
defparam \r_array_out[3][4]~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \i_array_out[3][2]~15 (
	.dataa(do_tdl3132),
	.datab(do_tdl3131),
	.datac(gnd),
	.datad(slb_1pt_0),
	.cin(gnd),
	.combout(\i_array_out[3][2]~15_combout ),
	.cout());
defparam \i_array_out[3][2]~15 .lut_mask = 16'hAACC;
defparam \i_array_out[3][2]~15 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux57~2 (
	.dataa(do_tdl3133),
	.datab(do_tdl3134),
	.datac(slb_last_0),
	.datad(scale_dft_o_en),
	.cin(gnd),
	.combout(\Mux57~2_combout ),
	.cout());
defparam \Mux57~2 .lut_mask = 16'hEFFE;
defparam \Mux57~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \i_array_out[3][4]~7 (
	.dataa(\i_array_out[3][2]~15_combout ),
	.datab(\Mux57~2_combout ),
	.datac(gnd),
	.datad(slb_1pt_1),
	.cin(gnd),
	.combout(\i_array_out[3][4]~7_combout ),
	.cout());
defparam \i_array_out[3][4]~7 .lut_mask = 16'hAACC;
defparam \i_array_out[3][4]~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux1~0 (
	.dataa(do_tdl0034),
	.datab(do_tdl0035),
	.datac(slb_last_0),
	.datad(scale_dft_o_en),
	.cin(gnd),
	.combout(\Mux1~0_combout ),
	.cout());
defparam \Mux1~0 .lut_mask = 16'hEFFE;
defparam \Mux1~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \r_array_out[0][5]~8 (
	.dataa(\Mux1~1_combout ),
	.datab(\Mux1~0_combout ),
	.datac(gnd),
	.datad(slb_1pt_1),
	.cin(gnd),
	.combout(\r_array_out[0][5]~8_combout ),
	.cout());
defparam \r_array_out[0][5]~8 .lut_mask = 16'hAACC;
defparam \r_array_out[0][5]~8 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux33~0 (
	.dataa(do_tdl0134),
	.datab(do_tdl0135),
	.datac(slb_last_0),
	.datad(scale_dft_o_en),
	.cin(gnd),
	.combout(\Mux33~0_combout ),
	.cout());
defparam \Mux33~0 .lut_mask = 16'hEFFE;
defparam \Mux33~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \i_array_out[0][5]~8 (
	.dataa(\Mux33~1_combout ),
	.datab(\Mux33~0_combout ),
	.datac(gnd),
	.datad(slb_1pt_1),
	.cin(gnd),
	.combout(\i_array_out[0][5]~8_combout ),
	.cout());
defparam \i_array_out[0][5]~8 .lut_mask = 16'hAACC;
defparam \i_array_out[0][5]~8 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux9~0 (
	.dataa(do_tdl1034),
	.datab(do_tdl1035),
	.datac(slb_last_0),
	.datad(scale_dft_o_en),
	.cin(gnd),
	.combout(\Mux9~0_combout ),
	.cout());
defparam \Mux9~0 .lut_mask = 16'hEFFE;
defparam \Mux9~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \r_array_out[1][5]~9 (
	.dataa(\Mux9~1_combout ),
	.datab(\Mux9~0_combout ),
	.datac(gnd),
	.datad(slb_1pt_1),
	.cin(gnd),
	.combout(\r_array_out[1][5]~9_combout ),
	.cout());
defparam \r_array_out[1][5]~9 .lut_mask = 16'hAACC;
defparam \r_array_out[1][5]~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux41~0 (
	.dataa(do_tdl1134),
	.datab(do_tdl1135),
	.datac(slb_last_0),
	.datad(scale_dft_o_en),
	.cin(gnd),
	.combout(\Mux41~0_combout ),
	.cout());
defparam \Mux41~0 .lut_mask = 16'hEFFE;
defparam \Mux41~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \i_array_out[1][5]~9 (
	.dataa(\Mux41~1_combout ),
	.datab(\Mux41~0_combout ),
	.datac(gnd),
	.datad(slb_1pt_1),
	.cin(gnd),
	.combout(\i_array_out[1][5]~9_combout ),
	.cout());
defparam \i_array_out[1][5]~9 .lut_mask = 16'hAACC;
defparam \i_array_out[1][5]~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux17~0 (
	.dataa(do_tdl2034),
	.datab(do_tdl2035),
	.datac(slb_last_0),
	.datad(scale_dft_o_en),
	.cin(gnd),
	.combout(\Mux17~0_combout ),
	.cout());
defparam \Mux17~0 .lut_mask = 16'hEFFE;
defparam \Mux17~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \r_array_out[2][5]~10 (
	.dataa(\Mux17~1_combout ),
	.datab(\Mux17~0_combout ),
	.datac(gnd),
	.datad(slb_1pt_1),
	.cin(gnd),
	.combout(\r_array_out[2][5]~10_combout ),
	.cout());
defparam \r_array_out[2][5]~10 .lut_mask = 16'hAACC;
defparam \r_array_out[2][5]~10 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux49~0 (
	.dataa(do_tdl2134),
	.datab(do_tdl2135),
	.datac(slb_last_0),
	.datad(scale_dft_o_en),
	.cin(gnd),
	.combout(\Mux49~0_combout ),
	.cout());
defparam \Mux49~0 .lut_mask = 16'hEFFE;
defparam \Mux49~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \i_array_out[2][5]~10 (
	.dataa(\Mux49~1_combout ),
	.datab(\Mux49~0_combout ),
	.datac(gnd),
	.datad(slb_1pt_1),
	.cin(gnd),
	.combout(\i_array_out[2][5]~10_combout ),
	.cout());
defparam \i_array_out[2][5]~10 .lut_mask = 16'hAACC;
defparam \i_array_out[2][5]~10 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux25~0 (
	.dataa(do_tdl3034),
	.datab(do_tdl3035),
	.datac(slb_last_0),
	.datad(scale_dft_o_en),
	.cin(gnd),
	.combout(\Mux25~0_combout ),
	.cout());
defparam \Mux25~0 .lut_mask = 16'hEFFE;
defparam \Mux25~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \r_array_out[3][5]~11 (
	.dataa(\Mux25~1_combout ),
	.datab(\Mux25~0_combout ),
	.datac(gnd),
	.datad(slb_1pt_1),
	.cin(gnd),
	.combout(\r_array_out[3][5]~11_combout ),
	.cout());
defparam \r_array_out[3][5]~11 .lut_mask = 16'hAACC;
defparam \r_array_out[3][5]~11 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux57~0 (
	.dataa(do_tdl3134),
	.datab(do_tdl3135),
	.datac(slb_last_0),
	.datad(scale_dft_o_en),
	.cin(gnd),
	.combout(\Mux57~0_combout ),
	.cout());
defparam \Mux57~0 .lut_mask = 16'hEFFE;
defparam \Mux57~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \i_array_out[3][5]~11 (
	.dataa(\Mux57~1_combout ),
	.datab(\Mux57~0_combout ),
	.datac(gnd),
	.datad(slb_1pt_1),
	.cin(gnd),
	.combout(\i_array_out[3][5]~11_combout ),
	.cout());
defparam \i_array_out[3][5]~11 .lut_mask = 16'hAACC;
defparam \i_array_out[3][5]~11 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux49~5 (
	.dataa(do_tdl2130),
	.datab(gnd),
	.datac(slb_last_0),
	.datad(scale_dft_o_en),
	.cin(gnd),
	.combout(\Mux49~5_combout ),
	.cout());
defparam \Mux49~5 .lut_mask = 16'hAFFF;
defparam \Mux49~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux41~5 (
	.dataa(do_tdl1130),
	.datab(gnd),
	.datac(slb_last_0),
	.datad(scale_dft_o_en),
	.cin(gnd),
	.combout(\Mux41~5_combout ),
	.cout());
defparam \Mux41~5 .lut_mask = 16'hAFFF;
defparam \Mux41~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux33~5 (
	.dataa(do_tdl0130),
	.datab(gnd),
	.datac(slb_last_0),
	.datad(scale_dft_o_en),
	.cin(gnd),
	.combout(\Mux33~5_combout ),
	.cout());
defparam \Mux33~5 .lut_mask = 16'hAFFF;
defparam \Mux33~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux57~5 (
	.dataa(do_tdl3130),
	.datab(gnd),
	.datac(slb_last_0),
	.datad(scale_dft_o_en),
	.cin(gnd),
	.combout(\Mux57~5_combout ),
	.cout());
defparam \Mux57~5 .lut_mask = 16'hAFFF;
defparam \Mux57~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux17~5 (
	.dataa(do_tdl2030),
	.datab(gnd),
	.datac(slb_last_0),
	.datad(scale_dft_o_en),
	.cin(gnd),
	.combout(\Mux17~5_combout ),
	.cout());
defparam \Mux17~5 .lut_mask = 16'hAFFF;
defparam \Mux17~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux9~5 (
	.dataa(do_tdl1030),
	.datab(gnd),
	.datac(slb_last_0),
	.datad(scale_dft_o_en),
	.cin(gnd),
	.combout(\Mux9~5_combout ),
	.cout());
defparam \Mux9~5 .lut_mask = 16'hAFFF;
defparam \Mux9~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux1~5 (
	.dataa(do_tdl0030),
	.datab(gnd),
	.datac(slb_last_0),
	.datad(scale_dft_o_en),
	.cin(gnd),
	.combout(\Mux1~5_combout ),
	.cout());
defparam \Mux1~5 .lut_mask = 16'hAFFF;
defparam \Mux1~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux25~5 (
	.dataa(do_tdl3030),
	.datab(gnd),
	.datac(slb_last_0),
	.datad(scale_dft_o_en),
	.cin(gnd),
	.combout(\Mux25~5_combout ),
	.cout());
defparam \Mux25~5 .lut_mask = 16'hAFFF;
defparam \Mux25~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \i_array_out[0][6]~16 (
	.dataa(scale_dft_o_en),
	.datab(slb_last_2),
	.datac(slb_last_0),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\i_array_out[0][6]~16_combout ),
	.cout());
defparam \i_array_out[0][6]~16 .lut_mask = 16'hFEFF;
defparam \i_array_out[0][6]~16 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \i_array_out[0][6]~17 (
	.dataa(scale_dft_o_en),
	.datab(slb_last_1),
	.datac(slb_last_2),
	.datad(gnd),
	.cin(gnd),
	.combout(\i_array_out[0][6]~17_combout ),
	.cout());
defparam \i_array_out[0][6]~17 .lut_mask = 16'hFEFE;
defparam \i_array_out[0][6]~17 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux0~0 (
	.dataa(\i_array_out[0][6]~16_combout ),
	.datab(do_tdl0037),
	.datac(\i_array_out[0][6]~17_combout ),
	.datad(\Mux1~0_combout ),
	.cin(gnd),
	.combout(\Mux0~0_combout ),
	.cout());
defparam \Mux0~0 .lut_mask = 16'hFFDE;
defparam \Mux0~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux0~1 (
	.dataa(do_tdl0033),
	.datab(\i_array_out[0][6]~16_combout ),
	.datac(\Mux0~0_combout ),
	.datad(do_tdl0036),
	.cin(gnd),
	.combout(\Mux0~1_combout ),
	.cout());
defparam \Mux0~1 .lut_mask = 16'hFFBE;
defparam \Mux0~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux32~0 (
	.dataa(\i_array_out[0][6]~16_combout ),
	.datab(do_tdl0137),
	.datac(\i_array_out[0][6]~17_combout ),
	.datad(\Mux33~0_combout ),
	.cin(gnd),
	.combout(\Mux32~0_combout ),
	.cout());
defparam \Mux32~0 .lut_mask = 16'hFFDE;
defparam \Mux32~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux32~1 (
	.dataa(do_tdl0133),
	.datab(\i_array_out[0][6]~16_combout ),
	.datac(\Mux32~0_combout ),
	.datad(do_tdl0136),
	.cin(gnd),
	.combout(\Mux32~1_combout ),
	.cout());
defparam \Mux32~1 .lut_mask = 16'hFFBE;
defparam \Mux32~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux8~0 (
	.dataa(\i_array_out[0][6]~16_combout ),
	.datab(do_tdl1037),
	.datac(\i_array_out[0][6]~17_combout ),
	.datad(\Mux9~0_combout ),
	.cin(gnd),
	.combout(\Mux8~0_combout ),
	.cout());
defparam \Mux8~0 .lut_mask = 16'hFFDE;
defparam \Mux8~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux8~1 (
	.dataa(do_tdl1033),
	.datab(\i_array_out[0][6]~16_combout ),
	.datac(\Mux8~0_combout ),
	.datad(do_tdl1036),
	.cin(gnd),
	.combout(\Mux8~1_combout ),
	.cout());
defparam \Mux8~1 .lut_mask = 16'hFFBE;
defparam \Mux8~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux40~0 (
	.dataa(\i_array_out[0][6]~16_combout ),
	.datab(do_tdl1137),
	.datac(\i_array_out[0][6]~17_combout ),
	.datad(\Mux41~0_combout ),
	.cin(gnd),
	.combout(\Mux40~0_combout ),
	.cout());
defparam \Mux40~0 .lut_mask = 16'hFFDE;
defparam \Mux40~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux40~1 (
	.dataa(do_tdl1133),
	.datab(\i_array_out[0][6]~16_combout ),
	.datac(\Mux40~0_combout ),
	.datad(do_tdl1136),
	.cin(gnd),
	.combout(\Mux40~1_combout ),
	.cout());
defparam \Mux40~1 .lut_mask = 16'hFFBE;
defparam \Mux40~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux16~0 (
	.dataa(\i_array_out[0][6]~16_combout ),
	.datab(do_tdl2037),
	.datac(\i_array_out[0][6]~17_combout ),
	.datad(\Mux17~0_combout ),
	.cin(gnd),
	.combout(\Mux16~0_combout ),
	.cout());
defparam \Mux16~0 .lut_mask = 16'hFFDE;
defparam \Mux16~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux16~1 (
	.dataa(do_tdl2033),
	.datab(\i_array_out[0][6]~16_combout ),
	.datac(\Mux16~0_combout ),
	.datad(do_tdl2036),
	.cin(gnd),
	.combout(\Mux16~1_combout ),
	.cout());
defparam \Mux16~1 .lut_mask = 16'hFFBE;
defparam \Mux16~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux48~0 (
	.dataa(\i_array_out[0][6]~16_combout ),
	.datab(do_tdl2137),
	.datac(\i_array_out[0][6]~17_combout ),
	.datad(\Mux49~0_combout ),
	.cin(gnd),
	.combout(\Mux48~0_combout ),
	.cout());
defparam \Mux48~0 .lut_mask = 16'hFFDE;
defparam \Mux48~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux48~1 (
	.dataa(do_tdl2133),
	.datab(\i_array_out[0][6]~16_combout ),
	.datac(\Mux48~0_combout ),
	.datad(do_tdl2136),
	.cin(gnd),
	.combout(\Mux48~1_combout ),
	.cout());
defparam \Mux48~1 .lut_mask = 16'hFFBE;
defparam \Mux48~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux24~0 (
	.dataa(\i_array_out[0][6]~16_combout ),
	.datab(do_tdl3037),
	.datac(\i_array_out[0][6]~17_combout ),
	.datad(\Mux25~0_combout ),
	.cin(gnd),
	.combout(\Mux24~0_combout ),
	.cout());
defparam \Mux24~0 .lut_mask = 16'hFFDE;
defparam \Mux24~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux24~1 (
	.dataa(do_tdl3033),
	.datab(\i_array_out[0][6]~16_combout ),
	.datac(\Mux24~0_combout ),
	.datad(do_tdl3036),
	.cin(gnd),
	.combout(\Mux24~1_combout ),
	.cout());
defparam \Mux24~1 .lut_mask = 16'hFFBE;
defparam \Mux24~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux56~0 (
	.dataa(\i_array_out[0][6]~16_combout ),
	.datab(do_tdl3137),
	.datac(\i_array_out[0][6]~17_combout ),
	.datad(\Mux57~0_combout ),
	.cin(gnd),
	.combout(\Mux56~0_combout ),
	.cout());
defparam \Mux56~0 .lut_mask = 16'hFFDE;
defparam \Mux56~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux56~1 (
	.dataa(do_tdl3133),
	.datab(\i_array_out[0][6]~16_combout ),
	.datac(\Mux56~0_combout ),
	.datad(do_tdl3136),
	.cin(gnd),
	.combout(\Mux56~1_combout ),
	.cout());
defparam \Mux56~1 .lut_mask = 16'hFFBE;
defparam \Mux56~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux1~3 (
	.dataa(\i_array_out[0][6]~16_combout ),
	.datab(do_tdl0036),
	.datac(\i_array_out[0][6]~17_combout ),
	.datad(\Mux1~2_combout ),
	.cin(gnd),
	.combout(\Mux1~3_combout ),
	.cout());
defparam \Mux1~3 .lut_mask = 16'hFFDE;
defparam \Mux1~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux1~4 (
	.dataa(do_tdl0032),
	.datab(\i_array_out[0][6]~16_combout ),
	.datac(\Mux1~3_combout ),
	.datad(do_tdl0035),
	.cin(gnd),
	.combout(\Mux1~4_combout ),
	.cout());
defparam \Mux1~4 .lut_mask = 16'hFFBE;
defparam \Mux1~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux33~3 (
	.dataa(\i_array_out[0][6]~16_combout ),
	.datab(do_tdl0136),
	.datac(\i_array_out[0][6]~17_combout ),
	.datad(\Mux33~2_combout ),
	.cin(gnd),
	.combout(\Mux33~3_combout ),
	.cout());
defparam \Mux33~3 .lut_mask = 16'hFFDE;
defparam \Mux33~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux33~4 (
	.dataa(do_tdl0132),
	.datab(\i_array_out[0][6]~16_combout ),
	.datac(\Mux33~3_combout ),
	.datad(do_tdl0135),
	.cin(gnd),
	.combout(\Mux33~4_combout ),
	.cout());
defparam \Mux33~4 .lut_mask = 16'hFFBE;
defparam \Mux33~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux9~3 (
	.dataa(\i_array_out[0][6]~16_combout ),
	.datab(do_tdl1036),
	.datac(\i_array_out[0][6]~17_combout ),
	.datad(\Mux9~2_combout ),
	.cin(gnd),
	.combout(\Mux9~3_combout ),
	.cout());
defparam \Mux9~3 .lut_mask = 16'hFFDE;
defparam \Mux9~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux9~4 (
	.dataa(do_tdl1032),
	.datab(\i_array_out[0][6]~16_combout ),
	.datac(\Mux9~3_combout ),
	.datad(do_tdl1035),
	.cin(gnd),
	.combout(\Mux9~4_combout ),
	.cout());
defparam \Mux9~4 .lut_mask = 16'hFFBE;
defparam \Mux9~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux41~3 (
	.dataa(\i_array_out[0][6]~16_combout ),
	.datab(do_tdl1136),
	.datac(\i_array_out[0][6]~17_combout ),
	.datad(\Mux41~2_combout ),
	.cin(gnd),
	.combout(\Mux41~3_combout ),
	.cout());
defparam \Mux41~3 .lut_mask = 16'hFFDE;
defparam \Mux41~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux41~4 (
	.dataa(do_tdl1132),
	.datab(\i_array_out[0][6]~16_combout ),
	.datac(\Mux41~3_combout ),
	.datad(do_tdl1135),
	.cin(gnd),
	.combout(\Mux41~4_combout ),
	.cout());
defparam \Mux41~4 .lut_mask = 16'hFFBE;
defparam \Mux41~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux17~3 (
	.dataa(\i_array_out[0][6]~16_combout ),
	.datab(do_tdl2036),
	.datac(\i_array_out[0][6]~17_combout ),
	.datad(\Mux17~2_combout ),
	.cin(gnd),
	.combout(\Mux17~3_combout ),
	.cout());
defparam \Mux17~3 .lut_mask = 16'hFFDE;
defparam \Mux17~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux17~4 (
	.dataa(do_tdl2032),
	.datab(\i_array_out[0][6]~16_combout ),
	.datac(\Mux17~3_combout ),
	.datad(do_tdl2035),
	.cin(gnd),
	.combout(\Mux17~4_combout ),
	.cout());
defparam \Mux17~4 .lut_mask = 16'hFFBE;
defparam \Mux17~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux49~3 (
	.dataa(\i_array_out[0][6]~17_combout ),
	.datab(do_tdl2132),
	.datac(\i_array_out[0][6]~16_combout ),
	.datad(\Mux49~2_combout ),
	.cin(gnd),
	.combout(\Mux49~3_combout ),
	.cout());
defparam \Mux49~3 .lut_mask = 16'hFFDE;
defparam \Mux49~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux49~4 (
	.dataa(do_tdl2136),
	.datab(\i_array_out[0][6]~17_combout ),
	.datac(\Mux49~3_combout ),
	.datad(do_tdl2135),
	.cin(gnd),
	.combout(\Mux49~4_combout ),
	.cout());
defparam \Mux49~4 .lut_mask = 16'hFFBE;
defparam \Mux49~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux25~3 (
	.dataa(\i_array_out[0][6]~17_combout ),
	.datab(do_tdl3032),
	.datac(\i_array_out[0][6]~16_combout ),
	.datad(\Mux25~2_combout ),
	.cin(gnd),
	.combout(\Mux25~3_combout ),
	.cout());
defparam \Mux25~3 .lut_mask = 16'hFFDE;
defparam \Mux25~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux25~4 (
	.dataa(do_tdl3036),
	.datab(\i_array_out[0][6]~17_combout ),
	.datac(\Mux25~3_combout ),
	.datad(do_tdl3035),
	.cin(gnd),
	.combout(\Mux25~4_combout ),
	.cout());
defparam \Mux25~4 .lut_mask = 16'hFFBE;
defparam \Mux25~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux57~3 (
	.dataa(\i_array_out[0][6]~17_combout ),
	.datab(do_tdl3132),
	.datac(\i_array_out[0][6]~16_combout ),
	.datad(\Mux57~2_combout ),
	.cin(gnd),
	.combout(\Mux57~3_combout ),
	.cout());
defparam \Mux57~3 .lut_mask = 16'hFFDE;
defparam \Mux57~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux57~4 (
	.dataa(do_tdl3136),
	.datab(\i_array_out[0][6]~17_combout ),
	.datac(\Mux57~3_combout ),
	.datad(do_tdl3135),
	.cin(gnd),
	.combout(\Mux57~4_combout ),
	.cout());
defparam \Mux57~4 .lut_mask = 16'hFFBE;
defparam \Mux57~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux54~2 (
	.dataa(scale_dft_o_en),
	.datab(slb_last_1),
	.datac(slb_last_2),
	.datad(\i_array_out[2][3]~2_combout ),
	.cin(gnd),
	.combout(\Mux54~2_combout ),
	.cout());
defparam \Mux54~2 .lut_mask = 16'hFF7F;
defparam \Mux54~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux46~2 (
	.dataa(scale_dft_o_en),
	.datab(slb_last_1),
	.datac(slb_last_2),
	.datad(\i_array_out[1][3]~1_combout ),
	.cin(gnd),
	.combout(\Mux46~2_combout ),
	.cout());
defparam \Mux46~2 .lut_mask = 16'hFF7F;
defparam \Mux46~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux38~2 (
	.dataa(scale_dft_o_en),
	.datab(slb_last_1),
	.datac(slb_last_2),
	.datad(\i_array_out[0][3]~0_combout ),
	.cin(gnd),
	.combout(\Mux38~2_combout ),
	.cout());
defparam \Mux38~2 .lut_mask = 16'hFF7F;
defparam \Mux38~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux62~2 (
	.dataa(scale_dft_o_en),
	.datab(slb_last_1),
	.datac(slb_last_2),
	.datad(\i_array_out[3][3]~3_combout ),
	.cin(gnd),
	.combout(\Mux62~2_combout ),
	.cout());
defparam \Mux62~2 .lut_mask = 16'hFF7F;
defparam \Mux62~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux7~0 (
	.dataa(scale_dft_o_en),
	.datab(slb_last_0),
	.datac(slb_last_1),
	.datad(slb_last_2),
	.cin(gnd),
	.combout(\Mux7~0_combout ),
	.cout());
defparam \Mux7~0 .lut_mask = 16'hFFFE;
defparam \Mux7~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux55~0 (
	.dataa(do_tdl2130),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mux7~0_combout ),
	.cin(gnd),
	.combout(\Mux55~0_combout ),
	.cout());
defparam \Mux55~0 .lut_mask = 16'hAAFF;
defparam \Mux55~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux47~0 (
	.dataa(do_tdl1130),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mux7~0_combout ),
	.cin(gnd),
	.combout(\Mux47~0_combout ),
	.cout());
defparam \Mux47~0 .lut_mask = 16'hAAFF;
defparam \Mux47~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux39~0 (
	.dataa(do_tdl0130),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mux7~0_combout ),
	.cin(gnd),
	.combout(\Mux39~0_combout ),
	.cout());
defparam \Mux39~0 .lut_mask = 16'hAAFF;
defparam \Mux39~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux63~0 (
	.dataa(do_tdl3130),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mux7~0_combout ),
	.cin(gnd),
	.combout(\Mux63~0_combout ),
	.cout());
defparam \Mux63~0 .lut_mask = 16'hAAFF;
defparam \Mux63~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux22~2 (
	.dataa(scale_dft_o_en),
	.datab(slb_last_1),
	.datac(slb_last_2),
	.datad(\r_array_out[2][3]~2_combout ),
	.cin(gnd),
	.combout(\Mux22~2_combout ),
	.cout());
defparam \Mux22~2 .lut_mask = 16'hFF7F;
defparam \Mux22~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux14~2 (
	.dataa(scale_dft_o_en),
	.datab(slb_last_1),
	.datac(slb_last_2),
	.datad(\r_array_out[1][3]~1_combout ),
	.cin(gnd),
	.combout(\Mux14~2_combout ),
	.cout());
defparam \Mux14~2 .lut_mask = 16'hFF7F;
defparam \Mux14~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux6~2 (
	.dataa(scale_dft_o_en),
	.datab(slb_last_1),
	.datac(slb_last_2),
	.datad(\r_array_out[0][3]~0_combout ),
	.cin(gnd),
	.combout(\Mux6~2_combout ),
	.cout());
defparam \Mux6~2 .lut_mask = 16'hFF7F;
defparam \Mux6~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux30~2 (
	.dataa(scale_dft_o_en),
	.datab(slb_last_1),
	.datac(slb_last_2),
	.datad(\r_array_out[3][3]~3_combout ),
	.cin(gnd),
	.combout(\Mux30~2_combout ),
	.cout());
defparam \Mux30~2 .lut_mask = 16'hFF7F;
defparam \Mux30~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux23~0 (
	.dataa(do_tdl2030),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mux7~0_combout ),
	.cin(gnd),
	.combout(\Mux23~0_combout ),
	.cout());
defparam \Mux23~0 .lut_mask = 16'hAAFF;
defparam \Mux23~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux15~0 (
	.dataa(do_tdl1030),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mux7~0_combout ),
	.cin(gnd),
	.combout(\Mux15~0_combout ),
	.cout());
defparam \Mux15~0 .lut_mask = 16'hAAFF;
defparam \Mux15~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux7~1 (
	.dataa(do_tdl0030),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mux7~0_combout ),
	.cin(gnd),
	.combout(\Mux7~1_combout ),
	.cout());
defparam \Mux7~1 .lut_mask = 16'hAAFF;
defparam \Mux7~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux31~0 (
	.dataa(do_tdl3030),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mux7~0_combout ),
	.cin(gnd),
	.combout(\Mux31~0_combout ),
	.cout());
defparam \Mux31~0 .lut_mask = 16'hAAFF;
defparam \Mux31~0 .sum_lutc_input = "datac";

endmodule

module fft_asj_fft_bfp_o_1pt_fft_120 (
	r_array_out_3_0,
	i_array_out_3_0,
	r_array_out_3_1,
	i_array_out_3_1,
	r_array_out_3_2,
	i_array_out_3_2,
	r_array_out_3_3,
	i_array_out_3_3,
	r_array_out_4_0,
	i_array_out_4_0,
	r_array_out_4_1,
	i_array_out_4_1,
	r_array_out_4_2,
	i_array_out_4_2,
	r_array_out_4_3,
	i_array_out_4_3,
	r_array_out_5_0,
	i_array_out_5_0,
	r_array_out_5_1,
	i_array_out_5_1,
	r_array_out_5_2,
	i_array_out_5_2,
	r_array_out_5_3,
	i_array_out_5_3,
	global_clock_enable,
	gain_lut_8pts_0,
	gain_lut_8pts_1,
	gain_lut_8pts_2,
	gain_lut_8pts_3,
	enable_op,
	r_array_out_7_0,
	i_array_out_7_0,
	r_array_out_7_1,
	i_array_out_7_1,
	r_array_out_7_2,
	i_array_out_7_2,
	r_array_out_7_3,
	i_array_out_7_3,
	r_array_out_6_0,
	i_array_out_6_0,
	r_array_out_6_1,
	i_array_out_6_1,
	r_array_out_6_2,
	i_array_out_6_2,
	r_array_out_6_3,
	i_array_out_6_3,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	r_array_out_3_0;
input 	i_array_out_3_0;
input 	r_array_out_3_1;
input 	i_array_out_3_1;
input 	r_array_out_3_2;
input 	i_array_out_3_2;
input 	r_array_out_3_3;
input 	i_array_out_3_3;
input 	r_array_out_4_0;
input 	i_array_out_4_0;
input 	r_array_out_4_1;
input 	i_array_out_4_1;
input 	r_array_out_4_2;
input 	i_array_out_4_2;
input 	r_array_out_4_3;
input 	i_array_out_4_3;
input 	r_array_out_5_0;
input 	i_array_out_5_0;
input 	r_array_out_5_1;
input 	i_array_out_5_1;
input 	r_array_out_5_2;
input 	i_array_out_5_2;
input 	r_array_out_5_3;
input 	i_array_out_5_3;
input 	global_clock_enable;
output 	gain_lut_8pts_0;
output 	gain_lut_8pts_1;
output 	gain_lut_8pts_2;
output 	gain_lut_8pts_3;
input 	enable_op;
input 	r_array_out_7_0;
input 	i_array_out_7_0;
input 	r_array_out_7_1;
input 	i_array_out_7_1;
input 	r_array_out_7_2;
input 	i_array_out_7_2;
input 	r_array_out_7_3;
input 	i_array_out_7_3;
input 	r_array_out_6_0;
input 	i_array_out_6_0;
input 	r_array_out_6_1;
input 	i_array_out_6_1;
input 	r_array_out_6_2;
input 	i_array_out_6_2;
input 	r_array_out_6_3;
input 	i_array_out_6_3;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \gain_lut_8pts~0_combout ;
wire \gain_lut_8pts~6_combout ;
wire \gain_lut_8pts~12_combout ;
wire \gain_lut_8pts~18_combout ;
wire \gain_lut_8pts~1_combout ;
wire \gain_lut_8pts~2_combout ;
wire \gain_lut_8pts~3_combout ;
wire \gain_lut_8pts~4_combout ;
wire \gain_lut_8pts~5_combout ;
wire \gain_lut_8pts~7_combout ;
wire \gain_lut_8pts~8_combout ;
wire \gain_lut_8pts~9_combout ;
wire \gain_lut_8pts~10_combout ;
wire \gain_lut_8pts~11_combout ;
wire \gain_lut_8pts~13_combout ;
wire \gain_lut_8pts~14_combout ;
wire \gain_lut_8pts~15_combout ;
wire \gain_lut_8pts~16_combout ;
wire \gain_lut_8pts~17_combout ;
wire \gain_lut_8pts~19_combout ;
wire \gain_lut_8pts~20_combout ;
wire \gain_lut_8pts~21_combout ;
wire \gain_lut_8pts~22_combout ;
wire \gain_lut_8pts~23_combout ;


cycloneiii_lcell_comb \gain_lut_8pts~0 (
	.dataa(r_array_out_7_0),
	.datab(r_array_out_3_0),
	.datac(i_array_out_7_0),
	.datad(i_array_out_3_0),
	.cin(gnd),
	.combout(\gain_lut_8pts~0_combout ),
	.cout());
defparam \gain_lut_8pts~0 .lut_mask = 16'h6996;
defparam \gain_lut_8pts~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \gain_lut_8pts~6 (
	.dataa(r_array_out_7_0),
	.datab(r_array_out_4_0),
	.datac(i_array_out_7_0),
	.datad(i_array_out_4_0),
	.cin(gnd),
	.combout(\gain_lut_8pts~6_combout ),
	.cout());
defparam \gain_lut_8pts~6 .lut_mask = 16'h6996;
defparam \gain_lut_8pts~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \gain_lut_8pts~12 (
	.dataa(r_array_out_7_0),
	.datab(r_array_out_5_0),
	.datac(i_array_out_7_0),
	.datad(i_array_out_5_0),
	.cin(gnd),
	.combout(\gain_lut_8pts~12_combout ),
	.cout());
defparam \gain_lut_8pts~12 .lut_mask = 16'h6996;
defparam \gain_lut_8pts~12 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \gain_lut_8pts~18 (
	.dataa(r_array_out_7_0),
	.datab(r_array_out_6_0),
	.datac(i_array_out_7_0),
	.datad(i_array_out_6_0),
	.cin(gnd),
	.combout(\gain_lut_8pts~18_combout ),
	.cout());
defparam \gain_lut_8pts~18 .lut_mask = 16'h6996;
defparam \gain_lut_8pts~18 .sum_lutc_input = "datac";

dffeas \gain_lut_8pts[0] (
	.clk(clk),
	.d(\gain_lut_8pts~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(gain_lut_8pts_0),
	.prn(vcc));
defparam \gain_lut_8pts[0] .is_wysiwyg = "true";
defparam \gain_lut_8pts[0] .power_up = "low";

dffeas \gain_lut_8pts[1] (
	.clk(clk),
	.d(\gain_lut_8pts~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(gain_lut_8pts_1),
	.prn(vcc));
defparam \gain_lut_8pts[1] .is_wysiwyg = "true";
defparam \gain_lut_8pts[1] .power_up = "low";

dffeas \gain_lut_8pts[2] (
	.clk(clk),
	.d(\gain_lut_8pts~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(gain_lut_8pts_2),
	.prn(vcc));
defparam \gain_lut_8pts[2] .is_wysiwyg = "true";
defparam \gain_lut_8pts[2] .power_up = "low";

dffeas \gain_lut_8pts[3] (
	.clk(clk),
	.d(\gain_lut_8pts~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(gain_lut_8pts_3),
	.prn(vcc));
defparam \gain_lut_8pts[3] .is_wysiwyg = "true";
defparam \gain_lut_8pts[3] .power_up = "low";

cycloneiii_lcell_comb \gain_lut_8pts~1 (
	.dataa(r_array_out_7_1),
	.datab(r_array_out_3_1),
	.datac(i_array_out_7_1),
	.datad(i_array_out_3_1),
	.cin(gnd),
	.combout(\gain_lut_8pts~1_combout ),
	.cout());
defparam \gain_lut_8pts~1 .lut_mask = 16'h6996;
defparam \gain_lut_8pts~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \gain_lut_8pts~2 (
	.dataa(r_array_out_7_2),
	.datab(r_array_out_3_2),
	.datac(i_array_out_7_2),
	.datad(i_array_out_3_2),
	.cin(gnd),
	.combout(\gain_lut_8pts~2_combout ),
	.cout());
defparam \gain_lut_8pts~2 .lut_mask = 16'h6996;
defparam \gain_lut_8pts~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \gain_lut_8pts~3 (
	.dataa(r_array_out_7_3),
	.datab(r_array_out_3_3),
	.datac(i_array_out_7_3),
	.datad(i_array_out_3_3),
	.cin(gnd),
	.combout(\gain_lut_8pts~3_combout ),
	.cout());
defparam \gain_lut_8pts~3 .lut_mask = 16'h6996;
defparam \gain_lut_8pts~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \gain_lut_8pts~4 (
	.dataa(\gain_lut_8pts~0_combout ),
	.datab(\gain_lut_8pts~1_combout ),
	.datac(\gain_lut_8pts~2_combout ),
	.datad(\gain_lut_8pts~3_combout ),
	.cin(gnd),
	.combout(\gain_lut_8pts~4_combout ),
	.cout());
defparam \gain_lut_8pts~4 .lut_mask = 16'hFFFE;
defparam \gain_lut_8pts~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \gain_lut_8pts~5 (
	.dataa(reset_n),
	.datab(enable_op),
	.datac(\gain_lut_8pts~4_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\gain_lut_8pts~5_combout ),
	.cout());
defparam \gain_lut_8pts~5 .lut_mask = 16'hFEFE;
defparam \gain_lut_8pts~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \gain_lut_8pts~7 (
	.dataa(r_array_out_7_1),
	.datab(r_array_out_4_1),
	.datac(i_array_out_7_1),
	.datad(i_array_out_4_1),
	.cin(gnd),
	.combout(\gain_lut_8pts~7_combout ),
	.cout());
defparam \gain_lut_8pts~7 .lut_mask = 16'h6996;
defparam \gain_lut_8pts~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \gain_lut_8pts~8 (
	.dataa(r_array_out_7_2),
	.datab(r_array_out_4_2),
	.datac(i_array_out_7_2),
	.datad(i_array_out_4_2),
	.cin(gnd),
	.combout(\gain_lut_8pts~8_combout ),
	.cout());
defparam \gain_lut_8pts~8 .lut_mask = 16'h6996;
defparam \gain_lut_8pts~8 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \gain_lut_8pts~9 (
	.dataa(r_array_out_7_3),
	.datab(r_array_out_4_3),
	.datac(i_array_out_7_3),
	.datad(i_array_out_4_3),
	.cin(gnd),
	.combout(\gain_lut_8pts~9_combout ),
	.cout());
defparam \gain_lut_8pts~9 .lut_mask = 16'h6996;
defparam \gain_lut_8pts~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \gain_lut_8pts~10 (
	.dataa(\gain_lut_8pts~6_combout ),
	.datab(\gain_lut_8pts~7_combout ),
	.datac(\gain_lut_8pts~8_combout ),
	.datad(\gain_lut_8pts~9_combout ),
	.cin(gnd),
	.combout(\gain_lut_8pts~10_combout ),
	.cout());
defparam \gain_lut_8pts~10 .lut_mask = 16'hFFFE;
defparam \gain_lut_8pts~10 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \gain_lut_8pts~11 (
	.dataa(reset_n),
	.datab(enable_op),
	.datac(\gain_lut_8pts~10_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\gain_lut_8pts~11_combout ),
	.cout());
defparam \gain_lut_8pts~11 .lut_mask = 16'hFEFE;
defparam \gain_lut_8pts~11 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \gain_lut_8pts~13 (
	.dataa(r_array_out_7_1),
	.datab(r_array_out_5_1),
	.datac(i_array_out_7_1),
	.datad(i_array_out_5_1),
	.cin(gnd),
	.combout(\gain_lut_8pts~13_combout ),
	.cout());
defparam \gain_lut_8pts~13 .lut_mask = 16'h6996;
defparam \gain_lut_8pts~13 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \gain_lut_8pts~14 (
	.dataa(r_array_out_7_2),
	.datab(r_array_out_5_2),
	.datac(i_array_out_7_2),
	.datad(i_array_out_5_2),
	.cin(gnd),
	.combout(\gain_lut_8pts~14_combout ),
	.cout());
defparam \gain_lut_8pts~14 .lut_mask = 16'h6996;
defparam \gain_lut_8pts~14 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \gain_lut_8pts~15 (
	.dataa(r_array_out_7_3),
	.datab(r_array_out_5_3),
	.datac(i_array_out_7_3),
	.datad(i_array_out_5_3),
	.cin(gnd),
	.combout(\gain_lut_8pts~15_combout ),
	.cout());
defparam \gain_lut_8pts~15 .lut_mask = 16'h6996;
defparam \gain_lut_8pts~15 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \gain_lut_8pts~16 (
	.dataa(\gain_lut_8pts~12_combout ),
	.datab(\gain_lut_8pts~13_combout ),
	.datac(\gain_lut_8pts~14_combout ),
	.datad(\gain_lut_8pts~15_combout ),
	.cin(gnd),
	.combout(\gain_lut_8pts~16_combout ),
	.cout());
defparam \gain_lut_8pts~16 .lut_mask = 16'hFFFE;
defparam \gain_lut_8pts~16 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \gain_lut_8pts~17 (
	.dataa(reset_n),
	.datab(enable_op),
	.datac(\gain_lut_8pts~16_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\gain_lut_8pts~17_combout ),
	.cout());
defparam \gain_lut_8pts~17 .lut_mask = 16'hFEFE;
defparam \gain_lut_8pts~17 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \gain_lut_8pts~19 (
	.dataa(r_array_out_7_1),
	.datab(r_array_out_6_1),
	.datac(i_array_out_7_1),
	.datad(i_array_out_6_1),
	.cin(gnd),
	.combout(\gain_lut_8pts~19_combout ),
	.cout());
defparam \gain_lut_8pts~19 .lut_mask = 16'h6996;
defparam \gain_lut_8pts~19 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \gain_lut_8pts~20 (
	.dataa(r_array_out_7_2),
	.datab(r_array_out_6_2),
	.datac(i_array_out_7_2),
	.datad(i_array_out_6_2),
	.cin(gnd),
	.combout(\gain_lut_8pts~20_combout ),
	.cout());
defparam \gain_lut_8pts~20 .lut_mask = 16'h6996;
defparam \gain_lut_8pts~20 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \gain_lut_8pts~21 (
	.dataa(r_array_out_7_3),
	.datab(r_array_out_6_3),
	.datac(i_array_out_7_3),
	.datad(i_array_out_6_3),
	.cin(gnd),
	.combout(\gain_lut_8pts~21_combout ),
	.cout());
defparam \gain_lut_8pts~21 .lut_mask = 16'h6996;
defparam \gain_lut_8pts~21 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \gain_lut_8pts~22 (
	.dataa(\gain_lut_8pts~18_combout ),
	.datab(\gain_lut_8pts~19_combout ),
	.datac(\gain_lut_8pts~20_combout ),
	.datad(\gain_lut_8pts~21_combout ),
	.cin(gnd),
	.combout(\gain_lut_8pts~22_combout ),
	.cout());
defparam \gain_lut_8pts~22 .lut_mask = 16'hFFFE;
defparam \gain_lut_8pts~22 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \gain_lut_8pts~23 (
	.dataa(reset_n),
	.datab(enable_op),
	.datac(\gain_lut_8pts~22_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\gain_lut_8pts~23_combout ),
	.cout());
defparam \gain_lut_8pts~23 .lut_mask = 16'hFEFE;
defparam \gain_lut_8pts~23 .sum_lutc_input = "datac";

endmodule

module fft_asj_fft_bfp_o_fft_120 (
	gain_out_4pts_0,
	gain_out_4pts_1,
	gain_out_4pts_2,
	gain_out_4pts_3,
	pipeline_dffe_11,
	pipeline_dffe_15,
	pipeline_dffe_111,
	pipeline_dffe_151,
	pipeline_dffe_112,
	pipeline_dffe_152,
	pipeline_dffe_12,
	pipeline_dffe_121,
	pipeline_dffe_122,
	pipeline_dffe_13,
	pipeline_dffe_131,
	pipeline_dffe_132,
	pipeline_dffe_14,
	pipeline_dffe_141,
	pipeline_dffe_142,
	global_clock_enable,
	slb_i_0,
	slb_i_1,
	slb_i_2,
	slb_i_3,
	Mux2,
	Mux1,
	reg_no_twiddle603,
	reg_no_twiddle607,
	reg_no_twiddle617,
	reg_no_twiddle613,
	real_out_3,
	real_out_7,
	real_out_31,
	real_out_71,
	real_out_32,
	real_out_72,
	reg_no_twiddle604,
	reg_no_twiddle614,
	real_out_4,
	real_out_41,
	real_out_42,
	reg_no_twiddle605,
	reg_no_twiddle615,
	real_out_5,
	real_out_51,
	real_out_52,
	reg_no_twiddle606,
	reg_no_twiddle616,
	real_out_6,
	real_out_61,
	real_out_62,
	blk_done_vec_2,
	tdl_arr_22,
	next_pass_vec_2,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	gain_out_4pts_0;
input 	gain_out_4pts_1;
input 	gain_out_4pts_2;
input 	gain_out_4pts_3;
input 	pipeline_dffe_11;
input 	pipeline_dffe_15;
input 	pipeline_dffe_111;
input 	pipeline_dffe_151;
input 	pipeline_dffe_112;
input 	pipeline_dffe_152;
input 	pipeline_dffe_12;
input 	pipeline_dffe_121;
input 	pipeline_dffe_122;
input 	pipeline_dffe_13;
input 	pipeline_dffe_131;
input 	pipeline_dffe_132;
input 	pipeline_dffe_14;
input 	pipeline_dffe_141;
input 	pipeline_dffe_142;
input 	global_clock_enable;
output 	slb_i_0;
output 	slb_i_1;
output 	slb_i_2;
output 	slb_i_3;
output 	Mux2;
output 	Mux1;
input 	reg_no_twiddle603;
input 	reg_no_twiddle607;
input 	reg_no_twiddle617;
input 	reg_no_twiddle613;
input 	real_out_3;
input 	real_out_7;
input 	real_out_31;
input 	real_out_71;
input 	real_out_32;
input 	real_out_72;
input 	reg_no_twiddle604;
input 	reg_no_twiddle614;
input 	real_out_4;
input 	real_out_41;
input 	real_out_42;
input 	reg_no_twiddle605;
input 	reg_no_twiddle615;
input 	real_out_5;
input 	real_out_51;
input 	real_out_52;
input 	reg_no_twiddle606;
input 	reg_no_twiddle616;
input 	real_out_6;
input 	real_out_61;
input 	real_out_62;
input 	blk_done_vec_2;
input 	tdl_arr_22;
input 	next_pass_vec_2;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \sdet.BLOCK_READY~q ;
wire \del_np_cnt[4]~q ;
wire \del_np_cnt[0]~q ;
wire \del_np_cnt[2]~q ;
wire \del_np_cnt[1]~q ;
wire \del_np_cnt[3]~q ;
wire \del_np_cnt[0]~6 ;
wire \del_np_cnt[0]~5_combout ;
wire \del_np_cnt[1]~8 ;
wire \del_np_cnt[1]~7_combout ;
wire \del_np_cnt[2]~10 ;
wire \del_np_cnt[2]~9_combout ;
wire \del_np_cnt[3]~12 ;
wire \del_np_cnt[3]~11_combout ;
wire \del_np_cnt[4]~13_combout ;
wire \gain_lut_8pts~0_combout ;
wire \gen_blk_float:gen_streaming:gen_cont:delay_next_pass|tdl_arr[8]~q ;
wire \Equal0~0_combout ;
wire \Selector1~0_combout ;
wire \gain_lut_8pts~6_combout ;
wire \gain_lut_8pts~12_combout ;
wire \gain_lut_8pts~18_combout ;
wire \sdet.IDLE~q ;
wire \Selector0~0_combout ;
wire \delay_next_pass_counter~2_combout ;
wire \gap_reg~0_combout ;
wire \gap_reg~q ;
wire \Selector1~1_combout ;
wire \Selector1~2_combout ;
wire \sdet.ENABLE~q ;
wire \sdet~7_combout ;
wire \sdet.DISABLE~q ;
wire \sdet~8_combout ;
wire \sdet.BLOCK_GAP~q ;
wire \en_gain_lut_8_pts~0_combout ;
wire \en_gain_lut_8_pts~1_combout ;
wire \en_gain_lut_8_pts~q ;
wire \gain_lut_8pts~1_combout ;
wire \gain_lut_8pts~2_combout ;
wire \gain_lut_8pts~3_combout ;
wire \gain_lut_8pts~4_combout ;
wire \gain_lut_8pts~5_combout ;
wire \gain_lut_8pts[0]~q ;
wire \gain_lut_blk~0_combout ;
wire \gain_lut_blk[0]~q ;
wire \Selector5~0_combout ;
wire \slb_i[3]~0_combout ;
wire \gain_lut_8pts~7_combout ;
wire \gain_lut_8pts~8_combout ;
wire \gain_lut_8pts~9_combout ;
wire \gain_lut_8pts~10_combout ;
wire \gain_lut_8pts~11_combout ;
wire \gain_lut_8pts[1]~q ;
wire \gain_lut_blk~1_combout ;
wire \gain_lut_blk[1]~q ;
wire \Selector4~0_combout ;
wire \gain_lut_8pts~13_combout ;
wire \gain_lut_8pts~14_combout ;
wire \gain_lut_8pts~15_combout ;
wire \gain_lut_8pts~16_combout ;
wire \gain_lut_8pts~17_combout ;
wire \gain_lut_8pts[2]~q ;
wire \gain_lut_blk~2_combout ;
wire \gain_lut_blk[2]~q ;
wire \Selector3~0_combout ;
wire \gain_lut_8pts~19_combout ;
wire \gain_lut_8pts~20_combout ;
wire \gain_lut_8pts~21_combout ;
wire \gain_lut_8pts~22_combout ;
wire \gain_lut_8pts~23_combout ;
wire \gain_lut_8pts[3]~q ;
wire \gain_lut_blk~3_combout ;
wire \gain_lut_blk[3]~q ;
wire \Selector2~0_combout ;


fft_asj_fft_tdl_bit_fft_120_1 \gen_blk_float:gen_streaming:gen_cont:delay_next_pass (
	.global_clock_enable(global_clock_enable),
	.tdl_arr_8(\gen_blk_float:gen_streaming:gen_cont:delay_next_pass|tdl_arr[8]~q ),
	.data_in(next_pass_vec_2),
	.clk(clk));

dffeas \sdet.BLOCK_READY (
	.clk(clk),
	.d(\Selector0~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sdet.BLOCK_READY~q ),
	.prn(vcc));
defparam \sdet.BLOCK_READY .is_wysiwyg = "true";
defparam \sdet.BLOCK_READY .power_up = "low";

dffeas \del_np_cnt[4] (
	.clk(clk),
	.d(\del_np_cnt[4]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\delay_next_pass_counter~2_combout ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\del_np_cnt[4]~q ),
	.prn(vcc));
defparam \del_np_cnt[4] .is_wysiwyg = "true";
defparam \del_np_cnt[4] .power_up = "low";

dffeas \del_np_cnt[0] (
	.clk(clk),
	.d(\del_np_cnt[0]~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\delay_next_pass_counter~2_combout ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\del_np_cnt[0]~q ),
	.prn(vcc));
defparam \del_np_cnt[0] .is_wysiwyg = "true";
defparam \del_np_cnt[0] .power_up = "low";

dffeas \del_np_cnt[2] (
	.clk(clk),
	.d(\del_np_cnt[2]~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\delay_next_pass_counter~2_combout ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\del_np_cnt[2]~q ),
	.prn(vcc));
defparam \del_np_cnt[2] .is_wysiwyg = "true";
defparam \del_np_cnt[2] .power_up = "low";

dffeas \del_np_cnt[1] (
	.clk(clk),
	.d(\del_np_cnt[1]~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\delay_next_pass_counter~2_combout ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\del_np_cnt[1]~q ),
	.prn(vcc));
defparam \del_np_cnt[1] .is_wysiwyg = "true";
defparam \del_np_cnt[1] .power_up = "low";

dffeas \del_np_cnt[3] (
	.clk(clk),
	.d(\del_np_cnt[3]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\delay_next_pass_counter~2_combout ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\del_np_cnt[3]~q ),
	.prn(vcc));
defparam \del_np_cnt[3] .is_wysiwyg = "true";
defparam \del_np_cnt[3] .power_up = "low";

cycloneiii_lcell_comb \del_np_cnt[0]~5 (
	.dataa(\del_np_cnt[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\del_np_cnt[0]~5_combout ),
	.cout(\del_np_cnt[0]~6 ));
defparam \del_np_cnt[0]~5 .lut_mask = 16'h55AA;
defparam \del_np_cnt[0]~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \del_np_cnt[1]~7 (
	.dataa(\del_np_cnt[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\del_np_cnt[0]~6 ),
	.combout(\del_np_cnt[1]~7_combout ),
	.cout(\del_np_cnt[1]~8 ));
defparam \del_np_cnt[1]~7 .lut_mask = 16'h5A5F;
defparam \del_np_cnt[1]~7 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \del_np_cnt[2]~9 (
	.dataa(\del_np_cnt[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\del_np_cnt[1]~8 ),
	.combout(\del_np_cnt[2]~9_combout ),
	.cout(\del_np_cnt[2]~10 ));
defparam \del_np_cnt[2]~9 .lut_mask = 16'h5AAF;
defparam \del_np_cnt[2]~9 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \del_np_cnt[3]~11 (
	.dataa(\del_np_cnt[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\del_np_cnt[2]~10 ),
	.combout(\del_np_cnt[3]~11_combout ),
	.cout(\del_np_cnt[3]~12 ));
defparam \del_np_cnt[3]~11 .lut_mask = 16'h5A5F;
defparam \del_np_cnt[3]~11 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \del_np_cnt[4]~13 (
	.dataa(\del_np_cnt[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\del_np_cnt[3]~12 ),
	.combout(\del_np_cnt[4]~13_combout ),
	.cout());
defparam \del_np_cnt[4]~13 .lut_mask = 16'h5A5A;
defparam \del_np_cnt[4]~13 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \gain_lut_8pts~0 (
	.dataa(reg_no_twiddle603),
	.datab(reg_no_twiddle607),
	.datac(reg_no_twiddle617),
	.datad(reg_no_twiddle613),
	.cin(gnd),
	.combout(\gain_lut_8pts~0_combout ),
	.cout());
defparam \gain_lut_8pts~0 .lut_mask = 16'h6996;
defparam \gain_lut_8pts~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Equal0~0 (
	.dataa(\del_np_cnt[0]~q ),
	.datab(\del_np_cnt[2]~q ),
	.datac(\del_np_cnt[1]~q ),
	.datad(\del_np_cnt[3]~q ),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
defparam \Equal0~0 .lut_mask = 16'hEFFF;
defparam \Equal0~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector1~0 (
	.dataa(\sdet.BLOCK_READY~q ),
	.datab(\del_np_cnt[4]~q ),
	.datac(\Equal0~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector1~0_combout ),
	.cout());
defparam \Selector1~0 .lut_mask = 16'hFEFE;
defparam \Selector1~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \gain_lut_8pts~6 (
	.dataa(reg_no_twiddle607),
	.datab(reg_no_twiddle604),
	.datac(reg_no_twiddle617),
	.datad(reg_no_twiddle614),
	.cin(gnd),
	.combout(\gain_lut_8pts~6_combout ),
	.cout());
defparam \gain_lut_8pts~6 .lut_mask = 16'h6996;
defparam \gain_lut_8pts~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \gain_lut_8pts~12 (
	.dataa(reg_no_twiddle607),
	.datab(reg_no_twiddle605),
	.datac(reg_no_twiddle617),
	.datad(reg_no_twiddle615),
	.cin(gnd),
	.combout(\gain_lut_8pts~12_combout ),
	.cout());
defparam \gain_lut_8pts~12 .lut_mask = 16'h6996;
defparam \gain_lut_8pts~12 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \gain_lut_8pts~18 (
	.dataa(reg_no_twiddle607),
	.datab(reg_no_twiddle606),
	.datac(reg_no_twiddle617),
	.datad(reg_no_twiddle616),
	.cin(gnd),
	.combout(\gain_lut_8pts~18_combout ),
	.cout());
defparam \gain_lut_8pts~18 .lut_mask = 16'h6996;
defparam \gain_lut_8pts~18 .sum_lutc_input = "datac";

dffeas \sdet.IDLE (
	.clk(clk),
	.d(reset_n),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sdet.IDLE~q ),
	.prn(vcc));
defparam \sdet.IDLE .is_wysiwyg = "true";
defparam \sdet.IDLE .power_up = "low";

cycloneiii_lcell_comb \Selector0~0 (
	.dataa(\sdet.BLOCK_READY~q ),
	.datab(\del_np_cnt[4]~q ),
	.datac(\Equal0~0_combout ),
	.datad(\sdet.IDLE~q ),
	.cin(gnd),
	.combout(\Selector0~0_combout ),
	.cout());
defparam \Selector0~0 .lut_mask = 16'hBFFF;
defparam \Selector0~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \delay_next_pass_counter~2 (
	.dataa(\sdet.DISABLE~q ),
	.datab(\sdet.BLOCK_READY~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_next_pass_counter~2_combout ),
	.cout());
defparam \delay_next_pass_counter~2 .lut_mask = 16'h7777;
defparam \delay_next_pass_counter~2 .sum_lutc_input = "datac";

dffeas \slb_i[0] (
	.clk(clk),
	.d(\Selector5~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\slb_i[3]~0_combout ),
	.q(slb_i_0),
	.prn(vcc));
defparam \slb_i[0] .is_wysiwyg = "true";
defparam \slb_i[0] .power_up = "low";

dffeas \slb_i[1] (
	.clk(clk),
	.d(\Selector4~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\slb_i[3]~0_combout ),
	.q(slb_i_1),
	.prn(vcc));
defparam \slb_i[1] .is_wysiwyg = "true";
defparam \slb_i[1] .power_up = "low";

dffeas \slb_i[2] (
	.clk(clk),
	.d(\Selector3~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\slb_i[3]~0_combout ),
	.q(slb_i_2),
	.prn(vcc));
defparam \slb_i[2] .is_wysiwyg = "true";
defparam \slb_i[2] .power_up = "low";

dffeas \slb_i[3] (
	.clk(clk),
	.d(\Selector2~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\slb_i[3]~0_combout ),
	.q(slb_i_3),
	.prn(vcc));
defparam \slb_i[3] .is_wysiwyg = "true";
defparam \slb_i[3] .power_up = "low";

cycloneiii_lcell_comb \Mux2~0 (
	.dataa(slb_i_0),
	.datab(slb_i_1),
	.datac(slb_i_2),
	.datad(slb_i_3),
	.cin(gnd),
	.combout(Mux2),
	.cout());
defparam \Mux2~0 .lut_mask = 16'hFBFF;
defparam \Mux2~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux1~0 (
	.dataa(slb_i_0),
	.datab(slb_i_1),
	.datac(slb_i_2),
	.datad(slb_i_3),
	.cin(gnd),
	.combout(Mux1),
	.cout());
defparam \Mux1~0 .lut_mask = 16'hEFFF;
defparam \Mux1~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \gap_reg~0 (
	.dataa(blk_done_vec_2),
	.datab(\gap_reg~q ),
	.datac(gnd),
	.datad(tdl_arr_22),
	.cin(gnd),
	.combout(\gap_reg~0_combout ),
	.cout());
defparam \gap_reg~0 .lut_mask = 16'hEEFF;
defparam \gap_reg~0 .sum_lutc_input = "datac";

dffeas gap_reg(
	.clk(clk),
	.d(\gap_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\gap_reg~q ),
	.prn(vcc));
defparam gap_reg.is_wysiwyg = "true";
defparam gap_reg.power_up = "low";

cycloneiii_lcell_comb \Selector1~1 (
	.dataa(\sdet.DISABLE~q ),
	.datab(\sdet.BLOCK_GAP~q ),
	.datac(gnd),
	.datad(\gap_reg~q ),
	.cin(gnd),
	.combout(\Selector1~1_combout ),
	.cout());
defparam \Selector1~1 .lut_mask = 16'hEEFF;
defparam \Selector1~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector1~2 (
	.dataa(\Selector1~0_combout ),
	.datab(\Selector1~1_combout ),
	.datac(\sdet.ENABLE~q ),
	.datad(\gen_blk_float:gen_streaming:gen_cont:delay_next_pass|tdl_arr[8]~q ),
	.cin(gnd),
	.combout(\Selector1~2_combout ),
	.cout());
defparam \Selector1~2 .lut_mask = 16'hFEFF;
defparam \Selector1~2 .sum_lutc_input = "datac";

dffeas \sdet.ENABLE (
	.clk(clk),
	.d(\Selector1~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sdet.ENABLE~q ),
	.prn(vcc));
defparam \sdet.ENABLE .is_wysiwyg = "true";
defparam \sdet.ENABLE .power_up = "low";

cycloneiii_lcell_comb \sdet~7 (
	.dataa(reset_n),
	.datab(\sdet.ENABLE~q ),
	.datac(\gen_blk_float:gen_streaming:gen_cont:delay_next_pass|tdl_arr[8]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\sdet~7_combout ),
	.cout());
defparam \sdet~7 .lut_mask = 16'hFEFE;
defparam \sdet~7 .sum_lutc_input = "datac";

dffeas \sdet.DISABLE (
	.clk(clk),
	.d(\sdet~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sdet.DISABLE~q ),
	.prn(vcc));
defparam \sdet.DISABLE .is_wysiwyg = "true";
defparam \sdet.DISABLE .power_up = "low";

cycloneiii_lcell_comb \sdet~8 (
	.dataa(reset_n),
	.datab(\gap_reg~q ),
	.datac(\sdet.DISABLE~q ),
	.datad(\sdet.BLOCK_GAP~q ),
	.cin(gnd),
	.combout(\sdet~8_combout ),
	.cout());
defparam \sdet~8 .lut_mask = 16'hFFFE;
defparam \sdet~8 .sum_lutc_input = "datac";

dffeas \sdet.BLOCK_GAP (
	.clk(clk),
	.d(\sdet~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sdet.BLOCK_GAP~q ),
	.prn(vcc));
defparam \sdet.BLOCK_GAP .is_wysiwyg = "true";
defparam \sdet.BLOCK_GAP .power_up = "low";

cycloneiii_lcell_comb \en_gain_lut_8_pts~0 (
	.dataa(\sdet.DISABLE~q ),
	.datab(\en_gain_lut_8_pts~q ),
	.datac(\sdet.BLOCK_GAP~q ),
	.datad(\gap_reg~q ),
	.cin(gnd),
	.combout(\en_gain_lut_8_pts~0_combout ),
	.cout());
defparam \en_gain_lut_8_pts~0 .lut_mask = 16'hACFF;
defparam \en_gain_lut_8_pts~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \en_gain_lut_8_pts~1 (
	.dataa(\sdet.ENABLE~q ),
	.datab(\en_gain_lut_8_pts~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\en_gain_lut_8_pts~1_combout ),
	.cout());
defparam \en_gain_lut_8_pts~1 .lut_mask = 16'hEEEE;
defparam \en_gain_lut_8_pts~1 .sum_lutc_input = "datac";

dffeas en_gain_lut_8_pts(
	.clk(clk),
	.d(\en_gain_lut_8_pts~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\en_gain_lut_8_pts~q ),
	.prn(vcc));
defparam en_gain_lut_8_pts.is_wysiwyg = "true";
defparam en_gain_lut_8_pts.power_up = "low";

cycloneiii_lcell_comb \gain_lut_8pts~1 (
	.dataa(pipeline_dffe_11),
	.datab(pipeline_dffe_15),
	.datac(real_out_3),
	.datad(real_out_7),
	.cin(gnd),
	.combout(\gain_lut_8pts~1_combout ),
	.cout());
defparam \gain_lut_8pts~1 .lut_mask = 16'h6996;
defparam \gain_lut_8pts~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \gain_lut_8pts~2 (
	.dataa(pipeline_dffe_111),
	.datab(pipeline_dffe_151),
	.datac(real_out_31),
	.datad(real_out_71),
	.cin(gnd),
	.combout(\gain_lut_8pts~2_combout ),
	.cout());
defparam \gain_lut_8pts~2 .lut_mask = 16'h6996;
defparam \gain_lut_8pts~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \gain_lut_8pts~3 (
	.dataa(pipeline_dffe_112),
	.datab(pipeline_dffe_152),
	.datac(real_out_32),
	.datad(real_out_72),
	.cin(gnd),
	.combout(\gain_lut_8pts~3_combout ),
	.cout());
defparam \gain_lut_8pts~3 .lut_mask = 16'h6996;
defparam \gain_lut_8pts~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \gain_lut_8pts~4 (
	.dataa(\gain_lut_8pts~0_combout ),
	.datab(\gain_lut_8pts~1_combout ),
	.datac(\gain_lut_8pts~2_combout ),
	.datad(\gain_lut_8pts~3_combout ),
	.cin(gnd),
	.combout(\gain_lut_8pts~4_combout ),
	.cout());
defparam \gain_lut_8pts~4 .lut_mask = 16'hFFFE;
defparam \gain_lut_8pts~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \gain_lut_8pts~5 (
	.dataa(reset_n),
	.datab(\en_gain_lut_8_pts~q ),
	.datac(\gain_lut_8pts~4_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\gain_lut_8pts~5_combout ),
	.cout());
defparam \gain_lut_8pts~5 .lut_mask = 16'hFEFE;
defparam \gain_lut_8pts~5 .sum_lutc_input = "datac";

dffeas \gain_lut_8pts[0] (
	.clk(clk),
	.d(\gain_lut_8pts~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\gain_lut_8pts[0]~q ),
	.prn(vcc));
defparam \gain_lut_8pts[0] .is_wysiwyg = "true";
defparam \gain_lut_8pts[0] .power_up = "low";

cycloneiii_lcell_comb \gain_lut_blk~0 (
	.dataa(\sdet.ENABLE~q ),
	.datab(\gain_lut_8pts[0]~q ),
	.datac(\gain_lut_blk[0]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\gain_lut_blk~0_combout ),
	.cout());
defparam \gain_lut_blk~0 .lut_mask = 16'hFEFE;
defparam \gain_lut_blk~0 .sum_lutc_input = "datac";

dffeas \gain_lut_blk[0] (
	.clk(clk),
	.d(\gain_lut_blk~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\gain_lut_blk[0]~q ),
	.prn(vcc));
defparam \gain_lut_blk[0] .is_wysiwyg = "true";
defparam \gain_lut_blk[0] .power_up = "low";

cycloneiii_lcell_comb \Selector5~0 (
	.dataa(\gain_lut_8pts[0]~q ),
	.datab(\gain_lut_blk[0]~q ),
	.datac(gain_out_4pts_0),
	.datad(\sdet.DISABLE~q ),
	.cin(gnd),
	.combout(\Selector5~0_combout ),
	.cout());
defparam \Selector5~0 .lut_mask = 16'hFEFF;
defparam \Selector5~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \slb_i[3]~0 (
	.dataa(global_clock_enable),
	.datab(\sdet.BLOCK_GAP~q ),
	.datac(\sdet.ENABLE~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\slb_i[3]~0_combout ),
	.cout());
defparam \slb_i[3]~0 .lut_mask = 16'hBFBF;
defparam \slb_i[3]~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \gain_lut_8pts~7 (
	.dataa(pipeline_dffe_15),
	.datab(pipeline_dffe_12),
	.datac(real_out_7),
	.datad(real_out_4),
	.cin(gnd),
	.combout(\gain_lut_8pts~7_combout ),
	.cout());
defparam \gain_lut_8pts~7 .lut_mask = 16'h6996;
defparam \gain_lut_8pts~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \gain_lut_8pts~8 (
	.dataa(pipeline_dffe_151),
	.datab(pipeline_dffe_121),
	.datac(real_out_71),
	.datad(real_out_41),
	.cin(gnd),
	.combout(\gain_lut_8pts~8_combout ),
	.cout());
defparam \gain_lut_8pts~8 .lut_mask = 16'h6996;
defparam \gain_lut_8pts~8 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \gain_lut_8pts~9 (
	.dataa(pipeline_dffe_152),
	.datab(pipeline_dffe_122),
	.datac(real_out_72),
	.datad(real_out_42),
	.cin(gnd),
	.combout(\gain_lut_8pts~9_combout ),
	.cout());
defparam \gain_lut_8pts~9 .lut_mask = 16'h6996;
defparam \gain_lut_8pts~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \gain_lut_8pts~10 (
	.dataa(\gain_lut_8pts~6_combout ),
	.datab(\gain_lut_8pts~7_combout ),
	.datac(\gain_lut_8pts~8_combout ),
	.datad(\gain_lut_8pts~9_combout ),
	.cin(gnd),
	.combout(\gain_lut_8pts~10_combout ),
	.cout());
defparam \gain_lut_8pts~10 .lut_mask = 16'hFFFE;
defparam \gain_lut_8pts~10 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \gain_lut_8pts~11 (
	.dataa(reset_n),
	.datab(\en_gain_lut_8_pts~q ),
	.datac(\gain_lut_8pts~10_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\gain_lut_8pts~11_combout ),
	.cout());
defparam \gain_lut_8pts~11 .lut_mask = 16'hFEFE;
defparam \gain_lut_8pts~11 .sum_lutc_input = "datac";

dffeas \gain_lut_8pts[1] (
	.clk(clk),
	.d(\gain_lut_8pts~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\gain_lut_8pts[1]~q ),
	.prn(vcc));
defparam \gain_lut_8pts[1] .is_wysiwyg = "true";
defparam \gain_lut_8pts[1] .power_up = "low";

cycloneiii_lcell_comb \gain_lut_blk~1 (
	.dataa(\sdet.ENABLE~q ),
	.datab(\gain_lut_8pts[1]~q ),
	.datac(\gain_lut_blk[1]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\gain_lut_blk~1_combout ),
	.cout());
defparam \gain_lut_blk~1 .lut_mask = 16'hFEFE;
defparam \gain_lut_blk~1 .sum_lutc_input = "datac";

dffeas \gain_lut_blk[1] (
	.clk(clk),
	.d(\gain_lut_blk~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\gain_lut_blk[1]~q ),
	.prn(vcc));
defparam \gain_lut_blk[1] .is_wysiwyg = "true";
defparam \gain_lut_blk[1] .power_up = "low";

cycloneiii_lcell_comb \Selector4~0 (
	.dataa(\gain_lut_8pts[1]~q ),
	.datab(\gain_lut_blk[1]~q ),
	.datac(gain_out_4pts_1),
	.datad(\sdet.DISABLE~q ),
	.cin(gnd),
	.combout(\Selector4~0_combout ),
	.cout());
defparam \Selector4~0 .lut_mask = 16'hFEFF;
defparam \Selector4~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \gain_lut_8pts~13 (
	.dataa(pipeline_dffe_15),
	.datab(pipeline_dffe_13),
	.datac(real_out_7),
	.datad(real_out_5),
	.cin(gnd),
	.combout(\gain_lut_8pts~13_combout ),
	.cout());
defparam \gain_lut_8pts~13 .lut_mask = 16'h6996;
defparam \gain_lut_8pts~13 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \gain_lut_8pts~14 (
	.dataa(pipeline_dffe_151),
	.datab(pipeline_dffe_131),
	.datac(real_out_71),
	.datad(real_out_51),
	.cin(gnd),
	.combout(\gain_lut_8pts~14_combout ),
	.cout());
defparam \gain_lut_8pts~14 .lut_mask = 16'h6996;
defparam \gain_lut_8pts~14 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \gain_lut_8pts~15 (
	.dataa(pipeline_dffe_152),
	.datab(pipeline_dffe_132),
	.datac(real_out_72),
	.datad(real_out_52),
	.cin(gnd),
	.combout(\gain_lut_8pts~15_combout ),
	.cout());
defparam \gain_lut_8pts~15 .lut_mask = 16'h6996;
defparam \gain_lut_8pts~15 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \gain_lut_8pts~16 (
	.dataa(\gain_lut_8pts~12_combout ),
	.datab(\gain_lut_8pts~13_combout ),
	.datac(\gain_lut_8pts~14_combout ),
	.datad(\gain_lut_8pts~15_combout ),
	.cin(gnd),
	.combout(\gain_lut_8pts~16_combout ),
	.cout());
defparam \gain_lut_8pts~16 .lut_mask = 16'hFFFE;
defparam \gain_lut_8pts~16 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \gain_lut_8pts~17 (
	.dataa(reset_n),
	.datab(\en_gain_lut_8_pts~q ),
	.datac(\gain_lut_8pts~16_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\gain_lut_8pts~17_combout ),
	.cout());
defparam \gain_lut_8pts~17 .lut_mask = 16'hFEFE;
defparam \gain_lut_8pts~17 .sum_lutc_input = "datac";

dffeas \gain_lut_8pts[2] (
	.clk(clk),
	.d(\gain_lut_8pts~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\gain_lut_8pts[2]~q ),
	.prn(vcc));
defparam \gain_lut_8pts[2] .is_wysiwyg = "true";
defparam \gain_lut_8pts[2] .power_up = "low";

cycloneiii_lcell_comb \gain_lut_blk~2 (
	.dataa(\sdet.ENABLE~q ),
	.datab(\gain_lut_8pts[2]~q ),
	.datac(\gain_lut_blk[2]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\gain_lut_blk~2_combout ),
	.cout());
defparam \gain_lut_blk~2 .lut_mask = 16'hFEFE;
defparam \gain_lut_blk~2 .sum_lutc_input = "datac";

dffeas \gain_lut_blk[2] (
	.clk(clk),
	.d(\gain_lut_blk~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\gain_lut_blk[2]~q ),
	.prn(vcc));
defparam \gain_lut_blk[2] .is_wysiwyg = "true";
defparam \gain_lut_blk[2] .power_up = "low";

cycloneiii_lcell_comb \Selector3~0 (
	.dataa(\gain_lut_8pts[2]~q ),
	.datab(\gain_lut_blk[2]~q ),
	.datac(gain_out_4pts_2),
	.datad(\sdet.DISABLE~q ),
	.cin(gnd),
	.combout(\Selector3~0_combout ),
	.cout());
defparam \Selector3~0 .lut_mask = 16'hFEFF;
defparam \Selector3~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \gain_lut_8pts~19 (
	.dataa(pipeline_dffe_15),
	.datab(pipeline_dffe_14),
	.datac(real_out_7),
	.datad(real_out_6),
	.cin(gnd),
	.combout(\gain_lut_8pts~19_combout ),
	.cout());
defparam \gain_lut_8pts~19 .lut_mask = 16'h6996;
defparam \gain_lut_8pts~19 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \gain_lut_8pts~20 (
	.dataa(pipeline_dffe_151),
	.datab(pipeline_dffe_141),
	.datac(real_out_71),
	.datad(real_out_61),
	.cin(gnd),
	.combout(\gain_lut_8pts~20_combout ),
	.cout());
defparam \gain_lut_8pts~20 .lut_mask = 16'h6996;
defparam \gain_lut_8pts~20 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \gain_lut_8pts~21 (
	.dataa(pipeline_dffe_152),
	.datab(pipeline_dffe_142),
	.datac(real_out_72),
	.datad(real_out_62),
	.cin(gnd),
	.combout(\gain_lut_8pts~21_combout ),
	.cout());
defparam \gain_lut_8pts~21 .lut_mask = 16'h6996;
defparam \gain_lut_8pts~21 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \gain_lut_8pts~22 (
	.dataa(\gain_lut_8pts~18_combout ),
	.datab(\gain_lut_8pts~19_combout ),
	.datac(\gain_lut_8pts~20_combout ),
	.datad(\gain_lut_8pts~21_combout ),
	.cin(gnd),
	.combout(\gain_lut_8pts~22_combout ),
	.cout());
defparam \gain_lut_8pts~22 .lut_mask = 16'hFFFE;
defparam \gain_lut_8pts~22 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \gain_lut_8pts~23 (
	.dataa(reset_n),
	.datab(\en_gain_lut_8_pts~q ),
	.datac(\gain_lut_8pts~22_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\gain_lut_8pts~23_combout ),
	.cout());
defparam \gain_lut_8pts~23 .lut_mask = 16'hFEFE;
defparam \gain_lut_8pts~23 .sum_lutc_input = "datac";

dffeas \gain_lut_8pts[3] (
	.clk(clk),
	.d(\gain_lut_8pts~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\gain_lut_8pts[3]~q ),
	.prn(vcc));
defparam \gain_lut_8pts[3] .is_wysiwyg = "true";
defparam \gain_lut_8pts[3] .power_up = "low";

cycloneiii_lcell_comb \gain_lut_blk~3 (
	.dataa(\sdet.ENABLE~q ),
	.datab(\gain_lut_8pts[3]~q ),
	.datac(\gain_lut_blk[3]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\gain_lut_blk~3_combout ),
	.cout());
defparam \gain_lut_blk~3 .lut_mask = 16'hFEFE;
defparam \gain_lut_blk~3 .sum_lutc_input = "datac";

dffeas \gain_lut_blk[3] (
	.clk(clk),
	.d(\gain_lut_blk~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\gain_lut_blk[3]~q ),
	.prn(vcc));
defparam \gain_lut_blk[3] .is_wysiwyg = "true";
defparam \gain_lut_blk[3] .power_up = "low";

cycloneiii_lcell_comb \Selector2~0 (
	.dataa(\gain_lut_8pts[3]~q ),
	.datab(\gain_lut_blk[3]~q ),
	.datac(gain_out_4pts_3),
	.datad(\sdet.DISABLE~q ),
	.cin(gnd),
	.combout(\Selector2~0_combout ),
	.cout());
defparam \Selector2~0 .lut_mask = 16'hFEFF;
defparam \Selector2~0 .sum_lutc_input = "datac";

endmodule

module fft_asj_fft_tdl_bit_fft_120_1 (
	global_clock_enable,
	tdl_arr_8,
	data_in,
	clk)/* synthesis synthesis_greybox=1 */;
input 	global_clock_enable;
output 	tdl_arr_8;
input 	data_in;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \tdl_arr[0]~q ;
wire \tdl_arr[1]~q ;
wire \tdl_arr[2]~q ;
wire \tdl_arr[3]~q ;
wire \tdl_arr[4]~q ;
wire \tdl_arr[5]~q ;
wire \tdl_arr[6]~q ;
wire \tdl_arr[7]~q ;


dffeas \tdl_arr[8] (
	.clk(clk),
	.d(\tdl_arr[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_8),
	.prn(vcc));
defparam \tdl_arr[8] .is_wysiwyg = "true";
defparam \tdl_arr[8] .power_up = "low";

dffeas \tdl_arr[0] (
	.clk(clk),
	.d(data_in),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0]~q ),
	.prn(vcc));
defparam \tdl_arr[0] .is_wysiwyg = "true";
defparam \tdl_arr[0] .power_up = "low";

dffeas \tdl_arr[1] (
	.clk(clk),
	.d(\tdl_arr[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[1]~q ),
	.prn(vcc));
defparam \tdl_arr[1] .is_wysiwyg = "true";
defparam \tdl_arr[1] .power_up = "low";

dffeas \tdl_arr[2] (
	.clk(clk),
	.d(\tdl_arr[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[2]~q ),
	.prn(vcc));
defparam \tdl_arr[2] .is_wysiwyg = "true";
defparam \tdl_arr[2] .power_up = "low";

dffeas \tdl_arr[3] (
	.clk(clk),
	.d(\tdl_arr[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[3]~q ),
	.prn(vcc));
defparam \tdl_arr[3] .is_wysiwyg = "true";
defparam \tdl_arr[3] .power_up = "low";

dffeas \tdl_arr[4] (
	.clk(clk),
	.d(\tdl_arr[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[4]~q ),
	.prn(vcc));
defparam \tdl_arr[4] .is_wysiwyg = "true";
defparam \tdl_arr[4] .power_up = "low";

dffeas \tdl_arr[5] (
	.clk(clk),
	.d(\tdl_arr[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[5]~q ),
	.prn(vcc));
defparam \tdl_arr[5] .is_wysiwyg = "true";
defparam \tdl_arr[5] .power_up = "low";

dffeas \tdl_arr[6] (
	.clk(clk),
	.d(\tdl_arr[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[6]~q ),
	.prn(vcc));
defparam \tdl_arr[6] .is_wysiwyg = "true";
defparam \tdl_arr[6] .power_up = "low";

dffeas \tdl_arr[7] (
	.clk(clk),
	.d(\tdl_arr[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[7]~q ),
	.prn(vcc));
defparam \tdl_arr[7] .is_wysiwyg = "true";
defparam \tdl_arr[7] .power_up = "low";

endmodule

module fft_asj_fft_cmult_can_fft_120 (
	pipeline_dffe_11,
	pipeline_dffe_15,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	pipeline_dffe_9,
	pipeline_dffe_8,
	pipeline_dffe_10,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_81,
	pipeline_dffe_91,
	pipeline_dffe_21,
	pipeline_dffe_31,
	pipeline_dffe_41,
	pipeline_dffe_51,
	pipeline_dffe_61,
	pipeline_dffe_71,
	pipeline_dffe_82,
	pipeline_dffe_92,
	global_clock_enable,
	real_out_3,
	real_out_7,
	real_out_4,
	real_out_5,
	real_out_6,
	real_out_1,
	real_out_0,
	real_out_2,
	twiddle_data000,
	twiddle_data001,
	twiddle_data002,
	twiddle_data003,
	twiddle_data004,
	twiddle_data005,
	twiddle_data006,
	twiddle_data007,
	twiddle_data010,
	twiddle_data011,
	twiddle_data012,
	twiddle_data013,
	twiddle_data014,
	twiddle_data015,
	twiddle_data016,
	twiddle_data017,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_11;
output 	pipeline_dffe_15;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
output 	pipeline_dffe_9;
output 	pipeline_dffe_8;
output 	pipeline_dffe_10;
input 	pipeline_dffe_2;
input 	pipeline_dffe_3;
input 	pipeline_dffe_4;
input 	pipeline_dffe_5;
input 	pipeline_dffe_6;
input 	pipeline_dffe_7;
input 	pipeline_dffe_81;
input 	pipeline_dffe_91;
input 	pipeline_dffe_21;
input 	pipeline_dffe_31;
input 	pipeline_dffe_41;
input 	pipeline_dffe_51;
input 	pipeline_dffe_61;
input 	pipeline_dffe_71;
input 	pipeline_dffe_82;
input 	pipeline_dffe_92;
input 	global_clock_enable;
output 	real_out_3;
output 	real_out_7;
output 	real_out_4;
output 	real_out_5;
output 	real_out_6;
output 	real_out_1;
output 	real_out_0;
output 	real_out_2;
input 	twiddle_data000;
input 	twiddle_data001;
input 	twiddle_data002;
input 	twiddle_data003;
input 	twiddle_data004;
input 	twiddle_data005;
input 	twiddle_data006;
input 	twiddle_data007;
input 	twiddle_data010;
input 	twiddle_data011;
input 	twiddle_data012;
input 	twiddle_data013;
input 	twiddle_data014;
input 	twiddle_data015;
input 	twiddle_data016;
input 	twiddle_data017;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \result_imag_1[11]~q ;
wire \result_imag_1[10]~q ;
wire \result_imag_1[9]~q ;
wire \result_imag_1[8]~q ;
wire \result_imag_1[7]~q ;
wire \result_imag_1[6]~q ;
wire \result_imag_1[5]~q ;
wire \result_imag_1[4]~q ;
wire \result_imag_1[3]~q ;
wire \result_imag_1[2]~q ;
wire \result_imag_1[1]~q ;
wire \result_imag_1[0]~q ;
wire \result_imag_1[15]~q ;
wire \result_imag_1[14]~q ;
wire \result_imag_1[13]~q ;
wire \result_imag_1[12]~q ;
wire \gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ;
wire \gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ;
wire \gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ;
wire \gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ;
wire \gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ;
wire \addresult_ac_bd[11]~q ;
wire \addresult_ac_bd[10]~q ;
wire \addresult_ac_bd[9]~q ;
wire \addresult_ac_bd[8]~q ;
wire \addresult_ac_bd[7]~q ;
wire \addresult_ac_bd[6]~q ;
wire \addresult_ac_bd[5]~q ;
wire \addresult_ac_bd[4]~q ;
wire \addresult_ac_bd[3]~q ;
wire \addresult_ac_bd[2]~q ;
wire \addresult_ac_bd[1]~q ;
wire \addresult_ac_bd[0]~q ;
wire \result_imag_1[0]~17 ;
wire \result_imag_1[0]~16_combout ;
wire \result_imag_1[1]~19 ;
wire \result_imag_1[1]~18_combout ;
wire \result_imag_1[2]~21 ;
wire \result_imag_1[2]~20_combout ;
wire \result_imag_1[3]~23 ;
wire \result_imag_1[3]~22_combout ;
wire \result_imag_1[4]~25 ;
wire \result_imag_1[4]~24_combout ;
wire \result_imag_1[5]~27 ;
wire \result_imag_1[5]~26_combout ;
wire \result_imag_1[6]~29 ;
wire \result_imag_1[6]~28_combout ;
wire \result_imag_1[7]~31 ;
wire \result_imag_1[7]~30_combout ;
wire \result_imag_1[8]~33 ;
wire \result_imag_1[8]~32_combout ;
wire \result_imag_1[9]~35 ;
wire \result_imag_1[9]~34_combout ;
wire \result_imag_1[10]~37 ;
wire \result_imag_1[10]~36_combout ;
wire \result_imag_1[11]~39 ;
wire \result_imag_1[11]~38_combout ;
wire \addresult_ac_bd[15]~q ;
wire \addresult_ac_bd[14]~q ;
wire \addresult_ac_bd[13]~q ;
wire \addresult_ac_bd[12]~q ;
wire \result_imag_1[12]~41 ;
wire \result_imag_1[12]~40_combout ;
wire \result_imag_1[13]~43 ;
wire \result_imag_1[13]~42_combout ;
wire \result_imag_1[14]~45 ;
wire \result_imag_1[14]~44_combout ;
wire \result_imag_1[15]~46_combout ;
wire \result_real_1_tmp[11]~q ;
wire \result_real_1_tmp[10]~q ;
wire \result_real_1_tmp[9]~q ;
wire \result_real_1_tmp[8]~q ;
wire \result_real_1_tmp[7]~q ;
wire \result_real_1_tmp[6]~q ;
wire \result_real_1_tmp[5]~q ;
wire \result_real_1_tmp[4]~q ;
wire \result_real_1_tmp[3]~q ;
wire \result_real_1_tmp[2]~q ;
wire \result_real_1_tmp[1]~q ;
wire \result_real_1_tmp[0]~q ;
wire \result_real_1_tmp[15]~q ;
wire \result_real_1_tmp[14]~q ;
wire \result_real_1_tmp[13]~q ;
wire \result_real_1_tmp[12]~q ;
wire \addresult_ac_bd[0]~17 ;
wire \addresult_ac_bd[0]~16_combout ;
wire \addresult_ac_bd[1]~19 ;
wire \addresult_ac_bd[1]~18_combout ;
wire \addresult_ac_bd[2]~21 ;
wire \addresult_ac_bd[2]~20_combout ;
wire \addresult_ac_bd[3]~23 ;
wire \addresult_ac_bd[3]~22_combout ;
wire \addresult_ac_bd[4]~25 ;
wire \addresult_ac_bd[4]~24_combout ;
wire \addresult_ac_bd[5]~27 ;
wire \addresult_ac_bd[5]~26_combout ;
wire \addresult_ac_bd[6]~29 ;
wire \addresult_ac_bd[6]~28_combout ;
wire \addresult_ac_bd[7]~31 ;
wire \addresult_ac_bd[7]~30_combout ;
wire \addresult_ac_bd[8]~33 ;
wire \addresult_ac_bd[8]~32_combout ;
wire \addresult_ac_bd[9]~35 ;
wire \addresult_ac_bd[9]~34_combout ;
wire \addresult_ac_bd[10]~37 ;
wire \addresult_ac_bd[10]~36_combout ;
wire \addresult_ac_bd[11]~39 ;
wire \addresult_ac_bd[11]~38_combout ;
wire \addresult_ac_bd[12]~41 ;
wire \addresult_ac_bd[12]~40_combout ;
wire \addresult_ac_bd[13]~43 ;
wire \addresult_ac_bd[13]~42_combout ;
wire \addresult_ac_bd[14]~45 ;
wire \addresult_ac_bd[14]~44_combout ;
wire \addresult_ac_bd[15]~46_combout ;
wire \result_real_1_tmp[0]~17 ;
wire \result_real_1_tmp[0]~16_combout ;
wire \result_real_1_tmp[1]~19 ;
wire \result_real_1_tmp[1]~18_combout ;
wire \result_real_1_tmp[2]~21 ;
wire \result_real_1_tmp[2]~20_combout ;
wire \result_real_1_tmp[3]~23 ;
wire \result_real_1_tmp[3]~22_combout ;
wire \result_real_1_tmp[4]~25 ;
wire \result_real_1_tmp[4]~24_combout ;
wire \result_real_1_tmp[5]~27 ;
wire \result_real_1_tmp[5]~26_combout ;
wire \result_real_1_tmp[6]~29 ;
wire \result_real_1_tmp[6]~28_combout ;
wire \result_real_1_tmp[7]~31 ;
wire \result_real_1_tmp[7]~30_combout ;
wire \result_real_1_tmp[8]~33 ;
wire \result_real_1_tmp[8]~32_combout ;
wire \result_real_1_tmp[9]~35 ;
wire \result_real_1_tmp[9]~34_combout ;
wire \result_real_1_tmp[10]~37 ;
wire \result_real_1_tmp[10]~36_combout ;
wire \result_real_1_tmp[11]~39 ;
wire \result_real_1_tmp[11]~38_combout ;
wire \result_real_1_tmp[12]~41 ;
wire \result_real_1_tmp[12]~40_combout ;
wire \result_real_1_tmp[13]~43 ;
wire \result_real_1_tmp[13]~42_combout ;
wire \result_real_1_tmp[14]~45 ;
wire \result_real_1_tmp[14]~44_combout ;
wire \result_real_1_tmp[15]~46_combout ;
wire \addresult_a_b[0]~q ;
wire \addresult_a_b[1]~q ;
wire \addresult_a_b[2]~q ;
wire \addresult_a_b[3]~q ;
wire \addresult_a_b[4]~q ;
wire \addresult_a_b[5]~q ;
wire \addresult_a_b[6]~q ;
wire \addresult_a_b[7]~q ;
wire \addresult_a_b[8]~q ;
wire \addresult_c_d[0]~q ;
wire \addresult_c_d[1]~q ;
wire \addresult_c_d[2]~q ;
wire \addresult_c_d[3]~q ;
wire \addresult_c_d[4]~q ;
wire \addresult_c_d[5]~q ;
wire \addresult_c_d[6]~q ;
wire \addresult_c_d[7]~q ;
wire \addresult_c_d[8]~q ;
wire \addresult_a_b[0]~10 ;
wire \addresult_a_b[0]~9_combout ;
wire \addresult_a_b[1]~12 ;
wire \addresult_a_b[1]~11_combout ;
wire \addresult_a_b[2]~14 ;
wire \addresult_a_b[2]~13_combout ;
wire \addresult_a_b[3]~16 ;
wire \addresult_a_b[3]~15_combout ;
wire \addresult_a_b[4]~18 ;
wire \addresult_a_b[4]~17_combout ;
wire \addresult_a_b[5]~20 ;
wire \addresult_a_b[5]~19_combout ;
wire \addresult_a_b[6]~22 ;
wire \addresult_a_b[6]~21_combout ;
wire \addresult_a_b[7]~24 ;
wire \addresult_a_b[7]~23_combout ;
wire \addresult_a_b[8]~25_combout ;
wire \addresult_c_d[0]~10 ;
wire \addresult_c_d[0]~9_combout ;
wire \addresult_c_d[1]~12 ;
wire \addresult_c_d[1]~11_combout ;
wire \addresult_c_d[2]~14 ;
wire \addresult_c_d[2]~13_combout ;
wire \addresult_c_d[3]~16 ;
wire \addresult_c_d[3]~15_combout ;
wire \addresult_c_d[4]~18 ;
wire \addresult_c_d[4]~17_combout ;
wire \addresult_c_d[5]~20 ;
wire \addresult_c_d[5]~19_combout ;
wire \addresult_c_d[6]~22 ;
wire \addresult_c_d[6]~21_combout ;
wire \addresult_c_d[7]~24 ;
wire \addresult_c_d[7]~23_combout ;
wire \addresult_c_d[8]~25_combout ;
wire \gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ;
wire \gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ;
wire \gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ;
wire \result_a_b_c_d_se[11]~q ;
wire \result_a_b_c_d_se[10]~q ;
wire \result_a_b_c_d_se[9]~q ;
wire \result_a_b_c_d_se[8]~q ;
wire \result_a_b_c_d_se[7]~q ;
wire \result_a_b_c_d_se[6]~q ;
wire \result_a_b_c_d_se[5]~q ;
wire \result_a_b_c_d_se[4]~q ;
wire \result_a_b_c_d_se[3]~q ;
wire \result_a_b_c_d_se[2]~q ;
wire \result_a_b_c_d_se[1]~q ;
wire \result_a_b_c_d_se[0]~q ;
wire \result_a_b_c_d_se[15]~q ;
wire \result_a_b_c_d_se[14]~q ;
wire \result_a_b_c_d_se[13]~q ;
wire \result_a_b_c_d_se[12]~q ;
wire \result_a_c_se[11]~q ;
wire \result_b_d_se[11]~q ;
wire \result_a_c_se[10]~q ;
wire \result_b_d_se[10]~q ;
wire \result_a_c_se[9]~q ;
wire \result_b_d_se[9]~q ;
wire \result_a_c_se[8]~q ;
wire \result_b_d_se[8]~q ;
wire \result_a_c_se[7]~q ;
wire \result_b_d_se[7]~q ;
wire \result_a_c_se[6]~q ;
wire \result_b_d_se[6]~q ;
wire \result_a_c_se[5]~q ;
wire \result_b_d_se[5]~q ;
wire \result_a_c_se[4]~q ;
wire \result_b_d_se[4]~q ;
wire \result_a_c_se[3]~q ;
wire \result_b_d_se[3]~q ;
wire \result_a_c_se[2]~q ;
wire \result_b_d_se[2]~q ;
wire \result_a_c_se[1]~q ;
wire \result_b_d_se[1]~q ;
wire \result_a_c_se[0]~q ;
wire \result_b_d_se[0]~q ;
wire \gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[11]~q ;
wire \gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[10]~q ;
wire \gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[9]~q ;
wire \gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[8]~q ;
wire \gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[7]~q ;
wire \gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[6]~q ;
wire \gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[5]~q ;
wire \gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[4]~q ;
wire \gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[3]~q ;
wire \gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[2]~q ;
wire \gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[1]~q ;
wire \gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[0]~q ;
wire \result_a_c_se[15]~q ;
wire \result_b_d_se[15]~q ;
wire \result_a_c_se[14]~q ;
wire \result_b_d_se[14]~q ;
wire \result_a_c_se[13]~q ;
wire \result_b_d_se[13]~q ;
wire \result_a_c_se[12]~q ;
wire \result_b_d_se[12]~q ;
wire \gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[15]~q ;
wire \gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[14]~q ;
wire \gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[13]~q ;
wire \gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[12]~q ;
wire \gen_dsp_only:m_ac|auto_generated|dffe3a[11]~q ;
wire \gen_dsp_only:m_bd|auto_generated|dffe3a[11]~q ;
wire \gen_dsp_only:m_ac|auto_generated|dffe3a[10]~q ;
wire \gen_dsp_only:m_bd|auto_generated|dffe3a[10]~q ;
wire \gen_dsp_only:m_ac|auto_generated|dffe3a[9]~q ;
wire \gen_dsp_only:m_bd|auto_generated|dffe3a[9]~q ;
wire \gen_dsp_only:m_ac|auto_generated|dffe3a[8]~q ;
wire \gen_dsp_only:m_bd|auto_generated|dffe3a[8]~q ;
wire \gen_dsp_only:m_ac|auto_generated|dffe3a[7]~q ;
wire \gen_dsp_only:m_bd|auto_generated|dffe3a[7]~q ;
wire \gen_dsp_only:m_ac|auto_generated|dffe3a[6]~q ;
wire \gen_dsp_only:m_bd|auto_generated|dffe3a[6]~q ;
wire \gen_dsp_only:m_ac|auto_generated|dffe3a[5]~q ;
wire \gen_dsp_only:m_bd|auto_generated|dffe3a[5]~q ;
wire \gen_dsp_only:m_ac|auto_generated|dffe3a[4]~q ;
wire \gen_dsp_only:m_bd|auto_generated|dffe3a[4]~q ;
wire \gen_dsp_only:m_ac|auto_generated|dffe3a[3]~q ;
wire \gen_dsp_only:m_bd|auto_generated|dffe3a[3]~q ;
wire \gen_dsp_only:m_ac|auto_generated|dffe3a[2]~q ;
wire \gen_dsp_only:m_bd|auto_generated|dffe3a[2]~q ;
wire \gen_dsp_only:m_ac|auto_generated|dffe3a[1]~q ;
wire \gen_dsp_only:m_bd|auto_generated|dffe3a[1]~q ;
wire \gen_dsp_only:m_ac|auto_generated|dffe3a[0]~q ;
wire \gen_dsp_only:m_bd|auto_generated|dffe3a[0]~q ;
wire \gen_dsp_only:m_ac|auto_generated|dffe3a[15]~q ;
wire \gen_dsp_only:m_bd|auto_generated|dffe3a[15]~q ;
wire \gen_dsp_only:m_ac|auto_generated|dffe3a[14]~q ;
wire \gen_dsp_only:m_bd|auto_generated|dffe3a[14]~q ;
wire \gen_dsp_only:m_ac|auto_generated|dffe3a[13]~q ;
wire \gen_dsp_only:m_bd|auto_generated|dffe3a[13]~q ;
wire \gen_dsp_only:m_ac|auto_generated|dffe3a[12]~q ;
wire \gen_dsp_only:m_bd|auto_generated|dffe3a[12]~q ;


fft_asj_fft_pround_fft_120_1 \gen_unsc:u1 (
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_14(pipeline_dffe_14),
	.result_imag_1_11(\result_imag_1[11]~q ),
	.result_imag_1_10(\result_imag_1[10]~q ),
	.result_imag_1_9(\result_imag_1[9]~q ),
	.result_imag_1_8(\result_imag_1[8]~q ),
	.result_imag_1_7(\result_imag_1[7]~q ),
	.result_imag_1_6(\result_imag_1[6]~q ),
	.result_imag_1_5(\result_imag_1[5]~q ),
	.result_imag_1_4(\result_imag_1[4]~q ),
	.result_imag_1_3(\result_imag_1[3]~q ),
	.result_imag_1_2(\result_imag_1[2]~q ),
	.result_imag_1_1(\result_imag_1[1]~q ),
	.result_imag_1_0(\result_imag_1[0]~q ),
	.result_imag_1_15(\result_imag_1[15]~q ),
	.result_imag_1_14(\result_imag_1[14]~q ),
	.result_imag_1_13(\result_imag_1[13]~q ),
	.result_imag_1_12(\result_imag_1[12]~q ),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_10(pipeline_dffe_10),
	.global_clock_enable(global_clock_enable),
	.clk(clk));

fft_asj_fft_pround_fft_120 \gen_unsc:u0 (
	.pipeline_dffe_11(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_15(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_12(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_13(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ),
	.pipeline_dffe_14(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ),
	.result_real_1_tmp_11(\result_real_1_tmp[11]~q ),
	.result_real_1_tmp_10(\result_real_1_tmp[10]~q ),
	.result_real_1_tmp_9(\result_real_1_tmp[9]~q ),
	.result_real_1_tmp_8(\result_real_1_tmp[8]~q ),
	.result_real_1_tmp_7(\result_real_1_tmp[7]~q ),
	.result_real_1_tmp_6(\result_real_1_tmp[6]~q ),
	.result_real_1_tmp_5(\result_real_1_tmp[5]~q ),
	.result_real_1_tmp_4(\result_real_1_tmp[4]~q ),
	.result_real_1_tmp_3(\result_real_1_tmp[3]~q ),
	.result_real_1_tmp_2(\result_real_1_tmp[2]~q ),
	.result_real_1_tmp_1(\result_real_1_tmp[1]~q ),
	.result_real_1_tmp_0(\result_real_1_tmp[0]~q ),
	.result_real_1_tmp_15(\result_real_1_tmp[15]~q ),
	.result_real_1_tmp_14(\result_real_1_tmp[14]~q ),
	.result_real_1_tmp_13(\result_real_1_tmp[13]~q ),
	.result_real_1_tmp_12(\result_real_1_tmp[12]~q ),
	.pipeline_dffe_9(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_8(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_10(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ),
	.global_clock_enable(global_clock_enable),
	.clk(clk));

fft_LPM_MULT_1 \gen_dsp_only:m_a_b_c_d (
	.dataa({\addresult_a_b[8]~q ,\addresult_a_b[7]~q ,\addresult_a_b[6]~q ,\addresult_a_b[5]~q ,\addresult_a_b[4]~q ,\addresult_a_b[3]~q ,\addresult_a_b[2]~q ,\addresult_a_b[1]~q ,\addresult_a_b[0]~q }),
	.datab({\addresult_c_d[8]~q ,\addresult_c_d[7]~q ,\addresult_c_d[6]~q ,\addresult_c_d[5]~q ,\addresult_c_d[4]~q ,\addresult_c_d[3]~q ,\addresult_c_d[2]~q ,\addresult_c_d[1]~q ,\addresult_c_d[0]~q }),
	.clken(global_clock_enable),
	.dffe3a_11(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[11]~q ),
	.dffe3a_10(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[10]~q ),
	.dffe3a_9(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[9]~q ),
	.dffe3a_8(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[8]~q ),
	.dffe3a_7(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[7]~q ),
	.dffe3a_6(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[6]~q ),
	.dffe3a_5(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[5]~q ),
	.dffe3a_4(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[4]~q ),
	.dffe3a_3(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[3]~q ),
	.dffe3a_2(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[2]~q ),
	.dffe3a_1(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[1]~q ),
	.dffe3a_0(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[0]~q ),
	.dffe3a_15(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[15]~q ),
	.dffe3a_14(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[14]~q ),
	.dffe3a_13(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[13]~q ),
	.dffe3a_12(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[12]~q ),
	.clock(clk));

fft_LPM_MULT_3 \gen_dsp_only:m_bd (
	.dataa({gnd,pipeline_dffe_92,pipeline_dffe_82,pipeline_dffe_71,pipeline_dffe_61,pipeline_dffe_51,pipeline_dffe_41,pipeline_dffe_31,pipeline_dffe_21}),
	.clken(global_clock_enable),
	.dffe3a_11(\gen_dsp_only:m_bd|auto_generated|dffe3a[11]~q ),
	.dffe3a_10(\gen_dsp_only:m_bd|auto_generated|dffe3a[10]~q ),
	.dffe3a_9(\gen_dsp_only:m_bd|auto_generated|dffe3a[9]~q ),
	.dffe3a_8(\gen_dsp_only:m_bd|auto_generated|dffe3a[8]~q ),
	.dffe3a_7(\gen_dsp_only:m_bd|auto_generated|dffe3a[7]~q ),
	.dffe3a_6(\gen_dsp_only:m_bd|auto_generated|dffe3a[6]~q ),
	.dffe3a_5(\gen_dsp_only:m_bd|auto_generated|dffe3a[5]~q ),
	.dffe3a_4(\gen_dsp_only:m_bd|auto_generated|dffe3a[4]~q ),
	.dffe3a_3(\gen_dsp_only:m_bd|auto_generated|dffe3a[3]~q ),
	.dffe3a_2(\gen_dsp_only:m_bd|auto_generated|dffe3a[2]~q ),
	.dffe3a_1(\gen_dsp_only:m_bd|auto_generated|dffe3a[1]~q ),
	.dffe3a_0(\gen_dsp_only:m_bd|auto_generated|dffe3a[0]~q ),
	.dffe3a_15(\gen_dsp_only:m_bd|auto_generated|dffe3a[15]~q ),
	.dffe3a_14(\gen_dsp_only:m_bd|auto_generated|dffe3a[14]~q ),
	.dffe3a_13(\gen_dsp_only:m_bd|auto_generated|dffe3a[13]~q ),
	.dffe3a_12(\gen_dsp_only:m_bd|auto_generated|dffe3a[12]~q ),
	.datab({gnd,twiddle_data017,twiddle_data016,twiddle_data015,twiddle_data014,twiddle_data013,twiddle_data012,twiddle_data011,twiddle_data010}),
	.clock(clk));

fft_LPM_MULT_2 \gen_dsp_only:m_ac (
	.dataa({gnd,pipeline_dffe_91,pipeline_dffe_81,pipeline_dffe_7,pipeline_dffe_6,pipeline_dffe_5,pipeline_dffe_4,pipeline_dffe_3,pipeline_dffe_2}),
	.clken(global_clock_enable),
	.dffe3a_11(\gen_dsp_only:m_ac|auto_generated|dffe3a[11]~q ),
	.dffe3a_10(\gen_dsp_only:m_ac|auto_generated|dffe3a[10]~q ),
	.dffe3a_9(\gen_dsp_only:m_ac|auto_generated|dffe3a[9]~q ),
	.dffe3a_8(\gen_dsp_only:m_ac|auto_generated|dffe3a[8]~q ),
	.dffe3a_7(\gen_dsp_only:m_ac|auto_generated|dffe3a[7]~q ),
	.dffe3a_6(\gen_dsp_only:m_ac|auto_generated|dffe3a[6]~q ),
	.dffe3a_5(\gen_dsp_only:m_ac|auto_generated|dffe3a[5]~q ),
	.dffe3a_4(\gen_dsp_only:m_ac|auto_generated|dffe3a[4]~q ),
	.dffe3a_3(\gen_dsp_only:m_ac|auto_generated|dffe3a[3]~q ),
	.dffe3a_2(\gen_dsp_only:m_ac|auto_generated|dffe3a[2]~q ),
	.dffe3a_1(\gen_dsp_only:m_ac|auto_generated|dffe3a[1]~q ),
	.dffe3a_0(\gen_dsp_only:m_ac|auto_generated|dffe3a[0]~q ),
	.dffe3a_15(\gen_dsp_only:m_ac|auto_generated|dffe3a[15]~q ),
	.dffe3a_14(\gen_dsp_only:m_ac|auto_generated|dffe3a[14]~q ),
	.dffe3a_13(\gen_dsp_only:m_ac|auto_generated|dffe3a[13]~q ),
	.dffe3a_12(\gen_dsp_only:m_ac|auto_generated|dffe3a[12]~q ),
	.datab({gnd,twiddle_data007,twiddle_data006,twiddle_data005,twiddle_data004,twiddle_data003,twiddle_data002,twiddle_data001,twiddle_data000}),
	.clock(clk));

dffeas \result_imag_1[11] (
	.clk(clk),
	.d(\result_imag_1[11]~38_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[11]~q ),
	.prn(vcc));
defparam \result_imag_1[11] .is_wysiwyg = "true";
defparam \result_imag_1[11] .power_up = "low";

dffeas \result_imag_1[10] (
	.clk(clk),
	.d(\result_imag_1[10]~36_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[10]~q ),
	.prn(vcc));
defparam \result_imag_1[10] .is_wysiwyg = "true";
defparam \result_imag_1[10] .power_up = "low";

dffeas \result_imag_1[9] (
	.clk(clk),
	.d(\result_imag_1[9]~34_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[9]~q ),
	.prn(vcc));
defparam \result_imag_1[9] .is_wysiwyg = "true";
defparam \result_imag_1[9] .power_up = "low";

dffeas \result_imag_1[8] (
	.clk(clk),
	.d(\result_imag_1[8]~32_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[8]~q ),
	.prn(vcc));
defparam \result_imag_1[8] .is_wysiwyg = "true";
defparam \result_imag_1[8] .power_up = "low";

dffeas \result_imag_1[7] (
	.clk(clk),
	.d(\result_imag_1[7]~30_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[7]~q ),
	.prn(vcc));
defparam \result_imag_1[7] .is_wysiwyg = "true";
defparam \result_imag_1[7] .power_up = "low";

dffeas \result_imag_1[6] (
	.clk(clk),
	.d(\result_imag_1[6]~28_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[6]~q ),
	.prn(vcc));
defparam \result_imag_1[6] .is_wysiwyg = "true";
defparam \result_imag_1[6] .power_up = "low";

dffeas \result_imag_1[5] (
	.clk(clk),
	.d(\result_imag_1[5]~26_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[5]~q ),
	.prn(vcc));
defparam \result_imag_1[5] .is_wysiwyg = "true";
defparam \result_imag_1[5] .power_up = "low";

dffeas \result_imag_1[4] (
	.clk(clk),
	.d(\result_imag_1[4]~24_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[4]~q ),
	.prn(vcc));
defparam \result_imag_1[4] .is_wysiwyg = "true";
defparam \result_imag_1[4] .power_up = "low";

dffeas \result_imag_1[3] (
	.clk(clk),
	.d(\result_imag_1[3]~22_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[3]~q ),
	.prn(vcc));
defparam \result_imag_1[3] .is_wysiwyg = "true";
defparam \result_imag_1[3] .power_up = "low";

dffeas \result_imag_1[2] (
	.clk(clk),
	.d(\result_imag_1[2]~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[2]~q ),
	.prn(vcc));
defparam \result_imag_1[2] .is_wysiwyg = "true";
defparam \result_imag_1[2] .power_up = "low";

dffeas \result_imag_1[1] (
	.clk(clk),
	.d(\result_imag_1[1]~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[1]~q ),
	.prn(vcc));
defparam \result_imag_1[1] .is_wysiwyg = "true";
defparam \result_imag_1[1] .power_up = "low";

dffeas \result_imag_1[0] (
	.clk(clk),
	.d(\result_imag_1[0]~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[0]~q ),
	.prn(vcc));
defparam \result_imag_1[0] .is_wysiwyg = "true";
defparam \result_imag_1[0] .power_up = "low";

dffeas \result_imag_1[15] (
	.clk(clk),
	.d(\result_imag_1[15]~46_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[15]~q ),
	.prn(vcc));
defparam \result_imag_1[15] .is_wysiwyg = "true";
defparam \result_imag_1[15] .power_up = "low";

dffeas \result_imag_1[14] (
	.clk(clk),
	.d(\result_imag_1[14]~44_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[14]~q ),
	.prn(vcc));
defparam \result_imag_1[14] .is_wysiwyg = "true";
defparam \result_imag_1[14] .power_up = "low";

dffeas \result_imag_1[13] (
	.clk(clk),
	.d(\result_imag_1[13]~42_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[13]~q ),
	.prn(vcc));
defparam \result_imag_1[13] .is_wysiwyg = "true";
defparam \result_imag_1[13] .power_up = "low";

dffeas \result_imag_1[12] (
	.clk(clk),
	.d(\result_imag_1[12]~40_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[12]~q ),
	.prn(vcc));
defparam \result_imag_1[12] .is_wysiwyg = "true";
defparam \result_imag_1[12] .power_up = "low";

dffeas \addresult_ac_bd[11] (
	.clk(clk),
	.d(\addresult_ac_bd[11]~38_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[11]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[11] .is_wysiwyg = "true";
defparam \addresult_ac_bd[11] .power_up = "low";

dffeas \addresult_ac_bd[10] (
	.clk(clk),
	.d(\addresult_ac_bd[10]~36_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[10]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[10] .is_wysiwyg = "true";
defparam \addresult_ac_bd[10] .power_up = "low";

dffeas \addresult_ac_bd[9] (
	.clk(clk),
	.d(\addresult_ac_bd[9]~34_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[9]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[9] .is_wysiwyg = "true";
defparam \addresult_ac_bd[9] .power_up = "low";

dffeas \addresult_ac_bd[8] (
	.clk(clk),
	.d(\addresult_ac_bd[8]~32_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[8]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[8] .is_wysiwyg = "true";
defparam \addresult_ac_bd[8] .power_up = "low";

dffeas \addresult_ac_bd[7] (
	.clk(clk),
	.d(\addresult_ac_bd[7]~30_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[7]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[7] .is_wysiwyg = "true";
defparam \addresult_ac_bd[7] .power_up = "low";

dffeas \addresult_ac_bd[6] (
	.clk(clk),
	.d(\addresult_ac_bd[6]~28_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[6]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[6] .is_wysiwyg = "true";
defparam \addresult_ac_bd[6] .power_up = "low";

dffeas \addresult_ac_bd[5] (
	.clk(clk),
	.d(\addresult_ac_bd[5]~26_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[5]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[5] .is_wysiwyg = "true";
defparam \addresult_ac_bd[5] .power_up = "low";

dffeas \addresult_ac_bd[4] (
	.clk(clk),
	.d(\addresult_ac_bd[4]~24_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[4]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[4] .is_wysiwyg = "true";
defparam \addresult_ac_bd[4] .power_up = "low";

dffeas \addresult_ac_bd[3] (
	.clk(clk),
	.d(\addresult_ac_bd[3]~22_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[3]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[3] .is_wysiwyg = "true";
defparam \addresult_ac_bd[3] .power_up = "low";

dffeas \addresult_ac_bd[2] (
	.clk(clk),
	.d(\addresult_ac_bd[2]~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[2]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[2] .is_wysiwyg = "true";
defparam \addresult_ac_bd[2] .power_up = "low";

dffeas \addresult_ac_bd[1] (
	.clk(clk),
	.d(\addresult_ac_bd[1]~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[1]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[1] .is_wysiwyg = "true";
defparam \addresult_ac_bd[1] .power_up = "low";

dffeas \addresult_ac_bd[0] (
	.clk(clk),
	.d(\addresult_ac_bd[0]~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[0]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[0] .is_wysiwyg = "true";
defparam \addresult_ac_bd[0] .power_up = "low";

cycloneiii_lcell_comb \result_imag_1[0]~16 (
	.dataa(\addresult_ac_bd[0]~q ),
	.datab(\result_a_b_c_d_se[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\result_imag_1[0]~16_combout ),
	.cout(\result_imag_1[0]~17 ));
defparam \result_imag_1[0]~16 .lut_mask = 16'h66DD;
defparam \result_imag_1[0]~16 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \result_imag_1[1]~18 (
	.dataa(\addresult_ac_bd[1]~q ),
	.datab(\result_a_b_c_d_se[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[0]~17 ),
	.combout(\result_imag_1[1]~18_combout ),
	.cout(\result_imag_1[1]~19 ));
defparam \result_imag_1[1]~18 .lut_mask = 16'h96BF;
defparam \result_imag_1[1]~18 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_imag_1[2]~20 (
	.dataa(\addresult_ac_bd[2]~q ),
	.datab(\result_a_b_c_d_se[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[1]~19 ),
	.combout(\result_imag_1[2]~20_combout ),
	.cout(\result_imag_1[2]~21 ));
defparam \result_imag_1[2]~20 .lut_mask = 16'h96DF;
defparam \result_imag_1[2]~20 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_imag_1[3]~22 (
	.dataa(\addresult_ac_bd[3]~q ),
	.datab(\result_a_b_c_d_se[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[2]~21 ),
	.combout(\result_imag_1[3]~22_combout ),
	.cout(\result_imag_1[3]~23 ));
defparam \result_imag_1[3]~22 .lut_mask = 16'h96BF;
defparam \result_imag_1[3]~22 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_imag_1[4]~24 (
	.dataa(\addresult_ac_bd[4]~q ),
	.datab(\result_a_b_c_d_se[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[3]~23 ),
	.combout(\result_imag_1[4]~24_combout ),
	.cout(\result_imag_1[4]~25 ));
defparam \result_imag_1[4]~24 .lut_mask = 16'h96DF;
defparam \result_imag_1[4]~24 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_imag_1[5]~26 (
	.dataa(\addresult_ac_bd[5]~q ),
	.datab(\result_a_b_c_d_se[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[4]~25 ),
	.combout(\result_imag_1[5]~26_combout ),
	.cout(\result_imag_1[5]~27 ));
defparam \result_imag_1[5]~26 .lut_mask = 16'h96BF;
defparam \result_imag_1[5]~26 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_imag_1[6]~28 (
	.dataa(\addresult_ac_bd[6]~q ),
	.datab(\result_a_b_c_d_se[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[5]~27 ),
	.combout(\result_imag_1[6]~28_combout ),
	.cout(\result_imag_1[6]~29 ));
defparam \result_imag_1[6]~28 .lut_mask = 16'h96DF;
defparam \result_imag_1[6]~28 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_imag_1[7]~30 (
	.dataa(\addresult_ac_bd[7]~q ),
	.datab(\result_a_b_c_d_se[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[6]~29 ),
	.combout(\result_imag_1[7]~30_combout ),
	.cout(\result_imag_1[7]~31 ));
defparam \result_imag_1[7]~30 .lut_mask = 16'h96BF;
defparam \result_imag_1[7]~30 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_imag_1[8]~32 (
	.dataa(\addresult_ac_bd[8]~q ),
	.datab(\result_a_b_c_d_se[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[7]~31 ),
	.combout(\result_imag_1[8]~32_combout ),
	.cout(\result_imag_1[8]~33 ));
defparam \result_imag_1[8]~32 .lut_mask = 16'h96DF;
defparam \result_imag_1[8]~32 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_imag_1[9]~34 (
	.dataa(\addresult_ac_bd[9]~q ),
	.datab(\result_a_b_c_d_se[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[8]~33 ),
	.combout(\result_imag_1[9]~34_combout ),
	.cout(\result_imag_1[9]~35 ));
defparam \result_imag_1[9]~34 .lut_mask = 16'h96BF;
defparam \result_imag_1[9]~34 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_imag_1[10]~36 (
	.dataa(\addresult_ac_bd[10]~q ),
	.datab(\result_a_b_c_d_se[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[9]~35 ),
	.combout(\result_imag_1[10]~36_combout ),
	.cout(\result_imag_1[10]~37 ));
defparam \result_imag_1[10]~36 .lut_mask = 16'h96DF;
defparam \result_imag_1[10]~36 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_imag_1[11]~38 (
	.dataa(\addresult_ac_bd[11]~q ),
	.datab(\result_a_b_c_d_se[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[10]~37 ),
	.combout(\result_imag_1[11]~38_combout ),
	.cout(\result_imag_1[11]~39 ));
defparam \result_imag_1[11]~38 .lut_mask = 16'h96BF;
defparam \result_imag_1[11]~38 .sum_lutc_input = "cin";

dffeas \addresult_ac_bd[15] (
	.clk(clk),
	.d(\addresult_ac_bd[15]~46_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[15]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[15] .is_wysiwyg = "true";
defparam \addresult_ac_bd[15] .power_up = "low";

dffeas \addresult_ac_bd[14] (
	.clk(clk),
	.d(\addresult_ac_bd[14]~44_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[14]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[14] .is_wysiwyg = "true";
defparam \addresult_ac_bd[14] .power_up = "low";

dffeas \addresult_ac_bd[13] (
	.clk(clk),
	.d(\addresult_ac_bd[13]~42_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[13]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[13] .is_wysiwyg = "true";
defparam \addresult_ac_bd[13] .power_up = "low";

dffeas \addresult_ac_bd[12] (
	.clk(clk),
	.d(\addresult_ac_bd[12]~40_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[12]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[12] .is_wysiwyg = "true";
defparam \addresult_ac_bd[12] .power_up = "low";

cycloneiii_lcell_comb \result_imag_1[12]~40 (
	.dataa(\addresult_ac_bd[12]~q ),
	.datab(\result_a_b_c_d_se[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[11]~39 ),
	.combout(\result_imag_1[12]~40_combout ),
	.cout(\result_imag_1[12]~41 ));
defparam \result_imag_1[12]~40 .lut_mask = 16'h96DF;
defparam \result_imag_1[12]~40 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_imag_1[13]~42 (
	.dataa(\addresult_ac_bd[13]~q ),
	.datab(\result_a_b_c_d_se[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[12]~41 ),
	.combout(\result_imag_1[13]~42_combout ),
	.cout(\result_imag_1[13]~43 ));
defparam \result_imag_1[13]~42 .lut_mask = 16'h96BF;
defparam \result_imag_1[13]~42 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_imag_1[14]~44 (
	.dataa(\addresult_ac_bd[14]~q ),
	.datab(\result_a_b_c_d_se[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[13]~43 ),
	.combout(\result_imag_1[14]~44_combout ),
	.cout(\result_imag_1[14]~45 ));
defparam \result_imag_1[14]~44 .lut_mask = 16'h96DF;
defparam \result_imag_1[14]~44 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_imag_1[15]~46 (
	.dataa(\addresult_ac_bd[15]~q ),
	.datab(\result_a_b_c_d_se[15]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\result_imag_1[14]~45 ),
	.combout(\result_imag_1[15]~46_combout ),
	.cout());
defparam \result_imag_1[15]~46 .lut_mask = 16'h9696;
defparam \result_imag_1[15]~46 .sum_lutc_input = "cin";

dffeas \result_real_1_tmp[11] (
	.clk(clk),
	.d(\result_real_1_tmp[11]~38_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[11]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[11] .is_wysiwyg = "true";
defparam \result_real_1_tmp[11] .power_up = "low";

dffeas \result_real_1_tmp[10] (
	.clk(clk),
	.d(\result_real_1_tmp[10]~36_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[10]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[10] .is_wysiwyg = "true";
defparam \result_real_1_tmp[10] .power_up = "low";

dffeas \result_real_1_tmp[9] (
	.clk(clk),
	.d(\result_real_1_tmp[9]~34_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[9]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[9] .is_wysiwyg = "true";
defparam \result_real_1_tmp[9] .power_up = "low";

dffeas \result_real_1_tmp[8] (
	.clk(clk),
	.d(\result_real_1_tmp[8]~32_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[8]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[8] .is_wysiwyg = "true";
defparam \result_real_1_tmp[8] .power_up = "low";

dffeas \result_real_1_tmp[7] (
	.clk(clk),
	.d(\result_real_1_tmp[7]~30_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[7]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[7] .is_wysiwyg = "true";
defparam \result_real_1_tmp[7] .power_up = "low";

dffeas \result_real_1_tmp[6] (
	.clk(clk),
	.d(\result_real_1_tmp[6]~28_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[6]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[6] .is_wysiwyg = "true";
defparam \result_real_1_tmp[6] .power_up = "low";

dffeas \result_real_1_tmp[5] (
	.clk(clk),
	.d(\result_real_1_tmp[5]~26_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[5]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[5] .is_wysiwyg = "true";
defparam \result_real_1_tmp[5] .power_up = "low";

dffeas \result_real_1_tmp[4] (
	.clk(clk),
	.d(\result_real_1_tmp[4]~24_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[4]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[4] .is_wysiwyg = "true";
defparam \result_real_1_tmp[4] .power_up = "low";

dffeas \result_real_1_tmp[3] (
	.clk(clk),
	.d(\result_real_1_tmp[3]~22_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[3]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[3] .is_wysiwyg = "true";
defparam \result_real_1_tmp[3] .power_up = "low";

dffeas \result_real_1_tmp[2] (
	.clk(clk),
	.d(\result_real_1_tmp[2]~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[2]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[2] .is_wysiwyg = "true";
defparam \result_real_1_tmp[2] .power_up = "low";

dffeas \result_real_1_tmp[1] (
	.clk(clk),
	.d(\result_real_1_tmp[1]~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[1]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[1] .is_wysiwyg = "true";
defparam \result_real_1_tmp[1] .power_up = "low";

dffeas \result_real_1_tmp[0] (
	.clk(clk),
	.d(\result_real_1_tmp[0]~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[0]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[0] .is_wysiwyg = "true";
defparam \result_real_1_tmp[0] .power_up = "low";

dffeas \result_real_1_tmp[15] (
	.clk(clk),
	.d(\result_real_1_tmp[15]~46_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[15]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[15] .is_wysiwyg = "true";
defparam \result_real_1_tmp[15] .power_up = "low";

dffeas \result_real_1_tmp[14] (
	.clk(clk),
	.d(\result_real_1_tmp[14]~44_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[14]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[14] .is_wysiwyg = "true";
defparam \result_real_1_tmp[14] .power_up = "low";

dffeas \result_real_1_tmp[13] (
	.clk(clk),
	.d(\result_real_1_tmp[13]~42_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[13]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[13] .is_wysiwyg = "true";
defparam \result_real_1_tmp[13] .power_up = "low";

dffeas \result_real_1_tmp[12] (
	.clk(clk),
	.d(\result_real_1_tmp[12]~40_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[12]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[12] .is_wysiwyg = "true";
defparam \result_real_1_tmp[12] .power_up = "low";

cycloneiii_lcell_comb \addresult_ac_bd[0]~16 (
	.dataa(\result_a_c_se[0]~q ),
	.datab(\result_b_d_se[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\addresult_ac_bd[0]~16_combout ),
	.cout(\addresult_ac_bd[0]~17 ));
defparam \addresult_ac_bd[0]~16 .lut_mask = 16'h66EE;
defparam \addresult_ac_bd[0]~16 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \addresult_ac_bd[1]~18 (
	.dataa(\result_a_c_se[1]~q ),
	.datab(\result_b_d_se[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[0]~17 ),
	.combout(\addresult_ac_bd[1]~18_combout ),
	.cout(\addresult_ac_bd[1]~19 ));
defparam \addresult_ac_bd[1]~18 .lut_mask = 16'h967F;
defparam \addresult_ac_bd[1]~18 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_ac_bd[2]~20 (
	.dataa(\result_a_c_se[2]~q ),
	.datab(\result_b_d_se[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[1]~19 ),
	.combout(\addresult_ac_bd[2]~20_combout ),
	.cout(\addresult_ac_bd[2]~21 ));
defparam \addresult_ac_bd[2]~20 .lut_mask = 16'h96EF;
defparam \addresult_ac_bd[2]~20 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_ac_bd[3]~22 (
	.dataa(\result_a_c_se[3]~q ),
	.datab(\result_b_d_se[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[2]~21 ),
	.combout(\addresult_ac_bd[3]~22_combout ),
	.cout(\addresult_ac_bd[3]~23 ));
defparam \addresult_ac_bd[3]~22 .lut_mask = 16'h967F;
defparam \addresult_ac_bd[3]~22 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_ac_bd[4]~24 (
	.dataa(\result_a_c_se[4]~q ),
	.datab(\result_b_d_se[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[3]~23 ),
	.combout(\addresult_ac_bd[4]~24_combout ),
	.cout(\addresult_ac_bd[4]~25 ));
defparam \addresult_ac_bd[4]~24 .lut_mask = 16'h96EF;
defparam \addresult_ac_bd[4]~24 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_ac_bd[5]~26 (
	.dataa(\result_a_c_se[5]~q ),
	.datab(\result_b_d_se[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[4]~25 ),
	.combout(\addresult_ac_bd[5]~26_combout ),
	.cout(\addresult_ac_bd[5]~27 ));
defparam \addresult_ac_bd[5]~26 .lut_mask = 16'h967F;
defparam \addresult_ac_bd[5]~26 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_ac_bd[6]~28 (
	.dataa(\result_a_c_se[6]~q ),
	.datab(\result_b_d_se[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[5]~27 ),
	.combout(\addresult_ac_bd[6]~28_combout ),
	.cout(\addresult_ac_bd[6]~29 ));
defparam \addresult_ac_bd[6]~28 .lut_mask = 16'h96EF;
defparam \addresult_ac_bd[6]~28 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_ac_bd[7]~30 (
	.dataa(\result_a_c_se[7]~q ),
	.datab(\result_b_d_se[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[6]~29 ),
	.combout(\addresult_ac_bd[7]~30_combout ),
	.cout(\addresult_ac_bd[7]~31 ));
defparam \addresult_ac_bd[7]~30 .lut_mask = 16'h967F;
defparam \addresult_ac_bd[7]~30 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_ac_bd[8]~32 (
	.dataa(\result_a_c_se[8]~q ),
	.datab(\result_b_d_se[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[7]~31 ),
	.combout(\addresult_ac_bd[8]~32_combout ),
	.cout(\addresult_ac_bd[8]~33 ));
defparam \addresult_ac_bd[8]~32 .lut_mask = 16'h96EF;
defparam \addresult_ac_bd[8]~32 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_ac_bd[9]~34 (
	.dataa(\result_a_c_se[9]~q ),
	.datab(\result_b_d_se[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[8]~33 ),
	.combout(\addresult_ac_bd[9]~34_combout ),
	.cout(\addresult_ac_bd[9]~35 ));
defparam \addresult_ac_bd[9]~34 .lut_mask = 16'h967F;
defparam \addresult_ac_bd[9]~34 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_ac_bd[10]~36 (
	.dataa(\result_a_c_se[10]~q ),
	.datab(\result_b_d_se[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[9]~35 ),
	.combout(\addresult_ac_bd[10]~36_combout ),
	.cout(\addresult_ac_bd[10]~37 ));
defparam \addresult_ac_bd[10]~36 .lut_mask = 16'h96EF;
defparam \addresult_ac_bd[10]~36 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_ac_bd[11]~38 (
	.dataa(\result_a_c_se[11]~q ),
	.datab(\result_b_d_se[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[10]~37 ),
	.combout(\addresult_ac_bd[11]~38_combout ),
	.cout(\addresult_ac_bd[11]~39 ));
defparam \addresult_ac_bd[11]~38 .lut_mask = 16'h967F;
defparam \addresult_ac_bd[11]~38 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_ac_bd[12]~40 (
	.dataa(\result_a_c_se[12]~q ),
	.datab(\result_b_d_se[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[11]~39 ),
	.combout(\addresult_ac_bd[12]~40_combout ),
	.cout(\addresult_ac_bd[12]~41 ));
defparam \addresult_ac_bd[12]~40 .lut_mask = 16'h96EF;
defparam \addresult_ac_bd[12]~40 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_ac_bd[13]~42 (
	.dataa(\result_a_c_se[13]~q ),
	.datab(\result_b_d_se[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[12]~41 ),
	.combout(\addresult_ac_bd[13]~42_combout ),
	.cout(\addresult_ac_bd[13]~43 ));
defparam \addresult_ac_bd[13]~42 .lut_mask = 16'h967F;
defparam \addresult_ac_bd[13]~42 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_ac_bd[14]~44 (
	.dataa(\result_a_c_se[14]~q ),
	.datab(\result_b_d_se[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[13]~43 ),
	.combout(\addresult_ac_bd[14]~44_combout ),
	.cout(\addresult_ac_bd[14]~45 ));
defparam \addresult_ac_bd[14]~44 .lut_mask = 16'h96EF;
defparam \addresult_ac_bd[14]~44 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_ac_bd[15]~46 (
	.dataa(\result_a_c_se[15]~q ),
	.datab(\result_b_d_se[15]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\addresult_ac_bd[14]~45 ),
	.combout(\addresult_ac_bd[15]~46_combout ),
	.cout());
defparam \addresult_ac_bd[15]~46 .lut_mask = 16'h9696;
defparam \addresult_ac_bd[15]~46 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_real_1_tmp[0]~16 (
	.dataa(\result_a_c_se[0]~q ),
	.datab(\result_b_d_se[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\result_real_1_tmp[0]~16_combout ),
	.cout(\result_real_1_tmp[0]~17 ));
defparam \result_real_1_tmp[0]~16 .lut_mask = 16'h66BB;
defparam \result_real_1_tmp[0]~16 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \result_real_1_tmp[1]~18 (
	.dataa(\result_a_c_se[1]~q ),
	.datab(\result_b_d_se[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[0]~17 ),
	.combout(\result_real_1_tmp[1]~18_combout ),
	.cout(\result_real_1_tmp[1]~19 ));
defparam \result_real_1_tmp[1]~18 .lut_mask = 16'h96DF;
defparam \result_real_1_tmp[1]~18 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_real_1_tmp[2]~20 (
	.dataa(\result_a_c_se[2]~q ),
	.datab(\result_b_d_se[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[1]~19 ),
	.combout(\result_real_1_tmp[2]~20_combout ),
	.cout(\result_real_1_tmp[2]~21 ));
defparam \result_real_1_tmp[2]~20 .lut_mask = 16'h96BF;
defparam \result_real_1_tmp[2]~20 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_real_1_tmp[3]~22 (
	.dataa(\result_a_c_se[3]~q ),
	.datab(\result_b_d_se[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[2]~21 ),
	.combout(\result_real_1_tmp[3]~22_combout ),
	.cout(\result_real_1_tmp[3]~23 ));
defparam \result_real_1_tmp[3]~22 .lut_mask = 16'h96DF;
defparam \result_real_1_tmp[3]~22 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_real_1_tmp[4]~24 (
	.dataa(\result_a_c_se[4]~q ),
	.datab(\result_b_d_se[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[3]~23 ),
	.combout(\result_real_1_tmp[4]~24_combout ),
	.cout(\result_real_1_tmp[4]~25 ));
defparam \result_real_1_tmp[4]~24 .lut_mask = 16'h96BF;
defparam \result_real_1_tmp[4]~24 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_real_1_tmp[5]~26 (
	.dataa(\result_a_c_se[5]~q ),
	.datab(\result_b_d_se[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[4]~25 ),
	.combout(\result_real_1_tmp[5]~26_combout ),
	.cout(\result_real_1_tmp[5]~27 ));
defparam \result_real_1_tmp[5]~26 .lut_mask = 16'h96DF;
defparam \result_real_1_tmp[5]~26 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_real_1_tmp[6]~28 (
	.dataa(\result_a_c_se[6]~q ),
	.datab(\result_b_d_se[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[5]~27 ),
	.combout(\result_real_1_tmp[6]~28_combout ),
	.cout(\result_real_1_tmp[6]~29 ));
defparam \result_real_1_tmp[6]~28 .lut_mask = 16'h96BF;
defparam \result_real_1_tmp[6]~28 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_real_1_tmp[7]~30 (
	.dataa(\result_a_c_se[7]~q ),
	.datab(\result_b_d_se[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[6]~29 ),
	.combout(\result_real_1_tmp[7]~30_combout ),
	.cout(\result_real_1_tmp[7]~31 ));
defparam \result_real_1_tmp[7]~30 .lut_mask = 16'h96DF;
defparam \result_real_1_tmp[7]~30 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_real_1_tmp[8]~32 (
	.dataa(\result_a_c_se[8]~q ),
	.datab(\result_b_d_se[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[7]~31 ),
	.combout(\result_real_1_tmp[8]~32_combout ),
	.cout(\result_real_1_tmp[8]~33 ));
defparam \result_real_1_tmp[8]~32 .lut_mask = 16'h96BF;
defparam \result_real_1_tmp[8]~32 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_real_1_tmp[9]~34 (
	.dataa(\result_a_c_se[9]~q ),
	.datab(\result_b_d_se[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[8]~33 ),
	.combout(\result_real_1_tmp[9]~34_combout ),
	.cout(\result_real_1_tmp[9]~35 ));
defparam \result_real_1_tmp[9]~34 .lut_mask = 16'h96DF;
defparam \result_real_1_tmp[9]~34 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_real_1_tmp[10]~36 (
	.dataa(\result_a_c_se[10]~q ),
	.datab(\result_b_d_se[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[9]~35 ),
	.combout(\result_real_1_tmp[10]~36_combout ),
	.cout(\result_real_1_tmp[10]~37 ));
defparam \result_real_1_tmp[10]~36 .lut_mask = 16'h96BF;
defparam \result_real_1_tmp[10]~36 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_real_1_tmp[11]~38 (
	.dataa(\result_a_c_se[11]~q ),
	.datab(\result_b_d_se[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[10]~37 ),
	.combout(\result_real_1_tmp[11]~38_combout ),
	.cout(\result_real_1_tmp[11]~39 ));
defparam \result_real_1_tmp[11]~38 .lut_mask = 16'h96DF;
defparam \result_real_1_tmp[11]~38 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_real_1_tmp[12]~40 (
	.dataa(\result_a_c_se[12]~q ),
	.datab(\result_b_d_se[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[11]~39 ),
	.combout(\result_real_1_tmp[12]~40_combout ),
	.cout(\result_real_1_tmp[12]~41 ));
defparam \result_real_1_tmp[12]~40 .lut_mask = 16'h96BF;
defparam \result_real_1_tmp[12]~40 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_real_1_tmp[13]~42 (
	.dataa(\result_a_c_se[13]~q ),
	.datab(\result_b_d_se[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[12]~41 ),
	.combout(\result_real_1_tmp[13]~42_combout ),
	.cout(\result_real_1_tmp[13]~43 ));
defparam \result_real_1_tmp[13]~42 .lut_mask = 16'h96DF;
defparam \result_real_1_tmp[13]~42 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_real_1_tmp[14]~44 (
	.dataa(\result_a_c_se[14]~q ),
	.datab(\result_b_d_se[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[13]~43 ),
	.combout(\result_real_1_tmp[14]~44_combout ),
	.cout(\result_real_1_tmp[14]~45 ));
defparam \result_real_1_tmp[14]~44 .lut_mask = 16'h96BF;
defparam \result_real_1_tmp[14]~44 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_real_1_tmp[15]~46 (
	.dataa(\result_a_c_se[15]~q ),
	.datab(\result_b_d_se[15]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\result_real_1_tmp[14]~45 ),
	.combout(\result_real_1_tmp[15]~46_combout ),
	.cout());
defparam \result_real_1_tmp[15]~46 .lut_mask = 16'h9696;
defparam \result_real_1_tmp[15]~46 .sum_lutc_input = "cin";

dffeas \addresult_a_b[0] (
	.clk(clk),
	.d(\addresult_a_b[0]~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_a_b[0]~q ),
	.prn(vcc));
defparam \addresult_a_b[0] .is_wysiwyg = "true";
defparam \addresult_a_b[0] .power_up = "low";

dffeas \addresult_a_b[1] (
	.clk(clk),
	.d(\addresult_a_b[1]~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_a_b[1]~q ),
	.prn(vcc));
defparam \addresult_a_b[1] .is_wysiwyg = "true";
defparam \addresult_a_b[1] .power_up = "low";

dffeas \addresult_a_b[2] (
	.clk(clk),
	.d(\addresult_a_b[2]~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_a_b[2]~q ),
	.prn(vcc));
defparam \addresult_a_b[2] .is_wysiwyg = "true";
defparam \addresult_a_b[2] .power_up = "low";

dffeas \addresult_a_b[3] (
	.clk(clk),
	.d(\addresult_a_b[3]~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_a_b[3]~q ),
	.prn(vcc));
defparam \addresult_a_b[3] .is_wysiwyg = "true";
defparam \addresult_a_b[3] .power_up = "low";

dffeas \addresult_a_b[4] (
	.clk(clk),
	.d(\addresult_a_b[4]~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_a_b[4]~q ),
	.prn(vcc));
defparam \addresult_a_b[4] .is_wysiwyg = "true";
defparam \addresult_a_b[4] .power_up = "low";

dffeas \addresult_a_b[5] (
	.clk(clk),
	.d(\addresult_a_b[5]~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_a_b[5]~q ),
	.prn(vcc));
defparam \addresult_a_b[5] .is_wysiwyg = "true";
defparam \addresult_a_b[5] .power_up = "low";

dffeas \addresult_a_b[6] (
	.clk(clk),
	.d(\addresult_a_b[6]~21_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_a_b[6]~q ),
	.prn(vcc));
defparam \addresult_a_b[6] .is_wysiwyg = "true";
defparam \addresult_a_b[6] .power_up = "low";

dffeas \addresult_a_b[7] (
	.clk(clk),
	.d(\addresult_a_b[7]~23_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_a_b[7]~q ),
	.prn(vcc));
defparam \addresult_a_b[7] .is_wysiwyg = "true";
defparam \addresult_a_b[7] .power_up = "low";

dffeas \addresult_a_b[8] (
	.clk(clk),
	.d(\addresult_a_b[8]~25_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_a_b[8]~q ),
	.prn(vcc));
defparam \addresult_a_b[8] .is_wysiwyg = "true";
defparam \addresult_a_b[8] .power_up = "low";

dffeas \addresult_c_d[0] (
	.clk(clk),
	.d(\addresult_c_d[0]~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_c_d[0]~q ),
	.prn(vcc));
defparam \addresult_c_d[0] .is_wysiwyg = "true";
defparam \addresult_c_d[0] .power_up = "low";

dffeas \addresult_c_d[1] (
	.clk(clk),
	.d(\addresult_c_d[1]~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_c_d[1]~q ),
	.prn(vcc));
defparam \addresult_c_d[1] .is_wysiwyg = "true";
defparam \addresult_c_d[1] .power_up = "low";

dffeas \addresult_c_d[2] (
	.clk(clk),
	.d(\addresult_c_d[2]~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_c_d[2]~q ),
	.prn(vcc));
defparam \addresult_c_d[2] .is_wysiwyg = "true";
defparam \addresult_c_d[2] .power_up = "low";

dffeas \addresult_c_d[3] (
	.clk(clk),
	.d(\addresult_c_d[3]~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_c_d[3]~q ),
	.prn(vcc));
defparam \addresult_c_d[3] .is_wysiwyg = "true";
defparam \addresult_c_d[3] .power_up = "low";

dffeas \addresult_c_d[4] (
	.clk(clk),
	.d(\addresult_c_d[4]~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_c_d[4]~q ),
	.prn(vcc));
defparam \addresult_c_d[4] .is_wysiwyg = "true";
defparam \addresult_c_d[4] .power_up = "low";

dffeas \addresult_c_d[5] (
	.clk(clk),
	.d(\addresult_c_d[5]~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_c_d[5]~q ),
	.prn(vcc));
defparam \addresult_c_d[5] .is_wysiwyg = "true";
defparam \addresult_c_d[5] .power_up = "low";

dffeas \addresult_c_d[6] (
	.clk(clk),
	.d(\addresult_c_d[6]~21_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_c_d[6]~q ),
	.prn(vcc));
defparam \addresult_c_d[6] .is_wysiwyg = "true";
defparam \addresult_c_d[6] .power_up = "low";

dffeas \addresult_c_d[7] (
	.clk(clk),
	.d(\addresult_c_d[7]~23_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_c_d[7]~q ),
	.prn(vcc));
defparam \addresult_c_d[7] .is_wysiwyg = "true";
defparam \addresult_c_d[7] .power_up = "low";

dffeas \addresult_c_d[8] (
	.clk(clk),
	.d(\addresult_c_d[8]~25_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_c_d[8]~q ),
	.prn(vcc));
defparam \addresult_c_d[8] .is_wysiwyg = "true";
defparam \addresult_c_d[8] .power_up = "low";

cycloneiii_lcell_comb \addresult_a_b[0]~9 (
	.dataa(pipeline_dffe_2),
	.datab(pipeline_dffe_21),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\addresult_a_b[0]~9_combout ),
	.cout(\addresult_a_b[0]~10 ));
defparam \addresult_a_b[0]~9 .lut_mask = 16'h66EE;
defparam \addresult_a_b[0]~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \addresult_a_b[1]~11 (
	.dataa(pipeline_dffe_3),
	.datab(pipeline_dffe_31),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_a_b[0]~10 ),
	.combout(\addresult_a_b[1]~11_combout ),
	.cout(\addresult_a_b[1]~12 ));
defparam \addresult_a_b[1]~11 .lut_mask = 16'h967F;
defparam \addresult_a_b[1]~11 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_a_b[2]~13 (
	.dataa(pipeline_dffe_4),
	.datab(pipeline_dffe_41),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_a_b[1]~12 ),
	.combout(\addresult_a_b[2]~13_combout ),
	.cout(\addresult_a_b[2]~14 ));
defparam \addresult_a_b[2]~13 .lut_mask = 16'h96EF;
defparam \addresult_a_b[2]~13 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_a_b[3]~15 (
	.dataa(pipeline_dffe_5),
	.datab(pipeline_dffe_51),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_a_b[2]~14 ),
	.combout(\addresult_a_b[3]~15_combout ),
	.cout(\addresult_a_b[3]~16 ));
defparam \addresult_a_b[3]~15 .lut_mask = 16'h967F;
defparam \addresult_a_b[3]~15 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_a_b[4]~17 (
	.dataa(pipeline_dffe_6),
	.datab(pipeline_dffe_61),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_a_b[3]~16 ),
	.combout(\addresult_a_b[4]~17_combout ),
	.cout(\addresult_a_b[4]~18 ));
defparam \addresult_a_b[4]~17 .lut_mask = 16'h96EF;
defparam \addresult_a_b[4]~17 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_a_b[5]~19 (
	.dataa(pipeline_dffe_7),
	.datab(pipeline_dffe_71),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_a_b[4]~18 ),
	.combout(\addresult_a_b[5]~19_combout ),
	.cout(\addresult_a_b[5]~20 ));
defparam \addresult_a_b[5]~19 .lut_mask = 16'h967F;
defparam \addresult_a_b[5]~19 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_a_b[6]~21 (
	.dataa(pipeline_dffe_81),
	.datab(pipeline_dffe_82),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_a_b[5]~20 ),
	.combout(\addresult_a_b[6]~21_combout ),
	.cout(\addresult_a_b[6]~22 ));
defparam \addresult_a_b[6]~21 .lut_mask = 16'h96EF;
defparam \addresult_a_b[6]~21 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_a_b[7]~23 (
	.dataa(pipeline_dffe_91),
	.datab(pipeline_dffe_92),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_a_b[6]~22 ),
	.combout(\addresult_a_b[7]~23_combout ),
	.cout(\addresult_a_b[7]~24 ));
defparam \addresult_a_b[7]~23 .lut_mask = 16'h967F;
defparam \addresult_a_b[7]~23 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_a_b[8]~25 (
	.dataa(pipeline_dffe_91),
	.datab(pipeline_dffe_92),
	.datac(gnd),
	.datad(gnd),
	.cin(\addresult_a_b[7]~24 ),
	.combout(\addresult_a_b[8]~25_combout ),
	.cout());
defparam \addresult_a_b[8]~25 .lut_mask = 16'h9696;
defparam \addresult_a_b[8]~25 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_c_d[0]~9 (
	.dataa(twiddle_data000),
	.datab(twiddle_data010),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\addresult_c_d[0]~9_combout ),
	.cout(\addresult_c_d[0]~10 ));
defparam \addresult_c_d[0]~9 .lut_mask = 16'h66EE;
defparam \addresult_c_d[0]~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \addresult_c_d[1]~11 (
	.dataa(twiddle_data001),
	.datab(twiddle_data011),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_c_d[0]~10 ),
	.combout(\addresult_c_d[1]~11_combout ),
	.cout(\addresult_c_d[1]~12 ));
defparam \addresult_c_d[1]~11 .lut_mask = 16'h967F;
defparam \addresult_c_d[1]~11 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_c_d[2]~13 (
	.dataa(twiddle_data002),
	.datab(twiddle_data012),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_c_d[1]~12 ),
	.combout(\addresult_c_d[2]~13_combout ),
	.cout(\addresult_c_d[2]~14 ));
defparam \addresult_c_d[2]~13 .lut_mask = 16'h96EF;
defparam \addresult_c_d[2]~13 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_c_d[3]~15 (
	.dataa(twiddle_data003),
	.datab(twiddle_data013),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_c_d[2]~14 ),
	.combout(\addresult_c_d[3]~15_combout ),
	.cout(\addresult_c_d[3]~16 ));
defparam \addresult_c_d[3]~15 .lut_mask = 16'h967F;
defparam \addresult_c_d[3]~15 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_c_d[4]~17 (
	.dataa(twiddle_data004),
	.datab(twiddle_data014),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_c_d[3]~16 ),
	.combout(\addresult_c_d[4]~17_combout ),
	.cout(\addresult_c_d[4]~18 ));
defparam \addresult_c_d[4]~17 .lut_mask = 16'h96EF;
defparam \addresult_c_d[4]~17 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_c_d[5]~19 (
	.dataa(twiddle_data005),
	.datab(twiddle_data015),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_c_d[4]~18 ),
	.combout(\addresult_c_d[5]~19_combout ),
	.cout(\addresult_c_d[5]~20 ));
defparam \addresult_c_d[5]~19 .lut_mask = 16'h967F;
defparam \addresult_c_d[5]~19 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_c_d[6]~21 (
	.dataa(twiddle_data006),
	.datab(twiddle_data016),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_c_d[5]~20 ),
	.combout(\addresult_c_d[6]~21_combout ),
	.cout(\addresult_c_d[6]~22 ));
defparam \addresult_c_d[6]~21 .lut_mask = 16'h96EF;
defparam \addresult_c_d[6]~21 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_c_d[7]~23 (
	.dataa(twiddle_data007),
	.datab(twiddle_data017),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_c_d[6]~22 ),
	.combout(\addresult_c_d[7]~23_combout ),
	.cout(\addresult_c_d[7]~24 ));
defparam \addresult_c_d[7]~23 .lut_mask = 16'h967F;
defparam \addresult_c_d[7]~23 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_c_d[8]~25 (
	.dataa(twiddle_data007),
	.datab(twiddle_data017),
	.datac(gnd),
	.datad(gnd),
	.cin(\addresult_c_d[7]~24 ),
	.combout(\addresult_c_d[8]~25_combout ),
	.cout());
defparam \addresult_c_d[8]~25 .lut_mask = 16'h9696;
defparam \addresult_c_d[8]~25 .sum_lutc_input = "cin";

dffeas \result_a_b_c_d_se[11] (
	.clk(clk),
	.d(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[11]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[11] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[11] .power_up = "low";

dffeas \result_a_b_c_d_se[10] (
	.clk(clk),
	.d(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[10]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[10] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[10] .power_up = "low";

dffeas \result_a_b_c_d_se[9] (
	.clk(clk),
	.d(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[9]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[9] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[9] .power_up = "low";

dffeas \result_a_b_c_d_se[8] (
	.clk(clk),
	.d(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[8]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[8] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[8] .power_up = "low";

dffeas \result_a_b_c_d_se[7] (
	.clk(clk),
	.d(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[7]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[7] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[7] .power_up = "low";

dffeas \result_a_b_c_d_se[6] (
	.clk(clk),
	.d(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[6]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[6] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[6] .power_up = "low";

dffeas \result_a_b_c_d_se[5] (
	.clk(clk),
	.d(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[5]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[5] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[5] .power_up = "low";

dffeas \result_a_b_c_d_se[4] (
	.clk(clk),
	.d(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[4]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[4] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[4] .power_up = "low";

dffeas \result_a_b_c_d_se[3] (
	.clk(clk),
	.d(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[3]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[3] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[3] .power_up = "low";

dffeas \result_a_b_c_d_se[2] (
	.clk(clk),
	.d(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[2]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[2] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[2] .power_up = "low";

dffeas \result_a_b_c_d_se[1] (
	.clk(clk),
	.d(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[1]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[1] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[1] .power_up = "low";

dffeas \result_a_b_c_d_se[0] (
	.clk(clk),
	.d(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[0]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[0] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[0] .power_up = "low";

dffeas \result_a_b_c_d_se[15] (
	.clk(clk),
	.d(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[15]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[15] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[15] .power_up = "low";

dffeas \result_a_b_c_d_se[14] (
	.clk(clk),
	.d(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[14]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[14] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[14] .power_up = "low";

dffeas \result_a_b_c_d_se[13] (
	.clk(clk),
	.d(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[13]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[13] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[13] .power_up = "low";

dffeas \result_a_b_c_d_se[12] (
	.clk(clk),
	.d(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[12]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[12] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[12] .power_up = "low";

dffeas \result_a_c_se[11] (
	.clk(clk),
	.d(\gen_dsp_only:m_ac|auto_generated|dffe3a[11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[11]~q ),
	.prn(vcc));
defparam \result_a_c_se[11] .is_wysiwyg = "true";
defparam \result_a_c_se[11] .power_up = "low";

dffeas \result_b_d_se[11] (
	.clk(clk),
	.d(\gen_dsp_only:m_bd|auto_generated|dffe3a[11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[11]~q ),
	.prn(vcc));
defparam \result_b_d_se[11] .is_wysiwyg = "true";
defparam \result_b_d_se[11] .power_up = "low";

dffeas \result_a_c_se[10] (
	.clk(clk),
	.d(\gen_dsp_only:m_ac|auto_generated|dffe3a[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[10]~q ),
	.prn(vcc));
defparam \result_a_c_se[10] .is_wysiwyg = "true";
defparam \result_a_c_se[10] .power_up = "low";

dffeas \result_b_d_se[10] (
	.clk(clk),
	.d(\gen_dsp_only:m_bd|auto_generated|dffe3a[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[10]~q ),
	.prn(vcc));
defparam \result_b_d_se[10] .is_wysiwyg = "true";
defparam \result_b_d_se[10] .power_up = "low";

dffeas \result_a_c_se[9] (
	.clk(clk),
	.d(\gen_dsp_only:m_ac|auto_generated|dffe3a[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[9]~q ),
	.prn(vcc));
defparam \result_a_c_se[9] .is_wysiwyg = "true";
defparam \result_a_c_se[9] .power_up = "low";

dffeas \result_b_d_se[9] (
	.clk(clk),
	.d(\gen_dsp_only:m_bd|auto_generated|dffe3a[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[9]~q ),
	.prn(vcc));
defparam \result_b_d_se[9] .is_wysiwyg = "true";
defparam \result_b_d_se[9] .power_up = "low";

dffeas \result_a_c_se[8] (
	.clk(clk),
	.d(\gen_dsp_only:m_ac|auto_generated|dffe3a[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[8]~q ),
	.prn(vcc));
defparam \result_a_c_se[8] .is_wysiwyg = "true";
defparam \result_a_c_se[8] .power_up = "low";

dffeas \result_b_d_se[8] (
	.clk(clk),
	.d(\gen_dsp_only:m_bd|auto_generated|dffe3a[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[8]~q ),
	.prn(vcc));
defparam \result_b_d_se[8] .is_wysiwyg = "true";
defparam \result_b_d_se[8] .power_up = "low";

dffeas \result_a_c_se[7] (
	.clk(clk),
	.d(\gen_dsp_only:m_ac|auto_generated|dffe3a[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[7]~q ),
	.prn(vcc));
defparam \result_a_c_se[7] .is_wysiwyg = "true";
defparam \result_a_c_se[7] .power_up = "low";

dffeas \result_b_d_se[7] (
	.clk(clk),
	.d(\gen_dsp_only:m_bd|auto_generated|dffe3a[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[7]~q ),
	.prn(vcc));
defparam \result_b_d_se[7] .is_wysiwyg = "true";
defparam \result_b_d_se[7] .power_up = "low";

dffeas \result_a_c_se[6] (
	.clk(clk),
	.d(\gen_dsp_only:m_ac|auto_generated|dffe3a[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[6]~q ),
	.prn(vcc));
defparam \result_a_c_se[6] .is_wysiwyg = "true";
defparam \result_a_c_se[6] .power_up = "low";

dffeas \result_b_d_se[6] (
	.clk(clk),
	.d(\gen_dsp_only:m_bd|auto_generated|dffe3a[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[6]~q ),
	.prn(vcc));
defparam \result_b_d_se[6] .is_wysiwyg = "true";
defparam \result_b_d_se[6] .power_up = "low";

dffeas \result_a_c_se[5] (
	.clk(clk),
	.d(\gen_dsp_only:m_ac|auto_generated|dffe3a[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[5]~q ),
	.prn(vcc));
defparam \result_a_c_se[5] .is_wysiwyg = "true";
defparam \result_a_c_se[5] .power_up = "low";

dffeas \result_b_d_se[5] (
	.clk(clk),
	.d(\gen_dsp_only:m_bd|auto_generated|dffe3a[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[5]~q ),
	.prn(vcc));
defparam \result_b_d_se[5] .is_wysiwyg = "true";
defparam \result_b_d_se[5] .power_up = "low";

dffeas \result_a_c_se[4] (
	.clk(clk),
	.d(\gen_dsp_only:m_ac|auto_generated|dffe3a[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[4]~q ),
	.prn(vcc));
defparam \result_a_c_se[4] .is_wysiwyg = "true";
defparam \result_a_c_se[4] .power_up = "low";

dffeas \result_b_d_se[4] (
	.clk(clk),
	.d(\gen_dsp_only:m_bd|auto_generated|dffe3a[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[4]~q ),
	.prn(vcc));
defparam \result_b_d_se[4] .is_wysiwyg = "true";
defparam \result_b_d_se[4] .power_up = "low";

dffeas \result_a_c_se[3] (
	.clk(clk),
	.d(\gen_dsp_only:m_ac|auto_generated|dffe3a[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[3]~q ),
	.prn(vcc));
defparam \result_a_c_se[3] .is_wysiwyg = "true";
defparam \result_a_c_se[3] .power_up = "low";

dffeas \result_b_d_se[3] (
	.clk(clk),
	.d(\gen_dsp_only:m_bd|auto_generated|dffe3a[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[3]~q ),
	.prn(vcc));
defparam \result_b_d_se[3] .is_wysiwyg = "true";
defparam \result_b_d_se[3] .power_up = "low";

dffeas \result_a_c_se[2] (
	.clk(clk),
	.d(\gen_dsp_only:m_ac|auto_generated|dffe3a[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[2]~q ),
	.prn(vcc));
defparam \result_a_c_se[2] .is_wysiwyg = "true";
defparam \result_a_c_se[2] .power_up = "low";

dffeas \result_b_d_se[2] (
	.clk(clk),
	.d(\gen_dsp_only:m_bd|auto_generated|dffe3a[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[2]~q ),
	.prn(vcc));
defparam \result_b_d_se[2] .is_wysiwyg = "true";
defparam \result_b_d_se[2] .power_up = "low";

dffeas \result_a_c_se[1] (
	.clk(clk),
	.d(\gen_dsp_only:m_ac|auto_generated|dffe3a[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[1]~q ),
	.prn(vcc));
defparam \result_a_c_se[1] .is_wysiwyg = "true";
defparam \result_a_c_se[1] .power_up = "low";

dffeas \result_b_d_se[1] (
	.clk(clk),
	.d(\gen_dsp_only:m_bd|auto_generated|dffe3a[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[1]~q ),
	.prn(vcc));
defparam \result_b_d_se[1] .is_wysiwyg = "true";
defparam \result_b_d_se[1] .power_up = "low";

dffeas \result_a_c_se[0] (
	.clk(clk),
	.d(\gen_dsp_only:m_ac|auto_generated|dffe3a[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[0]~q ),
	.prn(vcc));
defparam \result_a_c_se[0] .is_wysiwyg = "true";
defparam \result_a_c_se[0] .power_up = "low";

dffeas \result_b_d_se[0] (
	.clk(clk),
	.d(\gen_dsp_only:m_bd|auto_generated|dffe3a[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[0]~q ),
	.prn(vcc));
defparam \result_b_d_se[0] .is_wysiwyg = "true";
defparam \result_b_d_se[0] .power_up = "low";

dffeas \result_a_c_se[15] (
	.clk(clk),
	.d(\gen_dsp_only:m_ac|auto_generated|dffe3a[15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[15]~q ),
	.prn(vcc));
defparam \result_a_c_se[15] .is_wysiwyg = "true";
defparam \result_a_c_se[15] .power_up = "low";

dffeas \result_b_d_se[15] (
	.clk(clk),
	.d(\gen_dsp_only:m_bd|auto_generated|dffe3a[15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[15]~q ),
	.prn(vcc));
defparam \result_b_d_se[15] .is_wysiwyg = "true";
defparam \result_b_d_se[15] .power_up = "low";

dffeas \result_a_c_se[14] (
	.clk(clk),
	.d(\gen_dsp_only:m_ac|auto_generated|dffe3a[14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[14]~q ),
	.prn(vcc));
defparam \result_a_c_se[14] .is_wysiwyg = "true";
defparam \result_a_c_se[14] .power_up = "low";

dffeas \result_b_d_se[14] (
	.clk(clk),
	.d(\gen_dsp_only:m_bd|auto_generated|dffe3a[14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[14]~q ),
	.prn(vcc));
defparam \result_b_d_se[14] .is_wysiwyg = "true";
defparam \result_b_d_se[14] .power_up = "low";

dffeas \result_a_c_se[13] (
	.clk(clk),
	.d(\gen_dsp_only:m_ac|auto_generated|dffe3a[13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[13]~q ),
	.prn(vcc));
defparam \result_a_c_se[13] .is_wysiwyg = "true";
defparam \result_a_c_se[13] .power_up = "low";

dffeas \result_b_d_se[13] (
	.clk(clk),
	.d(\gen_dsp_only:m_bd|auto_generated|dffe3a[13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[13]~q ),
	.prn(vcc));
defparam \result_b_d_se[13] .is_wysiwyg = "true";
defparam \result_b_d_se[13] .power_up = "low";

dffeas \result_a_c_se[12] (
	.clk(clk),
	.d(\gen_dsp_only:m_ac|auto_generated|dffe3a[12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[12]~q ),
	.prn(vcc));
defparam \result_a_c_se[12] .is_wysiwyg = "true";
defparam \result_a_c_se[12] .power_up = "low";

dffeas \result_b_d_se[12] (
	.clk(clk),
	.d(\gen_dsp_only:m_bd|auto_generated|dffe3a[12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[12]~q ),
	.prn(vcc));
defparam \result_b_d_se[12] .is_wysiwyg = "true";
defparam \result_b_d_se[12] .power_up = "low";

dffeas \real_out[3] (
	.clk(clk),
	.d(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(real_out_3),
	.prn(vcc));
defparam \real_out[3] .is_wysiwyg = "true";
defparam \real_out[3] .power_up = "low";

dffeas \real_out[7] (
	.clk(clk),
	.d(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(real_out_7),
	.prn(vcc));
defparam \real_out[7] .is_wysiwyg = "true";
defparam \real_out[7] .power_up = "low";

dffeas \real_out[4] (
	.clk(clk),
	.d(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(real_out_4),
	.prn(vcc));
defparam \real_out[4] .is_wysiwyg = "true";
defparam \real_out[4] .power_up = "low";

dffeas \real_out[5] (
	.clk(clk),
	.d(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(real_out_5),
	.prn(vcc));
defparam \real_out[5] .is_wysiwyg = "true";
defparam \real_out[5] .power_up = "low";

dffeas \real_out[6] (
	.clk(clk),
	.d(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(real_out_6),
	.prn(vcc));
defparam \real_out[6] .is_wysiwyg = "true";
defparam \real_out[6] .power_up = "low";

dffeas \real_out[1] (
	.clk(clk),
	.d(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(real_out_1),
	.prn(vcc));
defparam \real_out[1] .is_wysiwyg = "true";
defparam \real_out[1] .power_up = "low";

dffeas \real_out[0] (
	.clk(clk),
	.d(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(real_out_0),
	.prn(vcc));
defparam \real_out[0] .is_wysiwyg = "true";
defparam \real_out[0] .power_up = "low";

dffeas \real_out[2] (
	.clk(clk),
	.d(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(real_out_2),
	.prn(vcc));
defparam \real_out[2] .is_wysiwyg = "true";
defparam \real_out[2] .power_up = "low";

endmodule

module fft_asj_fft_pround_fft_120 (
	pipeline_dffe_11,
	pipeline_dffe_15,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	result_real_1_tmp_11,
	result_real_1_tmp_10,
	result_real_1_tmp_9,
	result_real_1_tmp_8,
	result_real_1_tmp_7,
	result_real_1_tmp_6,
	result_real_1_tmp_5,
	result_real_1_tmp_4,
	result_real_1_tmp_3,
	result_real_1_tmp_2,
	result_real_1_tmp_1,
	result_real_1_tmp_0,
	result_real_1_tmp_15,
	result_real_1_tmp_14,
	result_real_1_tmp_13,
	result_real_1_tmp_12,
	pipeline_dffe_9,
	pipeline_dffe_8,
	pipeline_dffe_10,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_11;
output 	pipeline_dffe_15;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
input 	result_real_1_tmp_11;
input 	result_real_1_tmp_10;
input 	result_real_1_tmp_9;
input 	result_real_1_tmp_8;
input 	result_real_1_tmp_7;
input 	result_real_1_tmp_6;
input 	result_real_1_tmp_5;
input 	result_real_1_tmp_4;
input 	result_real_1_tmp_3;
input 	result_real_1_tmp_2;
input 	result_real_1_tmp_1;
input 	result_real_1_tmp_0;
input 	result_real_1_tmp_15;
input 	result_real_1_tmp_14;
input 	result_real_1_tmp_13;
input 	result_real_1_tmp_12;
output 	pipeline_dffe_9;
output 	pipeline_dffe_8;
output 	pipeline_dffe_10;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_LPM_ADD_SUB_1 \gbrnd:nev:gp:lpm_add_sub_component (
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_14(pipeline_dffe_14),
	.result_real_1_tmp_11(result_real_1_tmp_11),
	.result_real_1_tmp_10(result_real_1_tmp_10),
	.result_real_1_tmp_9(result_real_1_tmp_9),
	.result_real_1_tmp_8(result_real_1_tmp_8),
	.result_real_1_tmp_7(result_real_1_tmp_7),
	.result_real_1_tmp_6(result_real_1_tmp_6),
	.result_real_1_tmp_5(result_real_1_tmp_5),
	.result_real_1_tmp_4(result_real_1_tmp_4),
	.result_real_1_tmp_3(result_real_1_tmp_3),
	.result_real_1_tmp_2(result_real_1_tmp_2),
	.result_real_1_tmp_1(result_real_1_tmp_1),
	.result_real_1_tmp_0(result_real_1_tmp_0),
	.result_real_1_tmp_15(result_real_1_tmp_15),
	.result_real_1_tmp_14(result_real_1_tmp_14),
	.result_real_1_tmp_13(result_real_1_tmp_13),
	.result_real_1_tmp_12(result_real_1_tmp_12),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_10(pipeline_dffe_10),
	.clken(global_clock_enable),
	.clock(clk));

endmodule

module fft_LPM_ADD_SUB_1 (
	pipeline_dffe_11,
	pipeline_dffe_15,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	result_real_1_tmp_11,
	result_real_1_tmp_10,
	result_real_1_tmp_9,
	result_real_1_tmp_8,
	result_real_1_tmp_7,
	result_real_1_tmp_6,
	result_real_1_tmp_5,
	result_real_1_tmp_4,
	result_real_1_tmp_3,
	result_real_1_tmp_2,
	result_real_1_tmp_1,
	result_real_1_tmp_0,
	result_real_1_tmp_15,
	result_real_1_tmp_14,
	result_real_1_tmp_13,
	result_real_1_tmp_12,
	pipeline_dffe_9,
	pipeline_dffe_8,
	pipeline_dffe_10,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_11;
output 	pipeline_dffe_15;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
input 	result_real_1_tmp_11;
input 	result_real_1_tmp_10;
input 	result_real_1_tmp_9;
input 	result_real_1_tmp_8;
input 	result_real_1_tmp_7;
input 	result_real_1_tmp_6;
input 	result_real_1_tmp_5;
input 	result_real_1_tmp_4;
input 	result_real_1_tmp_3;
input 	result_real_1_tmp_2;
input 	result_real_1_tmp_1;
input 	result_real_1_tmp_0;
input 	result_real_1_tmp_15;
input 	result_real_1_tmp_14;
input 	result_real_1_tmp_13;
input 	result_real_1_tmp_12;
output 	pipeline_dffe_9;
output 	pipeline_dffe_8;
output 	pipeline_dffe_10;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_add_sub_dmj auto_generated(
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_14(pipeline_dffe_14),
	.result_real_1_tmp_11(result_real_1_tmp_11),
	.result_real_1_tmp_10(result_real_1_tmp_10),
	.result_real_1_tmp_9(result_real_1_tmp_9),
	.result_real_1_tmp_8(result_real_1_tmp_8),
	.result_real_1_tmp_7(result_real_1_tmp_7),
	.result_real_1_tmp_6(result_real_1_tmp_6),
	.result_real_1_tmp_5(result_real_1_tmp_5),
	.result_real_1_tmp_4(result_real_1_tmp_4),
	.result_real_1_tmp_3(result_real_1_tmp_3),
	.result_real_1_tmp_2(result_real_1_tmp_2),
	.result_real_1_tmp_1(result_real_1_tmp_1),
	.result_real_1_tmp_0(result_real_1_tmp_0),
	.result_real_1_tmp_15(result_real_1_tmp_15),
	.result_real_1_tmp_14(result_real_1_tmp_14),
	.result_real_1_tmp_13(result_real_1_tmp_13),
	.result_real_1_tmp_12(result_real_1_tmp_12),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_10(pipeline_dffe_10),
	.clken(clken),
	.clock(clock));

endmodule

module fft_add_sub_dmj (
	pipeline_dffe_11,
	pipeline_dffe_15,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	result_real_1_tmp_11,
	result_real_1_tmp_10,
	result_real_1_tmp_9,
	result_real_1_tmp_8,
	result_real_1_tmp_7,
	result_real_1_tmp_6,
	result_real_1_tmp_5,
	result_real_1_tmp_4,
	result_real_1_tmp_3,
	result_real_1_tmp_2,
	result_real_1_tmp_1,
	result_real_1_tmp_0,
	result_real_1_tmp_15,
	result_real_1_tmp_14,
	result_real_1_tmp_13,
	result_real_1_tmp_12,
	pipeline_dffe_9,
	pipeline_dffe_8,
	pipeline_dffe_10,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_11;
output 	pipeline_dffe_15;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
input 	result_real_1_tmp_11;
input 	result_real_1_tmp_10;
input 	result_real_1_tmp_9;
input 	result_real_1_tmp_8;
input 	result_real_1_tmp_7;
input 	result_real_1_tmp_6;
input 	result_real_1_tmp_5;
input 	result_real_1_tmp_4;
input 	result_real_1_tmp_3;
input 	result_real_1_tmp_2;
input 	result_real_1_tmp_1;
input 	result_real_1_tmp_0;
input 	result_real_1_tmp_15;
input 	result_real_1_tmp_14;
input 	result_real_1_tmp_13;
input 	result_real_1_tmp_12;
output 	pipeline_dffe_9;
output 	pipeline_dffe_8;
output 	pipeline_dffe_10;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~9_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~11_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~13_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~15_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~17_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~19_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~21_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~23_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~27 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~29 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~31 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~32_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~33 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~35 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~37 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~39 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~40_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~34_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~36_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~38_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~30_combout ;


dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_15),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_12),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_13),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_14),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .power_up = "low";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~9 (
	.dataa(result_real_1_tmp_15),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~9_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~9 .lut_mask = 16'h0055;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~11 (
	.dataa(result_real_1_tmp_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~9_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~11_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~11 .lut_mask = 16'h005F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~11 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~13 (
	.dataa(result_real_1_tmp_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~11_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~13_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~13 .lut_mask = 16'h00AF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~13 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~15 (
	.dataa(result_real_1_tmp_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~13_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~15_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~15 .lut_mask = 16'h005F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~15 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~17 (
	.dataa(result_real_1_tmp_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~15_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~17_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~17 .lut_mask = 16'h00AF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~17 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~19 (
	.dataa(result_real_1_tmp_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~17_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~19_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~19 .lut_mask = 16'h005F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~19 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~21 (
	.dataa(result_real_1_tmp_5),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~19_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~21_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~21 .lut_mask = 16'h00AF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~21 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~23 (
	.dataa(result_real_1_tmp_6),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~21_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~23_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~23 .lut_mask = 16'h005F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~23 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25 (
	.dataa(result_real_1_tmp_7),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~23_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25 .lut_mask = 16'h00AF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26 (
	.dataa(result_real_1_tmp_8),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25_cout ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~27 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28 (
	.dataa(result_real_1_tmp_9),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~27 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~29 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28 .lut_mask = 16'h5AAF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~30 (
	.dataa(result_real_1_tmp_10),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~29 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~30_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~31 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~30 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~30 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~32 (
	.dataa(result_real_1_tmp_11),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~31 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~32_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~33 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~32 .lut_mask = 16'h5AAF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~32 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~34 (
	.dataa(result_real_1_tmp_12),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~33 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~34_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~35 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~34 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~34 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~36 (
	.dataa(result_real_1_tmp_13),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~35 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~36_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~37 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~36 .lut_mask = 16'h5AAF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~36 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~38 (
	.dataa(result_real_1_tmp_14),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~37 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~38_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~39 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~38 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~38 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~40 (
	.dataa(result_real_1_tmp_15),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~39 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~40_combout ),
	.cout());
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~40 .lut_mask = 16'h5A5A;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~40 .sum_lutc_input = "cin";

endmodule

module fft_asj_fft_pround_fft_120_1 (
	pipeline_dffe_11,
	pipeline_dffe_15,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	result_imag_1_11,
	result_imag_1_10,
	result_imag_1_9,
	result_imag_1_8,
	result_imag_1_7,
	result_imag_1_6,
	result_imag_1_5,
	result_imag_1_4,
	result_imag_1_3,
	result_imag_1_2,
	result_imag_1_1,
	result_imag_1_0,
	result_imag_1_15,
	result_imag_1_14,
	result_imag_1_13,
	result_imag_1_12,
	pipeline_dffe_9,
	pipeline_dffe_8,
	pipeline_dffe_10,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_11;
output 	pipeline_dffe_15;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
input 	result_imag_1_11;
input 	result_imag_1_10;
input 	result_imag_1_9;
input 	result_imag_1_8;
input 	result_imag_1_7;
input 	result_imag_1_6;
input 	result_imag_1_5;
input 	result_imag_1_4;
input 	result_imag_1_3;
input 	result_imag_1_2;
input 	result_imag_1_1;
input 	result_imag_1_0;
input 	result_imag_1_15;
input 	result_imag_1_14;
input 	result_imag_1_13;
input 	result_imag_1_12;
output 	pipeline_dffe_9;
output 	pipeline_dffe_8;
output 	pipeline_dffe_10;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_LPM_ADD_SUB_2 \gbrnd:nev:gp:lpm_add_sub_component (
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_14(pipeline_dffe_14),
	.result_imag_1_11(result_imag_1_11),
	.result_imag_1_10(result_imag_1_10),
	.result_imag_1_9(result_imag_1_9),
	.result_imag_1_8(result_imag_1_8),
	.result_imag_1_7(result_imag_1_7),
	.result_imag_1_6(result_imag_1_6),
	.result_imag_1_5(result_imag_1_5),
	.result_imag_1_4(result_imag_1_4),
	.result_imag_1_3(result_imag_1_3),
	.result_imag_1_2(result_imag_1_2),
	.result_imag_1_1(result_imag_1_1),
	.result_imag_1_0(result_imag_1_0),
	.result_imag_1_15(result_imag_1_15),
	.result_imag_1_14(result_imag_1_14),
	.result_imag_1_13(result_imag_1_13),
	.result_imag_1_12(result_imag_1_12),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_10(pipeline_dffe_10),
	.clken(global_clock_enable),
	.clock(clk));

endmodule

module fft_LPM_ADD_SUB_2 (
	pipeline_dffe_11,
	pipeline_dffe_15,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	result_imag_1_11,
	result_imag_1_10,
	result_imag_1_9,
	result_imag_1_8,
	result_imag_1_7,
	result_imag_1_6,
	result_imag_1_5,
	result_imag_1_4,
	result_imag_1_3,
	result_imag_1_2,
	result_imag_1_1,
	result_imag_1_0,
	result_imag_1_15,
	result_imag_1_14,
	result_imag_1_13,
	result_imag_1_12,
	pipeline_dffe_9,
	pipeline_dffe_8,
	pipeline_dffe_10,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_11;
output 	pipeline_dffe_15;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
input 	result_imag_1_11;
input 	result_imag_1_10;
input 	result_imag_1_9;
input 	result_imag_1_8;
input 	result_imag_1_7;
input 	result_imag_1_6;
input 	result_imag_1_5;
input 	result_imag_1_4;
input 	result_imag_1_3;
input 	result_imag_1_2;
input 	result_imag_1_1;
input 	result_imag_1_0;
input 	result_imag_1_15;
input 	result_imag_1_14;
input 	result_imag_1_13;
input 	result_imag_1_12;
output 	pipeline_dffe_9;
output 	pipeline_dffe_8;
output 	pipeline_dffe_10;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_add_sub_dmj_1 auto_generated(
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_14(pipeline_dffe_14),
	.result_imag_1_11(result_imag_1_11),
	.result_imag_1_10(result_imag_1_10),
	.result_imag_1_9(result_imag_1_9),
	.result_imag_1_8(result_imag_1_8),
	.result_imag_1_7(result_imag_1_7),
	.result_imag_1_6(result_imag_1_6),
	.result_imag_1_5(result_imag_1_5),
	.result_imag_1_4(result_imag_1_4),
	.result_imag_1_3(result_imag_1_3),
	.result_imag_1_2(result_imag_1_2),
	.result_imag_1_1(result_imag_1_1),
	.result_imag_1_0(result_imag_1_0),
	.result_imag_1_15(result_imag_1_15),
	.result_imag_1_14(result_imag_1_14),
	.result_imag_1_13(result_imag_1_13),
	.result_imag_1_12(result_imag_1_12),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_10(pipeline_dffe_10),
	.clken(clken),
	.clock(clock));

endmodule

module fft_add_sub_dmj_1 (
	pipeline_dffe_11,
	pipeline_dffe_15,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	result_imag_1_11,
	result_imag_1_10,
	result_imag_1_9,
	result_imag_1_8,
	result_imag_1_7,
	result_imag_1_6,
	result_imag_1_5,
	result_imag_1_4,
	result_imag_1_3,
	result_imag_1_2,
	result_imag_1_1,
	result_imag_1_0,
	result_imag_1_15,
	result_imag_1_14,
	result_imag_1_13,
	result_imag_1_12,
	pipeline_dffe_9,
	pipeline_dffe_8,
	pipeline_dffe_10,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_11;
output 	pipeline_dffe_15;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
input 	result_imag_1_11;
input 	result_imag_1_10;
input 	result_imag_1_9;
input 	result_imag_1_8;
input 	result_imag_1_7;
input 	result_imag_1_6;
input 	result_imag_1_5;
input 	result_imag_1_4;
input 	result_imag_1_3;
input 	result_imag_1_2;
input 	result_imag_1_1;
input 	result_imag_1_0;
input 	result_imag_1_15;
input 	result_imag_1_14;
input 	result_imag_1_13;
input 	result_imag_1_12;
output 	pipeline_dffe_9;
output 	pipeline_dffe_8;
output 	pipeline_dffe_10;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~9_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~11_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~13_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~15_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~17_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~19_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~21_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~23_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~27 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~29 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~31 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~32_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~33 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~35 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~37 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~39 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~40_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~34_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~36_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~38_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~30_combout ;


dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_15),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_12),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_13),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_14),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .power_up = "low";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~9 (
	.dataa(result_imag_1_15),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~9_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~9 .lut_mask = 16'h0055;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~11 (
	.dataa(result_imag_1_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~9_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~11_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~11 .lut_mask = 16'h005F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~11 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~13 (
	.dataa(result_imag_1_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~11_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~13_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~13 .lut_mask = 16'h00AF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~13 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~15 (
	.dataa(result_imag_1_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~13_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~15_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~15 .lut_mask = 16'h005F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~15 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~17 (
	.dataa(result_imag_1_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~15_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~17_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~17 .lut_mask = 16'h00AF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~17 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~19 (
	.dataa(result_imag_1_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~17_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~19_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~19 .lut_mask = 16'h005F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~19 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~21 (
	.dataa(result_imag_1_5),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~19_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~21_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~21 .lut_mask = 16'h00AF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~21 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~23 (
	.dataa(result_imag_1_6),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~21_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~23_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~23 .lut_mask = 16'h005F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~23 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25 (
	.dataa(result_imag_1_7),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~23_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25 .lut_mask = 16'h00AF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26 (
	.dataa(result_imag_1_8),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25_cout ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~27 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28 (
	.dataa(result_imag_1_9),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~27 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~29 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28 .lut_mask = 16'h5AAF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~30 (
	.dataa(result_imag_1_10),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~29 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~30_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~31 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~30 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~30 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~32 (
	.dataa(result_imag_1_11),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~31 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~32_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~33 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~32 .lut_mask = 16'h5AAF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~32 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~34 (
	.dataa(result_imag_1_12),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~33 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~34_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~35 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~34 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~34 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~36 (
	.dataa(result_imag_1_13),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~35 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~36_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~37 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~36 .lut_mask = 16'h5AAF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~36 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~38 (
	.dataa(result_imag_1_14),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~37 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~38_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~39 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~38 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~38 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~40 (
	.dataa(result_imag_1_15),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~39 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~40_combout ),
	.cout());
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~40 .lut_mask = 16'h5A5A;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~40 .sum_lutc_input = "cin";

endmodule

module fft_LPM_MULT_1 (
	dataa,
	datab,
	clken,
	dffe3a_11,
	dffe3a_10,
	dffe3a_9,
	dffe3a_8,
	dffe3a_7,
	dffe3a_6,
	dffe3a_5,
	dffe3a_4,
	dffe3a_3,
	dffe3a_2,
	dffe3a_1,
	dffe3a_0,
	dffe3a_15,
	dffe3a_14,
	dffe3a_13,
	dffe3a_12,
	clock)/* synthesis synthesis_greybox=1 */;
input 	[8:0] dataa;
input 	[8:0] datab;
input 	clken;
output 	dffe3a_11;
output 	dffe3a_10;
output 	dffe3a_9;
output 	dffe3a_8;
output 	dffe3a_7;
output 	dffe3a_6;
output 	dffe3a_5;
output 	dffe3a_4;
output 	dffe3a_3;
output 	dffe3a_2;
output 	dffe3a_1;
output 	dffe3a_0;
output 	dffe3a_15;
output 	dffe3a_14;
output 	dffe3a_13;
output 	dffe3a_12;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_mult_4p01 auto_generated(
	.dataa({dataa[8],dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.datab({datab[8],datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.clken(clken),
	.dffe3a_11(dffe3a_11),
	.dffe3a_10(dffe3a_10),
	.dffe3a_9(dffe3a_9),
	.dffe3a_8(dffe3a_8),
	.dffe3a_7(dffe3a_7),
	.dffe3a_6(dffe3a_6),
	.dffe3a_5(dffe3a_5),
	.dffe3a_4(dffe3a_4),
	.dffe3a_3(dffe3a_3),
	.dffe3a_2(dffe3a_2),
	.dffe3a_1(dffe3a_1),
	.dffe3a_0(dffe3a_0),
	.dffe3a_15(dffe3a_15),
	.dffe3a_14(dffe3a_14),
	.dffe3a_13(dffe3a_13),
	.dffe3a_12(dffe3a_12),
	.clock(clock));

endmodule

module fft_mult_4p01 (
	dataa,
	datab,
	clken,
	dffe3a_11,
	dffe3a_10,
	dffe3a_9,
	dffe3a_8,
	dffe3a_7,
	dffe3a_6,
	dffe3a_5,
	dffe3a_4,
	dffe3a_3,
	dffe3a_2,
	dffe3a_1,
	dffe3a_0,
	dffe3a_15,
	dffe3a_14,
	dffe3a_13,
	dffe3a_12,
	clock)/* synthesis synthesis_greybox=1 */;
input 	[8:0] dataa;
input 	[8:0] datab;
input 	clken;
output 	dffe3a_11;
output 	dffe3a_10;
output 	dffe3a_9;
output 	dffe3a_8;
output 	dffe3a_7;
output 	dffe3a_6;
output 	dffe3a_5;
output 	dffe3a_4;
output 	dffe3a_3;
output 	dffe3a_2;
output 	dffe3a_1;
output 	dffe3a_0;
output 	dffe3a_15;
output 	dffe3a_14;
output 	dffe3a_13;
output 	dffe3a_12;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT16 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT17 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~dataout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT1 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT2 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT3 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT4 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT5 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT6 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT7 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT8 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT9 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT10 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT11 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT12 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT13 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT14 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT15 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT16 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT17 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT11 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT10 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT9 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT8 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT7 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT6 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT5 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT4 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT3 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT2 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT1 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~dataout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT15 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT14 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT13 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT12 ;

wire [35:0] \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus ;
wire [35:0] \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus ;

assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~dataout  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [0];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT1  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [1];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT2  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [2];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT3  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [3];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT4  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [4];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT5  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [5];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT6  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [6];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT7  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [7];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT8  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [8];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT9  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [9];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT10  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [10];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT11  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [11];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT12  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [12];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT13  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [13];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT14  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [14];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT15  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [15];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT16  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [16];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT17  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [17];

assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~dataout  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [0];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT1  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [1];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT2  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [2];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT3  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [3];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT4  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [4];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT5  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [5];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT6  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [6];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT7  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [7];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT8  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [8];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT9  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [9];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT10  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [10];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT11  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [11];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT12  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [12];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT13  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [13];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT14  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [14];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT15  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [15];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT16  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [16];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT17  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [17];

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[11] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT11 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_11),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[11] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[11] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[10] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT10 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_10),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[10] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[10] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[9] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT9 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_9),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[9] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[9] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[8] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT8 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_8),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[8] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[8] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[7] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT7 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_7),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[7] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[7] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[6] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT6 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_6),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[6] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[6] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[5] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT5 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_5),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[5] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[5] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[4] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT4 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_4),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[4] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[4] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[3] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT3 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_3),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[3] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[3] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[2] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT2 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_2),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[2] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[2] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[1] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT1 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_1),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[1] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[1] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[0] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~dataout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_0),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[0] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[0] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[15] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT15 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_15),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[15] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[15] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[14] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT14 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_14),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[14] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[14] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[13] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT13 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_13),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[13] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[13] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[12] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT12 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_12),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[12] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[12] .power_up = "low";

cycloneiii_mac_mult \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1 (
	.signa(vcc),
	.signb(vcc),
	.clk(clock),
	.aclr(gnd),
	.ena(clken),
	.dataa({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dataa[8],dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.datab({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,datab[8],datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.dataout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1 .dataa_clock = "0";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1 .dataa_width = 9;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1 .datab_clock = "0";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1 .datab_width = 9;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1 .signa_clock = "none";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1 .signb_clock = "none";

cycloneiii_mac_out \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2 (
	.clk(clock),
	.aclr(gnd),
	.ena(clken),
	.dataa({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT17 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT16 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT15 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT14 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT13 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT12 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT11 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT10 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT9 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT8 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT7 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT6 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT5 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT4 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT3 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT2 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT1 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~dataout }),
	.dataout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2 .dataa_width = 18;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2 .output_clock = "0";

endmodule

module fft_LPM_MULT_2 (
	dataa,
	clken,
	dffe3a_11,
	dffe3a_10,
	dffe3a_9,
	dffe3a_8,
	dffe3a_7,
	dffe3a_6,
	dffe3a_5,
	dffe3a_4,
	dffe3a_3,
	dffe3a_2,
	dffe3a_1,
	dffe3a_0,
	dffe3a_15,
	dffe3a_14,
	dffe3a_13,
	dffe3a_12,
	datab,
	clock)/* synthesis synthesis_greybox=1 */;
input 	[8:0] dataa;
input 	clken;
output 	dffe3a_11;
output 	dffe3a_10;
output 	dffe3a_9;
output 	dffe3a_8;
output 	dffe3a_7;
output 	dffe3a_6;
output 	dffe3a_5;
output 	dffe3a_4;
output 	dffe3a_3;
output 	dffe3a_2;
output 	dffe3a_1;
output 	dffe3a_0;
output 	dffe3a_15;
output 	dffe3a_14;
output 	dffe3a_13;
output 	dffe3a_12;
input 	[8:0] datab;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_mult_0p01 auto_generated(
	.dataa({dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.clken(clken),
	.dffe3a_11(dffe3a_11),
	.dffe3a_10(dffe3a_10),
	.dffe3a_9(dffe3a_9),
	.dffe3a_8(dffe3a_8),
	.dffe3a_7(dffe3a_7),
	.dffe3a_6(dffe3a_6),
	.dffe3a_5(dffe3a_5),
	.dffe3a_4(dffe3a_4),
	.dffe3a_3(dffe3a_3),
	.dffe3a_2(dffe3a_2),
	.dffe3a_1(dffe3a_1),
	.dffe3a_0(dffe3a_0),
	.dffe3a_15(dffe3a_15),
	.dffe3a_14(dffe3a_14),
	.dffe3a_13(dffe3a_13),
	.dffe3a_12(dffe3a_12),
	.datab({datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.clock(clock));

endmodule

module fft_mult_0p01 (
	dataa,
	clken,
	dffe3a_11,
	dffe3a_10,
	dffe3a_9,
	dffe3a_8,
	dffe3a_7,
	dffe3a_6,
	dffe3a_5,
	dffe3a_4,
	dffe3a_3,
	dffe3a_2,
	dffe3a_1,
	dffe3a_0,
	dffe3a_15,
	dffe3a_14,
	dffe3a_13,
	dffe3a_12,
	datab,
	clock)/* synthesis synthesis_greybox=1 */;
input 	[7:0] dataa;
input 	clken;
output 	dffe3a_11;
output 	dffe3a_10;
output 	dffe3a_9;
output 	dffe3a_8;
output 	dffe3a_7;
output 	dffe3a_6;
output 	dffe3a_5;
output 	dffe3a_4;
output 	dffe3a_3;
output 	dffe3a_2;
output 	dffe3a_1;
output 	dffe3a_0;
output 	dffe3a_15;
output 	dffe3a_14;
output 	dffe3a_13;
output 	dffe3a_12;
input 	[7:0] datab;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1~dataout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT1 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT2 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT3 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT4 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT5 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT6 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT7 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT8 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT9 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT10 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT11 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT12 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT13 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT14 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT15 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT11 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT10 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT9 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT8 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT7 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT6 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT5 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT4 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT3 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT2 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT1 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2~dataout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT15 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT14 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT13 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT12 ;

wire [35:0] \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2_DATAOUT_bus ;
wire [35:0] \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1_DATAOUT_bus ;

assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2~dataout  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2_DATAOUT_bus [0];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT1  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2_DATAOUT_bus [1];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT2  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2_DATAOUT_bus [2];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT3  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2_DATAOUT_bus [3];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT4  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2_DATAOUT_bus [4];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT5  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2_DATAOUT_bus [5];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT6  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2_DATAOUT_bus [6];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT7  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2_DATAOUT_bus [7];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT8  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2_DATAOUT_bus [8];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT9  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2_DATAOUT_bus [9];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT10  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2_DATAOUT_bus [10];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT11  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2_DATAOUT_bus [11];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT12  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2_DATAOUT_bus [12];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT13  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2_DATAOUT_bus [13];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT14  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2_DATAOUT_bus [14];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT15  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2_DATAOUT_bus [15];

assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1~dataout  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1_DATAOUT_bus [0];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT1  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1_DATAOUT_bus [1];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT2  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1_DATAOUT_bus [2];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT3  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1_DATAOUT_bus [3];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT4  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1_DATAOUT_bus [4];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT5  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1_DATAOUT_bus [5];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT6  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1_DATAOUT_bus [6];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT7  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1_DATAOUT_bus [7];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT8  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1_DATAOUT_bus [8];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT9  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1_DATAOUT_bus [9];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT10  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1_DATAOUT_bus [10];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT11  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1_DATAOUT_bus [11];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT12  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1_DATAOUT_bus [12];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT13  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1_DATAOUT_bus [13];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT14  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1_DATAOUT_bus [14];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT15  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1_DATAOUT_bus [15];

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|dffe3a[11] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT11 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_11),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|dffe3a[11] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|dffe3a[11] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|dffe3a[10] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT10 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_10),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|dffe3a[10] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|dffe3a[10] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|dffe3a[9] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT9 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_9),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|dffe3a[9] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|dffe3a[9] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|dffe3a[8] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT8 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_8),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|dffe3a[8] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|dffe3a[8] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|dffe3a[7] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT7 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_7),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|dffe3a[7] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|dffe3a[7] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|dffe3a[6] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT6 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_6),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|dffe3a[6] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|dffe3a[6] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|dffe3a[5] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT5 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_5),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|dffe3a[5] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|dffe3a[5] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|dffe3a[4] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT4 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_4),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|dffe3a[4] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|dffe3a[4] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|dffe3a[3] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT3 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_3),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|dffe3a[3] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|dffe3a[3] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|dffe3a[2] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT2 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_2),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|dffe3a[2] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|dffe3a[2] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|dffe3a[1] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT1 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_1),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|dffe3a[1] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|dffe3a[1] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|dffe3a[0] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2~dataout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_0),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|dffe3a[0] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|dffe3a[0] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|dffe3a[15] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT15 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_15),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|dffe3a[15] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|dffe3a[15] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|dffe3a[14] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT14 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_14),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|dffe3a[14] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|dffe3a[14] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|dffe3a[13] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT13 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_13),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|dffe3a[13] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|dffe3a[13] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|dffe3a[12] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT12 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_12),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|dffe3a[12] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|dffe3a[12] .power_up = "low";

cycloneiii_mac_mult \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1 (
	.signa(vcc),
	.signb(vcc),
	.clk(clock),
	.aclr(gnd),
	.ena(clken),
	.dataa({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.datab({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.dataout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1_DATAOUT_bus ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1 .dataa_clock = "0";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1 .dataa_width = 8;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1 .datab_clock = "0";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1 .datab_width = 8;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1 .signa_clock = "none";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1 .signb_clock = "none";

cycloneiii_mac_out \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2 (
	.clk(clock),
	.aclr(gnd),
	.ena(clken),
	.dataa({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT15 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT14 ,\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT13 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT12 ,\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT11 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT10 ,\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT9 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT8 ,\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT7 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT6 ,\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT5 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT4 ,\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT3 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT2 ,\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT1 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_mult1~dataout }),
	.dataout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2_DATAOUT_bus ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2 .dataa_width = 16;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_ac|auto_generated|mac_out2 .output_clock = "0";

endmodule

module fft_LPM_MULT_3 (
	dataa,
	clken,
	dffe3a_11,
	dffe3a_10,
	dffe3a_9,
	dffe3a_8,
	dffe3a_7,
	dffe3a_6,
	dffe3a_5,
	dffe3a_4,
	dffe3a_3,
	dffe3a_2,
	dffe3a_1,
	dffe3a_0,
	dffe3a_15,
	dffe3a_14,
	dffe3a_13,
	dffe3a_12,
	datab,
	clock)/* synthesis synthesis_greybox=1 */;
input 	[8:0] dataa;
input 	clken;
output 	dffe3a_11;
output 	dffe3a_10;
output 	dffe3a_9;
output 	dffe3a_8;
output 	dffe3a_7;
output 	dffe3a_6;
output 	dffe3a_5;
output 	dffe3a_4;
output 	dffe3a_3;
output 	dffe3a_2;
output 	dffe3a_1;
output 	dffe3a_0;
output 	dffe3a_15;
output 	dffe3a_14;
output 	dffe3a_13;
output 	dffe3a_12;
input 	[8:0] datab;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_mult_0p01_1 auto_generated(
	.dataa({dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.clken(clken),
	.dffe3a_11(dffe3a_11),
	.dffe3a_10(dffe3a_10),
	.dffe3a_9(dffe3a_9),
	.dffe3a_8(dffe3a_8),
	.dffe3a_7(dffe3a_7),
	.dffe3a_6(dffe3a_6),
	.dffe3a_5(dffe3a_5),
	.dffe3a_4(dffe3a_4),
	.dffe3a_3(dffe3a_3),
	.dffe3a_2(dffe3a_2),
	.dffe3a_1(dffe3a_1),
	.dffe3a_0(dffe3a_0),
	.dffe3a_15(dffe3a_15),
	.dffe3a_14(dffe3a_14),
	.dffe3a_13(dffe3a_13),
	.dffe3a_12(dffe3a_12),
	.datab({datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.clock(clock));

endmodule

module fft_mult_0p01_1 (
	dataa,
	clken,
	dffe3a_11,
	dffe3a_10,
	dffe3a_9,
	dffe3a_8,
	dffe3a_7,
	dffe3a_6,
	dffe3a_5,
	dffe3a_4,
	dffe3a_3,
	dffe3a_2,
	dffe3a_1,
	dffe3a_0,
	dffe3a_15,
	dffe3a_14,
	dffe3a_13,
	dffe3a_12,
	datab,
	clock)/* synthesis synthesis_greybox=1 */;
input 	[7:0] dataa;
input 	clken;
output 	dffe3a_11;
output 	dffe3a_10;
output 	dffe3a_9;
output 	dffe3a_8;
output 	dffe3a_7;
output 	dffe3a_6;
output 	dffe3a_5;
output 	dffe3a_4;
output 	dffe3a_3;
output 	dffe3a_2;
output 	dffe3a_1;
output 	dffe3a_0;
output 	dffe3a_15;
output 	dffe3a_14;
output 	dffe3a_13;
output 	dffe3a_12;
input 	[7:0] datab;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1~dataout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT1 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT2 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT3 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT4 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT5 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT6 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT7 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT8 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT9 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT10 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT11 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT12 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT13 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT14 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT15 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT11 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT10 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT9 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT8 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT7 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT6 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT5 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT4 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT3 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT2 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT1 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2~dataout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT15 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT14 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT13 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT12 ;

wire [35:0] \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2_DATAOUT_bus ;
wire [35:0] \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1_DATAOUT_bus ;

assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2~dataout  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2_DATAOUT_bus [0];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT1  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2_DATAOUT_bus [1];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT2  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2_DATAOUT_bus [2];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT3  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2_DATAOUT_bus [3];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT4  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2_DATAOUT_bus [4];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT5  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2_DATAOUT_bus [5];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT6  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2_DATAOUT_bus [6];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT7  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2_DATAOUT_bus [7];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT8  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2_DATAOUT_bus [8];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT9  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2_DATAOUT_bus [9];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT10  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2_DATAOUT_bus [10];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT11  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2_DATAOUT_bus [11];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT12  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2_DATAOUT_bus [12];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT13  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2_DATAOUT_bus [13];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT14  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2_DATAOUT_bus [14];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT15  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2_DATAOUT_bus [15];

assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1~dataout  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1_DATAOUT_bus [0];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT1  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1_DATAOUT_bus [1];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT2  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1_DATAOUT_bus [2];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT3  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1_DATAOUT_bus [3];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT4  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1_DATAOUT_bus [4];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT5  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1_DATAOUT_bus [5];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT6  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1_DATAOUT_bus [6];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT7  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1_DATAOUT_bus [7];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT8  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1_DATAOUT_bus [8];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT9  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1_DATAOUT_bus [9];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT10  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1_DATAOUT_bus [10];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT11  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1_DATAOUT_bus [11];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT12  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1_DATAOUT_bus [12];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT13  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1_DATAOUT_bus [13];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT14  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1_DATAOUT_bus [14];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT15  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1_DATAOUT_bus [15];

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|dffe3a[11] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT11 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_11),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|dffe3a[11] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|dffe3a[11] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|dffe3a[10] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT10 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_10),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|dffe3a[10] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|dffe3a[10] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|dffe3a[9] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT9 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_9),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|dffe3a[9] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|dffe3a[9] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|dffe3a[8] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT8 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_8),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|dffe3a[8] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|dffe3a[8] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|dffe3a[7] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT7 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_7),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|dffe3a[7] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|dffe3a[7] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|dffe3a[6] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT6 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_6),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|dffe3a[6] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|dffe3a[6] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|dffe3a[5] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT5 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_5),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|dffe3a[5] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|dffe3a[5] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|dffe3a[4] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT4 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_4),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|dffe3a[4] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|dffe3a[4] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|dffe3a[3] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT3 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_3),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|dffe3a[3] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|dffe3a[3] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|dffe3a[2] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT2 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_2),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|dffe3a[2] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|dffe3a[2] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|dffe3a[1] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT1 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_1),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|dffe3a[1] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|dffe3a[1] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|dffe3a[0] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2~dataout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_0),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|dffe3a[0] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|dffe3a[0] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|dffe3a[15] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT15 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_15),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|dffe3a[15] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|dffe3a[15] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|dffe3a[14] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT14 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_14),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|dffe3a[14] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|dffe3a[14] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|dffe3a[13] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT13 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_13),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|dffe3a[13] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|dffe3a[13] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|dffe3a[12] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT12 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_12),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|dffe3a[12] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|dffe3a[12] .power_up = "low";

cycloneiii_mac_mult \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1 (
	.signa(vcc),
	.signb(vcc),
	.clk(clock),
	.aclr(gnd),
	.ena(clken),
	.dataa({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.datab({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.dataout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1_DATAOUT_bus ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1 .dataa_clock = "0";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1 .dataa_width = 8;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1 .datab_clock = "0";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1 .datab_width = 8;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1 .signa_clock = "none";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1 .signb_clock = "none";

cycloneiii_mac_out \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2 (
	.clk(clock),
	.aclr(gnd),
	.ena(clken),
	.dataa({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT15 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT14 ,\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT13 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT12 ,\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT11 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT10 ,\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT9 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT8 ,\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT7 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT6 ,\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT5 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT4 ,\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT3 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT2 ,\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT1 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_mult1~dataout }),
	.dataout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2_DATAOUT_bus ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2 .dataa_width = 16;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm1|gen_dsp_only:m_bd|auto_generated|mac_out2 .output_clock = "0";

endmodule

module fft_asj_fft_cmult_can_fft_120_1 (
	pipeline_dffe_11,
	pipeline_dffe_15,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	pipeline_dffe_9,
	pipeline_dffe_8,
	pipeline_dffe_10,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_81,
	pipeline_dffe_91,
	pipeline_dffe_21,
	pipeline_dffe_31,
	pipeline_dffe_41,
	pipeline_dffe_51,
	pipeline_dffe_61,
	pipeline_dffe_71,
	pipeline_dffe_82,
	pipeline_dffe_92,
	global_clock_enable,
	real_out_3,
	real_out_7,
	real_out_4,
	real_out_5,
	real_out_6,
	real_out_1,
	real_out_0,
	real_out_2,
	twiddle_data100,
	twiddle_data101,
	twiddle_data102,
	twiddle_data103,
	twiddle_data104,
	twiddle_data105,
	twiddle_data106,
	twiddle_data107,
	twiddle_data110,
	twiddle_data111,
	twiddle_data112,
	twiddle_data113,
	twiddle_data114,
	twiddle_data115,
	twiddle_data116,
	twiddle_data117,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_11;
output 	pipeline_dffe_15;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
output 	pipeline_dffe_9;
output 	pipeline_dffe_8;
output 	pipeline_dffe_10;
input 	pipeline_dffe_2;
input 	pipeline_dffe_3;
input 	pipeline_dffe_4;
input 	pipeline_dffe_5;
input 	pipeline_dffe_6;
input 	pipeline_dffe_7;
input 	pipeline_dffe_81;
input 	pipeline_dffe_91;
input 	pipeline_dffe_21;
input 	pipeline_dffe_31;
input 	pipeline_dffe_41;
input 	pipeline_dffe_51;
input 	pipeline_dffe_61;
input 	pipeline_dffe_71;
input 	pipeline_dffe_82;
input 	pipeline_dffe_92;
input 	global_clock_enable;
output 	real_out_3;
output 	real_out_7;
output 	real_out_4;
output 	real_out_5;
output 	real_out_6;
output 	real_out_1;
output 	real_out_0;
output 	real_out_2;
input 	twiddle_data100;
input 	twiddle_data101;
input 	twiddle_data102;
input 	twiddle_data103;
input 	twiddle_data104;
input 	twiddle_data105;
input 	twiddle_data106;
input 	twiddle_data107;
input 	twiddle_data110;
input 	twiddle_data111;
input 	twiddle_data112;
input 	twiddle_data113;
input 	twiddle_data114;
input 	twiddle_data115;
input 	twiddle_data116;
input 	twiddle_data117;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \result_imag_1[11]~q ;
wire \result_imag_1[10]~q ;
wire \result_imag_1[9]~q ;
wire \result_imag_1[8]~q ;
wire \result_imag_1[7]~q ;
wire \result_imag_1[6]~q ;
wire \result_imag_1[5]~q ;
wire \result_imag_1[4]~q ;
wire \result_imag_1[3]~q ;
wire \result_imag_1[2]~q ;
wire \result_imag_1[1]~q ;
wire \result_imag_1[0]~q ;
wire \result_imag_1[15]~q ;
wire \result_imag_1[14]~q ;
wire \result_imag_1[13]~q ;
wire \result_imag_1[12]~q ;
wire \gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ;
wire \gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ;
wire \gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ;
wire \gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ;
wire \gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ;
wire \addresult_ac_bd[11]~q ;
wire \addresult_ac_bd[10]~q ;
wire \addresult_ac_bd[9]~q ;
wire \addresult_ac_bd[8]~q ;
wire \addresult_ac_bd[7]~q ;
wire \addresult_ac_bd[6]~q ;
wire \addresult_ac_bd[5]~q ;
wire \addresult_ac_bd[4]~q ;
wire \addresult_ac_bd[3]~q ;
wire \addresult_ac_bd[2]~q ;
wire \addresult_ac_bd[1]~q ;
wire \addresult_ac_bd[0]~q ;
wire \result_imag_1[0]~17 ;
wire \result_imag_1[0]~16_combout ;
wire \result_imag_1[1]~19 ;
wire \result_imag_1[1]~18_combout ;
wire \result_imag_1[2]~21 ;
wire \result_imag_1[2]~20_combout ;
wire \result_imag_1[3]~23 ;
wire \result_imag_1[3]~22_combout ;
wire \result_imag_1[4]~25 ;
wire \result_imag_1[4]~24_combout ;
wire \result_imag_1[5]~27 ;
wire \result_imag_1[5]~26_combout ;
wire \result_imag_1[6]~29 ;
wire \result_imag_1[6]~28_combout ;
wire \result_imag_1[7]~31 ;
wire \result_imag_1[7]~30_combout ;
wire \result_imag_1[8]~33 ;
wire \result_imag_1[8]~32_combout ;
wire \result_imag_1[9]~35 ;
wire \result_imag_1[9]~34_combout ;
wire \result_imag_1[10]~37 ;
wire \result_imag_1[10]~36_combout ;
wire \result_imag_1[11]~39 ;
wire \result_imag_1[11]~38_combout ;
wire \addresult_ac_bd[15]~q ;
wire \addresult_ac_bd[14]~q ;
wire \addresult_ac_bd[13]~q ;
wire \addresult_ac_bd[12]~q ;
wire \result_imag_1[12]~41 ;
wire \result_imag_1[12]~40_combout ;
wire \result_imag_1[13]~43 ;
wire \result_imag_1[13]~42_combout ;
wire \result_imag_1[14]~45 ;
wire \result_imag_1[14]~44_combout ;
wire \result_imag_1[15]~46_combout ;
wire \result_real_1_tmp[11]~q ;
wire \result_real_1_tmp[10]~q ;
wire \result_real_1_tmp[9]~q ;
wire \result_real_1_tmp[8]~q ;
wire \result_real_1_tmp[7]~q ;
wire \result_real_1_tmp[6]~q ;
wire \result_real_1_tmp[5]~q ;
wire \result_real_1_tmp[4]~q ;
wire \result_real_1_tmp[3]~q ;
wire \result_real_1_tmp[2]~q ;
wire \result_real_1_tmp[1]~q ;
wire \result_real_1_tmp[0]~q ;
wire \result_real_1_tmp[15]~q ;
wire \result_real_1_tmp[14]~q ;
wire \result_real_1_tmp[13]~q ;
wire \result_real_1_tmp[12]~q ;
wire \addresult_ac_bd[0]~17 ;
wire \addresult_ac_bd[0]~16_combout ;
wire \addresult_ac_bd[1]~19 ;
wire \addresult_ac_bd[1]~18_combout ;
wire \addresult_ac_bd[2]~21 ;
wire \addresult_ac_bd[2]~20_combout ;
wire \addresult_ac_bd[3]~23 ;
wire \addresult_ac_bd[3]~22_combout ;
wire \addresult_ac_bd[4]~25 ;
wire \addresult_ac_bd[4]~24_combout ;
wire \addresult_ac_bd[5]~27 ;
wire \addresult_ac_bd[5]~26_combout ;
wire \addresult_ac_bd[6]~29 ;
wire \addresult_ac_bd[6]~28_combout ;
wire \addresult_ac_bd[7]~31 ;
wire \addresult_ac_bd[7]~30_combout ;
wire \addresult_ac_bd[8]~33 ;
wire \addresult_ac_bd[8]~32_combout ;
wire \addresult_ac_bd[9]~35 ;
wire \addresult_ac_bd[9]~34_combout ;
wire \addresult_ac_bd[10]~37 ;
wire \addresult_ac_bd[10]~36_combout ;
wire \addresult_ac_bd[11]~39 ;
wire \addresult_ac_bd[11]~38_combout ;
wire \addresult_ac_bd[12]~41 ;
wire \addresult_ac_bd[12]~40_combout ;
wire \addresult_ac_bd[13]~43 ;
wire \addresult_ac_bd[13]~42_combout ;
wire \addresult_ac_bd[14]~45 ;
wire \addresult_ac_bd[14]~44_combout ;
wire \addresult_ac_bd[15]~46_combout ;
wire \result_real_1_tmp[0]~17 ;
wire \result_real_1_tmp[0]~16_combout ;
wire \result_real_1_tmp[1]~19 ;
wire \result_real_1_tmp[1]~18_combout ;
wire \result_real_1_tmp[2]~21 ;
wire \result_real_1_tmp[2]~20_combout ;
wire \result_real_1_tmp[3]~23 ;
wire \result_real_1_tmp[3]~22_combout ;
wire \result_real_1_tmp[4]~25 ;
wire \result_real_1_tmp[4]~24_combout ;
wire \result_real_1_tmp[5]~27 ;
wire \result_real_1_tmp[5]~26_combout ;
wire \result_real_1_tmp[6]~29 ;
wire \result_real_1_tmp[6]~28_combout ;
wire \result_real_1_tmp[7]~31 ;
wire \result_real_1_tmp[7]~30_combout ;
wire \result_real_1_tmp[8]~33 ;
wire \result_real_1_tmp[8]~32_combout ;
wire \result_real_1_tmp[9]~35 ;
wire \result_real_1_tmp[9]~34_combout ;
wire \result_real_1_tmp[10]~37 ;
wire \result_real_1_tmp[10]~36_combout ;
wire \result_real_1_tmp[11]~39 ;
wire \result_real_1_tmp[11]~38_combout ;
wire \result_real_1_tmp[12]~41 ;
wire \result_real_1_tmp[12]~40_combout ;
wire \result_real_1_tmp[13]~43 ;
wire \result_real_1_tmp[13]~42_combout ;
wire \result_real_1_tmp[14]~45 ;
wire \result_real_1_tmp[14]~44_combout ;
wire \result_real_1_tmp[15]~46_combout ;
wire \addresult_a_b[0]~q ;
wire \addresult_a_b[1]~q ;
wire \addresult_a_b[2]~q ;
wire \addresult_a_b[3]~q ;
wire \addresult_a_b[4]~q ;
wire \addresult_a_b[5]~q ;
wire \addresult_a_b[6]~q ;
wire \addresult_a_b[7]~q ;
wire \addresult_a_b[8]~q ;
wire \addresult_c_d[0]~q ;
wire \addresult_c_d[1]~q ;
wire \addresult_c_d[2]~q ;
wire \addresult_c_d[3]~q ;
wire \addresult_c_d[4]~q ;
wire \addresult_c_d[5]~q ;
wire \addresult_c_d[6]~q ;
wire \addresult_c_d[7]~q ;
wire \addresult_c_d[8]~q ;
wire \addresult_a_b[0]~10 ;
wire \addresult_a_b[0]~9_combout ;
wire \addresult_a_b[1]~12 ;
wire \addresult_a_b[1]~11_combout ;
wire \addresult_a_b[2]~14 ;
wire \addresult_a_b[2]~13_combout ;
wire \addresult_a_b[3]~16 ;
wire \addresult_a_b[3]~15_combout ;
wire \addresult_a_b[4]~18 ;
wire \addresult_a_b[4]~17_combout ;
wire \addresult_a_b[5]~20 ;
wire \addresult_a_b[5]~19_combout ;
wire \addresult_a_b[6]~22 ;
wire \addresult_a_b[6]~21_combout ;
wire \addresult_a_b[7]~24 ;
wire \addresult_a_b[7]~23_combout ;
wire \addresult_a_b[8]~25_combout ;
wire \addresult_c_d[0]~10 ;
wire \addresult_c_d[0]~9_combout ;
wire \addresult_c_d[1]~12 ;
wire \addresult_c_d[1]~11_combout ;
wire \addresult_c_d[2]~14 ;
wire \addresult_c_d[2]~13_combout ;
wire \addresult_c_d[3]~16 ;
wire \addresult_c_d[3]~15_combout ;
wire \addresult_c_d[4]~18 ;
wire \addresult_c_d[4]~17_combout ;
wire \addresult_c_d[5]~20 ;
wire \addresult_c_d[5]~19_combout ;
wire \addresult_c_d[6]~22 ;
wire \addresult_c_d[6]~21_combout ;
wire \addresult_c_d[7]~24 ;
wire \addresult_c_d[7]~23_combout ;
wire \addresult_c_d[8]~25_combout ;
wire \gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ;
wire \gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ;
wire \gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ;
wire \result_a_b_c_d_se[11]~q ;
wire \result_a_b_c_d_se[10]~q ;
wire \result_a_b_c_d_se[9]~q ;
wire \result_a_b_c_d_se[8]~q ;
wire \result_a_b_c_d_se[7]~q ;
wire \result_a_b_c_d_se[6]~q ;
wire \result_a_b_c_d_se[5]~q ;
wire \result_a_b_c_d_se[4]~q ;
wire \result_a_b_c_d_se[3]~q ;
wire \result_a_b_c_d_se[2]~q ;
wire \result_a_b_c_d_se[1]~q ;
wire \result_a_b_c_d_se[0]~q ;
wire \result_a_b_c_d_se[15]~q ;
wire \result_a_b_c_d_se[14]~q ;
wire \result_a_b_c_d_se[13]~q ;
wire \result_a_b_c_d_se[12]~q ;
wire \result_a_c_se[11]~q ;
wire \result_b_d_se[11]~q ;
wire \result_a_c_se[10]~q ;
wire \result_b_d_se[10]~q ;
wire \result_a_c_se[9]~q ;
wire \result_b_d_se[9]~q ;
wire \result_a_c_se[8]~q ;
wire \result_b_d_se[8]~q ;
wire \result_a_c_se[7]~q ;
wire \result_b_d_se[7]~q ;
wire \result_a_c_se[6]~q ;
wire \result_b_d_se[6]~q ;
wire \result_a_c_se[5]~q ;
wire \result_b_d_se[5]~q ;
wire \result_a_c_se[4]~q ;
wire \result_b_d_se[4]~q ;
wire \result_a_c_se[3]~q ;
wire \result_b_d_se[3]~q ;
wire \result_a_c_se[2]~q ;
wire \result_b_d_se[2]~q ;
wire \result_a_c_se[1]~q ;
wire \result_b_d_se[1]~q ;
wire \result_a_c_se[0]~q ;
wire \result_b_d_se[0]~q ;
wire \gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[11]~q ;
wire \gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[10]~q ;
wire \gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[9]~q ;
wire \gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[8]~q ;
wire \gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[7]~q ;
wire \gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[6]~q ;
wire \gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[5]~q ;
wire \gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[4]~q ;
wire \gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[3]~q ;
wire \gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[2]~q ;
wire \gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[1]~q ;
wire \gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[0]~q ;
wire \result_a_c_se[15]~q ;
wire \result_b_d_se[15]~q ;
wire \result_a_c_se[14]~q ;
wire \result_b_d_se[14]~q ;
wire \result_a_c_se[13]~q ;
wire \result_b_d_se[13]~q ;
wire \result_a_c_se[12]~q ;
wire \result_b_d_se[12]~q ;
wire \gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[15]~q ;
wire \gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[14]~q ;
wire \gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[13]~q ;
wire \gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[12]~q ;
wire \gen_dsp_only:m_ac|auto_generated|dffe3a[11]~q ;
wire \gen_dsp_only:m_bd|auto_generated|dffe3a[11]~q ;
wire \gen_dsp_only:m_ac|auto_generated|dffe3a[10]~q ;
wire \gen_dsp_only:m_bd|auto_generated|dffe3a[10]~q ;
wire \gen_dsp_only:m_ac|auto_generated|dffe3a[9]~q ;
wire \gen_dsp_only:m_bd|auto_generated|dffe3a[9]~q ;
wire \gen_dsp_only:m_ac|auto_generated|dffe3a[8]~q ;
wire \gen_dsp_only:m_bd|auto_generated|dffe3a[8]~q ;
wire \gen_dsp_only:m_ac|auto_generated|dffe3a[7]~q ;
wire \gen_dsp_only:m_bd|auto_generated|dffe3a[7]~q ;
wire \gen_dsp_only:m_ac|auto_generated|dffe3a[6]~q ;
wire \gen_dsp_only:m_bd|auto_generated|dffe3a[6]~q ;
wire \gen_dsp_only:m_ac|auto_generated|dffe3a[5]~q ;
wire \gen_dsp_only:m_bd|auto_generated|dffe3a[5]~q ;
wire \gen_dsp_only:m_ac|auto_generated|dffe3a[4]~q ;
wire \gen_dsp_only:m_bd|auto_generated|dffe3a[4]~q ;
wire \gen_dsp_only:m_ac|auto_generated|dffe3a[3]~q ;
wire \gen_dsp_only:m_bd|auto_generated|dffe3a[3]~q ;
wire \gen_dsp_only:m_ac|auto_generated|dffe3a[2]~q ;
wire \gen_dsp_only:m_bd|auto_generated|dffe3a[2]~q ;
wire \gen_dsp_only:m_ac|auto_generated|dffe3a[1]~q ;
wire \gen_dsp_only:m_bd|auto_generated|dffe3a[1]~q ;
wire \gen_dsp_only:m_ac|auto_generated|dffe3a[0]~q ;
wire \gen_dsp_only:m_bd|auto_generated|dffe3a[0]~q ;
wire \gen_dsp_only:m_ac|auto_generated|dffe3a[15]~q ;
wire \gen_dsp_only:m_bd|auto_generated|dffe3a[15]~q ;
wire \gen_dsp_only:m_ac|auto_generated|dffe3a[14]~q ;
wire \gen_dsp_only:m_bd|auto_generated|dffe3a[14]~q ;
wire \gen_dsp_only:m_ac|auto_generated|dffe3a[13]~q ;
wire \gen_dsp_only:m_bd|auto_generated|dffe3a[13]~q ;
wire \gen_dsp_only:m_ac|auto_generated|dffe3a[12]~q ;
wire \gen_dsp_only:m_bd|auto_generated|dffe3a[12]~q ;


fft_asj_fft_pround_fft_120_3 \gen_unsc:u1 (
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_14(pipeline_dffe_14),
	.result_imag_1_11(\result_imag_1[11]~q ),
	.result_imag_1_10(\result_imag_1[10]~q ),
	.result_imag_1_9(\result_imag_1[9]~q ),
	.result_imag_1_8(\result_imag_1[8]~q ),
	.result_imag_1_7(\result_imag_1[7]~q ),
	.result_imag_1_6(\result_imag_1[6]~q ),
	.result_imag_1_5(\result_imag_1[5]~q ),
	.result_imag_1_4(\result_imag_1[4]~q ),
	.result_imag_1_3(\result_imag_1[3]~q ),
	.result_imag_1_2(\result_imag_1[2]~q ),
	.result_imag_1_1(\result_imag_1[1]~q ),
	.result_imag_1_0(\result_imag_1[0]~q ),
	.result_imag_1_15(\result_imag_1[15]~q ),
	.result_imag_1_14(\result_imag_1[14]~q ),
	.result_imag_1_13(\result_imag_1[13]~q ),
	.result_imag_1_12(\result_imag_1[12]~q ),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_10(pipeline_dffe_10),
	.global_clock_enable(global_clock_enable),
	.clk(clk));

fft_asj_fft_pround_fft_120_2 \gen_unsc:u0 (
	.pipeline_dffe_11(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_15(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_12(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_13(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ),
	.pipeline_dffe_14(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ),
	.result_real_1_tmp_11(\result_real_1_tmp[11]~q ),
	.result_real_1_tmp_10(\result_real_1_tmp[10]~q ),
	.result_real_1_tmp_9(\result_real_1_tmp[9]~q ),
	.result_real_1_tmp_8(\result_real_1_tmp[8]~q ),
	.result_real_1_tmp_7(\result_real_1_tmp[7]~q ),
	.result_real_1_tmp_6(\result_real_1_tmp[6]~q ),
	.result_real_1_tmp_5(\result_real_1_tmp[5]~q ),
	.result_real_1_tmp_4(\result_real_1_tmp[4]~q ),
	.result_real_1_tmp_3(\result_real_1_tmp[3]~q ),
	.result_real_1_tmp_2(\result_real_1_tmp[2]~q ),
	.result_real_1_tmp_1(\result_real_1_tmp[1]~q ),
	.result_real_1_tmp_0(\result_real_1_tmp[0]~q ),
	.result_real_1_tmp_15(\result_real_1_tmp[15]~q ),
	.result_real_1_tmp_14(\result_real_1_tmp[14]~q ),
	.result_real_1_tmp_13(\result_real_1_tmp[13]~q ),
	.result_real_1_tmp_12(\result_real_1_tmp[12]~q ),
	.pipeline_dffe_9(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_8(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_10(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ),
	.global_clock_enable(global_clock_enable),
	.clk(clk));

fft_LPM_MULT_4 \gen_dsp_only:m_a_b_c_d (
	.dataa({\addresult_a_b[8]~q ,\addresult_a_b[7]~q ,\addresult_a_b[6]~q ,\addresult_a_b[5]~q ,\addresult_a_b[4]~q ,\addresult_a_b[3]~q ,\addresult_a_b[2]~q ,\addresult_a_b[1]~q ,\addresult_a_b[0]~q }),
	.datab({\addresult_c_d[8]~q ,\addresult_c_d[7]~q ,\addresult_c_d[6]~q ,\addresult_c_d[5]~q ,\addresult_c_d[4]~q ,\addresult_c_d[3]~q ,\addresult_c_d[2]~q ,\addresult_c_d[1]~q ,\addresult_c_d[0]~q }),
	.clken(global_clock_enable),
	.dffe3a_11(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[11]~q ),
	.dffe3a_10(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[10]~q ),
	.dffe3a_9(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[9]~q ),
	.dffe3a_8(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[8]~q ),
	.dffe3a_7(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[7]~q ),
	.dffe3a_6(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[6]~q ),
	.dffe3a_5(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[5]~q ),
	.dffe3a_4(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[4]~q ),
	.dffe3a_3(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[3]~q ),
	.dffe3a_2(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[2]~q ),
	.dffe3a_1(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[1]~q ),
	.dffe3a_0(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[0]~q ),
	.dffe3a_15(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[15]~q ),
	.dffe3a_14(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[14]~q ),
	.dffe3a_13(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[13]~q ),
	.dffe3a_12(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[12]~q ),
	.clock(clk));

fft_LPM_MULT_6 \gen_dsp_only:m_bd (
	.dataa({gnd,pipeline_dffe_92,pipeline_dffe_82,pipeline_dffe_71,pipeline_dffe_61,pipeline_dffe_51,pipeline_dffe_41,pipeline_dffe_31,pipeline_dffe_21}),
	.clken(global_clock_enable),
	.dffe3a_11(\gen_dsp_only:m_bd|auto_generated|dffe3a[11]~q ),
	.dffe3a_10(\gen_dsp_only:m_bd|auto_generated|dffe3a[10]~q ),
	.dffe3a_9(\gen_dsp_only:m_bd|auto_generated|dffe3a[9]~q ),
	.dffe3a_8(\gen_dsp_only:m_bd|auto_generated|dffe3a[8]~q ),
	.dffe3a_7(\gen_dsp_only:m_bd|auto_generated|dffe3a[7]~q ),
	.dffe3a_6(\gen_dsp_only:m_bd|auto_generated|dffe3a[6]~q ),
	.dffe3a_5(\gen_dsp_only:m_bd|auto_generated|dffe3a[5]~q ),
	.dffe3a_4(\gen_dsp_only:m_bd|auto_generated|dffe3a[4]~q ),
	.dffe3a_3(\gen_dsp_only:m_bd|auto_generated|dffe3a[3]~q ),
	.dffe3a_2(\gen_dsp_only:m_bd|auto_generated|dffe3a[2]~q ),
	.dffe3a_1(\gen_dsp_only:m_bd|auto_generated|dffe3a[1]~q ),
	.dffe3a_0(\gen_dsp_only:m_bd|auto_generated|dffe3a[0]~q ),
	.dffe3a_15(\gen_dsp_only:m_bd|auto_generated|dffe3a[15]~q ),
	.dffe3a_14(\gen_dsp_only:m_bd|auto_generated|dffe3a[14]~q ),
	.dffe3a_13(\gen_dsp_only:m_bd|auto_generated|dffe3a[13]~q ),
	.dffe3a_12(\gen_dsp_only:m_bd|auto_generated|dffe3a[12]~q ),
	.datab({gnd,twiddle_data117,twiddle_data116,twiddle_data115,twiddle_data114,twiddle_data113,twiddle_data112,twiddle_data111,twiddle_data110}),
	.clock(clk));

fft_LPM_MULT_5 \gen_dsp_only:m_ac (
	.dataa({gnd,pipeline_dffe_91,pipeline_dffe_81,pipeline_dffe_7,pipeline_dffe_6,pipeline_dffe_5,pipeline_dffe_4,pipeline_dffe_3,pipeline_dffe_2}),
	.clken(global_clock_enable),
	.dffe3a_11(\gen_dsp_only:m_ac|auto_generated|dffe3a[11]~q ),
	.dffe3a_10(\gen_dsp_only:m_ac|auto_generated|dffe3a[10]~q ),
	.dffe3a_9(\gen_dsp_only:m_ac|auto_generated|dffe3a[9]~q ),
	.dffe3a_8(\gen_dsp_only:m_ac|auto_generated|dffe3a[8]~q ),
	.dffe3a_7(\gen_dsp_only:m_ac|auto_generated|dffe3a[7]~q ),
	.dffe3a_6(\gen_dsp_only:m_ac|auto_generated|dffe3a[6]~q ),
	.dffe3a_5(\gen_dsp_only:m_ac|auto_generated|dffe3a[5]~q ),
	.dffe3a_4(\gen_dsp_only:m_ac|auto_generated|dffe3a[4]~q ),
	.dffe3a_3(\gen_dsp_only:m_ac|auto_generated|dffe3a[3]~q ),
	.dffe3a_2(\gen_dsp_only:m_ac|auto_generated|dffe3a[2]~q ),
	.dffe3a_1(\gen_dsp_only:m_ac|auto_generated|dffe3a[1]~q ),
	.dffe3a_0(\gen_dsp_only:m_ac|auto_generated|dffe3a[0]~q ),
	.dffe3a_15(\gen_dsp_only:m_ac|auto_generated|dffe3a[15]~q ),
	.dffe3a_14(\gen_dsp_only:m_ac|auto_generated|dffe3a[14]~q ),
	.dffe3a_13(\gen_dsp_only:m_ac|auto_generated|dffe3a[13]~q ),
	.dffe3a_12(\gen_dsp_only:m_ac|auto_generated|dffe3a[12]~q ),
	.datab({gnd,twiddle_data107,twiddle_data106,twiddle_data105,twiddle_data104,twiddle_data103,twiddle_data102,twiddle_data101,twiddle_data100}),
	.clock(clk));

dffeas \result_imag_1[11] (
	.clk(clk),
	.d(\result_imag_1[11]~38_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[11]~q ),
	.prn(vcc));
defparam \result_imag_1[11] .is_wysiwyg = "true";
defparam \result_imag_1[11] .power_up = "low";

dffeas \result_imag_1[10] (
	.clk(clk),
	.d(\result_imag_1[10]~36_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[10]~q ),
	.prn(vcc));
defparam \result_imag_1[10] .is_wysiwyg = "true";
defparam \result_imag_1[10] .power_up = "low";

dffeas \result_imag_1[9] (
	.clk(clk),
	.d(\result_imag_1[9]~34_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[9]~q ),
	.prn(vcc));
defparam \result_imag_1[9] .is_wysiwyg = "true";
defparam \result_imag_1[9] .power_up = "low";

dffeas \result_imag_1[8] (
	.clk(clk),
	.d(\result_imag_1[8]~32_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[8]~q ),
	.prn(vcc));
defparam \result_imag_1[8] .is_wysiwyg = "true";
defparam \result_imag_1[8] .power_up = "low";

dffeas \result_imag_1[7] (
	.clk(clk),
	.d(\result_imag_1[7]~30_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[7]~q ),
	.prn(vcc));
defparam \result_imag_1[7] .is_wysiwyg = "true";
defparam \result_imag_1[7] .power_up = "low";

dffeas \result_imag_1[6] (
	.clk(clk),
	.d(\result_imag_1[6]~28_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[6]~q ),
	.prn(vcc));
defparam \result_imag_1[6] .is_wysiwyg = "true";
defparam \result_imag_1[6] .power_up = "low";

dffeas \result_imag_1[5] (
	.clk(clk),
	.d(\result_imag_1[5]~26_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[5]~q ),
	.prn(vcc));
defparam \result_imag_1[5] .is_wysiwyg = "true";
defparam \result_imag_1[5] .power_up = "low";

dffeas \result_imag_1[4] (
	.clk(clk),
	.d(\result_imag_1[4]~24_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[4]~q ),
	.prn(vcc));
defparam \result_imag_1[4] .is_wysiwyg = "true";
defparam \result_imag_1[4] .power_up = "low";

dffeas \result_imag_1[3] (
	.clk(clk),
	.d(\result_imag_1[3]~22_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[3]~q ),
	.prn(vcc));
defparam \result_imag_1[3] .is_wysiwyg = "true";
defparam \result_imag_1[3] .power_up = "low";

dffeas \result_imag_1[2] (
	.clk(clk),
	.d(\result_imag_1[2]~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[2]~q ),
	.prn(vcc));
defparam \result_imag_1[2] .is_wysiwyg = "true";
defparam \result_imag_1[2] .power_up = "low";

dffeas \result_imag_1[1] (
	.clk(clk),
	.d(\result_imag_1[1]~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[1]~q ),
	.prn(vcc));
defparam \result_imag_1[1] .is_wysiwyg = "true";
defparam \result_imag_1[1] .power_up = "low";

dffeas \result_imag_1[0] (
	.clk(clk),
	.d(\result_imag_1[0]~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[0]~q ),
	.prn(vcc));
defparam \result_imag_1[0] .is_wysiwyg = "true";
defparam \result_imag_1[0] .power_up = "low";

dffeas \result_imag_1[15] (
	.clk(clk),
	.d(\result_imag_1[15]~46_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[15]~q ),
	.prn(vcc));
defparam \result_imag_1[15] .is_wysiwyg = "true";
defparam \result_imag_1[15] .power_up = "low";

dffeas \result_imag_1[14] (
	.clk(clk),
	.d(\result_imag_1[14]~44_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[14]~q ),
	.prn(vcc));
defparam \result_imag_1[14] .is_wysiwyg = "true";
defparam \result_imag_1[14] .power_up = "low";

dffeas \result_imag_1[13] (
	.clk(clk),
	.d(\result_imag_1[13]~42_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[13]~q ),
	.prn(vcc));
defparam \result_imag_1[13] .is_wysiwyg = "true";
defparam \result_imag_1[13] .power_up = "low";

dffeas \result_imag_1[12] (
	.clk(clk),
	.d(\result_imag_1[12]~40_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[12]~q ),
	.prn(vcc));
defparam \result_imag_1[12] .is_wysiwyg = "true";
defparam \result_imag_1[12] .power_up = "low";

dffeas \addresult_ac_bd[11] (
	.clk(clk),
	.d(\addresult_ac_bd[11]~38_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[11]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[11] .is_wysiwyg = "true";
defparam \addresult_ac_bd[11] .power_up = "low";

dffeas \addresult_ac_bd[10] (
	.clk(clk),
	.d(\addresult_ac_bd[10]~36_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[10]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[10] .is_wysiwyg = "true";
defparam \addresult_ac_bd[10] .power_up = "low";

dffeas \addresult_ac_bd[9] (
	.clk(clk),
	.d(\addresult_ac_bd[9]~34_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[9]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[9] .is_wysiwyg = "true";
defparam \addresult_ac_bd[9] .power_up = "low";

dffeas \addresult_ac_bd[8] (
	.clk(clk),
	.d(\addresult_ac_bd[8]~32_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[8]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[8] .is_wysiwyg = "true";
defparam \addresult_ac_bd[8] .power_up = "low";

dffeas \addresult_ac_bd[7] (
	.clk(clk),
	.d(\addresult_ac_bd[7]~30_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[7]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[7] .is_wysiwyg = "true";
defparam \addresult_ac_bd[7] .power_up = "low";

dffeas \addresult_ac_bd[6] (
	.clk(clk),
	.d(\addresult_ac_bd[6]~28_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[6]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[6] .is_wysiwyg = "true";
defparam \addresult_ac_bd[6] .power_up = "low";

dffeas \addresult_ac_bd[5] (
	.clk(clk),
	.d(\addresult_ac_bd[5]~26_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[5]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[5] .is_wysiwyg = "true";
defparam \addresult_ac_bd[5] .power_up = "low";

dffeas \addresult_ac_bd[4] (
	.clk(clk),
	.d(\addresult_ac_bd[4]~24_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[4]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[4] .is_wysiwyg = "true";
defparam \addresult_ac_bd[4] .power_up = "low";

dffeas \addresult_ac_bd[3] (
	.clk(clk),
	.d(\addresult_ac_bd[3]~22_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[3]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[3] .is_wysiwyg = "true";
defparam \addresult_ac_bd[3] .power_up = "low";

dffeas \addresult_ac_bd[2] (
	.clk(clk),
	.d(\addresult_ac_bd[2]~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[2]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[2] .is_wysiwyg = "true";
defparam \addresult_ac_bd[2] .power_up = "low";

dffeas \addresult_ac_bd[1] (
	.clk(clk),
	.d(\addresult_ac_bd[1]~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[1]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[1] .is_wysiwyg = "true";
defparam \addresult_ac_bd[1] .power_up = "low";

dffeas \addresult_ac_bd[0] (
	.clk(clk),
	.d(\addresult_ac_bd[0]~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[0]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[0] .is_wysiwyg = "true";
defparam \addresult_ac_bd[0] .power_up = "low";

cycloneiii_lcell_comb \result_imag_1[0]~16 (
	.dataa(\addresult_ac_bd[0]~q ),
	.datab(\result_a_b_c_d_se[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\result_imag_1[0]~16_combout ),
	.cout(\result_imag_1[0]~17 ));
defparam \result_imag_1[0]~16 .lut_mask = 16'h66DD;
defparam \result_imag_1[0]~16 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \result_imag_1[1]~18 (
	.dataa(\addresult_ac_bd[1]~q ),
	.datab(\result_a_b_c_d_se[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[0]~17 ),
	.combout(\result_imag_1[1]~18_combout ),
	.cout(\result_imag_1[1]~19 ));
defparam \result_imag_1[1]~18 .lut_mask = 16'h96BF;
defparam \result_imag_1[1]~18 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_imag_1[2]~20 (
	.dataa(\addresult_ac_bd[2]~q ),
	.datab(\result_a_b_c_d_se[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[1]~19 ),
	.combout(\result_imag_1[2]~20_combout ),
	.cout(\result_imag_1[2]~21 ));
defparam \result_imag_1[2]~20 .lut_mask = 16'h96DF;
defparam \result_imag_1[2]~20 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_imag_1[3]~22 (
	.dataa(\addresult_ac_bd[3]~q ),
	.datab(\result_a_b_c_d_se[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[2]~21 ),
	.combout(\result_imag_1[3]~22_combout ),
	.cout(\result_imag_1[3]~23 ));
defparam \result_imag_1[3]~22 .lut_mask = 16'h96BF;
defparam \result_imag_1[3]~22 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_imag_1[4]~24 (
	.dataa(\addresult_ac_bd[4]~q ),
	.datab(\result_a_b_c_d_se[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[3]~23 ),
	.combout(\result_imag_1[4]~24_combout ),
	.cout(\result_imag_1[4]~25 ));
defparam \result_imag_1[4]~24 .lut_mask = 16'h96DF;
defparam \result_imag_1[4]~24 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_imag_1[5]~26 (
	.dataa(\addresult_ac_bd[5]~q ),
	.datab(\result_a_b_c_d_se[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[4]~25 ),
	.combout(\result_imag_1[5]~26_combout ),
	.cout(\result_imag_1[5]~27 ));
defparam \result_imag_1[5]~26 .lut_mask = 16'h96BF;
defparam \result_imag_1[5]~26 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_imag_1[6]~28 (
	.dataa(\addresult_ac_bd[6]~q ),
	.datab(\result_a_b_c_d_se[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[5]~27 ),
	.combout(\result_imag_1[6]~28_combout ),
	.cout(\result_imag_1[6]~29 ));
defparam \result_imag_1[6]~28 .lut_mask = 16'h96DF;
defparam \result_imag_1[6]~28 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_imag_1[7]~30 (
	.dataa(\addresult_ac_bd[7]~q ),
	.datab(\result_a_b_c_d_se[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[6]~29 ),
	.combout(\result_imag_1[7]~30_combout ),
	.cout(\result_imag_1[7]~31 ));
defparam \result_imag_1[7]~30 .lut_mask = 16'h96BF;
defparam \result_imag_1[7]~30 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_imag_1[8]~32 (
	.dataa(\addresult_ac_bd[8]~q ),
	.datab(\result_a_b_c_d_se[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[7]~31 ),
	.combout(\result_imag_1[8]~32_combout ),
	.cout(\result_imag_1[8]~33 ));
defparam \result_imag_1[8]~32 .lut_mask = 16'h96DF;
defparam \result_imag_1[8]~32 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_imag_1[9]~34 (
	.dataa(\addresult_ac_bd[9]~q ),
	.datab(\result_a_b_c_d_se[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[8]~33 ),
	.combout(\result_imag_1[9]~34_combout ),
	.cout(\result_imag_1[9]~35 ));
defparam \result_imag_1[9]~34 .lut_mask = 16'h96BF;
defparam \result_imag_1[9]~34 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_imag_1[10]~36 (
	.dataa(\addresult_ac_bd[10]~q ),
	.datab(\result_a_b_c_d_se[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[9]~35 ),
	.combout(\result_imag_1[10]~36_combout ),
	.cout(\result_imag_1[10]~37 ));
defparam \result_imag_1[10]~36 .lut_mask = 16'h96DF;
defparam \result_imag_1[10]~36 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_imag_1[11]~38 (
	.dataa(\addresult_ac_bd[11]~q ),
	.datab(\result_a_b_c_d_se[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[10]~37 ),
	.combout(\result_imag_1[11]~38_combout ),
	.cout(\result_imag_1[11]~39 ));
defparam \result_imag_1[11]~38 .lut_mask = 16'h96BF;
defparam \result_imag_1[11]~38 .sum_lutc_input = "cin";

dffeas \addresult_ac_bd[15] (
	.clk(clk),
	.d(\addresult_ac_bd[15]~46_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[15]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[15] .is_wysiwyg = "true";
defparam \addresult_ac_bd[15] .power_up = "low";

dffeas \addresult_ac_bd[14] (
	.clk(clk),
	.d(\addresult_ac_bd[14]~44_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[14]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[14] .is_wysiwyg = "true";
defparam \addresult_ac_bd[14] .power_up = "low";

dffeas \addresult_ac_bd[13] (
	.clk(clk),
	.d(\addresult_ac_bd[13]~42_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[13]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[13] .is_wysiwyg = "true";
defparam \addresult_ac_bd[13] .power_up = "low";

dffeas \addresult_ac_bd[12] (
	.clk(clk),
	.d(\addresult_ac_bd[12]~40_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[12]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[12] .is_wysiwyg = "true";
defparam \addresult_ac_bd[12] .power_up = "low";

cycloneiii_lcell_comb \result_imag_1[12]~40 (
	.dataa(\addresult_ac_bd[12]~q ),
	.datab(\result_a_b_c_d_se[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[11]~39 ),
	.combout(\result_imag_1[12]~40_combout ),
	.cout(\result_imag_1[12]~41 ));
defparam \result_imag_1[12]~40 .lut_mask = 16'h96DF;
defparam \result_imag_1[12]~40 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_imag_1[13]~42 (
	.dataa(\addresult_ac_bd[13]~q ),
	.datab(\result_a_b_c_d_se[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[12]~41 ),
	.combout(\result_imag_1[13]~42_combout ),
	.cout(\result_imag_1[13]~43 ));
defparam \result_imag_1[13]~42 .lut_mask = 16'h96BF;
defparam \result_imag_1[13]~42 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_imag_1[14]~44 (
	.dataa(\addresult_ac_bd[14]~q ),
	.datab(\result_a_b_c_d_se[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[13]~43 ),
	.combout(\result_imag_1[14]~44_combout ),
	.cout(\result_imag_1[14]~45 ));
defparam \result_imag_1[14]~44 .lut_mask = 16'h96DF;
defparam \result_imag_1[14]~44 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_imag_1[15]~46 (
	.dataa(\addresult_ac_bd[15]~q ),
	.datab(\result_a_b_c_d_se[15]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\result_imag_1[14]~45 ),
	.combout(\result_imag_1[15]~46_combout ),
	.cout());
defparam \result_imag_1[15]~46 .lut_mask = 16'h9696;
defparam \result_imag_1[15]~46 .sum_lutc_input = "cin";

dffeas \result_real_1_tmp[11] (
	.clk(clk),
	.d(\result_real_1_tmp[11]~38_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[11]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[11] .is_wysiwyg = "true";
defparam \result_real_1_tmp[11] .power_up = "low";

dffeas \result_real_1_tmp[10] (
	.clk(clk),
	.d(\result_real_1_tmp[10]~36_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[10]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[10] .is_wysiwyg = "true";
defparam \result_real_1_tmp[10] .power_up = "low";

dffeas \result_real_1_tmp[9] (
	.clk(clk),
	.d(\result_real_1_tmp[9]~34_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[9]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[9] .is_wysiwyg = "true";
defparam \result_real_1_tmp[9] .power_up = "low";

dffeas \result_real_1_tmp[8] (
	.clk(clk),
	.d(\result_real_1_tmp[8]~32_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[8]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[8] .is_wysiwyg = "true";
defparam \result_real_1_tmp[8] .power_up = "low";

dffeas \result_real_1_tmp[7] (
	.clk(clk),
	.d(\result_real_1_tmp[7]~30_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[7]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[7] .is_wysiwyg = "true";
defparam \result_real_1_tmp[7] .power_up = "low";

dffeas \result_real_1_tmp[6] (
	.clk(clk),
	.d(\result_real_1_tmp[6]~28_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[6]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[6] .is_wysiwyg = "true";
defparam \result_real_1_tmp[6] .power_up = "low";

dffeas \result_real_1_tmp[5] (
	.clk(clk),
	.d(\result_real_1_tmp[5]~26_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[5]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[5] .is_wysiwyg = "true";
defparam \result_real_1_tmp[5] .power_up = "low";

dffeas \result_real_1_tmp[4] (
	.clk(clk),
	.d(\result_real_1_tmp[4]~24_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[4]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[4] .is_wysiwyg = "true";
defparam \result_real_1_tmp[4] .power_up = "low";

dffeas \result_real_1_tmp[3] (
	.clk(clk),
	.d(\result_real_1_tmp[3]~22_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[3]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[3] .is_wysiwyg = "true";
defparam \result_real_1_tmp[3] .power_up = "low";

dffeas \result_real_1_tmp[2] (
	.clk(clk),
	.d(\result_real_1_tmp[2]~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[2]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[2] .is_wysiwyg = "true";
defparam \result_real_1_tmp[2] .power_up = "low";

dffeas \result_real_1_tmp[1] (
	.clk(clk),
	.d(\result_real_1_tmp[1]~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[1]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[1] .is_wysiwyg = "true";
defparam \result_real_1_tmp[1] .power_up = "low";

dffeas \result_real_1_tmp[0] (
	.clk(clk),
	.d(\result_real_1_tmp[0]~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[0]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[0] .is_wysiwyg = "true";
defparam \result_real_1_tmp[0] .power_up = "low";

dffeas \result_real_1_tmp[15] (
	.clk(clk),
	.d(\result_real_1_tmp[15]~46_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[15]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[15] .is_wysiwyg = "true";
defparam \result_real_1_tmp[15] .power_up = "low";

dffeas \result_real_1_tmp[14] (
	.clk(clk),
	.d(\result_real_1_tmp[14]~44_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[14]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[14] .is_wysiwyg = "true";
defparam \result_real_1_tmp[14] .power_up = "low";

dffeas \result_real_1_tmp[13] (
	.clk(clk),
	.d(\result_real_1_tmp[13]~42_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[13]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[13] .is_wysiwyg = "true";
defparam \result_real_1_tmp[13] .power_up = "low";

dffeas \result_real_1_tmp[12] (
	.clk(clk),
	.d(\result_real_1_tmp[12]~40_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[12]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[12] .is_wysiwyg = "true";
defparam \result_real_1_tmp[12] .power_up = "low";

cycloneiii_lcell_comb \addresult_ac_bd[0]~16 (
	.dataa(\result_a_c_se[0]~q ),
	.datab(\result_b_d_se[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\addresult_ac_bd[0]~16_combout ),
	.cout(\addresult_ac_bd[0]~17 ));
defparam \addresult_ac_bd[0]~16 .lut_mask = 16'h66EE;
defparam \addresult_ac_bd[0]~16 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \addresult_ac_bd[1]~18 (
	.dataa(\result_a_c_se[1]~q ),
	.datab(\result_b_d_se[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[0]~17 ),
	.combout(\addresult_ac_bd[1]~18_combout ),
	.cout(\addresult_ac_bd[1]~19 ));
defparam \addresult_ac_bd[1]~18 .lut_mask = 16'h967F;
defparam \addresult_ac_bd[1]~18 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_ac_bd[2]~20 (
	.dataa(\result_a_c_se[2]~q ),
	.datab(\result_b_d_se[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[1]~19 ),
	.combout(\addresult_ac_bd[2]~20_combout ),
	.cout(\addresult_ac_bd[2]~21 ));
defparam \addresult_ac_bd[2]~20 .lut_mask = 16'h96EF;
defparam \addresult_ac_bd[2]~20 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_ac_bd[3]~22 (
	.dataa(\result_a_c_se[3]~q ),
	.datab(\result_b_d_se[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[2]~21 ),
	.combout(\addresult_ac_bd[3]~22_combout ),
	.cout(\addresult_ac_bd[3]~23 ));
defparam \addresult_ac_bd[3]~22 .lut_mask = 16'h967F;
defparam \addresult_ac_bd[3]~22 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_ac_bd[4]~24 (
	.dataa(\result_a_c_se[4]~q ),
	.datab(\result_b_d_se[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[3]~23 ),
	.combout(\addresult_ac_bd[4]~24_combout ),
	.cout(\addresult_ac_bd[4]~25 ));
defparam \addresult_ac_bd[4]~24 .lut_mask = 16'h96EF;
defparam \addresult_ac_bd[4]~24 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_ac_bd[5]~26 (
	.dataa(\result_a_c_se[5]~q ),
	.datab(\result_b_d_se[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[4]~25 ),
	.combout(\addresult_ac_bd[5]~26_combout ),
	.cout(\addresult_ac_bd[5]~27 ));
defparam \addresult_ac_bd[5]~26 .lut_mask = 16'h967F;
defparam \addresult_ac_bd[5]~26 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_ac_bd[6]~28 (
	.dataa(\result_a_c_se[6]~q ),
	.datab(\result_b_d_se[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[5]~27 ),
	.combout(\addresult_ac_bd[6]~28_combout ),
	.cout(\addresult_ac_bd[6]~29 ));
defparam \addresult_ac_bd[6]~28 .lut_mask = 16'h96EF;
defparam \addresult_ac_bd[6]~28 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_ac_bd[7]~30 (
	.dataa(\result_a_c_se[7]~q ),
	.datab(\result_b_d_se[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[6]~29 ),
	.combout(\addresult_ac_bd[7]~30_combout ),
	.cout(\addresult_ac_bd[7]~31 ));
defparam \addresult_ac_bd[7]~30 .lut_mask = 16'h967F;
defparam \addresult_ac_bd[7]~30 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_ac_bd[8]~32 (
	.dataa(\result_a_c_se[8]~q ),
	.datab(\result_b_d_se[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[7]~31 ),
	.combout(\addresult_ac_bd[8]~32_combout ),
	.cout(\addresult_ac_bd[8]~33 ));
defparam \addresult_ac_bd[8]~32 .lut_mask = 16'h96EF;
defparam \addresult_ac_bd[8]~32 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_ac_bd[9]~34 (
	.dataa(\result_a_c_se[9]~q ),
	.datab(\result_b_d_se[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[8]~33 ),
	.combout(\addresult_ac_bd[9]~34_combout ),
	.cout(\addresult_ac_bd[9]~35 ));
defparam \addresult_ac_bd[9]~34 .lut_mask = 16'h967F;
defparam \addresult_ac_bd[9]~34 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_ac_bd[10]~36 (
	.dataa(\result_a_c_se[10]~q ),
	.datab(\result_b_d_se[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[9]~35 ),
	.combout(\addresult_ac_bd[10]~36_combout ),
	.cout(\addresult_ac_bd[10]~37 ));
defparam \addresult_ac_bd[10]~36 .lut_mask = 16'h96EF;
defparam \addresult_ac_bd[10]~36 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_ac_bd[11]~38 (
	.dataa(\result_a_c_se[11]~q ),
	.datab(\result_b_d_se[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[10]~37 ),
	.combout(\addresult_ac_bd[11]~38_combout ),
	.cout(\addresult_ac_bd[11]~39 ));
defparam \addresult_ac_bd[11]~38 .lut_mask = 16'h967F;
defparam \addresult_ac_bd[11]~38 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_ac_bd[12]~40 (
	.dataa(\result_a_c_se[12]~q ),
	.datab(\result_b_d_se[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[11]~39 ),
	.combout(\addresult_ac_bd[12]~40_combout ),
	.cout(\addresult_ac_bd[12]~41 ));
defparam \addresult_ac_bd[12]~40 .lut_mask = 16'h96EF;
defparam \addresult_ac_bd[12]~40 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_ac_bd[13]~42 (
	.dataa(\result_a_c_se[13]~q ),
	.datab(\result_b_d_se[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[12]~41 ),
	.combout(\addresult_ac_bd[13]~42_combout ),
	.cout(\addresult_ac_bd[13]~43 ));
defparam \addresult_ac_bd[13]~42 .lut_mask = 16'h967F;
defparam \addresult_ac_bd[13]~42 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_ac_bd[14]~44 (
	.dataa(\result_a_c_se[14]~q ),
	.datab(\result_b_d_se[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[13]~43 ),
	.combout(\addresult_ac_bd[14]~44_combout ),
	.cout(\addresult_ac_bd[14]~45 ));
defparam \addresult_ac_bd[14]~44 .lut_mask = 16'h96EF;
defparam \addresult_ac_bd[14]~44 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_ac_bd[15]~46 (
	.dataa(\result_a_c_se[15]~q ),
	.datab(\result_b_d_se[15]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\addresult_ac_bd[14]~45 ),
	.combout(\addresult_ac_bd[15]~46_combout ),
	.cout());
defparam \addresult_ac_bd[15]~46 .lut_mask = 16'h9696;
defparam \addresult_ac_bd[15]~46 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_real_1_tmp[0]~16 (
	.dataa(\result_a_c_se[0]~q ),
	.datab(\result_b_d_se[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\result_real_1_tmp[0]~16_combout ),
	.cout(\result_real_1_tmp[0]~17 ));
defparam \result_real_1_tmp[0]~16 .lut_mask = 16'h66BB;
defparam \result_real_1_tmp[0]~16 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \result_real_1_tmp[1]~18 (
	.dataa(\result_a_c_se[1]~q ),
	.datab(\result_b_d_se[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[0]~17 ),
	.combout(\result_real_1_tmp[1]~18_combout ),
	.cout(\result_real_1_tmp[1]~19 ));
defparam \result_real_1_tmp[1]~18 .lut_mask = 16'h96DF;
defparam \result_real_1_tmp[1]~18 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_real_1_tmp[2]~20 (
	.dataa(\result_a_c_se[2]~q ),
	.datab(\result_b_d_se[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[1]~19 ),
	.combout(\result_real_1_tmp[2]~20_combout ),
	.cout(\result_real_1_tmp[2]~21 ));
defparam \result_real_1_tmp[2]~20 .lut_mask = 16'h96BF;
defparam \result_real_1_tmp[2]~20 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_real_1_tmp[3]~22 (
	.dataa(\result_a_c_se[3]~q ),
	.datab(\result_b_d_se[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[2]~21 ),
	.combout(\result_real_1_tmp[3]~22_combout ),
	.cout(\result_real_1_tmp[3]~23 ));
defparam \result_real_1_tmp[3]~22 .lut_mask = 16'h96DF;
defparam \result_real_1_tmp[3]~22 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_real_1_tmp[4]~24 (
	.dataa(\result_a_c_se[4]~q ),
	.datab(\result_b_d_se[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[3]~23 ),
	.combout(\result_real_1_tmp[4]~24_combout ),
	.cout(\result_real_1_tmp[4]~25 ));
defparam \result_real_1_tmp[4]~24 .lut_mask = 16'h96BF;
defparam \result_real_1_tmp[4]~24 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_real_1_tmp[5]~26 (
	.dataa(\result_a_c_se[5]~q ),
	.datab(\result_b_d_se[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[4]~25 ),
	.combout(\result_real_1_tmp[5]~26_combout ),
	.cout(\result_real_1_tmp[5]~27 ));
defparam \result_real_1_tmp[5]~26 .lut_mask = 16'h96DF;
defparam \result_real_1_tmp[5]~26 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_real_1_tmp[6]~28 (
	.dataa(\result_a_c_se[6]~q ),
	.datab(\result_b_d_se[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[5]~27 ),
	.combout(\result_real_1_tmp[6]~28_combout ),
	.cout(\result_real_1_tmp[6]~29 ));
defparam \result_real_1_tmp[6]~28 .lut_mask = 16'h96BF;
defparam \result_real_1_tmp[6]~28 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_real_1_tmp[7]~30 (
	.dataa(\result_a_c_se[7]~q ),
	.datab(\result_b_d_se[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[6]~29 ),
	.combout(\result_real_1_tmp[7]~30_combout ),
	.cout(\result_real_1_tmp[7]~31 ));
defparam \result_real_1_tmp[7]~30 .lut_mask = 16'h96DF;
defparam \result_real_1_tmp[7]~30 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_real_1_tmp[8]~32 (
	.dataa(\result_a_c_se[8]~q ),
	.datab(\result_b_d_se[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[7]~31 ),
	.combout(\result_real_1_tmp[8]~32_combout ),
	.cout(\result_real_1_tmp[8]~33 ));
defparam \result_real_1_tmp[8]~32 .lut_mask = 16'h96BF;
defparam \result_real_1_tmp[8]~32 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_real_1_tmp[9]~34 (
	.dataa(\result_a_c_se[9]~q ),
	.datab(\result_b_d_se[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[8]~33 ),
	.combout(\result_real_1_tmp[9]~34_combout ),
	.cout(\result_real_1_tmp[9]~35 ));
defparam \result_real_1_tmp[9]~34 .lut_mask = 16'h96DF;
defparam \result_real_1_tmp[9]~34 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_real_1_tmp[10]~36 (
	.dataa(\result_a_c_se[10]~q ),
	.datab(\result_b_d_se[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[9]~35 ),
	.combout(\result_real_1_tmp[10]~36_combout ),
	.cout(\result_real_1_tmp[10]~37 ));
defparam \result_real_1_tmp[10]~36 .lut_mask = 16'h96BF;
defparam \result_real_1_tmp[10]~36 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_real_1_tmp[11]~38 (
	.dataa(\result_a_c_se[11]~q ),
	.datab(\result_b_d_se[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[10]~37 ),
	.combout(\result_real_1_tmp[11]~38_combout ),
	.cout(\result_real_1_tmp[11]~39 ));
defparam \result_real_1_tmp[11]~38 .lut_mask = 16'h96DF;
defparam \result_real_1_tmp[11]~38 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_real_1_tmp[12]~40 (
	.dataa(\result_a_c_se[12]~q ),
	.datab(\result_b_d_se[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[11]~39 ),
	.combout(\result_real_1_tmp[12]~40_combout ),
	.cout(\result_real_1_tmp[12]~41 ));
defparam \result_real_1_tmp[12]~40 .lut_mask = 16'h96BF;
defparam \result_real_1_tmp[12]~40 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_real_1_tmp[13]~42 (
	.dataa(\result_a_c_se[13]~q ),
	.datab(\result_b_d_se[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[12]~41 ),
	.combout(\result_real_1_tmp[13]~42_combout ),
	.cout(\result_real_1_tmp[13]~43 ));
defparam \result_real_1_tmp[13]~42 .lut_mask = 16'h96DF;
defparam \result_real_1_tmp[13]~42 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_real_1_tmp[14]~44 (
	.dataa(\result_a_c_se[14]~q ),
	.datab(\result_b_d_se[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[13]~43 ),
	.combout(\result_real_1_tmp[14]~44_combout ),
	.cout(\result_real_1_tmp[14]~45 ));
defparam \result_real_1_tmp[14]~44 .lut_mask = 16'h96BF;
defparam \result_real_1_tmp[14]~44 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_real_1_tmp[15]~46 (
	.dataa(\result_a_c_se[15]~q ),
	.datab(\result_b_d_se[15]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\result_real_1_tmp[14]~45 ),
	.combout(\result_real_1_tmp[15]~46_combout ),
	.cout());
defparam \result_real_1_tmp[15]~46 .lut_mask = 16'h9696;
defparam \result_real_1_tmp[15]~46 .sum_lutc_input = "cin";

dffeas \addresult_a_b[0] (
	.clk(clk),
	.d(\addresult_a_b[0]~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_a_b[0]~q ),
	.prn(vcc));
defparam \addresult_a_b[0] .is_wysiwyg = "true";
defparam \addresult_a_b[0] .power_up = "low";

dffeas \addresult_a_b[1] (
	.clk(clk),
	.d(\addresult_a_b[1]~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_a_b[1]~q ),
	.prn(vcc));
defparam \addresult_a_b[1] .is_wysiwyg = "true";
defparam \addresult_a_b[1] .power_up = "low";

dffeas \addresult_a_b[2] (
	.clk(clk),
	.d(\addresult_a_b[2]~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_a_b[2]~q ),
	.prn(vcc));
defparam \addresult_a_b[2] .is_wysiwyg = "true";
defparam \addresult_a_b[2] .power_up = "low";

dffeas \addresult_a_b[3] (
	.clk(clk),
	.d(\addresult_a_b[3]~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_a_b[3]~q ),
	.prn(vcc));
defparam \addresult_a_b[3] .is_wysiwyg = "true";
defparam \addresult_a_b[3] .power_up = "low";

dffeas \addresult_a_b[4] (
	.clk(clk),
	.d(\addresult_a_b[4]~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_a_b[4]~q ),
	.prn(vcc));
defparam \addresult_a_b[4] .is_wysiwyg = "true";
defparam \addresult_a_b[4] .power_up = "low";

dffeas \addresult_a_b[5] (
	.clk(clk),
	.d(\addresult_a_b[5]~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_a_b[5]~q ),
	.prn(vcc));
defparam \addresult_a_b[5] .is_wysiwyg = "true";
defparam \addresult_a_b[5] .power_up = "low";

dffeas \addresult_a_b[6] (
	.clk(clk),
	.d(\addresult_a_b[6]~21_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_a_b[6]~q ),
	.prn(vcc));
defparam \addresult_a_b[6] .is_wysiwyg = "true";
defparam \addresult_a_b[6] .power_up = "low";

dffeas \addresult_a_b[7] (
	.clk(clk),
	.d(\addresult_a_b[7]~23_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_a_b[7]~q ),
	.prn(vcc));
defparam \addresult_a_b[7] .is_wysiwyg = "true";
defparam \addresult_a_b[7] .power_up = "low";

dffeas \addresult_a_b[8] (
	.clk(clk),
	.d(\addresult_a_b[8]~25_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_a_b[8]~q ),
	.prn(vcc));
defparam \addresult_a_b[8] .is_wysiwyg = "true";
defparam \addresult_a_b[8] .power_up = "low";

dffeas \addresult_c_d[0] (
	.clk(clk),
	.d(\addresult_c_d[0]~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_c_d[0]~q ),
	.prn(vcc));
defparam \addresult_c_d[0] .is_wysiwyg = "true";
defparam \addresult_c_d[0] .power_up = "low";

dffeas \addresult_c_d[1] (
	.clk(clk),
	.d(\addresult_c_d[1]~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_c_d[1]~q ),
	.prn(vcc));
defparam \addresult_c_d[1] .is_wysiwyg = "true";
defparam \addresult_c_d[1] .power_up = "low";

dffeas \addresult_c_d[2] (
	.clk(clk),
	.d(\addresult_c_d[2]~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_c_d[2]~q ),
	.prn(vcc));
defparam \addresult_c_d[2] .is_wysiwyg = "true";
defparam \addresult_c_d[2] .power_up = "low";

dffeas \addresult_c_d[3] (
	.clk(clk),
	.d(\addresult_c_d[3]~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_c_d[3]~q ),
	.prn(vcc));
defparam \addresult_c_d[3] .is_wysiwyg = "true";
defparam \addresult_c_d[3] .power_up = "low";

dffeas \addresult_c_d[4] (
	.clk(clk),
	.d(\addresult_c_d[4]~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_c_d[4]~q ),
	.prn(vcc));
defparam \addresult_c_d[4] .is_wysiwyg = "true";
defparam \addresult_c_d[4] .power_up = "low";

dffeas \addresult_c_d[5] (
	.clk(clk),
	.d(\addresult_c_d[5]~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_c_d[5]~q ),
	.prn(vcc));
defparam \addresult_c_d[5] .is_wysiwyg = "true";
defparam \addresult_c_d[5] .power_up = "low";

dffeas \addresult_c_d[6] (
	.clk(clk),
	.d(\addresult_c_d[6]~21_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_c_d[6]~q ),
	.prn(vcc));
defparam \addresult_c_d[6] .is_wysiwyg = "true";
defparam \addresult_c_d[6] .power_up = "low";

dffeas \addresult_c_d[7] (
	.clk(clk),
	.d(\addresult_c_d[7]~23_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_c_d[7]~q ),
	.prn(vcc));
defparam \addresult_c_d[7] .is_wysiwyg = "true";
defparam \addresult_c_d[7] .power_up = "low";

dffeas \addresult_c_d[8] (
	.clk(clk),
	.d(\addresult_c_d[8]~25_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_c_d[8]~q ),
	.prn(vcc));
defparam \addresult_c_d[8] .is_wysiwyg = "true";
defparam \addresult_c_d[8] .power_up = "low";

cycloneiii_lcell_comb \addresult_a_b[0]~9 (
	.dataa(pipeline_dffe_2),
	.datab(pipeline_dffe_21),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\addresult_a_b[0]~9_combout ),
	.cout(\addresult_a_b[0]~10 ));
defparam \addresult_a_b[0]~9 .lut_mask = 16'h66EE;
defparam \addresult_a_b[0]~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \addresult_a_b[1]~11 (
	.dataa(pipeline_dffe_3),
	.datab(pipeline_dffe_31),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_a_b[0]~10 ),
	.combout(\addresult_a_b[1]~11_combout ),
	.cout(\addresult_a_b[1]~12 ));
defparam \addresult_a_b[1]~11 .lut_mask = 16'h967F;
defparam \addresult_a_b[1]~11 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_a_b[2]~13 (
	.dataa(pipeline_dffe_4),
	.datab(pipeline_dffe_41),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_a_b[1]~12 ),
	.combout(\addresult_a_b[2]~13_combout ),
	.cout(\addresult_a_b[2]~14 ));
defparam \addresult_a_b[2]~13 .lut_mask = 16'h96EF;
defparam \addresult_a_b[2]~13 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_a_b[3]~15 (
	.dataa(pipeline_dffe_5),
	.datab(pipeline_dffe_51),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_a_b[2]~14 ),
	.combout(\addresult_a_b[3]~15_combout ),
	.cout(\addresult_a_b[3]~16 ));
defparam \addresult_a_b[3]~15 .lut_mask = 16'h967F;
defparam \addresult_a_b[3]~15 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_a_b[4]~17 (
	.dataa(pipeline_dffe_6),
	.datab(pipeline_dffe_61),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_a_b[3]~16 ),
	.combout(\addresult_a_b[4]~17_combout ),
	.cout(\addresult_a_b[4]~18 ));
defparam \addresult_a_b[4]~17 .lut_mask = 16'h96EF;
defparam \addresult_a_b[4]~17 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_a_b[5]~19 (
	.dataa(pipeline_dffe_7),
	.datab(pipeline_dffe_71),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_a_b[4]~18 ),
	.combout(\addresult_a_b[5]~19_combout ),
	.cout(\addresult_a_b[5]~20 ));
defparam \addresult_a_b[5]~19 .lut_mask = 16'h967F;
defparam \addresult_a_b[5]~19 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_a_b[6]~21 (
	.dataa(pipeline_dffe_81),
	.datab(pipeline_dffe_82),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_a_b[5]~20 ),
	.combout(\addresult_a_b[6]~21_combout ),
	.cout(\addresult_a_b[6]~22 ));
defparam \addresult_a_b[6]~21 .lut_mask = 16'h96EF;
defparam \addresult_a_b[6]~21 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_a_b[7]~23 (
	.dataa(pipeline_dffe_91),
	.datab(pipeline_dffe_92),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_a_b[6]~22 ),
	.combout(\addresult_a_b[7]~23_combout ),
	.cout(\addresult_a_b[7]~24 ));
defparam \addresult_a_b[7]~23 .lut_mask = 16'h967F;
defparam \addresult_a_b[7]~23 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_a_b[8]~25 (
	.dataa(pipeline_dffe_91),
	.datab(pipeline_dffe_92),
	.datac(gnd),
	.datad(gnd),
	.cin(\addresult_a_b[7]~24 ),
	.combout(\addresult_a_b[8]~25_combout ),
	.cout());
defparam \addresult_a_b[8]~25 .lut_mask = 16'h9696;
defparam \addresult_a_b[8]~25 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_c_d[0]~9 (
	.dataa(twiddle_data100),
	.datab(twiddle_data110),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\addresult_c_d[0]~9_combout ),
	.cout(\addresult_c_d[0]~10 ));
defparam \addresult_c_d[0]~9 .lut_mask = 16'h66EE;
defparam \addresult_c_d[0]~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \addresult_c_d[1]~11 (
	.dataa(twiddle_data101),
	.datab(twiddle_data111),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_c_d[0]~10 ),
	.combout(\addresult_c_d[1]~11_combout ),
	.cout(\addresult_c_d[1]~12 ));
defparam \addresult_c_d[1]~11 .lut_mask = 16'h967F;
defparam \addresult_c_d[1]~11 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_c_d[2]~13 (
	.dataa(twiddle_data102),
	.datab(twiddle_data112),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_c_d[1]~12 ),
	.combout(\addresult_c_d[2]~13_combout ),
	.cout(\addresult_c_d[2]~14 ));
defparam \addresult_c_d[2]~13 .lut_mask = 16'h96EF;
defparam \addresult_c_d[2]~13 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_c_d[3]~15 (
	.dataa(twiddle_data103),
	.datab(twiddle_data113),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_c_d[2]~14 ),
	.combout(\addresult_c_d[3]~15_combout ),
	.cout(\addresult_c_d[3]~16 ));
defparam \addresult_c_d[3]~15 .lut_mask = 16'h967F;
defparam \addresult_c_d[3]~15 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_c_d[4]~17 (
	.dataa(twiddle_data104),
	.datab(twiddle_data114),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_c_d[3]~16 ),
	.combout(\addresult_c_d[4]~17_combout ),
	.cout(\addresult_c_d[4]~18 ));
defparam \addresult_c_d[4]~17 .lut_mask = 16'h96EF;
defparam \addresult_c_d[4]~17 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_c_d[5]~19 (
	.dataa(twiddle_data105),
	.datab(twiddle_data115),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_c_d[4]~18 ),
	.combout(\addresult_c_d[5]~19_combout ),
	.cout(\addresult_c_d[5]~20 ));
defparam \addresult_c_d[5]~19 .lut_mask = 16'h967F;
defparam \addresult_c_d[5]~19 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_c_d[6]~21 (
	.dataa(twiddle_data106),
	.datab(twiddle_data116),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_c_d[5]~20 ),
	.combout(\addresult_c_d[6]~21_combout ),
	.cout(\addresult_c_d[6]~22 ));
defparam \addresult_c_d[6]~21 .lut_mask = 16'h96EF;
defparam \addresult_c_d[6]~21 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_c_d[7]~23 (
	.dataa(twiddle_data107),
	.datab(twiddle_data117),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_c_d[6]~22 ),
	.combout(\addresult_c_d[7]~23_combout ),
	.cout(\addresult_c_d[7]~24 ));
defparam \addresult_c_d[7]~23 .lut_mask = 16'h967F;
defparam \addresult_c_d[7]~23 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_c_d[8]~25 (
	.dataa(twiddle_data107),
	.datab(twiddle_data117),
	.datac(gnd),
	.datad(gnd),
	.cin(\addresult_c_d[7]~24 ),
	.combout(\addresult_c_d[8]~25_combout ),
	.cout());
defparam \addresult_c_d[8]~25 .lut_mask = 16'h9696;
defparam \addresult_c_d[8]~25 .sum_lutc_input = "cin";

dffeas \result_a_b_c_d_se[11] (
	.clk(clk),
	.d(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[11]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[11] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[11] .power_up = "low";

dffeas \result_a_b_c_d_se[10] (
	.clk(clk),
	.d(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[10]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[10] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[10] .power_up = "low";

dffeas \result_a_b_c_d_se[9] (
	.clk(clk),
	.d(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[9]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[9] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[9] .power_up = "low";

dffeas \result_a_b_c_d_se[8] (
	.clk(clk),
	.d(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[8]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[8] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[8] .power_up = "low";

dffeas \result_a_b_c_d_se[7] (
	.clk(clk),
	.d(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[7]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[7] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[7] .power_up = "low";

dffeas \result_a_b_c_d_se[6] (
	.clk(clk),
	.d(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[6]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[6] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[6] .power_up = "low";

dffeas \result_a_b_c_d_se[5] (
	.clk(clk),
	.d(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[5]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[5] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[5] .power_up = "low";

dffeas \result_a_b_c_d_se[4] (
	.clk(clk),
	.d(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[4]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[4] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[4] .power_up = "low";

dffeas \result_a_b_c_d_se[3] (
	.clk(clk),
	.d(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[3]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[3] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[3] .power_up = "low";

dffeas \result_a_b_c_d_se[2] (
	.clk(clk),
	.d(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[2]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[2] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[2] .power_up = "low";

dffeas \result_a_b_c_d_se[1] (
	.clk(clk),
	.d(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[1]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[1] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[1] .power_up = "low";

dffeas \result_a_b_c_d_se[0] (
	.clk(clk),
	.d(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[0]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[0] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[0] .power_up = "low";

dffeas \result_a_b_c_d_se[15] (
	.clk(clk),
	.d(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[15]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[15] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[15] .power_up = "low";

dffeas \result_a_b_c_d_se[14] (
	.clk(clk),
	.d(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[14]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[14] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[14] .power_up = "low";

dffeas \result_a_b_c_d_se[13] (
	.clk(clk),
	.d(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[13]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[13] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[13] .power_up = "low";

dffeas \result_a_b_c_d_se[12] (
	.clk(clk),
	.d(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[12]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[12] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[12] .power_up = "low";

dffeas \result_a_c_se[11] (
	.clk(clk),
	.d(\gen_dsp_only:m_ac|auto_generated|dffe3a[11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[11]~q ),
	.prn(vcc));
defparam \result_a_c_se[11] .is_wysiwyg = "true";
defparam \result_a_c_se[11] .power_up = "low";

dffeas \result_b_d_se[11] (
	.clk(clk),
	.d(\gen_dsp_only:m_bd|auto_generated|dffe3a[11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[11]~q ),
	.prn(vcc));
defparam \result_b_d_se[11] .is_wysiwyg = "true";
defparam \result_b_d_se[11] .power_up = "low";

dffeas \result_a_c_se[10] (
	.clk(clk),
	.d(\gen_dsp_only:m_ac|auto_generated|dffe3a[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[10]~q ),
	.prn(vcc));
defparam \result_a_c_se[10] .is_wysiwyg = "true";
defparam \result_a_c_se[10] .power_up = "low";

dffeas \result_b_d_se[10] (
	.clk(clk),
	.d(\gen_dsp_only:m_bd|auto_generated|dffe3a[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[10]~q ),
	.prn(vcc));
defparam \result_b_d_se[10] .is_wysiwyg = "true";
defparam \result_b_d_se[10] .power_up = "low";

dffeas \result_a_c_se[9] (
	.clk(clk),
	.d(\gen_dsp_only:m_ac|auto_generated|dffe3a[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[9]~q ),
	.prn(vcc));
defparam \result_a_c_se[9] .is_wysiwyg = "true";
defparam \result_a_c_se[9] .power_up = "low";

dffeas \result_b_d_se[9] (
	.clk(clk),
	.d(\gen_dsp_only:m_bd|auto_generated|dffe3a[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[9]~q ),
	.prn(vcc));
defparam \result_b_d_se[9] .is_wysiwyg = "true";
defparam \result_b_d_se[9] .power_up = "low";

dffeas \result_a_c_se[8] (
	.clk(clk),
	.d(\gen_dsp_only:m_ac|auto_generated|dffe3a[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[8]~q ),
	.prn(vcc));
defparam \result_a_c_se[8] .is_wysiwyg = "true";
defparam \result_a_c_se[8] .power_up = "low";

dffeas \result_b_d_se[8] (
	.clk(clk),
	.d(\gen_dsp_only:m_bd|auto_generated|dffe3a[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[8]~q ),
	.prn(vcc));
defparam \result_b_d_se[8] .is_wysiwyg = "true";
defparam \result_b_d_se[8] .power_up = "low";

dffeas \result_a_c_se[7] (
	.clk(clk),
	.d(\gen_dsp_only:m_ac|auto_generated|dffe3a[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[7]~q ),
	.prn(vcc));
defparam \result_a_c_se[7] .is_wysiwyg = "true";
defparam \result_a_c_se[7] .power_up = "low";

dffeas \result_b_d_se[7] (
	.clk(clk),
	.d(\gen_dsp_only:m_bd|auto_generated|dffe3a[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[7]~q ),
	.prn(vcc));
defparam \result_b_d_se[7] .is_wysiwyg = "true";
defparam \result_b_d_se[7] .power_up = "low";

dffeas \result_a_c_se[6] (
	.clk(clk),
	.d(\gen_dsp_only:m_ac|auto_generated|dffe3a[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[6]~q ),
	.prn(vcc));
defparam \result_a_c_se[6] .is_wysiwyg = "true";
defparam \result_a_c_se[6] .power_up = "low";

dffeas \result_b_d_se[6] (
	.clk(clk),
	.d(\gen_dsp_only:m_bd|auto_generated|dffe3a[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[6]~q ),
	.prn(vcc));
defparam \result_b_d_se[6] .is_wysiwyg = "true";
defparam \result_b_d_se[6] .power_up = "low";

dffeas \result_a_c_se[5] (
	.clk(clk),
	.d(\gen_dsp_only:m_ac|auto_generated|dffe3a[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[5]~q ),
	.prn(vcc));
defparam \result_a_c_se[5] .is_wysiwyg = "true";
defparam \result_a_c_se[5] .power_up = "low";

dffeas \result_b_d_se[5] (
	.clk(clk),
	.d(\gen_dsp_only:m_bd|auto_generated|dffe3a[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[5]~q ),
	.prn(vcc));
defparam \result_b_d_se[5] .is_wysiwyg = "true";
defparam \result_b_d_se[5] .power_up = "low";

dffeas \result_a_c_se[4] (
	.clk(clk),
	.d(\gen_dsp_only:m_ac|auto_generated|dffe3a[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[4]~q ),
	.prn(vcc));
defparam \result_a_c_se[4] .is_wysiwyg = "true";
defparam \result_a_c_se[4] .power_up = "low";

dffeas \result_b_d_se[4] (
	.clk(clk),
	.d(\gen_dsp_only:m_bd|auto_generated|dffe3a[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[4]~q ),
	.prn(vcc));
defparam \result_b_d_se[4] .is_wysiwyg = "true";
defparam \result_b_d_se[4] .power_up = "low";

dffeas \result_a_c_se[3] (
	.clk(clk),
	.d(\gen_dsp_only:m_ac|auto_generated|dffe3a[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[3]~q ),
	.prn(vcc));
defparam \result_a_c_se[3] .is_wysiwyg = "true";
defparam \result_a_c_se[3] .power_up = "low";

dffeas \result_b_d_se[3] (
	.clk(clk),
	.d(\gen_dsp_only:m_bd|auto_generated|dffe3a[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[3]~q ),
	.prn(vcc));
defparam \result_b_d_se[3] .is_wysiwyg = "true";
defparam \result_b_d_se[3] .power_up = "low";

dffeas \result_a_c_se[2] (
	.clk(clk),
	.d(\gen_dsp_only:m_ac|auto_generated|dffe3a[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[2]~q ),
	.prn(vcc));
defparam \result_a_c_se[2] .is_wysiwyg = "true";
defparam \result_a_c_se[2] .power_up = "low";

dffeas \result_b_d_se[2] (
	.clk(clk),
	.d(\gen_dsp_only:m_bd|auto_generated|dffe3a[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[2]~q ),
	.prn(vcc));
defparam \result_b_d_se[2] .is_wysiwyg = "true";
defparam \result_b_d_se[2] .power_up = "low";

dffeas \result_a_c_se[1] (
	.clk(clk),
	.d(\gen_dsp_only:m_ac|auto_generated|dffe3a[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[1]~q ),
	.prn(vcc));
defparam \result_a_c_se[1] .is_wysiwyg = "true";
defparam \result_a_c_se[1] .power_up = "low";

dffeas \result_b_d_se[1] (
	.clk(clk),
	.d(\gen_dsp_only:m_bd|auto_generated|dffe3a[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[1]~q ),
	.prn(vcc));
defparam \result_b_d_se[1] .is_wysiwyg = "true";
defparam \result_b_d_se[1] .power_up = "low";

dffeas \result_a_c_se[0] (
	.clk(clk),
	.d(\gen_dsp_only:m_ac|auto_generated|dffe3a[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[0]~q ),
	.prn(vcc));
defparam \result_a_c_se[0] .is_wysiwyg = "true";
defparam \result_a_c_se[0] .power_up = "low";

dffeas \result_b_d_se[0] (
	.clk(clk),
	.d(\gen_dsp_only:m_bd|auto_generated|dffe3a[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[0]~q ),
	.prn(vcc));
defparam \result_b_d_se[0] .is_wysiwyg = "true";
defparam \result_b_d_se[0] .power_up = "low";

dffeas \result_a_c_se[15] (
	.clk(clk),
	.d(\gen_dsp_only:m_ac|auto_generated|dffe3a[15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[15]~q ),
	.prn(vcc));
defparam \result_a_c_se[15] .is_wysiwyg = "true";
defparam \result_a_c_se[15] .power_up = "low";

dffeas \result_b_d_se[15] (
	.clk(clk),
	.d(\gen_dsp_only:m_bd|auto_generated|dffe3a[15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[15]~q ),
	.prn(vcc));
defparam \result_b_d_se[15] .is_wysiwyg = "true";
defparam \result_b_d_se[15] .power_up = "low";

dffeas \result_a_c_se[14] (
	.clk(clk),
	.d(\gen_dsp_only:m_ac|auto_generated|dffe3a[14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[14]~q ),
	.prn(vcc));
defparam \result_a_c_se[14] .is_wysiwyg = "true";
defparam \result_a_c_se[14] .power_up = "low";

dffeas \result_b_d_se[14] (
	.clk(clk),
	.d(\gen_dsp_only:m_bd|auto_generated|dffe3a[14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[14]~q ),
	.prn(vcc));
defparam \result_b_d_se[14] .is_wysiwyg = "true";
defparam \result_b_d_se[14] .power_up = "low";

dffeas \result_a_c_se[13] (
	.clk(clk),
	.d(\gen_dsp_only:m_ac|auto_generated|dffe3a[13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[13]~q ),
	.prn(vcc));
defparam \result_a_c_se[13] .is_wysiwyg = "true";
defparam \result_a_c_se[13] .power_up = "low";

dffeas \result_b_d_se[13] (
	.clk(clk),
	.d(\gen_dsp_only:m_bd|auto_generated|dffe3a[13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[13]~q ),
	.prn(vcc));
defparam \result_b_d_se[13] .is_wysiwyg = "true";
defparam \result_b_d_se[13] .power_up = "low";

dffeas \result_a_c_se[12] (
	.clk(clk),
	.d(\gen_dsp_only:m_ac|auto_generated|dffe3a[12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[12]~q ),
	.prn(vcc));
defparam \result_a_c_se[12] .is_wysiwyg = "true";
defparam \result_a_c_se[12] .power_up = "low";

dffeas \result_b_d_se[12] (
	.clk(clk),
	.d(\gen_dsp_only:m_bd|auto_generated|dffe3a[12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[12]~q ),
	.prn(vcc));
defparam \result_b_d_se[12] .is_wysiwyg = "true";
defparam \result_b_d_se[12] .power_up = "low";

dffeas \real_out[3] (
	.clk(clk),
	.d(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(real_out_3),
	.prn(vcc));
defparam \real_out[3] .is_wysiwyg = "true";
defparam \real_out[3] .power_up = "low";

dffeas \real_out[7] (
	.clk(clk),
	.d(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(real_out_7),
	.prn(vcc));
defparam \real_out[7] .is_wysiwyg = "true";
defparam \real_out[7] .power_up = "low";

dffeas \real_out[4] (
	.clk(clk),
	.d(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(real_out_4),
	.prn(vcc));
defparam \real_out[4] .is_wysiwyg = "true";
defparam \real_out[4] .power_up = "low";

dffeas \real_out[5] (
	.clk(clk),
	.d(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(real_out_5),
	.prn(vcc));
defparam \real_out[5] .is_wysiwyg = "true";
defparam \real_out[5] .power_up = "low";

dffeas \real_out[6] (
	.clk(clk),
	.d(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(real_out_6),
	.prn(vcc));
defparam \real_out[6] .is_wysiwyg = "true";
defparam \real_out[6] .power_up = "low";

dffeas \real_out[1] (
	.clk(clk),
	.d(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(real_out_1),
	.prn(vcc));
defparam \real_out[1] .is_wysiwyg = "true";
defparam \real_out[1] .power_up = "low";

dffeas \real_out[0] (
	.clk(clk),
	.d(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(real_out_0),
	.prn(vcc));
defparam \real_out[0] .is_wysiwyg = "true";
defparam \real_out[0] .power_up = "low";

dffeas \real_out[2] (
	.clk(clk),
	.d(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(real_out_2),
	.prn(vcc));
defparam \real_out[2] .is_wysiwyg = "true";
defparam \real_out[2] .power_up = "low";

endmodule

module fft_asj_fft_pround_fft_120_2 (
	pipeline_dffe_11,
	pipeline_dffe_15,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	result_real_1_tmp_11,
	result_real_1_tmp_10,
	result_real_1_tmp_9,
	result_real_1_tmp_8,
	result_real_1_tmp_7,
	result_real_1_tmp_6,
	result_real_1_tmp_5,
	result_real_1_tmp_4,
	result_real_1_tmp_3,
	result_real_1_tmp_2,
	result_real_1_tmp_1,
	result_real_1_tmp_0,
	result_real_1_tmp_15,
	result_real_1_tmp_14,
	result_real_1_tmp_13,
	result_real_1_tmp_12,
	pipeline_dffe_9,
	pipeline_dffe_8,
	pipeline_dffe_10,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_11;
output 	pipeline_dffe_15;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
input 	result_real_1_tmp_11;
input 	result_real_1_tmp_10;
input 	result_real_1_tmp_9;
input 	result_real_1_tmp_8;
input 	result_real_1_tmp_7;
input 	result_real_1_tmp_6;
input 	result_real_1_tmp_5;
input 	result_real_1_tmp_4;
input 	result_real_1_tmp_3;
input 	result_real_1_tmp_2;
input 	result_real_1_tmp_1;
input 	result_real_1_tmp_0;
input 	result_real_1_tmp_15;
input 	result_real_1_tmp_14;
input 	result_real_1_tmp_13;
input 	result_real_1_tmp_12;
output 	pipeline_dffe_9;
output 	pipeline_dffe_8;
output 	pipeline_dffe_10;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_LPM_ADD_SUB_3 \gbrnd:nev:gp:lpm_add_sub_component (
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_14(pipeline_dffe_14),
	.result_real_1_tmp_11(result_real_1_tmp_11),
	.result_real_1_tmp_10(result_real_1_tmp_10),
	.result_real_1_tmp_9(result_real_1_tmp_9),
	.result_real_1_tmp_8(result_real_1_tmp_8),
	.result_real_1_tmp_7(result_real_1_tmp_7),
	.result_real_1_tmp_6(result_real_1_tmp_6),
	.result_real_1_tmp_5(result_real_1_tmp_5),
	.result_real_1_tmp_4(result_real_1_tmp_4),
	.result_real_1_tmp_3(result_real_1_tmp_3),
	.result_real_1_tmp_2(result_real_1_tmp_2),
	.result_real_1_tmp_1(result_real_1_tmp_1),
	.result_real_1_tmp_0(result_real_1_tmp_0),
	.result_real_1_tmp_15(result_real_1_tmp_15),
	.result_real_1_tmp_14(result_real_1_tmp_14),
	.result_real_1_tmp_13(result_real_1_tmp_13),
	.result_real_1_tmp_12(result_real_1_tmp_12),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_10(pipeline_dffe_10),
	.clken(global_clock_enable),
	.clock(clk));

endmodule

module fft_LPM_ADD_SUB_3 (
	pipeline_dffe_11,
	pipeline_dffe_15,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	result_real_1_tmp_11,
	result_real_1_tmp_10,
	result_real_1_tmp_9,
	result_real_1_tmp_8,
	result_real_1_tmp_7,
	result_real_1_tmp_6,
	result_real_1_tmp_5,
	result_real_1_tmp_4,
	result_real_1_tmp_3,
	result_real_1_tmp_2,
	result_real_1_tmp_1,
	result_real_1_tmp_0,
	result_real_1_tmp_15,
	result_real_1_tmp_14,
	result_real_1_tmp_13,
	result_real_1_tmp_12,
	pipeline_dffe_9,
	pipeline_dffe_8,
	pipeline_dffe_10,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_11;
output 	pipeline_dffe_15;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
input 	result_real_1_tmp_11;
input 	result_real_1_tmp_10;
input 	result_real_1_tmp_9;
input 	result_real_1_tmp_8;
input 	result_real_1_tmp_7;
input 	result_real_1_tmp_6;
input 	result_real_1_tmp_5;
input 	result_real_1_tmp_4;
input 	result_real_1_tmp_3;
input 	result_real_1_tmp_2;
input 	result_real_1_tmp_1;
input 	result_real_1_tmp_0;
input 	result_real_1_tmp_15;
input 	result_real_1_tmp_14;
input 	result_real_1_tmp_13;
input 	result_real_1_tmp_12;
output 	pipeline_dffe_9;
output 	pipeline_dffe_8;
output 	pipeline_dffe_10;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_add_sub_dmj_2 auto_generated(
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_14(pipeline_dffe_14),
	.result_real_1_tmp_11(result_real_1_tmp_11),
	.result_real_1_tmp_10(result_real_1_tmp_10),
	.result_real_1_tmp_9(result_real_1_tmp_9),
	.result_real_1_tmp_8(result_real_1_tmp_8),
	.result_real_1_tmp_7(result_real_1_tmp_7),
	.result_real_1_tmp_6(result_real_1_tmp_6),
	.result_real_1_tmp_5(result_real_1_tmp_5),
	.result_real_1_tmp_4(result_real_1_tmp_4),
	.result_real_1_tmp_3(result_real_1_tmp_3),
	.result_real_1_tmp_2(result_real_1_tmp_2),
	.result_real_1_tmp_1(result_real_1_tmp_1),
	.result_real_1_tmp_0(result_real_1_tmp_0),
	.result_real_1_tmp_15(result_real_1_tmp_15),
	.result_real_1_tmp_14(result_real_1_tmp_14),
	.result_real_1_tmp_13(result_real_1_tmp_13),
	.result_real_1_tmp_12(result_real_1_tmp_12),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_10(pipeline_dffe_10),
	.clken(clken),
	.clock(clock));

endmodule

module fft_add_sub_dmj_2 (
	pipeline_dffe_11,
	pipeline_dffe_15,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	result_real_1_tmp_11,
	result_real_1_tmp_10,
	result_real_1_tmp_9,
	result_real_1_tmp_8,
	result_real_1_tmp_7,
	result_real_1_tmp_6,
	result_real_1_tmp_5,
	result_real_1_tmp_4,
	result_real_1_tmp_3,
	result_real_1_tmp_2,
	result_real_1_tmp_1,
	result_real_1_tmp_0,
	result_real_1_tmp_15,
	result_real_1_tmp_14,
	result_real_1_tmp_13,
	result_real_1_tmp_12,
	pipeline_dffe_9,
	pipeline_dffe_8,
	pipeline_dffe_10,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_11;
output 	pipeline_dffe_15;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
input 	result_real_1_tmp_11;
input 	result_real_1_tmp_10;
input 	result_real_1_tmp_9;
input 	result_real_1_tmp_8;
input 	result_real_1_tmp_7;
input 	result_real_1_tmp_6;
input 	result_real_1_tmp_5;
input 	result_real_1_tmp_4;
input 	result_real_1_tmp_3;
input 	result_real_1_tmp_2;
input 	result_real_1_tmp_1;
input 	result_real_1_tmp_0;
input 	result_real_1_tmp_15;
input 	result_real_1_tmp_14;
input 	result_real_1_tmp_13;
input 	result_real_1_tmp_12;
output 	pipeline_dffe_9;
output 	pipeline_dffe_8;
output 	pipeline_dffe_10;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~9_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~11_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~13_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~15_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~17_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~19_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~21_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~23_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~27 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~29 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~31 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~32_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~33 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~35 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~37 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~39 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~40_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~34_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~36_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~38_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~30_combout ;


dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_15),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_12),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_13),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_14),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .power_up = "low";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~9 (
	.dataa(result_real_1_tmp_15),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~9_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~9 .lut_mask = 16'h0055;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~11 (
	.dataa(result_real_1_tmp_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~9_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~11_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~11 .lut_mask = 16'h005F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~11 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~13 (
	.dataa(result_real_1_tmp_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~11_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~13_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~13 .lut_mask = 16'h00AF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~13 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~15 (
	.dataa(result_real_1_tmp_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~13_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~15_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~15 .lut_mask = 16'h005F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~15 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~17 (
	.dataa(result_real_1_tmp_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~15_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~17_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~17 .lut_mask = 16'h00AF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~17 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~19 (
	.dataa(result_real_1_tmp_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~17_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~19_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~19 .lut_mask = 16'h005F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~19 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~21 (
	.dataa(result_real_1_tmp_5),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~19_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~21_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~21 .lut_mask = 16'h00AF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~21 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~23 (
	.dataa(result_real_1_tmp_6),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~21_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~23_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~23 .lut_mask = 16'h005F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~23 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25 (
	.dataa(result_real_1_tmp_7),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~23_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25 .lut_mask = 16'h00AF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26 (
	.dataa(result_real_1_tmp_8),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25_cout ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~27 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28 (
	.dataa(result_real_1_tmp_9),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~27 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~29 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28 .lut_mask = 16'h5AAF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~30 (
	.dataa(result_real_1_tmp_10),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~29 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~30_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~31 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~30 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~30 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~32 (
	.dataa(result_real_1_tmp_11),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~31 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~32_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~33 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~32 .lut_mask = 16'h5AAF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~32 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~34 (
	.dataa(result_real_1_tmp_12),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~33 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~34_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~35 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~34 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~34 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~36 (
	.dataa(result_real_1_tmp_13),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~35 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~36_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~37 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~36 .lut_mask = 16'h5AAF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~36 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~38 (
	.dataa(result_real_1_tmp_14),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~37 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~38_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~39 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~38 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~38 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~40 (
	.dataa(result_real_1_tmp_15),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~39 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~40_combout ),
	.cout());
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~40 .lut_mask = 16'h5A5A;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~40 .sum_lutc_input = "cin";

endmodule

module fft_asj_fft_pround_fft_120_3 (
	pipeline_dffe_11,
	pipeline_dffe_15,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	result_imag_1_11,
	result_imag_1_10,
	result_imag_1_9,
	result_imag_1_8,
	result_imag_1_7,
	result_imag_1_6,
	result_imag_1_5,
	result_imag_1_4,
	result_imag_1_3,
	result_imag_1_2,
	result_imag_1_1,
	result_imag_1_0,
	result_imag_1_15,
	result_imag_1_14,
	result_imag_1_13,
	result_imag_1_12,
	pipeline_dffe_9,
	pipeline_dffe_8,
	pipeline_dffe_10,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_11;
output 	pipeline_dffe_15;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
input 	result_imag_1_11;
input 	result_imag_1_10;
input 	result_imag_1_9;
input 	result_imag_1_8;
input 	result_imag_1_7;
input 	result_imag_1_6;
input 	result_imag_1_5;
input 	result_imag_1_4;
input 	result_imag_1_3;
input 	result_imag_1_2;
input 	result_imag_1_1;
input 	result_imag_1_0;
input 	result_imag_1_15;
input 	result_imag_1_14;
input 	result_imag_1_13;
input 	result_imag_1_12;
output 	pipeline_dffe_9;
output 	pipeline_dffe_8;
output 	pipeline_dffe_10;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_LPM_ADD_SUB_4 \gbrnd:nev:gp:lpm_add_sub_component (
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_14(pipeline_dffe_14),
	.result_imag_1_11(result_imag_1_11),
	.result_imag_1_10(result_imag_1_10),
	.result_imag_1_9(result_imag_1_9),
	.result_imag_1_8(result_imag_1_8),
	.result_imag_1_7(result_imag_1_7),
	.result_imag_1_6(result_imag_1_6),
	.result_imag_1_5(result_imag_1_5),
	.result_imag_1_4(result_imag_1_4),
	.result_imag_1_3(result_imag_1_3),
	.result_imag_1_2(result_imag_1_2),
	.result_imag_1_1(result_imag_1_1),
	.result_imag_1_0(result_imag_1_0),
	.result_imag_1_15(result_imag_1_15),
	.result_imag_1_14(result_imag_1_14),
	.result_imag_1_13(result_imag_1_13),
	.result_imag_1_12(result_imag_1_12),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_10(pipeline_dffe_10),
	.clken(global_clock_enable),
	.clock(clk));

endmodule

module fft_LPM_ADD_SUB_4 (
	pipeline_dffe_11,
	pipeline_dffe_15,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	result_imag_1_11,
	result_imag_1_10,
	result_imag_1_9,
	result_imag_1_8,
	result_imag_1_7,
	result_imag_1_6,
	result_imag_1_5,
	result_imag_1_4,
	result_imag_1_3,
	result_imag_1_2,
	result_imag_1_1,
	result_imag_1_0,
	result_imag_1_15,
	result_imag_1_14,
	result_imag_1_13,
	result_imag_1_12,
	pipeline_dffe_9,
	pipeline_dffe_8,
	pipeline_dffe_10,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_11;
output 	pipeline_dffe_15;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
input 	result_imag_1_11;
input 	result_imag_1_10;
input 	result_imag_1_9;
input 	result_imag_1_8;
input 	result_imag_1_7;
input 	result_imag_1_6;
input 	result_imag_1_5;
input 	result_imag_1_4;
input 	result_imag_1_3;
input 	result_imag_1_2;
input 	result_imag_1_1;
input 	result_imag_1_0;
input 	result_imag_1_15;
input 	result_imag_1_14;
input 	result_imag_1_13;
input 	result_imag_1_12;
output 	pipeline_dffe_9;
output 	pipeline_dffe_8;
output 	pipeline_dffe_10;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_add_sub_dmj_3 auto_generated(
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_14(pipeline_dffe_14),
	.result_imag_1_11(result_imag_1_11),
	.result_imag_1_10(result_imag_1_10),
	.result_imag_1_9(result_imag_1_9),
	.result_imag_1_8(result_imag_1_8),
	.result_imag_1_7(result_imag_1_7),
	.result_imag_1_6(result_imag_1_6),
	.result_imag_1_5(result_imag_1_5),
	.result_imag_1_4(result_imag_1_4),
	.result_imag_1_3(result_imag_1_3),
	.result_imag_1_2(result_imag_1_2),
	.result_imag_1_1(result_imag_1_1),
	.result_imag_1_0(result_imag_1_0),
	.result_imag_1_15(result_imag_1_15),
	.result_imag_1_14(result_imag_1_14),
	.result_imag_1_13(result_imag_1_13),
	.result_imag_1_12(result_imag_1_12),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_10(pipeline_dffe_10),
	.clken(clken),
	.clock(clock));

endmodule

module fft_add_sub_dmj_3 (
	pipeline_dffe_11,
	pipeline_dffe_15,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	result_imag_1_11,
	result_imag_1_10,
	result_imag_1_9,
	result_imag_1_8,
	result_imag_1_7,
	result_imag_1_6,
	result_imag_1_5,
	result_imag_1_4,
	result_imag_1_3,
	result_imag_1_2,
	result_imag_1_1,
	result_imag_1_0,
	result_imag_1_15,
	result_imag_1_14,
	result_imag_1_13,
	result_imag_1_12,
	pipeline_dffe_9,
	pipeline_dffe_8,
	pipeline_dffe_10,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_11;
output 	pipeline_dffe_15;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
input 	result_imag_1_11;
input 	result_imag_1_10;
input 	result_imag_1_9;
input 	result_imag_1_8;
input 	result_imag_1_7;
input 	result_imag_1_6;
input 	result_imag_1_5;
input 	result_imag_1_4;
input 	result_imag_1_3;
input 	result_imag_1_2;
input 	result_imag_1_1;
input 	result_imag_1_0;
input 	result_imag_1_15;
input 	result_imag_1_14;
input 	result_imag_1_13;
input 	result_imag_1_12;
output 	pipeline_dffe_9;
output 	pipeline_dffe_8;
output 	pipeline_dffe_10;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~9_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~11_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~13_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~15_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~17_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~19_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~21_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~23_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~27 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~29 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~31 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~32_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~33 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~35 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~37 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~39 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~40_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~34_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~36_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~38_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~30_combout ;


dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_15),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_12),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_13),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_14),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .power_up = "low";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~9 (
	.dataa(result_imag_1_15),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~9_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~9 .lut_mask = 16'h0055;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~11 (
	.dataa(result_imag_1_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~9_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~11_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~11 .lut_mask = 16'h005F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~11 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~13 (
	.dataa(result_imag_1_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~11_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~13_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~13 .lut_mask = 16'h00AF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~13 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~15 (
	.dataa(result_imag_1_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~13_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~15_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~15 .lut_mask = 16'h005F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~15 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~17 (
	.dataa(result_imag_1_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~15_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~17_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~17 .lut_mask = 16'h00AF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~17 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~19 (
	.dataa(result_imag_1_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~17_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~19_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~19 .lut_mask = 16'h005F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~19 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~21 (
	.dataa(result_imag_1_5),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~19_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~21_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~21 .lut_mask = 16'h00AF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~21 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~23 (
	.dataa(result_imag_1_6),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~21_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~23_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~23 .lut_mask = 16'h005F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~23 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25 (
	.dataa(result_imag_1_7),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~23_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25 .lut_mask = 16'h00AF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26 (
	.dataa(result_imag_1_8),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25_cout ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~27 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28 (
	.dataa(result_imag_1_9),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~27 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~29 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28 .lut_mask = 16'h5AAF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~30 (
	.dataa(result_imag_1_10),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~29 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~30_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~31 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~30 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~30 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~32 (
	.dataa(result_imag_1_11),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~31 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~32_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~33 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~32 .lut_mask = 16'h5AAF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~32 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~34 (
	.dataa(result_imag_1_12),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~33 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~34_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~35 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~34 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~34 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~36 (
	.dataa(result_imag_1_13),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~35 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~36_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~37 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~36 .lut_mask = 16'h5AAF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~36 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~38 (
	.dataa(result_imag_1_14),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~37 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~38_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~39 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~38 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~38 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~40 (
	.dataa(result_imag_1_15),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~39 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~40_combout ),
	.cout());
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~40 .lut_mask = 16'h5A5A;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~40 .sum_lutc_input = "cin";

endmodule

module fft_LPM_MULT_4 (
	dataa,
	datab,
	clken,
	dffe3a_11,
	dffe3a_10,
	dffe3a_9,
	dffe3a_8,
	dffe3a_7,
	dffe3a_6,
	dffe3a_5,
	dffe3a_4,
	dffe3a_3,
	dffe3a_2,
	dffe3a_1,
	dffe3a_0,
	dffe3a_15,
	dffe3a_14,
	dffe3a_13,
	dffe3a_12,
	clock)/* synthesis synthesis_greybox=1 */;
input 	[8:0] dataa;
input 	[8:0] datab;
input 	clken;
output 	dffe3a_11;
output 	dffe3a_10;
output 	dffe3a_9;
output 	dffe3a_8;
output 	dffe3a_7;
output 	dffe3a_6;
output 	dffe3a_5;
output 	dffe3a_4;
output 	dffe3a_3;
output 	dffe3a_2;
output 	dffe3a_1;
output 	dffe3a_0;
output 	dffe3a_15;
output 	dffe3a_14;
output 	dffe3a_13;
output 	dffe3a_12;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_mult_4p01_1 auto_generated(
	.dataa({dataa[8],dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.datab({datab[8],datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.clken(clken),
	.dffe3a_11(dffe3a_11),
	.dffe3a_10(dffe3a_10),
	.dffe3a_9(dffe3a_9),
	.dffe3a_8(dffe3a_8),
	.dffe3a_7(dffe3a_7),
	.dffe3a_6(dffe3a_6),
	.dffe3a_5(dffe3a_5),
	.dffe3a_4(dffe3a_4),
	.dffe3a_3(dffe3a_3),
	.dffe3a_2(dffe3a_2),
	.dffe3a_1(dffe3a_1),
	.dffe3a_0(dffe3a_0),
	.dffe3a_15(dffe3a_15),
	.dffe3a_14(dffe3a_14),
	.dffe3a_13(dffe3a_13),
	.dffe3a_12(dffe3a_12),
	.clock(clock));

endmodule

module fft_mult_4p01_1 (
	dataa,
	datab,
	clken,
	dffe3a_11,
	dffe3a_10,
	dffe3a_9,
	dffe3a_8,
	dffe3a_7,
	dffe3a_6,
	dffe3a_5,
	dffe3a_4,
	dffe3a_3,
	dffe3a_2,
	dffe3a_1,
	dffe3a_0,
	dffe3a_15,
	dffe3a_14,
	dffe3a_13,
	dffe3a_12,
	clock)/* synthesis synthesis_greybox=1 */;
input 	[8:0] dataa;
input 	[8:0] datab;
input 	clken;
output 	dffe3a_11;
output 	dffe3a_10;
output 	dffe3a_9;
output 	dffe3a_8;
output 	dffe3a_7;
output 	dffe3a_6;
output 	dffe3a_5;
output 	dffe3a_4;
output 	dffe3a_3;
output 	dffe3a_2;
output 	dffe3a_1;
output 	dffe3a_0;
output 	dffe3a_15;
output 	dffe3a_14;
output 	dffe3a_13;
output 	dffe3a_12;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT16 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT17 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~dataout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT1 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT2 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT3 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT4 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT5 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT6 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT7 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT8 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT9 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT10 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT11 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT12 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT13 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT14 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT15 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT16 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT17 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT11 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT10 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT9 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT8 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT7 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT6 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT5 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT4 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT3 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT2 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT1 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~dataout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT15 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT14 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT13 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT12 ;

wire [35:0] \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus ;
wire [35:0] \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus ;

assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~dataout  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [0];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT1  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [1];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT2  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [2];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT3  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [3];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT4  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [4];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT5  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [5];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT6  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [6];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT7  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [7];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT8  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [8];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT9  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [9];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT10  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [10];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT11  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [11];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT12  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [12];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT13  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [13];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT14  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [14];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT15  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [15];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT16  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [16];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT17  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [17];

assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~dataout  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [0];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT1  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [1];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT2  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [2];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT3  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [3];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT4  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [4];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT5  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [5];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT6  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [6];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT7  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [7];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT8  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [8];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT9  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [9];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT10  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [10];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT11  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [11];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT12  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [12];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT13  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [13];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT14  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [14];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT15  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [15];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT16  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [16];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT17  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [17];

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[11] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT11 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_11),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[11] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[11] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[10] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT10 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_10),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[10] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[10] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[9] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT9 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_9),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[9] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[9] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[8] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT8 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_8),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[8] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[8] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[7] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT7 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_7),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[7] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[7] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[6] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT6 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_6),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[6] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[6] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[5] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT5 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_5),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[5] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[5] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[4] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT4 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_4),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[4] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[4] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[3] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT3 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_3),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[3] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[3] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[2] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT2 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_2),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[2] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[2] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[1] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT1 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_1),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[1] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[1] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[0] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~dataout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_0),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[0] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[0] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[15] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT15 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_15),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[15] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[15] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[14] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT14 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_14),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[14] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[14] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[13] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT13 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_13),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[13] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[13] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[12] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT12 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_12),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[12] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[12] .power_up = "low";

cycloneiii_mac_mult \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1 (
	.signa(vcc),
	.signb(vcc),
	.clk(clock),
	.aclr(gnd),
	.ena(clken),
	.dataa({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dataa[8],dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.datab({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,datab[8],datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.dataout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1 .dataa_clock = "0";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1 .dataa_width = 9;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1 .datab_clock = "0";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1 .datab_width = 9;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1 .signa_clock = "none";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1 .signb_clock = "none";

cycloneiii_mac_out \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2 (
	.clk(clock),
	.aclr(gnd),
	.ena(clken),
	.dataa({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT17 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT16 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT15 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT14 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT13 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT12 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT11 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT10 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT9 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT8 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT7 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT6 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT5 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT4 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT3 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT2 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT1 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~dataout }),
	.dataout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2 .dataa_width = 18;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2 .output_clock = "0";

endmodule

module fft_LPM_MULT_5 (
	dataa,
	clken,
	dffe3a_11,
	dffe3a_10,
	dffe3a_9,
	dffe3a_8,
	dffe3a_7,
	dffe3a_6,
	dffe3a_5,
	dffe3a_4,
	dffe3a_3,
	dffe3a_2,
	dffe3a_1,
	dffe3a_0,
	dffe3a_15,
	dffe3a_14,
	dffe3a_13,
	dffe3a_12,
	datab,
	clock)/* synthesis synthesis_greybox=1 */;
input 	[8:0] dataa;
input 	clken;
output 	dffe3a_11;
output 	dffe3a_10;
output 	dffe3a_9;
output 	dffe3a_8;
output 	dffe3a_7;
output 	dffe3a_6;
output 	dffe3a_5;
output 	dffe3a_4;
output 	dffe3a_3;
output 	dffe3a_2;
output 	dffe3a_1;
output 	dffe3a_0;
output 	dffe3a_15;
output 	dffe3a_14;
output 	dffe3a_13;
output 	dffe3a_12;
input 	[8:0] datab;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_mult_0p01_2 auto_generated(
	.dataa({dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.clken(clken),
	.dffe3a_11(dffe3a_11),
	.dffe3a_10(dffe3a_10),
	.dffe3a_9(dffe3a_9),
	.dffe3a_8(dffe3a_8),
	.dffe3a_7(dffe3a_7),
	.dffe3a_6(dffe3a_6),
	.dffe3a_5(dffe3a_5),
	.dffe3a_4(dffe3a_4),
	.dffe3a_3(dffe3a_3),
	.dffe3a_2(dffe3a_2),
	.dffe3a_1(dffe3a_1),
	.dffe3a_0(dffe3a_0),
	.dffe3a_15(dffe3a_15),
	.dffe3a_14(dffe3a_14),
	.dffe3a_13(dffe3a_13),
	.dffe3a_12(dffe3a_12),
	.datab({datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.clock(clock));

endmodule

module fft_mult_0p01_2 (
	dataa,
	clken,
	dffe3a_11,
	dffe3a_10,
	dffe3a_9,
	dffe3a_8,
	dffe3a_7,
	dffe3a_6,
	dffe3a_5,
	dffe3a_4,
	dffe3a_3,
	dffe3a_2,
	dffe3a_1,
	dffe3a_0,
	dffe3a_15,
	dffe3a_14,
	dffe3a_13,
	dffe3a_12,
	datab,
	clock)/* synthesis synthesis_greybox=1 */;
input 	[7:0] dataa;
input 	clken;
output 	dffe3a_11;
output 	dffe3a_10;
output 	dffe3a_9;
output 	dffe3a_8;
output 	dffe3a_7;
output 	dffe3a_6;
output 	dffe3a_5;
output 	dffe3a_4;
output 	dffe3a_3;
output 	dffe3a_2;
output 	dffe3a_1;
output 	dffe3a_0;
output 	dffe3a_15;
output 	dffe3a_14;
output 	dffe3a_13;
output 	dffe3a_12;
input 	[7:0] datab;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1~dataout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT1 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT2 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT3 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT4 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT5 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT6 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT7 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT8 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT9 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT10 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT11 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT12 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT13 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT14 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT15 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT11 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT10 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT9 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT8 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT7 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT6 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT5 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT4 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT3 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT2 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT1 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2~dataout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT15 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT14 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT13 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT12 ;

wire [35:0] \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2_DATAOUT_bus ;
wire [35:0] \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1_DATAOUT_bus ;

assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2~dataout  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2_DATAOUT_bus [0];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT1  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2_DATAOUT_bus [1];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT2  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2_DATAOUT_bus [2];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT3  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2_DATAOUT_bus [3];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT4  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2_DATAOUT_bus [4];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT5  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2_DATAOUT_bus [5];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT6  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2_DATAOUT_bus [6];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT7  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2_DATAOUT_bus [7];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT8  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2_DATAOUT_bus [8];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT9  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2_DATAOUT_bus [9];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT10  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2_DATAOUT_bus [10];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT11  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2_DATAOUT_bus [11];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT12  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2_DATAOUT_bus [12];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT13  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2_DATAOUT_bus [13];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT14  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2_DATAOUT_bus [14];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT15  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2_DATAOUT_bus [15];

assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1~dataout  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1_DATAOUT_bus [0];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT1  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1_DATAOUT_bus [1];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT2  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1_DATAOUT_bus [2];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT3  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1_DATAOUT_bus [3];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT4  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1_DATAOUT_bus [4];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT5  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1_DATAOUT_bus [5];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT6  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1_DATAOUT_bus [6];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT7  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1_DATAOUT_bus [7];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT8  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1_DATAOUT_bus [8];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT9  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1_DATAOUT_bus [9];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT10  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1_DATAOUT_bus [10];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT11  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1_DATAOUT_bus [11];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT12  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1_DATAOUT_bus [12];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT13  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1_DATAOUT_bus [13];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT14  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1_DATAOUT_bus [14];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT15  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1_DATAOUT_bus [15];

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|dffe3a[11] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT11 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_11),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|dffe3a[11] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|dffe3a[11] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|dffe3a[10] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT10 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_10),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|dffe3a[10] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|dffe3a[10] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|dffe3a[9] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT9 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_9),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|dffe3a[9] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|dffe3a[9] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|dffe3a[8] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT8 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_8),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|dffe3a[8] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|dffe3a[8] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|dffe3a[7] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT7 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_7),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|dffe3a[7] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|dffe3a[7] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|dffe3a[6] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT6 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_6),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|dffe3a[6] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|dffe3a[6] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|dffe3a[5] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT5 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_5),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|dffe3a[5] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|dffe3a[5] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|dffe3a[4] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT4 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_4),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|dffe3a[4] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|dffe3a[4] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|dffe3a[3] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT3 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_3),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|dffe3a[3] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|dffe3a[3] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|dffe3a[2] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT2 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_2),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|dffe3a[2] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|dffe3a[2] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|dffe3a[1] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT1 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_1),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|dffe3a[1] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|dffe3a[1] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|dffe3a[0] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2~dataout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_0),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|dffe3a[0] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|dffe3a[0] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|dffe3a[15] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT15 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_15),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|dffe3a[15] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|dffe3a[15] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|dffe3a[14] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT14 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_14),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|dffe3a[14] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|dffe3a[14] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|dffe3a[13] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT13 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_13),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|dffe3a[13] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|dffe3a[13] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|dffe3a[12] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT12 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_12),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|dffe3a[12] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|dffe3a[12] .power_up = "low";

cycloneiii_mac_mult \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1 (
	.signa(vcc),
	.signb(vcc),
	.clk(clock),
	.aclr(gnd),
	.ena(clken),
	.dataa({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.datab({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.dataout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1_DATAOUT_bus ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1 .dataa_clock = "0";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1 .dataa_width = 8;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1 .datab_clock = "0";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1 .datab_width = 8;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1 .signa_clock = "none";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1 .signb_clock = "none";

cycloneiii_mac_out \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2 (
	.clk(clock),
	.aclr(gnd),
	.ena(clken),
	.dataa({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT15 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT14 ,\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT13 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT12 ,\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT11 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT10 ,\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT9 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT8 ,\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT7 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT6 ,\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT5 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT4 ,\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT3 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT2 ,\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT1 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_mult1~dataout }),
	.dataout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2_DATAOUT_bus ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2 .dataa_width = 16;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_ac|auto_generated|mac_out2 .output_clock = "0";

endmodule

module fft_LPM_MULT_6 (
	dataa,
	clken,
	dffe3a_11,
	dffe3a_10,
	dffe3a_9,
	dffe3a_8,
	dffe3a_7,
	dffe3a_6,
	dffe3a_5,
	dffe3a_4,
	dffe3a_3,
	dffe3a_2,
	dffe3a_1,
	dffe3a_0,
	dffe3a_15,
	dffe3a_14,
	dffe3a_13,
	dffe3a_12,
	datab,
	clock)/* synthesis synthesis_greybox=1 */;
input 	[8:0] dataa;
input 	clken;
output 	dffe3a_11;
output 	dffe3a_10;
output 	dffe3a_9;
output 	dffe3a_8;
output 	dffe3a_7;
output 	dffe3a_6;
output 	dffe3a_5;
output 	dffe3a_4;
output 	dffe3a_3;
output 	dffe3a_2;
output 	dffe3a_1;
output 	dffe3a_0;
output 	dffe3a_15;
output 	dffe3a_14;
output 	dffe3a_13;
output 	dffe3a_12;
input 	[8:0] datab;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_mult_0p01_3 auto_generated(
	.dataa({dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.clken(clken),
	.dffe3a_11(dffe3a_11),
	.dffe3a_10(dffe3a_10),
	.dffe3a_9(dffe3a_9),
	.dffe3a_8(dffe3a_8),
	.dffe3a_7(dffe3a_7),
	.dffe3a_6(dffe3a_6),
	.dffe3a_5(dffe3a_5),
	.dffe3a_4(dffe3a_4),
	.dffe3a_3(dffe3a_3),
	.dffe3a_2(dffe3a_2),
	.dffe3a_1(dffe3a_1),
	.dffe3a_0(dffe3a_0),
	.dffe3a_15(dffe3a_15),
	.dffe3a_14(dffe3a_14),
	.dffe3a_13(dffe3a_13),
	.dffe3a_12(dffe3a_12),
	.datab({datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.clock(clock));

endmodule

module fft_mult_0p01_3 (
	dataa,
	clken,
	dffe3a_11,
	dffe3a_10,
	dffe3a_9,
	dffe3a_8,
	dffe3a_7,
	dffe3a_6,
	dffe3a_5,
	dffe3a_4,
	dffe3a_3,
	dffe3a_2,
	dffe3a_1,
	dffe3a_0,
	dffe3a_15,
	dffe3a_14,
	dffe3a_13,
	dffe3a_12,
	datab,
	clock)/* synthesis synthesis_greybox=1 */;
input 	[7:0] dataa;
input 	clken;
output 	dffe3a_11;
output 	dffe3a_10;
output 	dffe3a_9;
output 	dffe3a_8;
output 	dffe3a_7;
output 	dffe3a_6;
output 	dffe3a_5;
output 	dffe3a_4;
output 	dffe3a_3;
output 	dffe3a_2;
output 	dffe3a_1;
output 	dffe3a_0;
output 	dffe3a_15;
output 	dffe3a_14;
output 	dffe3a_13;
output 	dffe3a_12;
input 	[7:0] datab;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1~dataout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT1 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT2 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT3 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT4 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT5 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT6 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT7 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT8 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT9 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT10 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT11 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT12 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT13 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT14 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT15 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT11 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT10 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT9 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT8 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT7 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT6 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT5 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT4 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT3 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT2 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT1 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2~dataout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT15 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT14 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT13 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT12 ;

wire [35:0] \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2_DATAOUT_bus ;
wire [35:0] \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1_DATAOUT_bus ;

assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2~dataout  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2_DATAOUT_bus [0];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT1  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2_DATAOUT_bus [1];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT2  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2_DATAOUT_bus [2];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT3  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2_DATAOUT_bus [3];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT4  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2_DATAOUT_bus [4];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT5  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2_DATAOUT_bus [5];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT6  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2_DATAOUT_bus [6];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT7  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2_DATAOUT_bus [7];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT8  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2_DATAOUT_bus [8];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT9  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2_DATAOUT_bus [9];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT10  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2_DATAOUT_bus [10];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT11  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2_DATAOUT_bus [11];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT12  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2_DATAOUT_bus [12];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT13  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2_DATAOUT_bus [13];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT14  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2_DATAOUT_bus [14];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT15  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2_DATAOUT_bus [15];

assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1~dataout  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1_DATAOUT_bus [0];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT1  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1_DATAOUT_bus [1];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT2  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1_DATAOUT_bus [2];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT3  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1_DATAOUT_bus [3];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT4  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1_DATAOUT_bus [4];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT5  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1_DATAOUT_bus [5];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT6  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1_DATAOUT_bus [6];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT7  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1_DATAOUT_bus [7];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT8  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1_DATAOUT_bus [8];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT9  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1_DATAOUT_bus [9];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT10  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1_DATAOUT_bus [10];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT11  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1_DATAOUT_bus [11];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT12  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1_DATAOUT_bus [12];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT13  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1_DATAOUT_bus [13];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT14  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1_DATAOUT_bus [14];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT15  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1_DATAOUT_bus [15];

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|dffe3a[11] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT11 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_11),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|dffe3a[11] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|dffe3a[11] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|dffe3a[10] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT10 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_10),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|dffe3a[10] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|dffe3a[10] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|dffe3a[9] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT9 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_9),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|dffe3a[9] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|dffe3a[9] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|dffe3a[8] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT8 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_8),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|dffe3a[8] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|dffe3a[8] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|dffe3a[7] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT7 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_7),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|dffe3a[7] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|dffe3a[7] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|dffe3a[6] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT6 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_6),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|dffe3a[6] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|dffe3a[6] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|dffe3a[5] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT5 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_5),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|dffe3a[5] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|dffe3a[5] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|dffe3a[4] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT4 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_4),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|dffe3a[4] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|dffe3a[4] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|dffe3a[3] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT3 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_3),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|dffe3a[3] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|dffe3a[3] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|dffe3a[2] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT2 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_2),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|dffe3a[2] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|dffe3a[2] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|dffe3a[1] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT1 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_1),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|dffe3a[1] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|dffe3a[1] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|dffe3a[0] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2~dataout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_0),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|dffe3a[0] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|dffe3a[0] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|dffe3a[15] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT15 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_15),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|dffe3a[15] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|dffe3a[15] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|dffe3a[14] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT14 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_14),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|dffe3a[14] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|dffe3a[14] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|dffe3a[13] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT13 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_13),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|dffe3a[13] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|dffe3a[13] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|dffe3a[12] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT12 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_12),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|dffe3a[12] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|dffe3a[12] .power_up = "low";

cycloneiii_mac_mult \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1 (
	.signa(vcc),
	.signb(vcc),
	.clk(clock),
	.aclr(gnd),
	.ena(clken),
	.dataa({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.datab({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.dataout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1_DATAOUT_bus ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1 .dataa_clock = "0";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1 .dataa_width = 8;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1 .datab_clock = "0";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1 .datab_width = 8;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1 .signa_clock = "none";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1 .signb_clock = "none";

cycloneiii_mac_out \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2 (
	.clk(clock),
	.aclr(gnd),
	.ena(clken),
	.dataa({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT15 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT14 ,\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT13 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT12 ,\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT11 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT10 ,\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT9 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT8 ,\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT7 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT6 ,\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT5 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT4 ,\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT3 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT2 ,\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT1 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_mult1~dataout }),
	.dataout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2_DATAOUT_bus ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2 .dataa_width = 16;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm2|gen_dsp_only:m_bd|auto_generated|mac_out2 .output_clock = "0";

endmodule

module fft_asj_fft_cmult_can_fft_120_2 (
	pipeline_dffe_11,
	pipeline_dffe_15,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	pipeline_dffe_9,
	pipeline_dffe_8,
	pipeline_dffe_10,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_81,
	pipeline_dffe_91,
	pipeline_dffe_21,
	pipeline_dffe_31,
	pipeline_dffe_41,
	pipeline_dffe_51,
	pipeline_dffe_61,
	pipeline_dffe_71,
	pipeline_dffe_82,
	pipeline_dffe_92,
	global_clock_enable,
	real_out_3,
	real_out_7,
	real_out_4,
	real_out_5,
	real_out_6,
	real_out_1,
	real_out_0,
	real_out_2,
	twiddle_data200,
	twiddle_data201,
	twiddle_data202,
	twiddle_data203,
	twiddle_data204,
	twiddle_data205,
	twiddle_data206,
	twiddle_data207,
	twiddle_data210,
	twiddle_data211,
	twiddle_data212,
	twiddle_data213,
	twiddle_data214,
	twiddle_data215,
	twiddle_data216,
	twiddle_data217,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_11;
output 	pipeline_dffe_15;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
output 	pipeline_dffe_9;
output 	pipeline_dffe_8;
output 	pipeline_dffe_10;
input 	pipeline_dffe_2;
input 	pipeline_dffe_3;
input 	pipeline_dffe_4;
input 	pipeline_dffe_5;
input 	pipeline_dffe_6;
input 	pipeline_dffe_7;
input 	pipeline_dffe_81;
input 	pipeline_dffe_91;
input 	pipeline_dffe_21;
input 	pipeline_dffe_31;
input 	pipeline_dffe_41;
input 	pipeline_dffe_51;
input 	pipeline_dffe_61;
input 	pipeline_dffe_71;
input 	pipeline_dffe_82;
input 	pipeline_dffe_92;
input 	global_clock_enable;
output 	real_out_3;
output 	real_out_7;
output 	real_out_4;
output 	real_out_5;
output 	real_out_6;
output 	real_out_1;
output 	real_out_0;
output 	real_out_2;
input 	twiddle_data200;
input 	twiddle_data201;
input 	twiddle_data202;
input 	twiddle_data203;
input 	twiddle_data204;
input 	twiddle_data205;
input 	twiddle_data206;
input 	twiddle_data207;
input 	twiddle_data210;
input 	twiddle_data211;
input 	twiddle_data212;
input 	twiddle_data213;
input 	twiddle_data214;
input 	twiddle_data215;
input 	twiddle_data216;
input 	twiddle_data217;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \result_imag_1[11]~q ;
wire \result_imag_1[10]~q ;
wire \result_imag_1[9]~q ;
wire \result_imag_1[8]~q ;
wire \result_imag_1[7]~q ;
wire \result_imag_1[6]~q ;
wire \result_imag_1[5]~q ;
wire \result_imag_1[4]~q ;
wire \result_imag_1[3]~q ;
wire \result_imag_1[2]~q ;
wire \result_imag_1[1]~q ;
wire \result_imag_1[0]~q ;
wire \result_imag_1[15]~q ;
wire \result_imag_1[14]~q ;
wire \result_imag_1[13]~q ;
wire \result_imag_1[12]~q ;
wire \gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ;
wire \gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ;
wire \gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ;
wire \gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ;
wire \gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ;
wire \addresult_ac_bd[11]~q ;
wire \addresult_ac_bd[10]~q ;
wire \addresult_ac_bd[9]~q ;
wire \addresult_ac_bd[8]~q ;
wire \addresult_ac_bd[7]~q ;
wire \addresult_ac_bd[6]~q ;
wire \addresult_ac_bd[5]~q ;
wire \addresult_ac_bd[4]~q ;
wire \addresult_ac_bd[3]~q ;
wire \addresult_ac_bd[2]~q ;
wire \addresult_ac_bd[1]~q ;
wire \addresult_ac_bd[0]~q ;
wire \result_imag_1[0]~17 ;
wire \result_imag_1[0]~16_combout ;
wire \result_imag_1[1]~19 ;
wire \result_imag_1[1]~18_combout ;
wire \result_imag_1[2]~21 ;
wire \result_imag_1[2]~20_combout ;
wire \result_imag_1[3]~23 ;
wire \result_imag_1[3]~22_combout ;
wire \result_imag_1[4]~25 ;
wire \result_imag_1[4]~24_combout ;
wire \result_imag_1[5]~27 ;
wire \result_imag_1[5]~26_combout ;
wire \result_imag_1[6]~29 ;
wire \result_imag_1[6]~28_combout ;
wire \result_imag_1[7]~31 ;
wire \result_imag_1[7]~30_combout ;
wire \result_imag_1[8]~33 ;
wire \result_imag_1[8]~32_combout ;
wire \result_imag_1[9]~35 ;
wire \result_imag_1[9]~34_combout ;
wire \result_imag_1[10]~37 ;
wire \result_imag_1[10]~36_combout ;
wire \result_imag_1[11]~39 ;
wire \result_imag_1[11]~38_combout ;
wire \addresult_ac_bd[15]~q ;
wire \addresult_ac_bd[14]~q ;
wire \addresult_ac_bd[13]~q ;
wire \addresult_ac_bd[12]~q ;
wire \result_imag_1[12]~41 ;
wire \result_imag_1[12]~40_combout ;
wire \result_imag_1[13]~43 ;
wire \result_imag_1[13]~42_combout ;
wire \result_imag_1[14]~45 ;
wire \result_imag_1[14]~44_combout ;
wire \result_imag_1[15]~46_combout ;
wire \result_real_1_tmp[11]~q ;
wire \result_real_1_tmp[10]~q ;
wire \result_real_1_tmp[9]~q ;
wire \result_real_1_tmp[8]~q ;
wire \result_real_1_tmp[7]~q ;
wire \result_real_1_tmp[6]~q ;
wire \result_real_1_tmp[5]~q ;
wire \result_real_1_tmp[4]~q ;
wire \result_real_1_tmp[3]~q ;
wire \result_real_1_tmp[2]~q ;
wire \result_real_1_tmp[1]~q ;
wire \result_real_1_tmp[0]~q ;
wire \result_real_1_tmp[15]~q ;
wire \result_real_1_tmp[14]~q ;
wire \result_real_1_tmp[13]~q ;
wire \result_real_1_tmp[12]~q ;
wire \addresult_ac_bd[0]~17 ;
wire \addresult_ac_bd[0]~16_combout ;
wire \addresult_ac_bd[1]~19 ;
wire \addresult_ac_bd[1]~18_combout ;
wire \addresult_ac_bd[2]~21 ;
wire \addresult_ac_bd[2]~20_combout ;
wire \addresult_ac_bd[3]~23 ;
wire \addresult_ac_bd[3]~22_combout ;
wire \addresult_ac_bd[4]~25 ;
wire \addresult_ac_bd[4]~24_combout ;
wire \addresult_ac_bd[5]~27 ;
wire \addresult_ac_bd[5]~26_combout ;
wire \addresult_ac_bd[6]~29 ;
wire \addresult_ac_bd[6]~28_combout ;
wire \addresult_ac_bd[7]~31 ;
wire \addresult_ac_bd[7]~30_combout ;
wire \addresult_ac_bd[8]~33 ;
wire \addresult_ac_bd[8]~32_combout ;
wire \addresult_ac_bd[9]~35 ;
wire \addresult_ac_bd[9]~34_combout ;
wire \addresult_ac_bd[10]~37 ;
wire \addresult_ac_bd[10]~36_combout ;
wire \addresult_ac_bd[11]~39 ;
wire \addresult_ac_bd[11]~38_combout ;
wire \addresult_ac_bd[12]~41 ;
wire \addresult_ac_bd[12]~40_combout ;
wire \addresult_ac_bd[13]~43 ;
wire \addresult_ac_bd[13]~42_combout ;
wire \addresult_ac_bd[14]~45 ;
wire \addresult_ac_bd[14]~44_combout ;
wire \addresult_ac_bd[15]~46_combout ;
wire \result_real_1_tmp[0]~17 ;
wire \result_real_1_tmp[0]~16_combout ;
wire \result_real_1_tmp[1]~19 ;
wire \result_real_1_tmp[1]~18_combout ;
wire \result_real_1_tmp[2]~21 ;
wire \result_real_1_tmp[2]~20_combout ;
wire \result_real_1_tmp[3]~23 ;
wire \result_real_1_tmp[3]~22_combout ;
wire \result_real_1_tmp[4]~25 ;
wire \result_real_1_tmp[4]~24_combout ;
wire \result_real_1_tmp[5]~27 ;
wire \result_real_1_tmp[5]~26_combout ;
wire \result_real_1_tmp[6]~29 ;
wire \result_real_1_tmp[6]~28_combout ;
wire \result_real_1_tmp[7]~31 ;
wire \result_real_1_tmp[7]~30_combout ;
wire \result_real_1_tmp[8]~33 ;
wire \result_real_1_tmp[8]~32_combout ;
wire \result_real_1_tmp[9]~35 ;
wire \result_real_1_tmp[9]~34_combout ;
wire \result_real_1_tmp[10]~37 ;
wire \result_real_1_tmp[10]~36_combout ;
wire \result_real_1_tmp[11]~39 ;
wire \result_real_1_tmp[11]~38_combout ;
wire \result_real_1_tmp[12]~41 ;
wire \result_real_1_tmp[12]~40_combout ;
wire \result_real_1_tmp[13]~43 ;
wire \result_real_1_tmp[13]~42_combout ;
wire \result_real_1_tmp[14]~45 ;
wire \result_real_1_tmp[14]~44_combout ;
wire \result_real_1_tmp[15]~46_combout ;
wire \addresult_a_b[0]~q ;
wire \addresult_a_b[1]~q ;
wire \addresult_a_b[2]~q ;
wire \addresult_a_b[3]~q ;
wire \addresult_a_b[4]~q ;
wire \addresult_a_b[5]~q ;
wire \addresult_a_b[6]~q ;
wire \addresult_a_b[7]~q ;
wire \addresult_a_b[8]~q ;
wire \addresult_c_d[0]~q ;
wire \addresult_c_d[1]~q ;
wire \addresult_c_d[2]~q ;
wire \addresult_c_d[3]~q ;
wire \addresult_c_d[4]~q ;
wire \addresult_c_d[5]~q ;
wire \addresult_c_d[6]~q ;
wire \addresult_c_d[7]~q ;
wire \addresult_c_d[8]~q ;
wire \addresult_a_b[0]~10 ;
wire \addresult_a_b[0]~9_combout ;
wire \addresult_a_b[1]~12 ;
wire \addresult_a_b[1]~11_combout ;
wire \addresult_a_b[2]~14 ;
wire \addresult_a_b[2]~13_combout ;
wire \addresult_a_b[3]~16 ;
wire \addresult_a_b[3]~15_combout ;
wire \addresult_a_b[4]~18 ;
wire \addresult_a_b[4]~17_combout ;
wire \addresult_a_b[5]~20 ;
wire \addresult_a_b[5]~19_combout ;
wire \addresult_a_b[6]~22 ;
wire \addresult_a_b[6]~21_combout ;
wire \addresult_a_b[7]~24 ;
wire \addresult_a_b[7]~23_combout ;
wire \addresult_a_b[8]~25_combout ;
wire \addresult_c_d[0]~10 ;
wire \addresult_c_d[0]~9_combout ;
wire \addresult_c_d[1]~12 ;
wire \addresult_c_d[1]~11_combout ;
wire \addresult_c_d[2]~14 ;
wire \addresult_c_d[2]~13_combout ;
wire \addresult_c_d[3]~16 ;
wire \addresult_c_d[3]~15_combout ;
wire \addresult_c_d[4]~18 ;
wire \addresult_c_d[4]~17_combout ;
wire \addresult_c_d[5]~20 ;
wire \addresult_c_d[5]~19_combout ;
wire \addresult_c_d[6]~22 ;
wire \addresult_c_d[6]~21_combout ;
wire \addresult_c_d[7]~24 ;
wire \addresult_c_d[7]~23_combout ;
wire \addresult_c_d[8]~25_combout ;
wire \gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ;
wire \gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ;
wire \gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ;
wire \result_a_b_c_d_se[11]~q ;
wire \result_a_b_c_d_se[10]~q ;
wire \result_a_b_c_d_se[9]~q ;
wire \result_a_b_c_d_se[8]~q ;
wire \result_a_b_c_d_se[7]~q ;
wire \result_a_b_c_d_se[6]~q ;
wire \result_a_b_c_d_se[5]~q ;
wire \result_a_b_c_d_se[4]~q ;
wire \result_a_b_c_d_se[3]~q ;
wire \result_a_b_c_d_se[2]~q ;
wire \result_a_b_c_d_se[1]~q ;
wire \result_a_b_c_d_se[0]~q ;
wire \result_a_b_c_d_se[15]~q ;
wire \result_a_b_c_d_se[14]~q ;
wire \result_a_b_c_d_se[13]~q ;
wire \result_a_b_c_d_se[12]~q ;
wire \result_a_c_se[11]~q ;
wire \result_b_d_se[11]~q ;
wire \result_a_c_se[10]~q ;
wire \result_b_d_se[10]~q ;
wire \result_a_c_se[9]~q ;
wire \result_b_d_se[9]~q ;
wire \result_a_c_se[8]~q ;
wire \result_b_d_se[8]~q ;
wire \result_a_c_se[7]~q ;
wire \result_b_d_se[7]~q ;
wire \result_a_c_se[6]~q ;
wire \result_b_d_se[6]~q ;
wire \result_a_c_se[5]~q ;
wire \result_b_d_se[5]~q ;
wire \result_a_c_se[4]~q ;
wire \result_b_d_se[4]~q ;
wire \result_a_c_se[3]~q ;
wire \result_b_d_se[3]~q ;
wire \result_a_c_se[2]~q ;
wire \result_b_d_se[2]~q ;
wire \result_a_c_se[1]~q ;
wire \result_b_d_se[1]~q ;
wire \result_a_c_se[0]~q ;
wire \result_b_d_se[0]~q ;
wire \gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[11]~q ;
wire \gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[10]~q ;
wire \gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[9]~q ;
wire \gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[8]~q ;
wire \gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[7]~q ;
wire \gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[6]~q ;
wire \gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[5]~q ;
wire \gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[4]~q ;
wire \gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[3]~q ;
wire \gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[2]~q ;
wire \gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[1]~q ;
wire \gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[0]~q ;
wire \result_a_c_se[15]~q ;
wire \result_b_d_se[15]~q ;
wire \result_a_c_se[14]~q ;
wire \result_b_d_se[14]~q ;
wire \result_a_c_se[13]~q ;
wire \result_b_d_se[13]~q ;
wire \result_a_c_se[12]~q ;
wire \result_b_d_se[12]~q ;
wire \gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[15]~q ;
wire \gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[14]~q ;
wire \gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[13]~q ;
wire \gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[12]~q ;
wire \gen_dsp_only:m_ac|auto_generated|dffe3a[11]~q ;
wire \gen_dsp_only:m_bd|auto_generated|dffe3a[11]~q ;
wire \gen_dsp_only:m_ac|auto_generated|dffe3a[10]~q ;
wire \gen_dsp_only:m_bd|auto_generated|dffe3a[10]~q ;
wire \gen_dsp_only:m_ac|auto_generated|dffe3a[9]~q ;
wire \gen_dsp_only:m_bd|auto_generated|dffe3a[9]~q ;
wire \gen_dsp_only:m_ac|auto_generated|dffe3a[8]~q ;
wire \gen_dsp_only:m_bd|auto_generated|dffe3a[8]~q ;
wire \gen_dsp_only:m_ac|auto_generated|dffe3a[7]~q ;
wire \gen_dsp_only:m_bd|auto_generated|dffe3a[7]~q ;
wire \gen_dsp_only:m_ac|auto_generated|dffe3a[6]~q ;
wire \gen_dsp_only:m_bd|auto_generated|dffe3a[6]~q ;
wire \gen_dsp_only:m_ac|auto_generated|dffe3a[5]~q ;
wire \gen_dsp_only:m_bd|auto_generated|dffe3a[5]~q ;
wire \gen_dsp_only:m_ac|auto_generated|dffe3a[4]~q ;
wire \gen_dsp_only:m_bd|auto_generated|dffe3a[4]~q ;
wire \gen_dsp_only:m_ac|auto_generated|dffe3a[3]~q ;
wire \gen_dsp_only:m_bd|auto_generated|dffe3a[3]~q ;
wire \gen_dsp_only:m_ac|auto_generated|dffe3a[2]~q ;
wire \gen_dsp_only:m_bd|auto_generated|dffe3a[2]~q ;
wire \gen_dsp_only:m_ac|auto_generated|dffe3a[1]~q ;
wire \gen_dsp_only:m_bd|auto_generated|dffe3a[1]~q ;
wire \gen_dsp_only:m_ac|auto_generated|dffe3a[0]~q ;
wire \gen_dsp_only:m_bd|auto_generated|dffe3a[0]~q ;
wire \gen_dsp_only:m_ac|auto_generated|dffe3a[15]~q ;
wire \gen_dsp_only:m_bd|auto_generated|dffe3a[15]~q ;
wire \gen_dsp_only:m_ac|auto_generated|dffe3a[14]~q ;
wire \gen_dsp_only:m_bd|auto_generated|dffe3a[14]~q ;
wire \gen_dsp_only:m_ac|auto_generated|dffe3a[13]~q ;
wire \gen_dsp_only:m_bd|auto_generated|dffe3a[13]~q ;
wire \gen_dsp_only:m_ac|auto_generated|dffe3a[12]~q ;
wire \gen_dsp_only:m_bd|auto_generated|dffe3a[12]~q ;


fft_asj_fft_pround_fft_120_5 \gen_unsc:u1 (
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_14(pipeline_dffe_14),
	.result_imag_1_11(\result_imag_1[11]~q ),
	.result_imag_1_10(\result_imag_1[10]~q ),
	.result_imag_1_9(\result_imag_1[9]~q ),
	.result_imag_1_8(\result_imag_1[8]~q ),
	.result_imag_1_7(\result_imag_1[7]~q ),
	.result_imag_1_6(\result_imag_1[6]~q ),
	.result_imag_1_5(\result_imag_1[5]~q ),
	.result_imag_1_4(\result_imag_1[4]~q ),
	.result_imag_1_3(\result_imag_1[3]~q ),
	.result_imag_1_2(\result_imag_1[2]~q ),
	.result_imag_1_1(\result_imag_1[1]~q ),
	.result_imag_1_0(\result_imag_1[0]~q ),
	.result_imag_1_15(\result_imag_1[15]~q ),
	.result_imag_1_14(\result_imag_1[14]~q ),
	.result_imag_1_13(\result_imag_1[13]~q ),
	.result_imag_1_12(\result_imag_1[12]~q ),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_10(pipeline_dffe_10),
	.global_clock_enable(global_clock_enable),
	.clk(clk));

fft_asj_fft_pround_fft_120_4 \gen_unsc:u0 (
	.pipeline_dffe_11(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_15(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_12(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_13(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ),
	.pipeline_dffe_14(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ),
	.result_real_1_tmp_11(\result_real_1_tmp[11]~q ),
	.result_real_1_tmp_10(\result_real_1_tmp[10]~q ),
	.result_real_1_tmp_9(\result_real_1_tmp[9]~q ),
	.result_real_1_tmp_8(\result_real_1_tmp[8]~q ),
	.result_real_1_tmp_7(\result_real_1_tmp[7]~q ),
	.result_real_1_tmp_6(\result_real_1_tmp[6]~q ),
	.result_real_1_tmp_5(\result_real_1_tmp[5]~q ),
	.result_real_1_tmp_4(\result_real_1_tmp[4]~q ),
	.result_real_1_tmp_3(\result_real_1_tmp[3]~q ),
	.result_real_1_tmp_2(\result_real_1_tmp[2]~q ),
	.result_real_1_tmp_1(\result_real_1_tmp[1]~q ),
	.result_real_1_tmp_0(\result_real_1_tmp[0]~q ),
	.result_real_1_tmp_15(\result_real_1_tmp[15]~q ),
	.result_real_1_tmp_14(\result_real_1_tmp[14]~q ),
	.result_real_1_tmp_13(\result_real_1_tmp[13]~q ),
	.result_real_1_tmp_12(\result_real_1_tmp[12]~q ),
	.pipeline_dffe_9(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_8(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_10(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ),
	.global_clock_enable(global_clock_enable),
	.clk(clk));

fft_LPM_MULT_7 \gen_dsp_only:m_a_b_c_d (
	.dataa({\addresult_a_b[8]~q ,\addresult_a_b[7]~q ,\addresult_a_b[6]~q ,\addresult_a_b[5]~q ,\addresult_a_b[4]~q ,\addresult_a_b[3]~q ,\addresult_a_b[2]~q ,\addresult_a_b[1]~q ,\addresult_a_b[0]~q }),
	.datab({\addresult_c_d[8]~q ,\addresult_c_d[7]~q ,\addresult_c_d[6]~q ,\addresult_c_d[5]~q ,\addresult_c_d[4]~q ,\addresult_c_d[3]~q ,\addresult_c_d[2]~q ,\addresult_c_d[1]~q ,\addresult_c_d[0]~q }),
	.clken(global_clock_enable),
	.dffe3a_11(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[11]~q ),
	.dffe3a_10(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[10]~q ),
	.dffe3a_9(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[9]~q ),
	.dffe3a_8(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[8]~q ),
	.dffe3a_7(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[7]~q ),
	.dffe3a_6(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[6]~q ),
	.dffe3a_5(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[5]~q ),
	.dffe3a_4(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[4]~q ),
	.dffe3a_3(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[3]~q ),
	.dffe3a_2(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[2]~q ),
	.dffe3a_1(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[1]~q ),
	.dffe3a_0(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[0]~q ),
	.dffe3a_15(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[15]~q ),
	.dffe3a_14(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[14]~q ),
	.dffe3a_13(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[13]~q ),
	.dffe3a_12(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[12]~q ),
	.clock(clk));

fft_LPM_MULT_9 \gen_dsp_only:m_bd (
	.dataa({gnd,pipeline_dffe_92,pipeline_dffe_82,pipeline_dffe_71,pipeline_dffe_61,pipeline_dffe_51,pipeline_dffe_41,pipeline_dffe_31,pipeline_dffe_21}),
	.clken(global_clock_enable),
	.dffe3a_11(\gen_dsp_only:m_bd|auto_generated|dffe3a[11]~q ),
	.dffe3a_10(\gen_dsp_only:m_bd|auto_generated|dffe3a[10]~q ),
	.dffe3a_9(\gen_dsp_only:m_bd|auto_generated|dffe3a[9]~q ),
	.dffe3a_8(\gen_dsp_only:m_bd|auto_generated|dffe3a[8]~q ),
	.dffe3a_7(\gen_dsp_only:m_bd|auto_generated|dffe3a[7]~q ),
	.dffe3a_6(\gen_dsp_only:m_bd|auto_generated|dffe3a[6]~q ),
	.dffe3a_5(\gen_dsp_only:m_bd|auto_generated|dffe3a[5]~q ),
	.dffe3a_4(\gen_dsp_only:m_bd|auto_generated|dffe3a[4]~q ),
	.dffe3a_3(\gen_dsp_only:m_bd|auto_generated|dffe3a[3]~q ),
	.dffe3a_2(\gen_dsp_only:m_bd|auto_generated|dffe3a[2]~q ),
	.dffe3a_1(\gen_dsp_only:m_bd|auto_generated|dffe3a[1]~q ),
	.dffe3a_0(\gen_dsp_only:m_bd|auto_generated|dffe3a[0]~q ),
	.dffe3a_15(\gen_dsp_only:m_bd|auto_generated|dffe3a[15]~q ),
	.dffe3a_14(\gen_dsp_only:m_bd|auto_generated|dffe3a[14]~q ),
	.dffe3a_13(\gen_dsp_only:m_bd|auto_generated|dffe3a[13]~q ),
	.dffe3a_12(\gen_dsp_only:m_bd|auto_generated|dffe3a[12]~q ),
	.datab({gnd,twiddle_data217,twiddle_data216,twiddle_data215,twiddle_data214,twiddle_data213,twiddle_data212,twiddle_data211,twiddle_data210}),
	.clock(clk));

fft_LPM_MULT_8 \gen_dsp_only:m_ac (
	.dataa({gnd,pipeline_dffe_91,pipeline_dffe_81,pipeline_dffe_7,pipeline_dffe_6,pipeline_dffe_5,pipeline_dffe_4,pipeline_dffe_3,pipeline_dffe_2}),
	.clken(global_clock_enable),
	.dffe3a_11(\gen_dsp_only:m_ac|auto_generated|dffe3a[11]~q ),
	.dffe3a_10(\gen_dsp_only:m_ac|auto_generated|dffe3a[10]~q ),
	.dffe3a_9(\gen_dsp_only:m_ac|auto_generated|dffe3a[9]~q ),
	.dffe3a_8(\gen_dsp_only:m_ac|auto_generated|dffe3a[8]~q ),
	.dffe3a_7(\gen_dsp_only:m_ac|auto_generated|dffe3a[7]~q ),
	.dffe3a_6(\gen_dsp_only:m_ac|auto_generated|dffe3a[6]~q ),
	.dffe3a_5(\gen_dsp_only:m_ac|auto_generated|dffe3a[5]~q ),
	.dffe3a_4(\gen_dsp_only:m_ac|auto_generated|dffe3a[4]~q ),
	.dffe3a_3(\gen_dsp_only:m_ac|auto_generated|dffe3a[3]~q ),
	.dffe3a_2(\gen_dsp_only:m_ac|auto_generated|dffe3a[2]~q ),
	.dffe3a_1(\gen_dsp_only:m_ac|auto_generated|dffe3a[1]~q ),
	.dffe3a_0(\gen_dsp_only:m_ac|auto_generated|dffe3a[0]~q ),
	.dffe3a_15(\gen_dsp_only:m_ac|auto_generated|dffe3a[15]~q ),
	.dffe3a_14(\gen_dsp_only:m_ac|auto_generated|dffe3a[14]~q ),
	.dffe3a_13(\gen_dsp_only:m_ac|auto_generated|dffe3a[13]~q ),
	.dffe3a_12(\gen_dsp_only:m_ac|auto_generated|dffe3a[12]~q ),
	.datab({gnd,twiddle_data207,twiddle_data206,twiddle_data205,twiddle_data204,twiddle_data203,twiddle_data202,twiddle_data201,twiddle_data200}),
	.clock(clk));

dffeas \result_imag_1[11] (
	.clk(clk),
	.d(\result_imag_1[11]~38_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[11]~q ),
	.prn(vcc));
defparam \result_imag_1[11] .is_wysiwyg = "true";
defparam \result_imag_1[11] .power_up = "low";

dffeas \result_imag_1[10] (
	.clk(clk),
	.d(\result_imag_1[10]~36_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[10]~q ),
	.prn(vcc));
defparam \result_imag_1[10] .is_wysiwyg = "true";
defparam \result_imag_1[10] .power_up = "low";

dffeas \result_imag_1[9] (
	.clk(clk),
	.d(\result_imag_1[9]~34_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[9]~q ),
	.prn(vcc));
defparam \result_imag_1[9] .is_wysiwyg = "true";
defparam \result_imag_1[9] .power_up = "low";

dffeas \result_imag_1[8] (
	.clk(clk),
	.d(\result_imag_1[8]~32_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[8]~q ),
	.prn(vcc));
defparam \result_imag_1[8] .is_wysiwyg = "true";
defparam \result_imag_1[8] .power_up = "low";

dffeas \result_imag_1[7] (
	.clk(clk),
	.d(\result_imag_1[7]~30_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[7]~q ),
	.prn(vcc));
defparam \result_imag_1[7] .is_wysiwyg = "true";
defparam \result_imag_1[7] .power_up = "low";

dffeas \result_imag_1[6] (
	.clk(clk),
	.d(\result_imag_1[6]~28_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[6]~q ),
	.prn(vcc));
defparam \result_imag_1[6] .is_wysiwyg = "true";
defparam \result_imag_1[6] .power_up = "low";

dffeas \result_imag_1[5] (
	.clk(clk),
	.d(\result_imag_1[5]~26_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[5]~q ),
	.prn(vcc));
defparam \result_imag_1[5] .is_wysiwyg = "true";
defparam \result_imag_1[5] .power_up = "low";

dffeas \result_imag_1[4] (
	.clk(clk),
	.d(\result_imag_1[4]~24_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[4]~q ),
	.prn(vcc));
defparam \result_imag_1[4] .is_wysiwyg = "true";
defparam \result_imag_1[4] .power_up = "low";

dffeas \result_imag_1[3] (
	.clk(clk),
	.d(\result_imag_1[3]~22_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[3]~q ),
	.prn(vcc));
defparam \result_imag_1[3] .is_wysiwyg = "true";
defparam \result_imag_1[3] .power_up = "low";

dffeas \result_imag_1[2] (
	.clk(clk),
	.d(\result_imag_1[2]~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[2]~q ),
	.prn(vcc));
defparam \result_imag_1[2] .is_wysiwyg = "true";
defparam \result_imag_1[2] .power_up = "low";

dffeas \result_imag_1[1] (
	.clk(clk),
	.d(\result_imag_1[1]~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[1]~q ),
	.prn(vcc));
defparam \result_imag_1[1] .is_wysiwyg = "true";
defparam \result_imag_1[1] .power_up = "low";

dffeas \result_imag_1[0] (
	.clk(clk),
	.d(\result_imag_1[0]~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[0]~q ),
	.prn(vcc));
defparam \result_imag_1[0] .is_wysiwyg = "true";
defparam \result_imag_1[0] .power_up = "low";

dffeas \result_imag_1[15] (
	.clk(clk),
	.d(\result_imag_1[15]~46_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[15]~q ),
	.prn(vcc));
defparam \result_imag_1[15] .is_wysiwyg = "true";
defparam \result_imag_1[15] .power_up = "low";

dffeas \result_imag_1[14] (
	.clk(clk),
	.d(\result_imag_1[14]~44_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[14]~q ),
	.prn(vcc));
defparam \result_imag_1[14] .is_wysiwyg = "true";
defparam \result_imag_1[14] .power_up = "low";

dffeas \result_imag_1[13] (
	.clk(clk),
	.d(\result_imag_1[13]~42_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[13]~q ),
	.prn(vcc));
defparam \result_imag_1[13] .is_wysiwyg = "true";
defparam \result_imag_1[13] .power_up = "low";

dffeas \result_imag_1[12] (
	.clk(clk),
	.d(\result_imag_1[12]~40_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[12]~q ),
	.prn(vcc));
defparam \result_imag_1[12] .is_wysiwyg = "true";
defparam \result_imag_1[12] .power_up = "low";

dffeas \addresult_ac_bd[11] (
	.clk(clk),
	.d(\addresult_ac_bd[11]~38_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[11]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[11] .is_wysiwyg = "true";
defparam \addresult_ac_bd[11] .power_up = "low";

dffeas \addresult_ac_bd[10] (
	.clk(clk),
	.d(\addresult_ac_bd[10]~36_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[10]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[10] .is_wysiwyg = "true";
defparam \addresult_ac_bd[10] .power_up = "low";

dffeas \addresult_ac_bd[9] (
	.clk(clk),
	.d(\addresult_ac_bd[9]~34_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[9]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[9] .is_wysiwyg = "true";
defparam \addresult_ac_bd[9] .power_up = "low";

dffeas \addresult_ac_bd[8] (
	.clk(clk),
	.d(\addresult_ac_bd[8]~32_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[8]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[8] .is_wysiwyg = "true";
defparam \addresult_ac_bd[8] .power_up = "low";

dffeas \addresult_ac_bd[7] (
	.clk(clk),
	.d(\addresult_ac_bd[7]~30_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[7]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[7] .is_wysiwyg = "true";
defparam \addresult_ac_bd[7] .power_up = "low";

dffeas \addresult_ac_bd[6] (
	.clk(clk),
	.d(\addresult_ac_bd[6]~28_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[6]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[6] .is_wysiwyg = "true";
defparam \addresult_ac_bd[6] .power_up = "low";

dffeas \addresult_ac_bd[5] (
	.clk(clk),
	.d(\addresult_ac_bd[5]~26_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[5]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[5] .is_wysiwyg = "true";
defparam \addresult_ac_bd[5] .power_up = "low";

dffeas \addresult_ac_bd[4] (
	.clk(clk),
	.d(\addresult_ac_bd[4]~24_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[4]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[4] .is_wysiwyg = "true";
defparam \addresult_ac_bd[4] .power_up = "low";

dffeas \addresult_ac_bd[3] (
	.clk(clk),
	.d(\addresult_ac_bd[3]~22_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[3]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[3] .is_wysiwyg = "true";
defparam \addresult_ac_bd[3] .power_up = "low";

dffeas \addresult_ac_bd[2] (
	.clk(clk),
	.d(\addresult_ac_bd[2]~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[2]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[2] .is_wysiwyg = "true";
defparam \addresult_ac_bd[2] .power_up = "low";

dffeas \addresult_ac_bd[1] (
	.clk(clk),
	.d(\addresult_ac_bd[1]~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[1]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[1] .is_wysiwyg = "true";
defparam \addresult_ac_bd[1] .power_up = "low";

dffeas \addresult_ac_bd[0] (
	.clk(clk),
	.d(\addresult_ac_bd[0]~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[0]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[0] .is_wysiwyg = "true";
defparam \addresult_ac_bd[0] .power_up = "low";

cycloneiii_lcell_comb \result_imag_1[0]~16 (
	.dataa(\addresult_ac_bd[0]~q ),
	.datab(\result_a_b_c_d_se[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\result_imag_1[0]~16_combout ),
	.cout(\result_imag_1[0]~17 ));
defparam \result_imag_1[0]~16 .lut_mask = 16'h66DD;
defparam \result_imag_1[0]~16 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \result_imag_1[1]~18 (
	.dataa(\addresult_ac_bd[1]~q ),
	.datab(\result_a_b_c_d_se[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[0]~17 ),
	.combout(\result_imag_1[1]~18_combout ),
	.cout(\result_imag_1[1]~19 ));
defparam \result_imag_1[1]~18 .lut_mask = 16'h96BF;
defparam \result_imag_1[1]~18 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_imag_1[2]~20 (
	.dataa(\addresult_ac_bd[2]~q ),
	.datab(\result_a_b_c_d_se[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[1]~19 ),
	.combout(\result_imag_1[2]~20_combout ),
	.cout(\result_imag_1[2]~21 ));
defparam \result_imag_1[2]~20 .lut_mask = 16'h96DF;
defparam \result_imag_1[2]~20 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_imag_1[3]~22 (
	.dataa(\addresult_ac_bd[3]~q ),
	.datab(\result_a_b_c_d_se[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[2]~21 ),
	.combout(\result_imag_1[3]~22_combout ),
	.cout(\result_imag_1[3]~23 ));
defparam \result_imag_1[3]~22 .lut_mask = 16'h96BF;
defparam \result_imag_1[3]~22 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_imag_1[4]~24 (
	.dataa(\addresult_ac_bd[4]~q ),
	.datab(\result_a_b_c_d_se[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[3]~23 ),
	.combout(\result_imag_1[4]~24_combout ),
	.cout(\result_imag_1[4]~25 ));
defparam \result_imag_1[4]~24 .lut_mask = 16'h96DF;
defparam \result_imag_1[4]~24 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_imag_1[5]~26 (
	.dataa(\addresult_ac_bd[5]~q ),
	.datab(\result_a_b_c_d_se[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[4]~25 ),
	.combout(\result_imag_1[5]~26_combout ),
	.cout(\result_imag_1[5]~27 ));
defparam \result_imag_1[5]~26 .lut_mask = 16'h96BF;
defparam \result_imag_1[5]~26 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_imag_1[6]~28 (
	.dataa(\addresult_ac_bd[6]~q ),
	.datab(\result_a_b_c_d_se[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[5]~27 ),
	.combout(\result_imag_1[6]~28_combout ),
	.cout(\result_imag_1[6]~29 ));
defparam \result_imag_1[6]~28 .lut_mask = 16'h96DF;
defparam \result_imag_1[6]~28 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_imag_1[7]~30 (
	.dataa(\addresult_ac_bd[7]~q ),
	.datab(\result_a_b_c_d_se[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[6]~29 ),
	.combout(\result_imag_1[7]~30_combout ),
	.cout(\result_imag_1[7]~31 ));
defparam \result_imag_1[7]~30 .lut_mask = 16'h96BF;
defparam \result_imag_1[7]~30 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_imag_1[8]~32 (
	.dataa(\addresult_ac_bd[8]~q ),
	.datab(\result_a_b_c_d_se[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[7]~31 ),
	.combout(\result_imag_1[8]~32_combout ),
	.cout(\result_imag_1[8]~33 ));
defparam \result_imag_1[8]~32 .lut_mask = 16'h96DF;
defparam \result_imag_1[8]~32 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_imag_1[9]~34 (
	.dataa(\addresult_ac_bd[9]~q ),
	.datab(\result_a_b_c_d_se[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[8]~33 ),
	.combout(\result_imag_1[9]~34_combout ),
	.cout(\result_imag_1[9]~35 ));
defparam \result_imag_1[9]~34 .lut_mask = 16'h96BF;
defparam \result_imag_1[9]~34 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_imag_1[10]~36 (
	.dataa(\addresult_ac_bd[10]~q ),
	.datab(\result_a_b_c_d_se[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[9]~35 ),
	.combout(\result_imag_1[10]~36_combout ),
	.cout(\result_imag_1[10]~37 ));
defparam \result_imag_1[10]~36 .lut_mask = 16'h96DF;
defparam \result_imag_1[10]~36 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_imag_1[11]~38 (
	.dataa(\addresult_ac_bd[11]~q ),
	.datab(\result_a_b_c_d_se[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[10]~37 ),
	.combout(\result_imag_1[11]~38_combout ),
	.cout(\result_imag_1[11]~39 ));
defparam \result_imag_1[11]~38 .lut_mask = 16'h96BF;
defparam \result_imag_1[11]~38 .sum_lutc_input = "cin";

dffeas \addresult_ac_bd[15] (
	.clk(clk),
	.d(\addresult_ac_bd[15]~46_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[15]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[15] .is_wysiwyg = "true";
defparam \addresult_ac_bd[15] .power_up = "low";

dffeas \addresult_ac_bd[14] (
	.clk(clk),
	.d(\addresult_ac_bd[14]~44_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[14]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[14] .is_wysiwyg = "true";
defparam \addresult_ac_bd[14] .power_up = "low";

dffeas \addresult_ac_bd[13] (
	.clk(clk),
	.d(\addresult_ac_bd[13]~42_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[13]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[13] .is_wysiwyg = "true";
defparam \addresult_ac_bd[13] .power_up = "low";

dffeas \addresult_ac_bd[12] (
	.clk(clk),
	.d(\addresult_ac_bd[12]~40_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[12]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[12] .is_wysiwyg = "true";
defparam \addresult_ac_bd[12] .power_up = "low";

cycloneiii_lcell_comb \result_imag_1[12]~40 (
	.dataa(\addresult_ac_bd[12]~q ),
	.datab(\result_a_b_c_d_se[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[11]~39 ),
	.combout(\result_imag_1[12]~40_combout ),
	.cout(\result_imag_1[12]~41 ));
defparam \result_imag_1[12]~40 .lut_mask = 16'h96DF;
defparam \result_imag_1[12]~40 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_imag_1[13]~42 (
	.dataa(\addresult_ac_bd[13]~q ),
	.datab(\result_a_b_c_d_se[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[12]~41 ),
	.combout(\result_imag_1[13]~42_combout ),
	.cout(\result_imag_1[13]~43 ));
defparam \result_imag_1[13]~42 .lut_mask = 16'h96BF;
defparam \result_imag_1[13]~42 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_imag_1[14]~44 (
	.dataa(\addresult_ac_bd[14]~q ),
	.datab(\result_a_b_c_d_se[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[13]~43 ),
	.combout(\result_imag_1[14]~44_combout ),
	.cout(\result_imag_1[14]~45 ));
defparam \result_imag_1[14]~44 .lut_mask = 16'h96DF;
defparam \result_imag_1[14]~44 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_imag_1[15]~46 (
	.dataa(\addresult_ac_bd[15]~q ),
	.datab(\result_a_b_c_d_se[15]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\result_imag_1[14]~45 ),
	.combout(\result_imag_1[15]~46_combout ),
	.cout());
defparam \result_imag_1[15]~46 .lut_mask = 16'h9696;
defparam \result_imag_1[15]~46 .sum_lutc_input = "cin";

dffeas \result_real_1_tmp[11] (
	.clk(clk),
	.d(\result_real_1_tmp[11]~38_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[11]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[11] .is_wysiwyg = "true";
defparam \result_real_1_tmp[11] .power_up = "low";

dffeas \result_real_1_tmp[10] (
	.clk(clk),
	.d(\result_real_1_tmp[10]~36_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[10]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[10] .is_wysiwyg = "true";
defparam \result_real_1_tmp[10] .power_up = "low";

dffeas \result_real_1_tmp[9] (
	.clk(clk),
	.d(\result_real_1_tmp[9]~34_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[9]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[9] .is_wysiwyg = "true";
defparam \result_real_1_tmp[9] .power_up = "low";

dffeas \result_real_1_tmp[8] (
	.clk(clk),
	.d(\result_real_1_tmp[8]~32_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[8]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[8] .is_wysiwyg = "true";
defparam \result_real_1_tmp[8] .power_up = "low";

dffeas \result_real_1_tmp[7] (
	.clk(clk),
	.d(\result_real_1_tmp[7]~30_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[7]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[7] .is_wysiwyg = "true";
defparam \result_real_1_tmp[7] .power_up = "low";

dffeas \result_real_1_tmp[6] (
	.clk(clk),
	.d(\result_real_1_tmp[6]~28_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[6]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[6] .is_wysiwyg = "true";
defparam \result_real_1_tmp[6] .power_up = "low";

dffeas \result_real_1_tmp[5] (
	.clk(clk),
	.d(\result_real_1_tmp[5]~26_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[5]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[5] .is_wysiwyg = "true";
defparam \result_real_1_tmp[5] .power_up = "low";

dffeas \result_real_1_tmp[4] (
	.clk(clk),
	.d(\result_real_1_tmp[4]~24_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[4]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[4] .is_wysiwyg = "true";
defparam \result_real_1_tmp[4] .power_up = "low";

dffeas \result_real_1_tmp[3] (
	.clk(clk),
	.d(\result_real_1_tmp[3]~22_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[3]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[3] .is_wysiwyg = "true";
defparam \result_real_1_tmp[3] .power_up = "low";

dffeas \result_real_1_tmp[2] (
	.clk(clk),
	.d(\result_real_1_tmp[2]~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[2]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[2] .is_wysiwyg = "true";
defparam \result_real_1_tmp[2] .power_up = "low";

dffeas \result_real_1_tmp[1] (
	.clk(clk),
	.d(\result_real_1_tmp[1]~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[1]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[1] .is_wysiwyg = "true";
defparam \result_real_1_tmp[1] .power_up = "low";

dffeas \result_real_1_tmp[0] (
	.clk(clk),
	.d(\result_real_1_tmp[0]~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[0]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[0] .is_wysiwyg = "true";
defparam \result_real_1_tmp[0] .power_up = "low";

dffeas \result_real_1_tmp[15] (
	.clk(clk),
	.d(\result_real_1_tmp[15]~46_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[15]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[15] .is_wysiwyg = "true";
defparam \result_real_1_tmp[15] .power_up = "low";

dffeas \result_real_1_tmp[14] (
	.clk(clk),
	.d(\result_real_1_tmp[14]~44_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[14]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[14] .is_wysiwyg = "true";
defparam \result_real_1_tmp[14] .power_up = "low";

dffeas \result_real_1_tmp[13] (
	.clk(clk),
	.d(\result_real_1_tmp[13]~42_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[13]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[13] .is_wysiwyg = "true";
defparam \result_real_1_tmp[13] .power_up = "low";

dffeas \result_real_1_tmp[12] (
	.clk(clk),
	.d(\result_real_1_tmp[12]~40_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[12]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[12] .is_wysiwyg = "true";
defparam \result_real_1_tmp[12] .power_up = "low";

cycloneiii_lcell_comb \addresult_ac_bd[0]~16 (
	.dataa(\result_a_c_se[0]~q ),
	.datab(\result_b_d_se[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\addresult_ac_bd[0]~16_combout ),
	.cout(\addresult_ac_bd[0]~17 ));
defparam \addresult_ac_bd[0]~16 .lut_mask = 16'h66EE;
defparam \addresult_ac_bd[0]~16 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \addresult_ac_bd[1]~18 (
	.dataa(\result_a_c_se[1]~q ),
	.datab(\result_b_d_se[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[0]~17 ),
	.combout(\addresult_ac_bd[1]~18_combout ),
	.cout(\addresult_ac_bd[1]~19 ));
defparam \addresult_ac_bd[1]~18 .lut_mask = 16'h967F;
defparam \addresult_ac_bd[1]~18 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_ac_bd[2]~20 (
	.dataa(\result_a_c_se[2]~q ),
	.datab(\result_b_d_se[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[1]~19 ),
	.combout(\addresult_ac_bd[2]~20_combout ),
	.cout(\addresult_ac_bd[2]~21 ));
defparam \addresult_ac_bd[2]~20 .lut_mask = 16'h96EF;
defparam \addresult_ac_bd[2]~20 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_ac_bd[3]~22 (
	.dataa(\result_a_c_se[3]~q ),
	.datab(\result_b_d_se[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[2]~21 ),
	.combout(\addresult_ac_bd[3]~22_combout ),
	.cout(\addresult_ac_bd[3]~23 ));
defparam \addresult_ac_bd[3]~22 .lut_mask = 16'h967F;
defparam \addresult_ac_bd[3]~22 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_ac_bd[4]~24 (
	.dataa(\result_a_c_se[4]~q ),
	.datab(\result_b_d_se[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[3]~23 ),
	.combout(\addresult_ac_bd[4]~24_combout ),
	.cout(\addresult_ac_bd[4]~25 ));
defparam \addresult_ac_bd[4]~24 .lut_mask = 16'h96EF;
defparam \addresult_ac_bd[4]~24 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_ac_bd[5]~26 (
	.dataa(\result_a_c_se[5]~q ),
	.datab(\result_b_d_se[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[4]~25 ),
	.combout(\addresult_ac_bd[5]~26_combout ),
	.cout(\addresult_ac_bd[5]~27 ));
defparam \addresult_ac_bd[5]~26 .lut_mask = 16'h967F;
defparam \addresult_ac_bd[5]~26 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_ac_bd[6]~28 (
	.dataa(\result_a_c_se[6]~q ),
	.datab(\result_b_d_se[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[5]~27 ),
	.combout(\addresult_ac_bd[6]~28_combout ),
	.cout(\addresult_ac_bd[6]~29 ));
defparam \addresult_ac_bd[6]~28 .lut_mask = 16'h96EF;
defparam \addresult_ac_bd[6]~28 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_ac_bd[7]~30 (
	.dataa(\result_a_c_se[7]~q ),
	.datab(\result_b_d_se[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[6]~29 ),
	.combout(\addresult_ac_bd[7]~30_combout ),
	.cout(\addresult_ac_bd[7]~31 ));
defparam \addresult_ac_bd[7]~30 .lut_mask = 16'h967F;
defparam \addresult_ac_bd[7]~30 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_ac_bd[8]~32 (
	.dataa(\result_a_c_se[8]~q ),
	.datab(\result_b_d_se[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[7]~31 ),
	.combout(\addresult_ac_bd[8]~32_combout ),
	.cout(\addresult_ac_bd[8]~33 ));
defparam \addresult_ac_bd[8]~32 .lut_mask = 16'h96EF;
defparam \addresult_ac_bd[8]~32 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_ac_bd[9]~34 (
	.dataa(\result_a_c_se[9]~q ),
	.datab(\result_b_d_se[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[8]~33 ),
	.combout(\addresult_ac_bd[9]~34_combout ),
	.cout(\addresult_ac_bd[9]~35 ));
defparam \addresult_ac_bd[9]~34 .lut_mask = 16'h967F;
defparam \addresult_ac_bd[9]~34 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_ac_bd[10]~36 (
	.dataa(\result_a_c_se[10]~q ),
	.datab(\result_b_d_se[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[9]~35 ),
	.combout(\addresult_ac_bd[10]~36_combout ),
	.cout(\addresult_ac_bd[10]~37 ));
defparam \addresult_ac_bd[10]~36 .lut_mask = 16'h96EF;
defparam \addresult_ac_bd[10]~36 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_ac_bd[11]~38 (
	.dataa(\result_a_c_se[11]~q ),
	.datab(\result_b_d_se[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[10]~37 ),
	.combout(\addresult_ac_bd[11]~38_combout ),
	.cout(\addresult_ac_bd[11]~39 ));
defparam \addresult_ac_bd[11]~38 .lut_mask = 16'h967F;
defparam \addresult_ac_bd[11]~38 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_ac_bd[12]~40 (
	.dataa(\result_a_c_se[12]~q ),
	.datab(\result_b_d_se[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[11]~39 ),
	.combout(\addresult_ac_bd[12]~40_combout ),
	.cout(\addresult_ac_bd[12]~41 ));
defparam \addresult_ac_bd[12]~40 .lut_mask = 16'h96EF;
defparam \addresult_ac_bd[12]~40 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_ac_bd[13]~42 (
	.dataa(\result_a_c_se[13]~q ),
	.datab(\result_b_d_se[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[12]~41 ),
	.combout(\addresult_ac_bd[13]~42_combout ),
	.cout(\addresult_ac_bd[13]~43 ));
defparam \addresult_ac_bd[13]~42 .lut_mask = 16'h967F;
defparam \addresult_ac_bd[13]~42 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_ac_bd[14]~44 (
	.dataa(\result_a_c_se[14]~q ),
	.datab(\result_b_d_se[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[13]~43 ),
	.combout(\addresult_ac_bd[14]~44_combout ),
	.cout(\addresult_ac_bd[14]~45 ));
defparam \addresult_ac_bd[14]~44 .lut_mask = 16'h96EF;
defparam \addresult_ac_bd[14]~44 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_ac_bd[15]~46 (
	.dataa(\result_a_c_se[15]~q ),
	.datab(\result_b_d_se[15]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\addresult_ac_bd[14]~45 ),
	.combout(\addresult_ac_bd[15]~46_combout ),
	.cout());
defparam \addresult_ac_bd[15]~46 .lut_mask = 16'h9696;
defparam \addresult_ac_bd[15]~46 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_real_1_tmp[0]~16 (
	.dataa(\result_a_c_se[0]~q ),
	.datab(\result_b_d_se[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\result_real_1_tmp[0]~16_combout ),
	.cout(\result_real_1_tmp[0]~17 ));
defparam \result_real_1_tmp[0]~16 .lut_mask = 16'h66BB;
defparam \result_real_1_tmp[0]~16 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \result_real_1_tmp[1]~18 (
	.dataa(\result_a_c_se[1]~q ),
	.datab(\result_b_d_se[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[0]~17 ),
	.combout(\result_real_1_tmp[1]~18_combout ),
	.cout(\result_real_1_tmp[1]~19 ));
defparam \result_real_1_tmp[1]~18 .lut_mask = 16'h96DF;
defparam \result_real_1_tmp[1]~18 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_real_1_tmp[2]~20 (
	.dataa(\result_a_c_se[2]~q ),
	.datab(\result_b_d_se[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[1]~19 ),
	.combout(\result_real_1_tmp[2]~20_combout ),
	.cout(\result_real_1_tmp[2]~21 ));
defparam \result_real_1_tmp[2]~20 .lut_mask = 16'h96BF;
defparam \result_real_1_tmp[2]~20 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_real_1_tmp[3]~22 (
	.dataa(\result_a_c_se[3]~q ),
	.datab(\result_b_d_se[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[2]~21 ),
	.combout(\result_real_1_tmp[3]~22_combout ),
	.cout(\result_real_1_tmp[3]~23 ));
defparam \result_real_1_tmp[3]~22 .lut_mask = 16'h96DF;
defparam \result_real_1_tmp[3]~22 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_real_1_tmp[4]~24 (
	.dataa(\result_a_c_se[4]~q ),
	.datab(\result_b_d_se[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[3]~23 ),
	.combout(\result_real_1_tmp[4]~24_combout ),
	.cout(\result_real_1_tmp[4]~25 ));
defparam \result_real_1_tmp[4]~24 .lut_mask = 16'h96BF;
defparam \result_real_1_tmp[4]~24 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_real_1_tmp[5]~26 (
	.dataa(\result_a_c_se[5]~q ),
	.datab(\result_b_d_se[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[4]~25 ),
	.combout(\result_real_1_tmp[5]~26_combout ),
	.cout(\result_real_1_tmp[5]~27 ));
defparam \result_real_1_tmp[5]~26 .lut_mask = 16'h96DF;
defparam \result_real_1_tmp[5]~26 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_real_1_tmp[6]~28 (
	.dataa(\result_a_c_se[6]~q ),
	.datab(\result_b_d_se[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[5]~27 ),
	.combout(\result_real_1_tmp[6]~28_combout ),
	.cout(\result_real_1_tmp[6]~29 ));
defparam \result_real_1_tmp[6]~28 .lut_mask = 16'h96BF;
defparam \result_real_1_tmp[6]~28 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_real_1_tmp[7]~30 (
	.dataa(\result_a_c_se[7]~q ),
	.datab(\result_b_d_se[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[6]~29 ),
	.combout(\result_real_1_tmp[7]~30_combout ),
	.cout(\result_real_1_tmp[7]~31 ));
defparam \result_real_1_tmp[7]~30 .lut_mask = 16'h96DF;
defparam \result_real_1_tmp[7]~30 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_real_1_tmp[8]~32 (
	.dataa(\result_a_c_se[8]~q ),
	.datab(\result_b_d_se[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[7]~31 ),
	.combout(\result_real_1_tmp[8]~32_combout ),
	.cout(\result_real_1_tmp[8]~33 ));
defparam \result_real_1_tmp[8]~32 .lut_mask = 16'h96BF;
defparam \result_real_1_tmp[8]~32 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_real_1_tmp[9]~34 (
	.dataa(\result_a_c_se[9]~q ),
	.datab(\result_b_d_se[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[8]~33 ),
	.combout(\result_real_1_tmp[9]~34_combout ),
	.cout(\result_real_1_tmp[9]~35 ));
defparam \result_real_1_tmp[9]~34 .lut_mask = 16'h96DF;
defparam \result_real_1_tmp[9]~34 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_real_1_tmp[10]~36 (
	.dataa(\result_a_c_se[10]~q ),
	.datab(\result_b_d_se[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[9]~35 ),
	.combout(\result_real_1_tmp[10]~36_combout ),
	.cout(\result_real_1_tmp[10]~37 ));
defparam \result_real_1_tmp[10]~36 .lut_mask = 16'h96BF;
defparam \result_real_1_tmp[10]~36 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_real_1_tmp[11]~38 (
	.dataa(\result_a_c_se[11]~q ),
	.datab(\result_b_d_se[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[10]~37 ),
	.combout(\result_real_1_tmp[11]~38_combout ),
	.cout(\result_real_1_tmp[11]~39 ));
defparam \result_real_1_tmp[11]~38 .lut_mask = 16'h96DF;
defparam \result_real_1_tmp[11]~38 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_real_1_tmp[12]~40 (
	.dataa(\result_a_c_se[12]~q ),
	.datab(\result_b_d_se[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[11]~39 ),
	.combout(\result_real_1_tmp[12]~40_combout ),
	.cout(\result_real_1_tmp[12]~41 ));
defparam \result_real_1_tmp[12]~40 .lut_mask = 16'h96BF;
defparam \result_real_1_tmp[12]~40 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_real_1_tmp[13]~42 (
	.dataa(\result_a_c_se[13]~q ),
	.datab(\result_b_d_se[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[12]~41 ),
	.combout(\result_real_1_tmp[13]~42_combout ),
	.cout(\result_real_1_tmp[13]~43 ));
defparam \result_real_1_tmp[13]~42 .lut_mask = 16'h96DF;
defparam \result_real_1_tmp[13]~42 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_real_1_tmp[14]~44 (
	.dataa(\result_a_c_se[14]~q ),
	.datab(\result_b_d_se[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[13]~43 ),
	.combout(\result_real_1_tmp[14]~44_combout ),
	.cout(\result_real_1_tmp[14]~45 ));
defparam \result_real_1_tmp[14]~44 .lut_mask = 16'h96BF;
defparam \result_real_1_tmp[14]~44 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \result_real_1_tmp[15]~46 (
	.dataa(\result_a_c_se[15]~q ),
	.datab(\result_b_d_se[15]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\result_real_1_tmp[14]~45 ),
	.combout(\result_real_1_tmp[15]~46_combout ),
	.cout());
defparam \result_real_1_tmp[15]~46 .lut_mask = 16'h9696;
defparam \result_real_1_tmp[15]~46 .sum_lutc_input = "cin";

dffeas \addresult_a_b[0] (
	.clk(clk),
	.d(\addresult_a_b[0]~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_a_b[0]~q ),
	.prn(vcc));
defparam \addresult_a_b[0] .is_wysiwyg = "true";
defparam \addresult_a_b[0] .power_up = "low";

dffeas \addresult_a_b[1] (
	.clk(clk),
	.d(\addresult_a_b[1]~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_a_b[1]~q ),
	.prn(vcc));
defparam \addresult_a_b[1] .is_wysiwyg = "true";
defparam \addresult_a_b[1] .power_up = "low";

dffeas \addresult_a_b[2] (
	.clk(clk),
	.d(\addresult_a_b[2]~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_a_b[2]~q ),
	.prn(vcc));
defparam \addresult_a_b[2] .is_wysiwyg = "true";
defparam \addresult_a_b[2] .power_up = "low";

dffeas \addresult_a_b[3] (
	.clk(clk),
	.d(\addresult_a_b[3]~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_a_b[3]~q ),
	.prn(vcc));
defparam \addresult_a_b[3] .is_wysiwyg = "true";
defparam \addresult_a_b[3] .power_up = "low";

dffeas \addresult_a_b[4] (
	.clk(clk),
	.d(\addresult_a_b[4]~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_a_b[4]~q ),
	.prn(vcc));
defparam \addresult_a_b[4] .is_wysiwyg = "true";
defparam \addresult_a_b[4] .power_up = "low";

dffeas \addresult_a_b[5] (
	.clk(clk),
	.d(\addresult_a_b[5]~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_a_b[5]~q ),
	.prn(vcc));
defparam \addresult_a_b[5] .is_wysiwyg = "true";
defparam \addresult_a_b[5] .power_up = "low";

dffeas \addresult_a_b[6] (
	.clk(clk),
	.d(\addresult_a_b[6]~21_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_a_b[6]~q ),
	.prn(vcc));
defparam \addresult_a_b[6] .is_wysiwyg = "true";
defparam \addresult_a_b[6] .power_up = "low";

dffeas \addresult_a_b[7] (
	.clk(clk),
	.d(\addresult_a_b[7]~23_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_a_b[7]~q ),
	.prn(vcc));
defparam \addresult_a_b[7] .is_wysiwyg = "true";
defparam \addresult_a_b[7] .power_up = "low";

dffeas \addresult_a_b[8] (
	.clk(clk),
	.d(\addresult_a_b[8]~25_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_a_b[8]~q ),
	.prn(vcc));
defparam \addresult_a_b[8] .is_wysiwyg = "true";
defparam \addresult_a_b[8] .power_up = "low";

dffeas \addresult_c_d[0] (
	.clk(clk),
	.d(\addresult_c_d[0]~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_c_d[0]~q ),
	.prn(vcc));
defparam \addresult_c_d[0] .is_wysiwyg = "true";
defparam \addresult_c_d[0] .power_up = "low";

dffeas \addresult_c_d[1] (
	.clk(clk),
	.d(\addresult_c_d[1]~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_c_d[1]~q ),
	.prn(vcc));
defparam \addresult_c_d[1] .is_wysiwyg = "true";
defparam \addresult_c_d[1] .power_up = "low";

dffeas \addresult_c_d[2] (
	.clk(clk),
	.d(\addresult_c_d[2]~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_c_d[2]~q ),
	.prn(vcc));
defparam \addresult_c_d[2] .is_wysiwyg = "true";
defparam \addresult_c_d[2] .power_up = "low";

dffeas \addresult_c_d[3] (
	.clk(clk),
	.d(\addresult_c_d[3]~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_c_d[3]~q ),
	.prn(vcc));
defparam \addresult_c_d[3] .is_wysiwyg = "true";
defparam \addresult_c_d[3] .power_up = "low";

dffeas \addresult_c_d[4] (
	.clk(clk),
	.d(\addresult_c_d[4]~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_c_d[4]~q ),
	.prn(vcc));
defparam \addresult_c_d[4] .is_wysiwyg = "true";
defparam \addresult_c_d[4] .power_up = "low";

dffeas \addresult_c_d[5] (
	.clk(clk),
	.d(\addresult_c_d[5]~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_c_d[5]~q ),
	.prn(vcc));
defparam \addresult_c_d[5] .is_wysiwyg = "true";
defparam \addresult_c_d[5] .power_up = "low";

dffeas \addresult_c_d[6] (
	.clk(clk),
	.d(\addresult_c_d[6]~21_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_c_d[6]~q ),
	.prn(vcc));
defparam \addresult_c_d[6] .is_wysiwyg = "true";
defparam \addresult_c_d[6] .power_up = "low";

dffeas \addresult_c_d[7] (
	.clk(clk),
	.d(\addresult_c_d[7]~23_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_c_d[7]~q ),
	.prn(vcc));
defparam \addresult_c_d[7] .is_wysiwyg = "true";
defparam \addresult_c_d[7] .power_up = "low";

dffeas \addresult_c_d[8] (
	.clk(clk),
	.d(\addresult_c_d[8]~25_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_c_d[8]~q ),
	.prn(vcc));
defparam \addresult_c_d[8] .is_wysiwyg = "true";
defparam \addresult_c_d[8] .power_up = "low";

cycloneiii_lcell_comb \addresult_a_b[0]~9 (
	.dataa(pipeline_dffe_2),
	.datab(pipeline_dffe_21),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\addresult_a_b[0]~9_combout ),
	.cout(\addresult_a_b[0]~10 ));
defparam \addresult_a_b[0]~9 .lut_mask = 16'h66EE;
defparam \addresult_a_b[0]~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \addresult_a_b[1]~11 (
	.dataa(pipeline_dffe_3),
	.datab(pipeline_dffe_31),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_a_b[0]~10 ),
	.combout(\addresult_a_b[1]~11_combout ),
	.cout(\addresult_a_b[1]~12 ));
defparam \addresult_a_b[1]~11 .lut_mask = 16'h967F;
defparam \addresult_a_b[1]~11 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_a_b[2]~13 (
	.dataa(pipeline_dffe_4),
	.datab(pipeline_dffe_41),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_a_b[1]~12 ),
	.combout(\addresult_a_b[2]~13_combout ),
	.cout(\addresult_a_b[2]~14 ));
defparam \addresult_a_b[2]~13 .lut_mask = 16'h96EF;
defparam \addresult_a_b[2]~13 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_a_b[3]~15 (
	.dataa(pipeline_dffe_5),
	.datab(pipeline_dffe_51),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_a_b[2]~14 ),
	.combout(\addresult_a_b[3]~15_combout ),
	.cout(\addresult_a_b[3]~16 ));
defparam \addresult_a_b[3]~15 .lut_mask = 16'h967F;
defparam \addresult_a_b[3]~15 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_a_b[4]~17 (
	.dataa(pipeline_dffe_6),
	.datab(pipeline_dffe_61),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_a_b[3]~16 ),
	.combout(\addresult_a_b[4]~17_combout ),
	.cout(\addresult_a_b[4]~18 ));
defparam \addresult_a_b[4]~17 .lut_mask = 16'h96EF;
defparam \addresult_a_b[4]~17 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_a_b[5]~19 (
	.dataa(pipeline_dffe_7),
	.datab(pipeline_dffe_71),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_a_b[4]~18 ),
	.combout(\addresult_a_b[5]~19_combout ),
	.cout(\addresult_a_b[5]~20 ));
defparam \addresult_a_b[5]~19 .lut_mask = 16'h967F;
defparam \addresult_a_b[5]~19 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_a_b[6]~21 (
	.dataa(pipeline_dffe_81),
	.datab(pipeline_dffe_82),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_a_b[5]~20 ),
	.combout(\addresult_a_b[6]~21_combout ),
	.cout(\addresult_a_b[6]~22 ));
defparam \addresult_a_b[6]~21 .lut_mask = 16'h96EF;
defparam \addresult_a_b[6]~21 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_a_b[7]~23 (
	.dataa(pipeline_dffe_91),
	.datab(pipeline_dffe_92),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_a_b[6]~22 ),
	.combout(\addresult_a_b[7]~23_combout ),
	.cout(\addresult_a_b[7]~24 ));
defparam \addresult_a_b[7]~23 .lut_mask = 16'h967F;
defparam \addresult_a_b[7]~23 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_a_b[8]~25 (
	.dataa(pipeline_dffe_91),
	.datab(pipeline_dffe_92),
	.datac(gnd),
	.datad(gnd),
	.cin(\addresult_a_b[7]~24 ),
	.combout(\addresult_a_b[8]~25_combout ),
	.cout());
defparam \addresult_a_b[8]~25 .lut_mask = 16'h9696;
defparam \addresult_a_b[8]~25 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_c_d[0]~9 (
	.dataa(twiddle_data200),
	.datab(twiddle_data210),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\addresult_c_d[0]~9_combout ),
	.cout(\addresult_c_d[0]~10 ));
defparam \addresult_c_d[0]~9 .lut_mask = 16'h66EE;
defparam \addresult_c_d[0]~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \addresult_c_d[1]~11 (
	.dataa(twiddle_data201),
	.datab(twiddle_data211),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_c_d[0]~10 ),
	.combout(\addresult_c_d[1]~11_combout ),
	.cout(\addresult_c_d[1]~12 ));
defparam \addresult_c_d[1]~11 .lut_mask = 16'h967F;
defparam \addresult_c_d[1]~11 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_c_d[2]~13 (
	.dataa(twiddle_data202),
	.datab(twiddle_data212),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_c_d[1]~12 ),
	.combout(\addresult_c_d[2]~13_combout ),
	.cout(\addresult_c_d[2]~14 ));
defparam \addresult_c_d[2]~13 .lut_mask = 16'h96EF;
defparam \addresult_c_d[2]~13 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_c_d[3]~15 (
	.dataa(twiddle_data203),
	.datab(twiddle_data213),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_c_d[2]~14 ),
	.combout(\addresult_c_d[3]~15_combout ),
	.cout(\addresult_c_d[3]~16 ));
defparam \addresult_c_d[3]~15 .lut_mask = 16'h967F;
defparam \addresult_c_d[3]~15 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_c_d[4]~17 (
	.dataa(twiddle_data204),
	.datab(twiddle_data214),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_c_d[3]~16 ),
	.combout(\addresult_c_d[4]~17_combout ),
	.cout(\addresult_c_d[4]~18 ));
defparam \addresult_c_d[4]~17 .lut_mask = 16'h96EF;
defparam \addresult_c_d[4]~17 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_c_d[5]~19 (
	.dataa(twiddle_data205),
	.datab(twiddle_data215),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_c_d[4]~18 ),
	.combout(\addresult_c_d[5]~19_combout ),
	.cout(\addresult_c_d[5]~20 ));
defparam \addresult_c_d[5]~19 .lut_mask = 16'h967F;
defparam \addresult_c_d[5]~19 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_c_d[6]~21 (
	.dataa(twiddle_data206),
	.datab(twiddle_data216),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_c_d[5]~20 ),
	.combout(\addresult_c_d[6]~21_combout ),
	.cout(\addresult_c_d[6]~22 ));
defparam \addresult_c_d[6]~21 .lut_mask = 16'h96EF;
defparam \addresult_c_d[6]~21 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_c_d[7]~23 (
	.dataa(twiddle_data207),
	.datab(twiddle_data217),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_c_d[6]~22 ),
	.combout(\addresult_c_d[7]~23_combout ),
	.cout(\addresult_c_d[7]~24 ));
defparam \addresult_c_d[7]~23 .lut_mask = 16'h967F;
defparam \addresult_c_d[7]~23 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \addresult_c_d[8]~25 (
	.dataa(twiddle_data207),
	.datab(twiddle_data217),
	.datac(gnd),
	.datad(gnd),
	.cin(\addresult_c_d[7]~24 ),
	.combout(\addresult_c_d[8]~25_combout ),
	.cout());
defparam \addresult_c_d[8]~25 .lut_mask = 16'h9696;
defparam \addresult_c_d[8]~25 .sum_lutc_input = "cin";

dffeas \result_a_b_c_d_se[11] (
	.clk(clk),
	.d(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[11]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[11] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[11] .power_up = "low";

dffeas \result_a_b_c_d_se[10] (
	.clk(clk),
	.d(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[10]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[10] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[10] .power_up = "low";

dffeas \result_a_b_c_d_se[9] (
	.clk(clk),
	.d(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[9]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[9] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[9] .power_up = "low";

dffeas \result_a_b_c_d_se[8] (
	.clk(clk),
	.d(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[8]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[8] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[8] .power_up = "low";

dffeas \result_a_b_c_d_se[7] (
	.clk(clk),
	.d(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[7]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[7] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[7] .power_up = "low";

dffeas \result_a_b_c_d_se[6] (
	.clk(clk),
	.d(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[6]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[6] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[6] .power_up = "low";

dffeas \result_a_b_c_d_se[5] (
	.clk(clk),
	.d(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[5]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[5] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[5] .power_up = "low";

dffeas \result_a_b_c_d_se[4] (
	.clk(clk),
	.d(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[4]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[4] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[4] .power_up = "low";

dffeas \result_a_b_c_d_se[3] (
	.clk(clk),
	.d(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[3]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[3] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[3] .power_up = "low";

dffeas \result_a_b_c_d_se[2] (
	.clk(clk),
	.d(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[2]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[2] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[2] .power_up = "low";

dffeas \result_a_b_c_d_se[1] (
	.clk(clk),
	.d(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[1]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[1] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[1] .power_up = "low";

dffeas \result_a_b_c_d_se[0] (
	.clk(clk),
	.d(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[0]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[0] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[0] .power_up = "low";

dffeas \result_a_b_c_d_se[15] (
	.clk(clk),
	.d(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[15]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[15] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[15] .power_up = "low";

dffeas \result_a_b_c_d_se[14] (
	.clk(clk),
	.d(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[14]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[14] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[14] .power_up = "low";

dffeas \result_a_b_c_d_se[13] (
	.clk(clk),
	.d(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[13]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[13] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[13] .power_up = "low";

dffeas \result_a_b_c_d_se[12] (
	.clk(clk),
	.d(\gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[12]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[12] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[12] .power_up = "low";

dffeas \result_a_c_se[11] (
	.clk(clk),
	.d(\gen_dsp_only:m_ac|auto_generated|dffe3a[11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[11]~q ),
	.prn(vcc));
defparam \result_a_c_se[11] .is_wysiwyg = "true";
defparam \result_a_c_se[11] .power_up = "low";

dffeas \result_b_d_se[11] (
	.clk(clk),
	.d(\gen_dsp_only:m_bd|auto_generated|dffe3a[11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[11]~q ),
	.prn(vcc));
defparam \result_b_d_se[11] .is_wysiwyg = "true";
defparam \result_b_d_se[11] .power_up = "low";

dffeas \result_a_c_se[10] (
	.clk(clk),
	.d(\gen_dsp_only:m_ac|auto_generated|dffe3a[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[10]~q ),
	.prn(vcc));
defparam \result_a_c_se[10] .is_wysiwyg = "true";
defparam \result_a_c_se[10] .power_up = "low";

dffeas \result_b_d_se[10] (
	.clk(clk),
	.d(\gen_dsp_only:m_bd|auto_generated|dffe3a[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[10]~q ),
	.prn(vcc));
defparam \result_b_d_se[10] .is_wysiwyg = "true";
defparam \result_b_d_se[10] .power_up = "low";

dffeas \result_a_c_se[9] (
	.clk(clk),
	.d(\gen_dsp_only:m_ac|auto_generated|dffe3a[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[9]~q ),
	.prn(vcc));
defparam \result_a_c_se[9] .is_wysiwyg = "true";
defparam \result_a_c_se[9] .power_up = "low";

dffeas \result_b_d_se[9] (
	.clk(clk),
	.d(\gen_dsp_only:m_bd|auto_generated|dffe3a[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[9]~q ),
	.prn(vcc));
defparam \result_b_d_se[9] .is_wysiwyg = "true";
defparam \result_b_d_se[9] .power_up = "low";

dffeas \result_a_c_se[8] (
	.clk(clk),
	.d(\gen_dsp_only:m_ac|auto_generated|dffe3a[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[8]~q ),
	.prn(vcc));
defparam \result_a_c_se[8] .is_wysiwyg = "true";
defparam \result_a_c_se[8] .power_up = "low";

dffeas \result_b_d_se[8] (
	.clk(clk),
	.d(\gen_dsp_only:m_bd|auto_generated|dffe3a[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[8]~q ),
	.prn(vcc));
defparam \result_b_d_se[8] .is_wysiwyg = "true";
defparam \result_b_d_se[8] .power_up = "low";

dffeas \result_a_c_se[7] (
	.clk(clk),
	.d(\gen_dsp_only:m_ac|auto_generated|dffe3a[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[7]~q ),
	.prn(vcc));
defparam \result_a_c_se[7] .is_wysiwyg = "true";
defparam \result_a_c_se[7] .power_up = "low";

dffeas \result_b_d_se[7] (
	.clk(clk),
	.d(\gen_dsp_only:m_bd|auto_generated|dffe3a[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[7]~q ),
	.prn(vcc));
defparam \result_b_d_se[7] .is_wysiwyg = "true";
defparam \result_b_d_se[7] .power_up = "low";

dffeas \result_a_c_se[6] (
	.clk(clk),
	.d(\gen_dsp_only:m_ac|auto_generated|dffe3a[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[6]~q ),
	.prn(vcc));
defparam \result_a_c_se[6] .is_wysiwyg = "true";
defparam \result_a_c_se[6] .power_up = "low";

dffeas \result_b_d_se[6] (
	.clk(clk),
	.d(\gen_dsp_only:m_bd|auto_generated|dffe3a[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[6]~q ),
	.prn(vcc));
defparam \result_b_d_se[6] .is_wysiwyg = "true";
defparam \result_b_d_se[6] .power_up = "low";

dffeas \result_a_c_se[5] (
	.clk(clk),
	.d(\gen_dsp_only:m_ac|auto_generated|dffe3a[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[5]~q ),
	.prn(vcc));
defparam \result_a_c_se[5] .is_wysiwyg = "true";
defparam \result_a_c_se[5] .power_up = "low";

dffeas \result_b_d_se[5] (
	.clk(clk),
	.d(\gen_dsp_only:m_bd|auto_generated|dffe3a[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[5]~q ),
	.prn(vcc));
defparam \result_b_d_se[5] .is_wysiwyg = "true";
defparam \result_b_d_se[5] .power_up = "low";

dffeas \result_a_c_se[4] (
	.clk(clk),
	.d(\gen_dsp_only:m_ac|auto_generated|dffe3a[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[4]~q ),
	.prn(vcc));
defparam \result_a_c_se[4] .is_wysiwyg = "true";
defparam \result_a_c_se[4] .power_up = "low";

dffeas \result_b_d_se[4] (
	.clk(clk),
	.d(\gen_dsp_only:m_bd|auto_generated|dffe3a[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[4]~q ),
	.prn(vcc));
defparam \result_b_d_se[4] .is_wysiwyg = "true";
defparam \result_b_d_se[4] .power_up = "low";

dffeas \result_a_c_se[3] (
	.clk(clk),
	.d(\gen_dsp_only:m_ac|auto_generated|dffe3a[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[3]~q ),
	.prn(vcc));
defparam \result_a_c_se[3] .is_wysiwyg = "true";
defparam \result_a_c_se[3] .power_up = "low";

dffeas \result_b_d_se[3] (
	.clk(clk),
	.d(\gen_dsp_only:m_bd|auto_generated|dffe3a[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[3]~q ),
	.prn(vcc));
defparam \result_b_d_se[3] .is_wysiwyg = "true";
defparam \result_b_d_se[3] .power_up = "low";

dffeas \result_a_c_se[2] (
	.clk(clk),
	.d(\gen_dsp_only:m_ac|auto_generated|dffe3a[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[2]~q ),
	.prn(vcc));
defparam \result_a_c_se[2] .is_wysiwyg = "true";
defparam \result_a_c_se[2] .power_up = "low";

dffeas \result_b_d_se[2] (
	.clk(clk),
	.d(\gen_dsp_only:m_bd|auto_generated|dffe3a[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[2]~q ),
	.prn(vcc));
defparam \result_b_d_se[2] .is_wysiwyg = "true";
defparam \result_b_d_se[2] .power_up = "low";

dffeas \result_a_c_se[1] (
	.clk(clk),
	.d(\gen_dsp_only:m_ac|auto_generated|dffe3a[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[1]~q ),
	.prn(vcc));
defparam \result_a_c_se[1] .is_wysiwyg = "true";
defparam \result_a_c_se[1] .power_up = "low";

dffeas \result_b_d_se[1] (
	.clk(clk),
	.d(\gen_dsp_only:m_bd|auto_generated|dffe3a[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[1]~q ),
	.prn(vcc));
defparam \result_b_d_se[1] .is_wysiwyg = "true";
defparam \result_b_d_se[1] .power_up = "low";

dffeas \result_a_c_se[0] (
	.clk(clk),
	.d(\gen_dsp_only:m_ac|auto_generated|dffe3a[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[0]~q ),
	.prn(vcc));
defparam \result_a_c_se[0] .is_wysiwyg = "true";
defparam \result_a_c_se[0] .power_up = "low";

dffeas \result_b_d_se[0] (
	.clk(clk),
	.d(\gen_dsp_only:m_bd|auto_generated|dffe3a[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[0]~q ),
	.prn(vcc));
defparam \result_b_d_se[0] .is_wysiwyg = "true";
defparam \result_b_d_se[0] .power_up = "low";

dffeas \result_a_c_se[15] (
	.clk(clk),
	.d(\gen_dsp_only:m_ac|auto_generated|dffe3a[15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[15]~q ),
	.prn(vcc));
defparam \result_a_c_se[15] .is_wysiwyg = "true";
defparam \result_a_c_se[15] .power_up = "low";

dffeas \result_b_d_se[15] (
	.clk(clk),
	.d(\gen_dsp_only:m_bd|auto_generated|dffe3a[15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[15]~q ),
	.prn(vcc));
defparam \result_b_d_se[15] .is_wysiwyg = "true";
defparam \result_b_d_se[15] .power_up = "low";

dffeas \result_a_c_se[14] (
	.clk(clk),
	.d(\gen_dsp_only:m_ac|auto_generated|dffe3a[14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[14]~q ),
	.prn(vcc));
defparam \result_a_c_se[14] .is_wysiwyg = "true";
defparam \result_a_c_se[14] .power_up = "low";

dffeas \result_b_d_se[14] (
	.clk(clk),
	.d(\gen_dsp_only:m_bd|auto_generated|dffe3a[14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[14]~q ),
	.prn(vcc));
defparam \result_b_d_se[14] .is_wysiwyg = "true";
defparam \result_b_d_se[14] .power_up = "low";

dffeas \result_a_c_se[13] (
	.clk(clk),
	.d(\gen_dsp_only:m_ac|auto_generated|dffe3a[13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[13]~q ),
	.prn(vcc));
defparam \result_a_c_se[13] .is_wysiwyg = "true";
defparam \result_a_c_se[13] .power_up = "low";

dffeas \result_b_d_se[13] (
	.clk(clk),
	.d(\gen_dsp_only:m_bd|auto_generated|dffe3a[13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[13]~q ),
	.prn(vcc));
defparam \result_b_d_se[13] .is_wysiwyg = "true";
defparam \result_b_d_se[13] .power_up = "low";

dffeas \result_a_c_se[12] (
	.clk(clk),
	.d(\gen_dsp_only:m_ac|auto_generated|dffe3a[12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[12]~q ),
	.prn(vcc));
defparam \result_a_c_se[12] .is_wysiwyg = "true";
defparam \result_a_c_se[12] .power_up = "low";

dffeas \result_b_d_se[12] (
	.clk(clk),
	.d(\gen_dsp_only:m_bd|auto_generated|dffe3a[12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[12]~q ),
	.prn(vcc));
defparam \result_b_d_se[12] .is_wysiwyg = "true";
defparam \result_b_d_se[12] .power_up = "low";

dffeas \real_out[3] (
	.clk(clk),
	.d(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(real_out_3),
	.prn(vcc));
defparam \real_out[3] .is_wysiwyg = "true";
defparam \real_out[3] .power_up = "low";

dffeas \real_out[7] (
	.clk(clk),
	.d(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(real_out_7),
	.prn(vcc));
defparam \real_out[7] .is_wysiwyg = "true";
defparam \real_out[7] .power_up = "low";

dffeas \real_out[4] (
	.clk(clk),
	.d(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(real_out_4),
	.prn(vcc));
defparam \real_out[4] .is_wysiwyg = "true";
defparam \real_out[4] .power_up = "low";

dffeas \real_out[5] (
	.clk(clk),
	.d(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(real_out_5),
	.prn(vcc));
defparam \real_out[5] .is_wysiwyg = "true";
defparam \real_out[5] .power_up = "low";

dffeas \real_out[6] (
	.clk(clk),
	.d(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(real_out_6),
	.prn(vcc));
defparam \real_out[6] .is_wysiwyg = "true";
defparam \real_out[6] .power_up = "low";

dffeas \real_out[1] (
	.clk(clk),
	.d(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(real_out_1),
	.prn(vcc));
defparam \real_out[1] .is_wysiwyg = "true";
defparam \real_out[1] .power_up = "low";

dffeas \real_out[0] (
	.clk(clk),
	.d(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(real_out_0),
	.prn(vcc));
defparam \real_out[0] .is_wysiwyg = "true";
defparam \real_out[0] .power_up = "low";

dffeas \real_out[2] (
	.clk(clk),
	.d(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(real_out_2),
	.prn(vcc));
defparam \real_out[2] .is_wysiwyg = "true";
defparam \real_out[2] .power_up = "low";

endmodule

module fft_asj_fft_pround_fft_120_4 (
	pipeline_dffe_11,
	pipeline_dffe_15,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	result_real_1_tmp_11,
	result_real_1_tmp_10,
	result_real_1_tmp_9,
	result_real_1_tmp_8,
	result_real_1_tmp_7,
	result_real_1_tmp_6,
	result_real_1_tmp_5,
	result_real_1_tmp_4,
	result_real_1_tmp_3,
	result_real_1_tmp_2,
	result_real_1_tmp_1,
	result_real_1_tmp_0,
	result_real_1_tmp_15,
	result_real_1_tmp_14,
	result_real_1_tmp_13,
	result_real_1_tmp_12,
	pipeline_dffe_9,
	pipeline_dffe_8,
	pipeline_dffe_10,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_11;
output 	pipeline_dffe_15;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
input 	result_real_1_tmp_11;
input 	result_real_1_tmp_10;
input 	result_real_1_tmp_9;
input 	result_real_1_tmp_8;
input 	result_real_1_tmp_7;
input 	result_real_1_tmp_6;
input 	result_real_1_tmp_5;
input 	result_real_1_tmp_4;
input 	result_real_1_tmp_3;
input 	result_real_1_tmp_2;
input 	result_real_1_tmp_1;
input 	result_real_1_tmp_0;
input 	result_real_1_tmp_15;
input 	result_real_1_tmp_14;
input 	result_real_1_tmp_13;
input 	result_real_1_tmp_12;
output 	pipeline_dffe_9;
output 	pipeline_dffe_8;
output 	pipeline_dffe_10;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_LPM_ADD_SUB_5 \gbrnd:nev:gp:lpm_add_sub_component (
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_14(pipeline_dffe_14),
	.result_real_1_tmp_11(result_real_1_tmp_11),
	.result_real_1_tmp_10(result_real_1_tmp_10),
	.result_real_1_tmp_9(result_real_1_tmp_9),
	.result_real_1_tmp_8(result_real_1_tmp_8),
	.result_real_1_tmp_7(result_real_1_tmp_7),
	.result_real_1_tmp_6(result_real_1_tmp_6),
	.result_real_1_tmp_5(result_real_1_tmp_5),
	.result_real_1_tmp_4(result_real_1_tmp_4),
	.result_real_1_tmp_3(result_real_1_tmp_3),
	.result_real_1_tmp_2(result_real_1_tmp_2),
	.result_real_1_tmp_1(result_real_1_tmp_1),
	.result_real_1_tmp_0(result_real_1_tmp_0),
	.result_real_1_tmp_15(result_real_1_tmp_15),
	.result_real_1_tmp_14(result_real_1_tmp_14),
	.result_real_1_tmp_13(result_real_1_tmp_13),
	.result_real_1_tmp_12(result_real_1_tmp_12),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_10(pipeline_dffe_10),
	.clken(global_clock_enable),
	.clock(clk));

endmodule

module fft_LPM_ADD_SUB_5 (
	pipeline_dffe_11,
	pipeline_dffe_15,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	result_real_1_tmp_11,
	result_real_1_tmp_10,
	result_real_1_tmp_9,
	result_real_1_tmp_8,
	result_real_1_tmp_7,
	result_real_1_tmp_6,
	result_real_1_tmp_5,
	result_real_1_tmp_4,
	result_real_1_tmp_3,
	result_real_1_tmp_2,
	result_real_1_tmp_1,
	result_real_1_tmp_0,
	result_real_1_tmp_15,
	result_real_1_tmp_14,
	result_real_1_tmp_13,
	result_real_1_tmp_12,
	pipeline_dffe_9,
	pipeline_dffe_8,
	pipeline_dffe_10,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_11;
output 	pipeline_dffe_15;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
input 	result_real_1_tmp_11;
input 	result_real_1_tmp_10;
input 	result_real_1_tmp_9;
input 	result_real_1_tmp_8;
input 	result_real_1_tmp_7;
input 	result_real_1_tmp_6;
input 	result_real_1_tmp_5;
input 	result_real_1_tmp_4;
input 	result_real_1_tmp_3;
input 	result_real_1_tmp_2;
input 	result_real_1_tmp_1;
input 	result_real_1_tmp_0;
input 	result_real_1_tmp_15;
input 	result_real_1_tmp_14;
input 	result_real_1_tmp_13;
input 	result_real_1_tmp_12;
output 	pipeline_dffe_9;
output 	pipeline_dffe_8;
output 	pipeline_dffe_10;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_add_sub_dmj_4 auto_generated(
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_14(pipeline_dffe_14),
	.result_real_1_tmp_11(result_real_1_tmp_11),
	.result_real_1_tmp_10(result_real_1_tmp_10),
	.result_real_1_tmp_9(result_real_1_tmp_9),
	.result_real_1_tmp_8(result_real_1_tmp_8),
	.result_real_1_tmp_7(result_real_1_tmp_7),
	.result_real_1_tmp_6(result_real_1_tmp_6),
	.result_real_1_tmp_5(result_real_1_tmp_5),
	.result_real_1_tmp_4(result_real_1_tmp_4),
	.result_real_1_tmp_3(result_real_1_tmp_3),
	.result_real_1_tmp_2(result_real_1_tmp_2),
	.result_real_1_tmp_1(result_real_1_tmp_1),
	.result_real_1_tmp_0(result_real_1_tmp_0),
	.result_real_1_tmp_15(result_real_1_tmp_15),
	.result_real_1_tmp_14(result_real_1_tmp_14),
	.result_real_1_tmp_13(result_real_1_tmp_13),
	.result_real_1_tmp_12(result_real_1_tmp_12),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_10(pipeline_dffe_10),
	.clken(clken),
	.clock(clock));

endmodule

module fft_add_sub_dmj_4 (
	pipeline_dffe_11,
	pipeline_dffe_15,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	result_real_1_tmp_11,
	result_real_1_tmp_10,
	result_real_1_tmp_9,
	result_real_1_tmp_8,
	result_real_1_tmp_7,
	result_real_1_tmp_6,
	result_real_1_tmp_5,
	result_real_1_tmp_4,
	result_real_1_tmp_3,
	result_real_1_tmp_2,
	result_real_1_tmp_1,
	result_real_1_tmp_0,
	result_real_1_tmp_15,
	result_real_1_tmp_14,
	result_real_1_tmp_13,
	result_real_1_tmp_12,
	pipeline_dffe_9,
	pipeline_dffe_8,
	pipeline_dffe_10,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_11;
output 	pipeline_dffe_15;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
input 	result_real_1_tmp_11;
input 	result_real_1_tmp_10;
input 	result_real_1_tmp_9;
input 	result_real_1_tmp_8;
input 	result_real_1_tmp_7;
input 	result_real_1_tmp_6;
input 	result_real_1_tmp_5;
input 	result_real_1_tmp_4;
input 	result_real_1_tmp_3;
input 	result_real_1_tmp_2;
input 	result_real_1_tmp_1;
input 	result_real_1_tmp_0;
input 	result_real_1_tmp_15;
input 	result_real_1_tmp_14;
input 	result_real_1_tmp_13;
input 	result_real_1_tmp_12;
output 	pipeline_dffe_9;
output 	pipeline_dffe_8;
output 	pipeline_dffe_10;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~9_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~11_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~13_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~15_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~17_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~19_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~21_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~23_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~27 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~29 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~31 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~32_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~33 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~35 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~37 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~39 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~40_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~34_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~36_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~38_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~30_combout ;


dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_15),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_12),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_13),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_14),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .power_up = "low";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~9 (
	.dataa(result_real_1_tmp_15),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~9_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~9 .lut_mask = 16'h0055;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~11 (
	.dataa(result_real_1_tmp_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~9_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~11_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~11 .lut_mask = 16'h005F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~11 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~13 (
	.dataa(result_real_1_tmp_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~11_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~13_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~13 .lut_mask = 16'h00AF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~13 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~15 (
	.dataa(result_real_1_tmp_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~13_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~15_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~15 .lut_mask = 16'h005F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~15 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~17 (
	.dataa(result_real_1_tmp_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~15_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~17_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~17 .lut_mask = 16'h00AF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~17 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~19 (
	.dataa(result_real_1_tmp_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~17_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~19_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~19 .lut_mask = 16'h005F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~19 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~21 (
	.dataa(result_real_1_tmp_5),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~19_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~21_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~21 .lut_mask = 16'h00AF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~21 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~23 (
	.dataa(result_real_1_tmp_6),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~21_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~23_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~23 .lut_mask = 16'h005F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~23 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25 (
	.dataa(result_real_1_tmp_7),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~23_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25 .lut_mask = 16'h00AF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26 (
	.dataa(result_real_1_tmp_8),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25_cout ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~27 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28 (
	.dataa(result_real_1_tmp_9),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~27 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~29 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28 .lut_mask = 16'h5AAF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~30 (
	.dataa(result_real_1_tmp_10),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~29 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~30_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~31 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~30 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~30 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~32 (
	.dataa(result_real_1_tmp_11),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~31 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~32_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~33 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~32 .lut_mask = 16'h5AAF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~32 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~34 (
	.dataa(result_real_1_tmp_12),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~33 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~34_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~35 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~34 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~34 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~36 (
	.dataa(result_real_1_tmp_13),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~35 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~36_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~37 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~36 .lut_mask = 16'h5AAF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~36 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~38 (
	.dataa(result_real_1_tmp_14),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~37 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~38_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~39 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~38 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~38 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~40 (
	.dataa(result_real_1_tmp_15),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~39 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~40_combout ),
	.cout());
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~40 .lut_mask = 16'h5A5A;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~40 .sum_lutc_input = "cin";

endmodule

module fft_asj_fft_pround_fft_120_5 (
	pipeline_dffe_11,
	pipeline_dffe_15,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	result_imag_1_11,
	result_imag_1_10,
	result_imag_1_9,
	result_imag_1_8,
	result_imag_1_7,
	result_imag_1_6,
	result_imag_1_5,
	result_imag_1_4,
	result_imag_1_3,
	result_imag_1_2,
	result_imag_1_1,
	result_imag_1_0,
	result_imag_1_15,
	result_imag_1_14,
	result_imag_1_13,
	result_imag_1_12,
	pipeline_dffe_9,
	pipeline_dffe_8,
	pipeline_dffe_10,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_11;
output 	pipeline_dffe_15;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
input 	result_imag_1_11;
input 	result_imag_1_10;
input 	result_imag_1_9;
input 	result_imag_1_8;
input 	result_imag_1_7;
input 	result_imag_1_6;
input 	result_imag_1_5;
input 	result_imag_1_4;
input 	result_imag_1_3;
input 	result_imag_1_2;
input 	result_imag_1_1;
input 	result_imag_1_0;
input 	result_imag_1_15;
input 	result_imag_1_14;
input 	result_imag_1_13;
input 	result_imag_1_12;
output 	pipeline_dffe_9;
output 	pipeline_dffe_8;
output 	pipeline_dffe_10;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_LPM_ADD_SUB_6 \gbrnd:nev:gp:lpm_add_sub_component (
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_14(pipeline_dffe_14),
	.result_imag_1_11(result_imag_1_11),
	.result_imag_1_10(result_imag_1_10),
	.result_imag_1_9(result_imag_1_9),
	.result_imag_1_8(result_imag_1_8),
	.result_imag_1_7(result_imag_1_7),
	.result_imag_1_6(result_imag_1_6),
	.result_imag_1_5(result_imag_1_5),
	.result_imag_1_4(result_imag_1_4),
	.result_imag_1_3(result_imag_1_3),
	.result_imag_1_2(result_imag_1_2),
	.result_imag_1_1(result_imag_1_1),
	.result_imag_1_0(result_imag_1_0),
	.result_imag_1_15(result_imag_1_15),
	.result_imag_1_14(result_imag_1_14),
	.result_imag_1_13(result_imag_1_13),
	.result_imag_1_12(result_imag_1_12),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_10(pipeline_dffe_10),
	.clken(global_clock_enable),
	.clock(clk));

endmodule

module fft_LPM_ADD_SUB_6 (
	pipeline_dffe_11,
	pipeline_dffe_15,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	result_imag_1_11,
	result_imag_1_10,
	result_imag_1_9,
	result_imag_1_8,
	result_imag_1_7,
	result_imag_1_6,
	result_imag_1_5,
	result_imag_1_4,
	result_imag_1_3,
	result_imag_1_2,
	result_imag_1_1,
	result_imag_1_0,
	result_imag_1_15,
	result_imag_1_14,
	result_imag_1_13,
	result_imag_1_12,
	pipeline_dffe_9,
	pipeline_dffe_8,
	pipeline_dffe_10,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_11;
output 	pipeline_dffe_15;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
input 	result_imag_1_11;
input 	result_imag_1_10;
input 	result_imag_1_9;
input 	result_imag_1_8;
input 	result_imag_1_7;
input 	result_imag_1_6;
input 	result_imag_1_5;
input 	result_imag_1_4;
input 	result_imag_1_3;
input 	result_imag_1_2;
input 	result_imag_1_1;
input 	result_imag_1_0;
input 	result_imag_1_15;
input 	result_imag_1_14;
input 	result_imag_1_13;
input 	result_imag_1_12;
output 	pipeline_dffe_9;
output 	pipeline_dffe_8;
output 	pipeline_dffe_10;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_add_sub_dmj_5 auto_generated(
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_14(pipeline_dffe_14),
	.result_imag_1_11(result_imag_1_11),
	.result_imag_1_10(result_imag_1_10),
	.result_imag_1_9(result_imag_1_9),
	.result_imag_1_8(result_imag_1_8),
	.result_imag_1_7(result_imag_1_7),
	.result_imag_1_6(result_imag_1_6),
	.result_imag_1_5(result_imag_1_5),
	.result_imag_1_4(result_imag_1_4),
	.result_imag_1_3(result_imag_1_3),
	.result_imag_1_2(result_imag_1_2),
	.result_imag_1_1(result_imag_1_1),
	.result_imag_1_0(result_imag_1_0),
	.result_imag_1_15(result_imag_1_15),
	.result_imag_1_14(result_imag_1_14),
	.result_imag_1_13(result_imag_1_13),
	.result_imag_1_12(result_imag_1_12),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_10(pipeline_dffe_10),
	.clken(clken),
	.clock(clock));

endmodule

module fft_add_sub_dmj_5 (
	pipeline_dffe_11,
	pipeline_dffe_15,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	result_imag_1_11,
	result_imag_1_10,
	result_imag_1_9,
	result_imag_1_8,
	result_imag_1_7,
	result_imag_1_6,
	result_imag_1_5,
	result_imag_1_4,
	result_imag_1_3,
	result_imag_1_2,
	result_imag_1_1,
	result_imag_1_0,
	result_imag_1_15,
	result_imag_1_14,
	result_imag_1_13,
	result_imag_1_12,
	pipeline_dffe_9,
	pipeline_dffe_8,
	pipeline_dffe_10,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_11;
output 	pipeline_dffe_15;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
input 	result_imag_1_11;
input 	result_imag_1_10;
input 	result_imag_1_9;
input 	result_imag_1_8;
input 	result_imag_1_7;
input 	result_imag_1_6;
input 	result_imag_1_5;
input 	result_imag_1_4;
input 	result_imag_1_3;
input 	result_imag_1_2;
input 	result_imag_1_1;
input 	result_imag_1_0;
input 	result_imag_1_15;
input 	result_imag_1_14;
input 	result_imag_1_13;
input 	result_imag_1_12;
output 	pipeline_dffe_9;
output 	pipeline_dffe_8;
output 	pipeline_dffe_10;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~9_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~11_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~13_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~15_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~17_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~19_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~21_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~23_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~27 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~29 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~31 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~32_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~33 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~35 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~37 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~39 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~40_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~34_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~36_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~38_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~30_combout ;


dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_15),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_12),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_13),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_14),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .power_up = "low";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~9 (
	.dataa(result_imag_1_15),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~9_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~9 .lut_mask = 16'h0055;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~11 (
	.dataa(result_imag_1_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~9_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~11_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~11 .lut_mask = 16'h005F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~11 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~13 (
	.dataa(result_imag_1_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~11_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~13_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~13 .lut_mask = 16'h00AF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~13 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~15 (
	.dataa(result_imag_1_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~13_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~15_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~15 .lut_mask = 16'h005F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~15 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~17 (
	.dataa(result_imag_1_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~15_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~17_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~17 .lut_mask = 16'h00AF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~17 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~19 (
	.dataa(result_imag_1_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~17_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~19_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~19 .lut_mask = 16'h005F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~19 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~21 (
	.dataa(result_imag_1_5),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~19_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~21_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~21 .lut_mask = 16'h00AF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~21 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~23 (
	.dataa(result_imag_1_6),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~21_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~23_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~23 .lut_mask = 16'h005F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~23 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25 (
	.dataa(result_imag_1_7),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~23_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25 .lut_mask = 16'h00AF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26 (
	.dataa(result_imag_1_8),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25_cout ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~27 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28 (
	.dataa(result_imag_1_9),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~27 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~29 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28 .lut_mask = 16'h5AAF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~30 (
	.dataa(result_imag_1_10),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~29 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~30_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~31 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~30 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~30 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~32 (
	.dataa(result_imag_1_11),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~31 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~32_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~33 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~32 .lut_mask = 16'h5AAF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~32 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~34 (
	.dataa(result_imag_1_12),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~33 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~34_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~35 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~34 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~34 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~36 (
	.dataa(result_imag_1_13),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~35 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~36_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~37 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~36 .lut_mask = 16'h5AAF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~36 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~38 (
	.dataa(result_imag_1_14),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~37 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~38_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~39 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~38 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~38 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~40 (
	.dataa(result_imag_1_15),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~39 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~40_combout ),
	.cout());
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~40 .lut_mask = 16'h5A5A;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~40 .sum_lutc_input = "cin";

endmodule

module fft_LPM_MULT_7 (
	dataa,
	datab,
	clken,
	dffe3a_11,
	dffe3a_10,
	dffe3a_9,
	dffe3a_8,
	dffe3a_7,
	dffe3a_6,
	dffe3a_5,
	dffe3a_4,
	dffe3a_3,
	dffe3a_2,
	dffe3a_1,
	dffe3a_0,
	dffe3a_15,
	dffe3a_14,
	dffe3a_13,
	dffe3a_12,
	clock)/* synthesis synthesis_greybox=1 */;
input 	[8:0] dataa;
input 	[8:0] datab;
input 	clken;
output 	dffe3a_11;
output 	dffe3a_10;
output 	dffe3a_9;
output 	dffe3a_8;
output 	dffe3a_7;
output 	dffe3a_6;
output 	dffe3a_5;
output 	dffe3a_4;
output 	dffe3a_3;
output 	dffe3a_2;
output 	dffe3a_1;
output 	dffe3a_0;
output 	dffe3a_15;
output 	dffe3a_14;
output 	dffe3a_13;
output 	dffe3a_12;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_mult_4p01_2 auto_generated(
	.dataa({dataa[8],dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.datab({datab[8],datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.clken(clken),
	.dffe3a_11(dffe3a_11),
	.dffe3a_10(dffe3a_10),
	.dffe3a_9(dffe3a_9),
	.dffe3a_8(dffe3a_8),
	.dffe3a_7(dffe3a_7),
	.dffe3a_6(dffe3a_6),
	.dffe3a_5(dffe3a_5),
	.dffe3a_4(dffe3a_4),
	.dffe3a_3(dffe3a_3),
	.dffe3a_2(dffe3a_2),
	.dffe3a_1(dffe3a_1),
	.dffe3a_0(dffe3a_0),
	.dffe3a_15(dffe3a_15),
	.dffe3a_14(dffe3a_14),
	.dffe3a_13(dffe3a_13),
	.dffe3a_12(dffe3a_12),
	.clock(clock));

endmodule

module fft_mult_4p01_2 (
	dataa,
	datab,
	clken,
	dffe3a_11,
	dffe3a_10,
	dffe3a_9,
	dffe3a_8,
	dffe3a_7,
	dffe3a_6,
	dffe3a_5,
	dffe3a_4,
	dffe3a_3,
	dffe3a_2,
	dffe3a_1,
	dffe3a_0,
	dffe3a_15,
	dffe3a_14,
	dffe3a_13,
	dffe3a_12,
	clock)/* synthesis synthesis_greybox=1 */;
input 	[8:0] dataa;
input 	[8:0] datab;
input 	clken;
output 	dffe3a_11;
output 	dffe3a_10;
output 	dffe3a_9;
output 	dffe3a_8;
output 	dffe3a_7;
output 	dffe3a_6;
output 	dffe3a_5;
output 	dffe3a_4;
output 	dffe3a_3;
output 	dffe3a_2;
output 	dffe3a_1;
output 	dffe3a_0;
output 	dffe3a_15;
output 	dffe3a_14;
output 	dffe3a_13;
output 	dffe3a_12;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT16 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT17 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~dataout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT1 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT2 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT3 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT4 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT5 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT6 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT7 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT8 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT9 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT10 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT11 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT12 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT13 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT14 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT15 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT16 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT17 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT11 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT10 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT9 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT8 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT7 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT6 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT5 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT4 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT3 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT2 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT1 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~dataout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT15 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT14 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT13 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT12 ;

wire [35:0] \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus ;
wire [35:0] \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus ;

assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~dataout  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [0];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT1  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [1];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT2  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [2];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT3  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [3];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT4  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [4];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT5  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [5];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT6  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [6];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT7  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [7];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT8  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [8];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT9  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [9];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT10  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [10];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT11  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [11];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT12  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [12];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT13  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [13];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT14  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [14];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT15  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [15];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT16  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [16];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT17  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [17];

assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~dataout  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [0];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT1  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [1];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT2  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [2];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT3  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [3];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT4  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [4];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT5  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [5];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT6  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [6];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT7  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [7];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT8  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [8];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT9  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [9];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT10  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [10];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT11  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [11];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT12  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [12];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT13  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [13];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT14  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [14];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT15  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [15];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT16  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [16];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT17  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [17];

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[11] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT11 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_11),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[11] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[11] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[10] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT10 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_10),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[10] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[10] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[9] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT9 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_9),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[9] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[9] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[8] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT8 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_8),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[8] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[8] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[7] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT7 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_7),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[7] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[7] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[6] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT6 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_6),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[6] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[6] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[5] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT5 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_5),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[5] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[5] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[4] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT4 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_4),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[4] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[4] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[3] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT3 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_3),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[3] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[3] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[2] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT2 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_2),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[2] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[2] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[1] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT1 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_1),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[1] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[1] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[0] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~dataout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_0),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[0] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[0] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[15] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT15 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_15),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[15] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[15] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[14] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT14 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_14),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[14] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[14] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[13] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT13 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_13),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[13] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[13] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[12] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2~DATAOUT12 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_12),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[12] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|dffe3a[12] .power_up = "low";

cycloneiii_mac_mult \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1 (
	.signa(vcc),
	.signb(vcc),
	.clk(clock),
	.aclr(gnd),
	.ena(clken),
	.dataa({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dataa[8],dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.datab({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,datab[8],datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.dataout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1 .dataa_clock = "0";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1 .dataa_width = 9;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1 .datab_clock = "0";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1 .datab_width = 9;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1 .signa_clock = "none";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1 .signb_clock = "none";

cycloneiii_mac_out \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2 (
	.clk(clock),
	.aclr(gnd),
	.ena(clken),
	.dataa({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT17 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT16 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT15 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT14 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT13 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT12 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT11 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT10 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT9 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT8 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT7 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT6 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT5 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT4 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT3 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT2 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT1 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_mult1~dataout }),
	.dataout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2 .dataa_width = 18;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_a_b_c_d|auto_generated|mac_out2 .output_clock = "0";

endmodule

module fft_LPM_MULT_8 (
	dataa,
	clken,
	dffe3a_11,
	dffe3a_10,
	dffe3a_9,
	dffe3a_8,
	dffe3a_7,
	dffe3a_6,
	dffe3a_5,
	dffe3a_4,
	dffe3a_3,
	dffe3a_2,
	dffe3a_1,
	dffe3a_0,
	dffe3a_15,
	dffe3a_14,
	dffe3a_13,
	dffe3a_12,
	datab,
	clock)/* synthesis synthesis_greybox=1 */;
input 	[8:0] dataa;
input 	clken;
output 	dffe3a_11;
output 	dffe3a_10;
output 	dffe3a_9;
output 	dffe3a_8;
output 	dffe3a_7;
output 	dffe3a_6;
output 	dffe3a_5;
output 	dffe3a_4;
output 	dffe3a_3;
output 	dffe3a_2;
output 	dffe3a_1;
output 	dffe3a_0;
output 	dffe3a_15;
output 	dffe3a_14;
output 	dffe3a_13;
output 	dffe3a_12;
input 	[8:0] datab;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_mult_0p01_4 auto_generated(
	.dataa({dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.clken(clken),
	.dffe3a_11(dffe3a_11),
	.dffe3a_10(dffe3a_10),
	.dffe3a_9(dffe3a_9),
	.dffe3a_8(dffe3a_8),
	.dffe3a_7(dffe3a_7),
	.dffe3a_6(dffe3a_6),
	.dffe3a_5(dffe3a_5),
	.dffe3a_4(dffe3a_4),
	.dffe3a_3(dffe3a_3),
	.dffe3a_2(dffe3a_2),
	.dffe3a_1(dffe3a_1),
	.dffe3a_0(dffe3a_0),
	.dffe3a_15(dffe3a_15),
	.dffe3a_14(dffe3a_14),
	.dffe3a_13(dffe3a_13),
	.dffe3a_12(dffe3a_12),
	.datab({datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.clock(clock));

endmodule

module fft_mult_0p01_4 (
	dataa,
	clken,
	dffe3a_11,
	dffe3a_10,
	dffe3a_9,
	dffe3a_8,
	dffe3a_7,
	dffe3a_6,
	dffe3a_5,
	dffe3a_4,
	dffe3a_3,
	dffe3a_2,
	dffe3a_1,
	dffe3a_0,
	dffe3a_15,
	dffe3a_14,
	dffe3a_13,
	dffe3a_12,
	datab,
	clock)/* synthesis synthesis_greybox=1 */;
input 	[7:0] dataa;
input 	clken;
output 	dffe3a_11;
output 	dffe3a_10;
output 	dffe3a_9;
output 	dffe3a_8;
output 	dffe3a_7;
output 	dffe3a_6;
output 	dffe3a_5;
output 	dffe3a_4;
output 	dffe3a_3;
output 	dffe3a_2;
output 	dffe3a_1;
output 	dffe3a_0;
output 	dffe3a_15;
output 	dffe3a_14;
output 	dffe3a_13;
output 	dffe3a_12;
input 	[7:0] datab;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1~dataout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT1 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT2 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT3 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT4 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT5 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT6 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT7 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT8 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT9 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT10 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT11 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT12 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT13 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT14 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT15 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT11 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT10 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT9 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT8 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT7 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT6 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT5 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT4 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT3 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT2 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT1 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2~dataout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT15 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT14 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT13 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT12 ;

wire [35:0] \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2_DATAOUT_bus ;
wire [35:0] \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1_DATAOUT_bus ;

assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2~dataout  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2_DATAOUT_bus [0];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT1  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2_DATAOUT_bus [1];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT2  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2_DATAOUT_bus [2];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT3  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2_DATAOUT_bus [3];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT4  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2_DATAOUT_bus [4];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT5  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2_DATAOUT_bus [5];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT6  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2_DATAOUT_bus [6];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT7  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2_DATAOUT_bus [7];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT8  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2_DATAOUT_bus [8];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT9  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2_DATAOUT_bus [9];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT10  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2_DATAOUT_bus [10];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT11  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2_DATAOUT_bus [11];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT12  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2_DATAOUT_bus [12];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT13  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2_DATAOUT_bus [13];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT14  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2_DATAOUT_bus [14];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT15  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2_DATAOUT_bus [15];

assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1~dataout  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1_DATAOUT_bus [0];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT1  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1_DATAOUT_bus [1];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT2  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1_DATAOUT_bus [2];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT3  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1_DATAOUT_bus [3];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT4  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1_DATAOUT_bus [4];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT5  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1_DATAOUT_bus [5];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT6  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1_DATAOUT_bus [6];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT7  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1_DATAOUT_bus [7];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT8  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1_DATAOUT_bus [8];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT9  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1_DATAOUT_bus [9];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT10  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1_DATAOUT_bus [10];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT11  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1_DATAOUT_bus [11];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT12  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1_DATAOUT_bus [12];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT13  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1_DATAOUT_bus [13];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT14  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1_DATAOUT_bus [14];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT15  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1_DATAOUT_bus [15];

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|dffe3a[11] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT11 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_11),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|dffe3a[11] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|dffe3a[11] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|dffe3a[10] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT10 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_10),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|dffe3a[10] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|dffe3a[10] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|dffe3a[9] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT9 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_9),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|dffe3a[9] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|dffe3a[9] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|dffe3a[8] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT8 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_8),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|dffe3a[8] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|dffe3a[8] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|dffe3a[7] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT7 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_7),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|dffe3a[7] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|dffe3a[7] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|dffe3a[6] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT6 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_6),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|dffe3a[6] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|dffe3a[6] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|dffe3a[5] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT5 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_5),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|dffe3a[5] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|dffe3a[5] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|dffe3a[4] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT4 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_4),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|dffe3a[4] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|dffe3a[4] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|dffe3a[3] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT3 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_3),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|dffe3a[3] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|dffe3a[3] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|dffe3a[2] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT2 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_2),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|dffe3a[2] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|dffe3a[2] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|dffe3a[1] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT1 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_1),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|dffe3a[1] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|dffe3a[1] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|dffe3a[0] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2~dataout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_0),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|dffe3a[0] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|dffe3a[0] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|dffe3a[15] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT15 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_15),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|dffe3a[15] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|dffe3a[15] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|dffe3a[14] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT14 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_14),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|dffe3a[14] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|dffe3a[14] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|dffe3a[13] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT13 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_13),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|dffe3a[13] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|dffe3a[13] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|dffe3a[12] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2~DATAOUT12 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_12),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|dffe3a[12] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|dffe3a[12] .power_up = "low";

cycloneiii_mac_mult \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1 (
	.signa(vcc),
	.signb(vcc),
	.clk(clock),
	.aclr(gnd),
	.ena(clken),
	.dataa({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.datab({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.dataout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1_DATAOUT_bus ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1 .dataa_clock = "0";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1 .dataa_width = 8;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1 .datab_clock = "0";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1 .datab_width = 8;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1 .signa_clock = "none";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1 .signb_clock = "none";

cycloneiii_mac_out \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2 (
	.clk(clock),
	.aclr(gnd),
	.ena(clken),
	.dataa({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT15 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT14 ,\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT13 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT12 ,\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT11 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT10 ,\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT9 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT8 ,\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT7 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT6 ,\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT5 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT4 ,\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT3 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT2 ,\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1~DATAOUT1 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_mult1~dataout }),
	.dataout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2_DATAOUT_bus ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2 .dataa_width = 16;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_ac|auto_generated|mac_out2 .output_clock = "0";

endmodule

module fft_LPM_MULT_9 (
	dataa,
	clken,
	dffe3a_11,
	dffe3a_10,
	dffe3a_9,
	dffe3a_8,
	dffe3a_7,
	dffe3a_6,
	dffe3a_5,
	dffe3a_4,
	dffe3a_3,
	dffe3a_2,
	dffe3a_1,
	dffe3a_0,
	dffe3a_15,
	dffe3a_14,
	dffe3a_13,
	dffe3a_12,
	datab,
	clock)/* synthesis synthesis_greybox=1 */;
input 	[8:0] dataa;
input 	clken;
output 	dffe3a_11;
output 	dffe3a_10;
output 	dffe3a_9;
output 	dffe3a_8;
output 	dffe3a_7;
output 	dffe3a_6;
output 	dffe3a_5;
output 	dffe3a_4;
output 	dffe3a_3;
output 	dffe3a_2;
output 	dffe3a_1;
output 	dffe3a_0;
output 	dffe3a_15;
output 	dffe3a_14;
output 	dffe3a_13;
output 	dffe3a_12;
input 	[8:0] datab;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_mult_0p01_5 auto_generated(
	.dataa({dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.clken(clken),
	.dffe3a_11(dffe3a_11),
	.dffe3a_10(dffe3a_10),
	.dffe3a_9(dffe3a_9),
	.dffe3a_8(dffe3a_8),
	.dffe3a_7(dffe3a_7),
	.dffe3a_6(dffe3a_6),
	.dffe3a_5(dffe3a_5),
	.dffe3a_4(dffe3a_4),
	.dffe3a_3(dffe3a_3),
	.dffe3a_2(dffe3a_2),
	.dffe3a_1(dffe3a_1),
	.dffe3a_0(dffe3a_0),
	.dffe3a_15(dffe3a_15),
	.dffe3a_14(dffe3a_14),
	.dffe3a_13(dffe3a_13),
	.dffe3a_12(dffe3a_12),
	.datab({datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.clock(clock));

endmodule

module fft_mult_0p01_5 (
	dataa,
	clken,
	dffe3a_11,
	dffe3a_10,
	dffe3a_9,
	dffe3a_8,
	dffe3a_7,
	dffe3a_6,
	dffe3a_5,
	dffe3a_4,
	dffe3a_3,
	dffe3a_2,
	dffe3a_1,
	dffe3a_0,
	dffe3a_15,
	dffe3a_14,
	dffe3a_13,
	dffe3a_12,
	datab,
	clock)/* synthesis synthesis_greybox=1 */;
input 	[7:0] dataa;
input 	clken;
output 	dffe3a_11;
output 	dffe3a_10;
output 	dffe3a_9;
output 	dffe3a_8;
output 	dffe3a_7;
output 	dffe3a_6;
output 	dffe3a_5;
output 	dffe3a_4;
output 	dffe3a_3;
output 	dffe3a_2;
output 	dffe3a_1;
output 	dffe3a_0;
output 	dffe3a_15;
output 	dffe3a_14;
output 	dffe3a_13;
output 	dffe3a_12;
input 	[7:0] datab;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1~dataout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT1 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT2 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT3 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT4 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT5 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT6 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT7 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT8 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT9 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT10 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT11 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT12 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT13 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT14 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT15 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT11 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT10 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT9 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT8 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT7 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT6 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT5 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT4 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT3 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT2 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT1 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2~dataout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT15 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT14 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT13 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT12 ;

wire [35:0] \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2_DATAOUT_bus ;
wire [35:0] \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1_DATAOUT_bus ;

assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2~dataout  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2_DATAOUT_bus [0];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT1  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2_DATAOUT_bus [1];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT2  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2_DATAOUT_bus [2];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT3  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2_DATAOUT_bus [3];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT4  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2_DATAOUT_bus [4];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT5  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2_DATAOUT_bus [5];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT6  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2_DATAOUT_bus [6];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT7  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2_DATAOUT_bus [7];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT8  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2_DATAOUT_bus [8];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT9  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2_DATAOUT_bus [9];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT10  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2_DATAOUT_bus [10];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT11  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2_DATAOUT_bus [11];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT12  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2_DATAOUT_bus [12];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT13  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2_DATAOUT_bus [13];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT14  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2_DATAOUT_bus [14];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT15  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2_DATAOUT_bus [15];

assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1~dataout  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1_DATAOUT_bus [0];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT1  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1_DATAOUT_bus [1];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT2  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1_DATAOUT_bus [2];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT3  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1_DATAOUT_bus [3];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT4  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1_DATAOUT_bus [4];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT5  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1_DATAOUT_bus [5];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT6  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1_DATAOUT_bus [6];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT7  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1_DATAOUT_bus [7];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT8  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1_DATAOUT_bus [8];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT9  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1_DATAOUT_bus [9];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT10  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1_DATAOUT_bus [10];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT11  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1_DATAOUT_bus [11];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT12  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1_DATAOUT_bus [12];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT13  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1_DATAOUT_bus [13];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT14  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1_DATAOUT_bus [14];
assign \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT15  = \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1_DATAOUT_bus [15];

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|dffe3a[11] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT11 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_11),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|dffe3a[11] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|dffe3a[11] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|dffe3a[10] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT10 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_10),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|dffe3a[10] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|dffe3a[10] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|dffe3a[9] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT9 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_9),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|dffe3a[9] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|dffe3a[9] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|dffe3a[8] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT8 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_8),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|dffe3a[8] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|dffe3a[8] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|dffe3a[7] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT7 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_7),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|dffe3a[7] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|dffe3a[7] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|dffe3a[6] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT6 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_6),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|dffe3a[6] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|dffe3a[6] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|dffe3a[5] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT5 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_5),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|dffe3a[5] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|dffe3a[5] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|dffe3a[4] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT4 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_4),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|dffe3a[4] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|dffe3a[4] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|dffe3a[3] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT3 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_3),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|dffe3a[3] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|dffe3a[3] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|dffe3a[2] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT2 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_2),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|dffe3a[2] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|dffe3a[2] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|dffe3a[1] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT1 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_1),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|dffe3a[1] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|dffe3a[1] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|dffe3a[0] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2~dataout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_0),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|dffe3a[0] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|dffe3a[0] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|dffe3a[15] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT15 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_15),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|dffe3a[15] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|dffe3a[15] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|dffe3a[14] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT14 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_14),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|dffe3a[14] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|dffe3a[14] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|dffe3a[13] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT13 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_13),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|dffe3a[13] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|dffe3a[13] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|dffe3a[12] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2~DATAOUT12 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_12),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|dffe3a[12] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|dffe3a[12] .power_up = "low";

cycloneiii_mac_mult \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1 (
	.signa(vcc),
	.signb(vcc),
	.clk(clock),
	.aclr(gnd),
	.ena(clken),
	.dataa({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.datab({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.dataout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1_DATAOUT_bus ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1 .dataa_clock = "0";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1 .dataa_width = 8;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1 .datab_clock = "0";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1 .datab_width = 8;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1 .signa_clock = "none";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1 .signb_clock = "none";

cycloneiii_mac_out \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2 (
	.clk(clock),
	.aclr(gnd),
	.ena(clken),
	.dataa({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT15 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT14 ,\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT13 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT12 ,\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT11 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT10 ,\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT9 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT8 ,\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT7 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT6 ,\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT5 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT4 ,\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT3 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT2 ,\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1~DATAOUT1 ,
\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_mult1~dataout }),
	.dataout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2_DATAOUT_bus ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2 .dataa_width = 16;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_da0:gen_canonic:cm3|gen_dsp_only:m_bd|auto_generated|mac_out2 .output_clock = "0";

endmodule

module fft_asj_fft_pround_fft_120_6 (
	pipeline_dffe_6,
	pipeline_dffe_5,
	pipeline_dffe_4,
	pipeline_dffe_3,
	pipeline_dffe_2,
	pipeline_dffe_9,
	pipeline_dffe_8,
	pipeline_dffe_7,
	butterfly_st2006,
	butterfly_st2005,
	butterfly_st2004,
	butterfly_st2003,
	butterfly_st2002,
	butterfly_st2001,
	butterfly_st2000,
	butterfly_st2009,
	butterfly_st2008,
	butterfly_st2007,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_6;
output 	pipeline_dffe_5;
output 	pipeline_dffe_4;
output 	pipeline_dffe_3;
output 	pipeline_dffe_2;
output 	pipeline_dffe_9;
output 	pipeline_dffe_8;
output 	pipeline_dffe_7;
input 	butterfly_st2006;
input 	butterfly_st2005;
input 	butterfly_st2004;
input 	butterfly_st2003;
input 	butterfly_st2002;
input 	butterfly_st2001;
input 	butterfly_st2000;
input 	butterfly_st2009;
input 	butterfly_st2008;
input 	butterfly_st2007;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_LPM_ADD_SUB_7 \gbrnd:nev:gp:lpm_add_sub_component (
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_7(pipeline_dffe_7),
	.butterfly_st2006(butterfly_st2006),
	.butterfly_st2005(butterfly_st2005),
	.butterfly_st2004(butterfly_st2004),
	.butterfly_st2003(butterfly_st2003),
	.butterfly_st2002(butterfly_st2002),
	.butterfly_st2001(butterfly_st2001),
	.butterfly_st2000(butterfly_st2000),
	.butterfly_st2009(butterfly_st2009),
	.butterfly_st2008(butterfly_st2008),
	.butterfly_st2007(butterfly_st2007),
	.clken(global_clock_enable),
	.clock(clk));

endmodule

module fft_LPM_ADD_SUB_7 (
	pipeline_dffe_6,
	pipeline_dffe_5,
	pipeline_dffe_4,
	pipeline_dffe_3,
	pipeline_dffe_2,
	pipeline_dffe_9,
	pipeline_dffe_8,
	pipeline_dffe_7,
	butterfly_st2006,
	butterfly_st2005,
	butterfly_st2004,
	butterfly_st2003,
	butterfly_st2002,
	butterfly_st2001,
	butterfly_st2000,
	butterfly_st2009,
	butterfly_st2008,
	butterfly_st2007,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_6;
output 	pipeline_dffe_5;
output 	pipeline_dffe_4;
output 	pipeline_dffe_3;
output 	pipeline_dffe_2;
output 	pipeline_dffe_9;
output 	pipeline_dffe_8;
output 	pipeline_dffe_7;
input 	butterfly_st2006;
input 	butterfly_st2005;
input 	butterfly_st2004;
input 	butterfly_st2003;
input 	butterfly_st2002;
input 	butterfly_st2001;
input 	butterfly_st2000;
input 	butterfly_st2009;
input 	butterfly_st2008;
input 	butterfly_st2007;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_add_sub_7mj auto_generated(
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_7(pipeline_dffe_7),
	.butterfly_st2006(butterfly_st2006),
	.butterfly_st2005(butterfly_st2005),
	.butterfly_st2004(butterfly_st2004),
	.butterfly_st2003(butterfly_st2003),
	.butterfly_st2002(butterfly_st2002),
	.butterfly_st2001(butterfly_st2001),
	.butterfly_st2000(butterfly_st2000),
	.butterfly_st2009(butterfly_st2009),
	.butterfly_st2008(butterfly_st2008),
	.butterfly_st2007(butterfly_st2007),
	.clken(clken),
	.clock(clock));

endmodule

module fft_add_sub_7mj (
	pipeline_dffe_6,
	pipeline_dffe_5,
	pipeline_dffe_4,
	pipeline_dffe_3,
	pipeline_dffe_2,
	pipeline_dffe_9,
	pipeline_dffe_8,
	pipeline_dffe_7,
	butterfly_st2006,
	butterfly_st2005,
	butterfly_st2004,
	butterfly_st2003,
	butterfly_st2002,
	butterfly_st2001,
	butterfly_st2000,
	butterfly_st2009,
	butterfly_st2008,
	butterfly_st2007,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_6;
output 	pipeline_dffe_5;
output 	pipeline_dffe_4;
output 	pipeline_dffe_3;
output 	pipeline_dffe_2;
output 	pipeline_dffe_9;
output 	pipeline_dffe_8;
output 	pipeline_dffe_7;
input 	butterfly_st2006;
input 	butterfly_st2005;
input 	butterfly_st2004;
input 	butterfly_st2003;
input 	butterfly_st2002;
input 	butterfly_st2001;
input 	butterfly_st2000;
input 	butterfly_st2009;
input 	butterfly_st2008;
input 	butterfly_st2007;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~17 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~19 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~21 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~23 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~25 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~27 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24_combout ;


dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .power_up = "low";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9 (
	.dataa(butterfly_st2009),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9 .lut_mask = 16'h0055;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 (
	.dataa(butterfly_st2000),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 .lut_mask = 16'h005F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 (
	.dataa(butterfly_st2001),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 .lut_mask = 16'h00AF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14 (
	.dataa(butterfly_st2002),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16 (
	.dataa(butterfly_st2003),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~17 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16 .lut_mask = 16'h5AAF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18 (
	.dataa(butterfly_st2004),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~17 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~19 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20 (
	.dataa(butterfly_st2005),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~19 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~21 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20 .lut_mask = 16'h5AAF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22 (
	.dataa(butterfly_st2006),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~21 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~23 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24 (
	.dataa(butterfly_st2007),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~23 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~25 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24 .lut_mask = 16'h5AAF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26 (
	.dataa(butterfly_st2008),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~25 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~27 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28 (
	.dataa(butterfly_st2009),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~27 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28_combout ),
	.cout());
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28 .lut_mask = 16'h5A5A;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28 .sum_lutc_input = "cin";

endmodule

module fft_asj_fft_pround_fft_120_7 (
	pipeline_dffe_9,
	pipeline_dffe_8,
	pipeline_dffe_7,
	pipeline_dffe_6,
	pipeline_dffe_5,
	pipeline_dffe_4,
	pipeline_dffe_3,
	pipeline_dffe_2,
	butterfly_st2019,
	butterfly_st2018,
	butterfly_st2017,
	butterfly_st2016,
	butterfly_st2015,
	butterfly_st2014,
	butterfly_st2013,
	butterfly_st2012,
	butterfly_st2011,
	butterfly_st2010,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_9;
output 	pipeline_dffe_8;
output 	pipeline_dffe_7;
output 	pipeline_dffe_6;
output 	pipeline_dffe_5;
output 	pipeline_dffe_4;
output 	pipeline_dffe_3;
output 	pipeline_dffe_2;
input 	butterfly_st2019;
input 	butterfly_st2018;
input 	butterfly_st2017;
input 	butterfly_st2016;
input 	butterfly_st2015;
input 	butterfly_st2014;
input 	butterfly_st2013;
input 	butterfly_st2012;
input 	butterfly_st2011;
input 	butterfly_st2010;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_LPM_ADD_SUB_8 \gbrnd:nev:gp:lpm_add_sub_component (
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_2(pipeline_dffe_2),
	.butterfly_st2019(butterfly_st2019),
	.butterfly_st2018(butterfly_st2018),
	.butterfly_st2017(butterfly_st2017),
	.butterfly_st2016(butterfly_st2016),
	.butterfly_st2015(butterfly_st2015),
	.butterfly_st2014(butterfly_st2014),
	.butterfly_st2013(butterfly_st2013),
	.butterfly_st2012(butterfly_st2012),
	.butterfly_st2011(butterfly_st2011),
	.butterfly_st2010(butterfly_st2010),
	.clken(global_clock_enable),
	.clock(clk));

endmodule

module fft_LPM_ADD_SUB_8 (
	pipeline_dffe_9,
	pipeline_dffe_8,
	pipeline_dffe_7,
	pipeline_dffe_6,
	pipeline_dffe_5,
	pipeline_dffe_4,
	pipeline_dffe_3,
	pipeline_dffe_2,
	butterfly_st2019,
	butterfly_st2018,
	butterfly_st2017,
	butterfly_st2016,
	butterfly_st2015,
	butterfly_st2014,
	butterfly_st2013,
	butterfly_st2012,
	butterfly_st2011,
	butterfly_st2010,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_9;
output 	pipeline_dffe_8;
output 	pipeline_dffe_7;
output 	pipeline_dffe_6;
output 	pipeline_dffe_5;
output 	pipeline_dffe_4;
output 	pipeline_dffe_3;
output 	pipeline_dffe_2;
input 	butterfly_st2019;
input 	butterfly_st2018;
input 	butterfly_st2017;
input 	butterfly_st2016;
input 	butterfly_st2015;
input 	butterfly_st2014;
input 	butterfly_st2013;
input 	butterfly_st2012;
input 	butterfly_st2011;
input 	butterfly_st2010;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_add_sub_7mj_1 auto_generated(
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_2(pipeline_dffe_2),
	.butterfly_st2019(butterfly_st2019),
	.butterfly_st2018(butterfly_st2018),
	.butterfly_st2017(butterfly_st2017),
	.butterfly_st2016(butterfly_st2016),
	.butterfly_st2015(butterfly_st2015),
	.butterfly_st2014(butterfly_st2014),
	.butterfly_st2013(butterfly_st2013),
	.butterfly_st2012(butterfly_st2012),
	.butterfly_st2011(butterfly_st2011),
	.butterfly_st2010(butterfly_st2010),
	.clken(clken),
	.clock(clock));

endmodule

module fft_add_sub_7mj_1 (
	pipeline_dffe_9,
	pipeline_dffe_8,
	pipeline_dffe_7,
	pipeline_dffe_6,
	pipeline_dffe_5,
	pipeline_dffe_4,
	pipeline_dffe_3,
	pipeline_dffe_2,
	butterfly_st2019,
	butterfly_st2018,
	butterfly_st2017,
	butterfly_st2016,
	butterfly_st2015,
	butterfly_st2014,
	butterfly_st2013,
	butterfly_st2012,
	butterfly_st2011,
	butterfly_st2010,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_9;
output 	pipeline_dffe_8;
output 	pipeline_dffe_7;
output 	pipeline_dffe_6;
output 	pipeline_dffe_5;
output 	pipeline_dffe_4;
output 	pipeline_dffe_3;
output 	pipeline_dffe_2;
input 	butterfly_st2019;
input 	butterfly_st2018;
input 	butterfly_st2017;
input 	butterfly_st2016;
input 	butterfly_st2015;
input 	butterfly_st2014;
input 	butterfly_st2013;
input 	butterfly_st2012;
input 	butterfly_st2011;
input 	butterfly_st2010;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~17 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~19 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~21 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~23 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~25 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~27 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14_combout ;


dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .power_up = "low";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9 (
	.dataa(butterfly_st2019),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9 .lut_mask = 16'h0055;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 (
	.dataa(butterfly_st2010),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 .lut_mask = 16'h005F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 (
	.dataa(butterfly_st2011),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 .lut_mask = 16'h00AF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14 (
	.dataa(butterfly_st2012),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16 (
	.dataa(butterfly_st2013),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~17 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16 .lut_mask = 16'h5AAF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18 (
	.dataa(butterfly_st2014),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~17 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~19 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20 (
	.dataa(butterfly_st2015),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~19 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~21 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20 .lut_mask = 16'h5AAF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22 (
	.dataa(butterfly_st2016),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~21 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~23 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24 (
	.dataa(butterfly_st2017),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~23 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~25 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24 .lut_mask = 16'h5AAF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26 (
	.dataa(butterfly_st2018),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~25 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~27 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28 (
	.dataa(butterfly_st2019),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~27 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28_combout ),
	.cout());
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28 .lut_mask = 16'h5A5A;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28 .sum_lutc_input = "cin";

endmodule

module fft_asj_fft_pround_fft_120_8 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	butterfly_st2102,
	butterfly_st2101,
	butterfly_st2100,
	butterfly_st2109,
	butterfly_st2103,
	butterfly_st2104,
	butterfly_st2105,
	butterfly_st2106,
	butterfly_st2107,
	butterfly_st2108,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	butterfly_st2102;
input 	butterfly_st2101;
input 	butterfly_st2100;
input 	butterfly_st2109;
input 	butterfly_st2103;
input 	butterfly_st2104;
input 	butterfly_st2105;
input 	butterfly_st2106;
input 	butterfly_st2107;
input 	butterfly_st2108;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_LPM_ADD_SUB_9 \gbrnd:nev:gp:lpm_add_sub_component (
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.butterfly_st2102(butterfly_st2102),
	.butterfly_st2101(butterfly_st2101),
	.butterfly_st2100(butterfly_st2100),
	.butterfly_st2109(butterfly_st2109),
	.butterfly_st2103(butterfly_st2103),
	.butterfly_st2104(butterfly_st2104),
	.butterfly_st2105(butterfly_st2105),
	.butterfly_st2106(butterfly_st2106),
	.butterfly_st2107(butterfly_st2107),
	.butterfly_st2108(butterfly_st2108),
	.clken(global_clock_enable),
	.clock(clk));

endmodule

module fft_LPM_ADD_SUB_9 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	butterfly_st2102,
	butterfly_st2101,
	butterfly_st2100,
	butterfly_st2109,
	butterfly_st2103,
	butterfly_st2104,
	butterfly_st2105,
	butterfly_st2106,
	butterfly_st2107,
	butterfly_st2108,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	butterfly_st2102;
input 	butterfly_st2101;
input 	butterfly_st2100;
input 	butterfly_st2109;
input 	butterfly_st2103;
input 	butterfly_st2104;
input 	butterfly_st2105;
input 	butterfly_st2106;
input 	butterfly_st2107;
input 	butterfly_st2108;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_add_sub_7mj_2 auto_generated(
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.butterfly_st2102(butterfly_st2102),
	.butterfly_st2101(butterfly_st2101),
	.butterfly_st2100(butterfly_st2100),
	.butterfly_st2109(butterfly_st2109),
	.butterfly_st2103(butterfly_st2103),
	.butterfly_st2104(butterfly_st2104),
	.butterfly_st2105(butterfly_st2105),
	.butterfly_st2106(butterfly_st2106),
	.butterfly_st2107(butterfly_st2107),
	.butterfly_st2108(butterfly_st2108),
	.clken(clken),
	.clock(clock));

endmodule

module fft_add_sub_7mj_2 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	butterfly_st2102,
	butterfly_st2101,
	butterfly_st2100,
	butterfly_st2109,
	butterfly_st2103,
	butterfly_st2104,
	butterfly_st2105,
	butterfly_st2106,
	butterfly_st2107,
	butterfly_st2108,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	butterfly_st2102;
input 	butterfly_st2101;
input 	butterfly_st2100;
input 	butterfly_st2109;
input 	butterfly_st2103;
input 	butterfly_st2104;
input 	butterfly_st2105;
input 	butterfly_st2106;
input 	butterfly_st2107;
input 	butterfly_st2108;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~17 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~19 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~21 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~23 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~25 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~27 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28_combout ;


dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .power_up = "low";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9 (
	.dataa(butterfly_st2109),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9 .lut_mask = 16'h0055;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 (
	.dataa(butterfly_st2100),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 .lut_mask = 16'h005F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 (
	.dataa(butterfly_st2101),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 .lut_mask = 16'h00AF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14 (
	.dataa(butterfly_st2102),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16 (
	.dataa(butterfly_st2103),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~17 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16 .lut_mask = 16'h5AAF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18 (
	.dataa(butterfly_st2104),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~17 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~19 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20 (
	.dataa(butterfly_st2105),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~19 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~21 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20 .lut_mask = 16'h5AAF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22 (
	.dataa(butterfly_st2106),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~21 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~23 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24 (
	.dataa(butterfly_st2107),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~23 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~25 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24 .lut_mask = 16'h5AAF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26 (
	.dataa(butterfly_st2108),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~25 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~27 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28 (
	.dataa(butterfly_st2109),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~27 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28_combout ),
	.cout());
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28 .lut_mask = 16'h5A5A;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28 .sum_lutc_input = "cin";

endmodule

module fft_asj_fft_pround_fft_120_9 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	butterfly_st2112,
	butterfly_st2111,
	butterfly_st2110,
	butterfly_st2119,
	butterfly_st2113,
	butterfly_st2114,
	butterfly_st2115,
	butterfly_st2116,
	butterfly_st2117,
	butterfly_st2118,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	butterfly_st2112;
input 	butterfly_st2111;
input 	butterfly_st2110;
input 	butterfly_st2119;
input 	butterfly_st2113;
input 	butterfly_st2114;
input 	butterfly_st2115;
input 	butterfly_st2116;
input 	butterfly_st2117;
input 	butterfly_st2118;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_LPM_ADD_SUB_10 \gbrnd:nev:gp:lpm_add_sub_component (
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.butterfly_st2112(butterfly_st2112),
	.butterfly_st2111(butterfly_st2111),
	.butterfly_st2110(butterfly_st2110),
	.butterfly_st2119(butterfly_st2119),
	.butterfly_st2113(butterfly_st2113),
	.butterfly_st2114(butterfly_st2114),
	.butterfly_st2115(butterfly_st2115),
	.butterfly_st2116(butterfly_st2116),
	.butterfly_st2117(butterfly_st2117),
	.butterfly_st2118(butterfly_st2118),
	.clken(global_clock_enable),
	.clock(clk));

endmodule

module fft_LPM_ADD_SUB_10 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	butterfly_st2112,
	butterfly_st2111,
	butterfly_st2110,
	butterfly_st2119,
	butterfly_st2113,
	butterfly_st2114,
	butterfly_st2115,
	butterfly_st2116,
	butterfly_st2117,
	butterfly_st2118,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	butterfly_st2112;
input 	butterfly_st2111;
input 	butterfly_st2110;
input 	butterfly_st2119;
input 	butterfly_st2113;
input 	butterfly_st2114;
input 	butterfly_st2115;
input 	butterfly_st2116;
input 	butterfly_st2117;
input 	butterfly_st2118;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_add_sub_7mj_3 auto_generated(
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.butterfly_st2112(butterfly_st2112),
	.butterfly_st2111(butterfly_st2111),
	.butterfly_st2110(butterfly_st2110),
	.butterfly_st2119(butterfly_st2119),
	.butterfly_st2113(butterfly_st2113),
	.butterfly_st2114(butterfly_st2114),
	.butterfly_st2115(butterfly_st2115),
	.butterfly_st2116(butterfly_st2116),
	.butterfly_st2117(butterfly_st2117),
	.butterfly_st2118(butterfly_st2118),
	.clken(clken),
	.clock(clock));

endmodule

module fft_add_sub_7mj_3 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	butterfly_st2112,
	butterfly_st2111,
	butterfly_st2110,
	butterfly_st2119,
	butterfly_st2113,
	butterfly_st2114,
	butterfly_st2115,
	butterfly_st2116,
	butterfly_st2117,
	butterfly_st2118,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	butterfly_st2112;
input 	butterfly_st2111;
input 	butterfly_st2110;
input 	butterfly_st2119;
input 	butterfly_st2113;
input 	butterfly_st2114;
input 	butterfly_st2115;
input 	butterfly_st2116;
input 	butterfly_st2117;
input 	butterfly_st2118;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~17 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~19 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~21 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~23 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~25 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~27 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28_combout ;


dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .power_up = "low";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9 (
	.dataa(butterfly_st2119),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9 .lut_mask = 16'h0055;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 (
	.dataa(butterfly_st2110),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 .lut_mask = 16'h005F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 (
	.dataa(butterfly_st2111),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 .lut_mask = 16'h00AF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14 (
	.dataa(butterfly_st2112),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16 (
	.dataa(butterfly_st2113),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~17 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16 .lut_mask = 16'h5AAF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18 (
	.dataa(butterfly_st2114),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~17 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~19 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20 (
	.dataa(butterfly_st2115),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~19 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~21 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20 .lut_mask = 16'h5AAF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22 (
	.dataa(butterfly_st2116),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~21 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~23 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24 (
	.dataa(butterfly_st2117),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~23 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~25 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24 .lut_mask = 16'h5AAF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26 (
	.dataa(butterfly_st2118),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~25 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~27 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28 (
	.dataa(butterfly_st2119),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~27 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28_combout ),
	.cout());
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28 .lut_mask = 16'h5A5A;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28 .sum_lutc_input = "cin";

endmodule

module fft_asj_fft_pround_fft_120_10 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	butterfly_st2202,
	butterfly_st2201,
	butterfly_st2200,
	butterfly_st2209,
	butterfly_st2203,
	butterfly_st2204,
	butterfly_st2205,
	butterfly_st2206,
	butterfly_st2207,
	butterfly_st2208,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	butterfly_st2202;
input 	butterfly_st2201;
input 	butterfly_st2200;
input 	butterfly_st2209;
input 	butterfly_st2203;
input 	butterfly_st2204;
input 	butterfly_st2205;
input 	butterfly_st2206;
input 	butterfly_st2207;
input 	butterfly_st2208;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_LPM_ADD_SUB_11 \gbrnd:nev:gp:lpm_add_sub_component (
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.butterfly_st2202(butterfly_st2202),
	.butterfly_st2201(butterfly_st2201),
	.butterfly_st2200(butterfly_st2200),
	.butterfly_st2209(butterfly_st2209),
	.butterfly_st2203(butterfly_st2203),
	.butterfly_st2204(butterfly_st2204),
	.butterfly_st2205(butterfly_st2205),
	.butterfly_st2206(butterfly_st2206),
	.butterfly_st2207(butterfly_st2207),
	.butterfly_st2208(butterfly_st2208),
	.clken(global_clock_enable),
	.clock(clk));

endmodule

module fft_LPM_ADD_SUB_11 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	butterfly_st2202,
	butterfly_st2201,
	butterfly_st2200,
	butterfly_st2209,
	butterfly_st2203,
	butterfly_st2204,
	butterfly_st2205,
	butterfly_st2206,
	butterfly_st2207,
	butterfly_st2208,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	butterfly_st2202;
input 	butterfly_st2201;
input 	butterfly_st2200;
input 	butterfly_st2209;
input 	butterfly_st2203;
input 	butterfly_st2204;
input 	butterfly_st2205;
input 	butterfly_st2206;
input 	butterfly_st2207;
input 	butterfly_st2208;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_add_sub_7mj_4 auto_generated(
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.butterfly_st2202(butterfly_st2202),
	.butterfly_st2201(butterfly_st2201),
	.butterfly_st2200(butterfly_st2200),
	.butterfly_st2209(butterfly_st2209),
	.butterfly_st2203(butterfly_st2203),
	.butterfly_st2204(butterfly_st2204),
	.butterfly_st2205(butterfly_st2205),
	.butterfly_st2206(butterfly_st2206),
	.butterfly_st2207(butterfly_st2207),
	.butterfly_st2208(butterfly_st2208),
	.clken(clken),
	.clock(clock));

endmodule

module fft_add_sub_7mj_4 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	butterfly_st2202,
	butterfly_st2201,
	butterfly_st2200,
	butterfly_st2209,
	butterfly_st2203,
	butterfly_st2204,
	butterfly_st2205,
	butterfly_st2206,
	butterfly_st2207,
	butterfly_st2208,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	butterfly_st2202;
input 	butterfly_st2201;
input 	butterfly_st2200;
input 	butterfly_st2209;
input 	butterfly_st2203;
input 	butterfly_st2204;
input 	butterfly_st2205;
input 	butterfly_st2206;
input 	butterfly_st2207;
input 	butterfly_st2208;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~17 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~19 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~21 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~23 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~25 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~27 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28_combout ;


dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .power_up = "low";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9 (
	.dataa(butterfly_st2209),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9 .lut_mask = 16'h0055;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 (
	.dataa(butterfly_st2200),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 .lut_mask = 16'h005F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 (
	.dataa(butterfly_st2201),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 .lut_mask = 16'h00AF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14 (
	.dataa(butterfly_st2202),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16 (
	.dataa(butterfly_st2203),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~17 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16 .lut_mask = 16'h5AAF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18 (
	.dataa(butterfly_st2204),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~17 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~19 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20 (
	.dataa(butterfly_st2205),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~19 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~21 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20 .lut_mask = 16'h5AAF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22 (
	.dataa(butterfly_st2206),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~21 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~23 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24 (
	.dataa(butterfly_st2207),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~23 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~25 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24 .lut_mask = 16'h5AAF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26 (
	.dataa(butterfly_st2208),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~25 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~27 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28 (
	.dataa(butterfly_st2209),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~27 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28_combout ),
	.cout());
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28 .lut_mask = 16'h5A5A;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28 .sum_lutc_input = "cin";

endmodule

module fft_asj_fft_pround_fft_120_11 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	butterfly_st2212,
	butterfly_st2211,
	butterfly_st2210,
	butterfly_st2219,
	butterfly_st2213,
	butterfly_st2214,
	butterfly_st2215,
	butterfly_st2216,
	butterfly_st2217,
	butterfly_st2218,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	butterfly_st2212;
input 	butterfly_st2211;
input 	butterfly_st2210;
input 	butterfly_st2219;
input 	butterfly_st2213;
input 	butterfly_st2214;
input 	butterfly_st2215;
input 	butterfly_st2216;
input 	butterfly_st2217;
input 	butterfly_st2218;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_LPM_ADD_SUB_12 \gbrnd:nev:gp:lpm_add_sub_component (
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.butterfly_st2212(butterfly_st2212),
	.butterfly_st2211(butterfly_st2211),
	.butterfly_st2210(butterfly_st2210),
	.butterfly_st2219(butterfly_st2219),
	.butterfly_st2213(butterfly_st2213),
	.butterfly_st2214(butterfly_st2214),
	.butterfly_st2215(butterfly_st2215),
	.butterfly_st2216(butterfly_st2216),
	.butterfly_st2217(butterfly_st2217),
	.butterfly_st2218(butterfly_st2218),
	.clken(global_clock_enable),
	.clock(clk));

endmodule

module fft_LPM_ADD_SUB_12 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	butterfly_st2212,
	butterfly_st2211,
	butterfly_st2210,
	butterfly_st2219,
	butterfly_st2213,
	butterfly_st2214,
	butterfly_st2215,
	butterfly_st2216,
	butterfly_st2217,
	butterfly_st2218,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	butterfly_st2212;
input 	butterfly_st2211;
input 	butterfly_st2210;
input 	butterfly_st2219;
input 	butterfly_st2213;
input 	butterfly_st2214;
input 	butterfly_st2215;
input 	butterfly_st2216;
input 	butterfly_st2217;
input 	butterfly_st2218;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_add_sub_7mj_5 auto_generated(
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.butterfly_st2212(butterfly_st2212),
	.butterfly_st2211(butterfly_st2211),
	.butterfly_st2210(butterfly_st2210),
	.butterfly_st2219(butterfly_st2219),
	.butterfly_st2213(butterfly_st2213),
	.butterfly_st2214(butterfly_st2214),
	.butterfly_st2215(butterfly_st2215),
	.butterfly_st2216(butterfly_st2216),
	.butterfly_st2217(butterfly_st2217),
	.butterfly_st2218(butterfly_st2218),
	.clken(clken),
	.clock(clock));

endmodule

module fft_add_sub_7mj_5 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	butterfly_st2212,
	butterfly_st2211,
	butterfly_st2210,
	butterfly_st2219,
	butterfly_st2213,
	butterfly_st2214,
	butterfly_st2215,
	butterfly_st2216,
	butterfly_st2217,
	butterfly_st2218,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	butterfly_st2212;
input 	butterfly_st2211;
input 	butterfly_st2210;
input 	butterfly_st2219;
input 	butterfly_st2213;
input 	butterfly_st2214;
input 	butterfly_st2215;
input 	butterfly_st2216;
input 	butterfly_st2217;
input 	butterfly_st2218;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~17 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~19 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~21 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~23 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~25 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~27 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28_combout ;


dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .power_up = "low";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9 (
	.dataa(butterfly_st2219),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9 .lut_mask = 16'h0055;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 (
	.dataa(butterfly_st2210),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 .lut_mask = 16'h005F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 (
	.dataa(butterfly_st2211),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 .lut_mask = 16'h00AF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14 (
	.dataa(butterfly_st2212),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16 (
	.dataa(butterfly_st2213),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~17 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16 .lut_mask = 16'h5AAF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18 (
	.dataa(butterfly_st2214),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~17 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~19 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20 (
	.dataa(butterfly_st2215),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~19 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~21 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20 .lut_mask = 16'h5AAF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22 (
	.dataa(butterfly_st2216),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~21 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~23 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24 (
	.dataa(butterfly_st2217),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~23 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~25 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24 .lut_mask = 16'h5AAF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26 (
	.dataa(butterfly_st2218),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~25 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~27 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28 (
	.dataa(butterfly_st2219),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~27 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28_combout ),
	.cout());
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28 .lut_mask = 16'h5A5A;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28 .sum_lutc_input = "cin";

endmodule

module fft_asj_fft_pround_fft_120_12 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	butterfly_st2302,
	butterfly_st2301,
	butterfly_st2300,
	butterfly_st2309,
	butterfly_st2303,
	butterfly_st2304,
	butterfly_st2305,
	butterfly_st2306,
	butterfly_st2307,
	butterfly_st2308,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	butterfly_st2302;
input 	butterfly_st2301;
input 	butterfly_st2300;
input 	butterfly_st2309;
input 	butterfly_st2303;
input 	butterfly_st2304;
input 	butterfly_st2305;
input 	butterfly_st2306;
input 	butterfly_st2307;
input 	butterfly_st2308;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_LPM_ADD_SUB_13 \gbrnd:nev:gp:lpm_add_sub_component (
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.butterfly_st2302(butterfly_st2302),
	.butterfly_st2301(butterfly_st2301),
	.butterfly_st2300(butterfly_st2300),
	.butterfly_st2309(butterfly_st2309),
	.butterfly_st2303(butterfly_st2303),
	.butterfly_st2304(butterfly_st2304),
	.butterfly_st2305(butterfly_st2305),
	.butterfly_st2306(butterfly_st2306),
	.butterfly_st2307(butterfly_st2307),
	.butterfly_st2308(butterfly_st2308),
	.clken(global_clock_enable),
	.clock(clk));

endmodule

module fft_LPM_ADD_SUB_13 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	butterfly_st2302,
	butterfly_st2301,
	butterfly_st2300,
	butterfly_st2309,
	butterfly_st2303,
	butterfly_st2304,
	butterfly_st2305,
	butterfly_st2306,
	butterfly_st2307,
	butterfly_st2308,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	butterfly_st2302;
input 	butterfly_st2301;
input 	butterfly_st2300;
input 	butterfly_st2309;
input 	butterfly_st2303;
input 	butterfly_st2304;
input 	butterfly_st2305;
input 	butterfly_st2306;
input 	butterfly_st2307;
input 	butterfly_st2308;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_add_sub_7mj_6 auto_generated(
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.butterfly_st2302(butterfly_st2302),
	.butterfly_st2301(butterfly_st2301),
	.butterfly_st2300(butterfly_st2300),
	.butterfly_st2309(butterfly_st2309),
	.butterfly_st2303(butterfly_st2303),
	.butterfly_st2304(butterfly_st2304),
	.butterfly_st2305(butterfly_st2305),
	.butterfly_st2306(butterfly_st2306),
	.butterfly_st2307(butterfly_st2307),
	.butterfly_st2308(butterfly_st2308),
	.clken(clken),
	.clock(clock));

endmodule

module fft_add_sub_7mj_6 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	butterfly_st2302,
	butterfly_st2301,
	butterfly_st2300,
	butterfly_st2309,
	butterfly_st2303,
	butterfly_st2304,
	butterfly_st2305,
	butterfly_st2306,
	butterfly_st2307,
	butterfly_st2308,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	butterfly_st2302;
input 	butterfly_st2301;
input 	butterfly_st2300;
input 	butterfly_st2309;
input 	butterfly_st2303;
input 	butterfly_st2304;
input 	butterfly_st2305;
input 	butterfly_st2306;
input 	butterfly_st2307;
input 	butterfly_st2308;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~17 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~19 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~21 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~23 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~25 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~27 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28_combout ;


dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .power_up = "low";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9 (
	.dataa(butterfly_st2309),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9 .lut_mask = 16'h0055;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 (
	.dataa(butterfly_st2300),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 .lut_mask = 16'h005F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 (
	.dataa(butterfly_st2301),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 .lut_mask = 16'h00AF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14 (
	.dataa(butterfly_st2302),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16 (
	.dataa(butterfly_st2303),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~17 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16 .lut_mask = 16'h5AAF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18 (
	.dataa(butterfly_st2304),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~17 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~19 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20 (
	.dataa(butterfly_st2305),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~19 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~21 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20 .lut_mask = 16'h5AAF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22 (
	.dataa(butterfly_st2306),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~21 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~23 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24 (
	.dataa(butterfly_st2307),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~23 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~25 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24 .lut_mask = 16'h5AAF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26 (
	.dataa(butterfly_st2308),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~25 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~27 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28 (
	.dataa(butterfly_st2309),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~27 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28_combout ),
	.cout());
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28 .lut_mask = 16'h5A5A;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28 .sum_lutc_input = "cin";

endmodule

module fft_asj_fft_pround_fft_120_13 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	butterfly_st2312,
	butterfly_st2311,
	butterfly_st2310,
	butterfly_st2319,
	butterfly_st2313,
	butterfly_st2314,
	butterfly_st2315,
	butterfly_st2316,
	butterfly_st2317,
	butterfly_st2318,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	butterfly_st2312;
input 	butterfly_st2311;
input 	butterfly_st2310;
input 	butterfly_st2319;
input 	butterfly_st2313;
input 	butterfly_st2314;
input 	butterfly_st2315;
input 	butterfly_st2316;
input 	butterfly_st2317;
input 	butterfly_st2318;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_LPM_ADD_SUB_14 \gbrnd:nev:gp:lpm_add_sub_component (
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.butterfly_st2312(butterfly_st2312),
	.butterfly_st2311(butterfly_st2311),
	.butterfly_st2310(butterfly_st2310),
	.butterfly_st2319(butterfly_st2319),
	.butterfly_st2313(butterfly_st2313),
	.butterfly_st2314(butterfly_st2314),
	.butterfly_st2315(butterfly_st2315),
	.butterfly_st2316(butterfly_st2316),
	.butterfly_st2317(butterfly_st2317),
	.butterfly_st2318(butterfly_st2318),
	.clken(global_clock_enable),
	.clock(clk));

endmodule

module fft_LPM_ADD_SUB_14 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	butterfly_st2312,
	butterfly_st2311,
	butterfly_st2310,
	butterfly_st2319,
	butterfly_st2313,
	butterfly_st2314,
	butterfly_st2315,
	butterfly_st2316,
	butterfly_st2317,
	butterfly_st2318,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	butterfly_st2312;
input 	butterfly_st2311;
input 	butterfly_st2310;
input 	butterfly_st2319;
input 	butterfly_st2313;
input 	butterfly_st2314;
input 	butterfly_st2315;
input 	butterfly_st2316;
input 	butterfly_st2317;
input 	butterfly_st2318;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_add_sub_7mj_7 auto_generated(
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.butterfly_st2312(butterfly_st2312),
	.butterfly_st2311(butterfly_st2311),
	.butterfly_st2310(butterfly_st2310),
	.butterfly_st2319(butterfly_st2319),
	.butterfly_st2313(butterfly_st2313),
	.butterfly_st2314(butterfly_st2314),
	.butterfly_st2315(butterfly_st2315),
	.butterfly_st2316(butterfly_st2316),
	.butterfly_st2317(butterfly_st2317),
	.butterfly_st2318(butterfly_st2318),
	.clken(clken),
	.clock(clock));

endmodule

module fft_add_sub_7mj_7 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	butterfly_st2312,
	butterfly_st2311,
	butterfly_st2310,
	butterfly_st2319,
	butterfly_st2313,
	butterfly_st2314,
	butterfly_st2315,
	butterfly_st2316,
	butterfly_st2317,
	butterfly_st2318,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	butterfly_st2312;
input 	butterfly_st2311;
input 	butterfly_st2310;
input 	butterfly_st2319;
input 	butterfly_st2313;
input 	butterfly_st2314;
input 	butterfly_st2315;
input 	butterfly_st2316;
input 	butterfly_st2317;
input 	butterfly_st2318;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~17 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~19 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~21 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~23 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~25 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~27 ;
wire \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28_combout ;


dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .power_up = "low";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9 (
	.dataa(butterfly_st2319),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9 .lut_mask = 16'h0055;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 (
	.dataa(butterfly_st2310),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 .lut_mask = 16'h005F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 (
	.dataa(butterfly_st2311),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 .lut_mask = 16'h00AF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14 (
	.dataa(butterfly_st2312),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16 (
	.dataa(butterfly_st2313),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~17 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16 .lut_mask = 16'h5AAF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18 (
	.dataa(butterfly_st2314),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~17 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~19 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20 (
	.dataa(butterfly_st2315),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~19 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~21 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20 .lut_mask = 16'h5AAF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22 (
	.dataa(butterfly_st2316),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~21 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~23 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24 (
	.dataa(butterfly_st2317),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~23 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~25 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24 .lut_mask = 16'h5AAF;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26 (
	.dataa(butterfly_st2318),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~25 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~27 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28 (
	.dataa(butterfly_st2319),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~27 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28_combout ),
	.cout());
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28 .lut_mask = 16'h5A5A;
defparam \asj_fft_sglstream_fft_120_inst|gen_dft_2:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28 .sum_lutc_input = "cin";

endmodule

module fft_asj_fft_tdl_bit_fft_120_2 (
	global_clock_enable,
	data_in,
	tdl_arr_4,
	tdl_arr_3,
	tdl_arr_22,
	tdl_arr_25,
	clk)/* synthesis synthesis_greybox=1 */;
input 	global_clock_enable;
input 	data_in;
output 	tdl_arr_4;
output 	tdl_arr_3;
output 	tdl_arr_22;
output 	tdl_arr_25;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \tdl_arr[0]~q ;
wire \tdl_arr[1]~q ;
wire \tdl_arr[2]~q ;
wire \tdl_arr[5]~q ;
wire \tdl_arr[6]~q ;
wire \tdl_arr[7]~q ;
wire \tdl_arr[8]~q ;
wire \tdl_arr[9]~q ;
wire \tdl_arr[10]~q ;
wire \tdl_arr[11]~q ;
wire \tdl_arr[12]~q ;
wire \tdl_arr[13]~q ;
wire \tdl_arr[14]~q ;
wire \tdl_arr[15]~q ;
wire \tdl_arr[16]~q ;
wire \tdl_arr[17]~q ;
wire \tdl_arr[18]~q ;
wire \tdl_arr[19]~q ;
wire \tdl_arr[20]~q ;
wire \tdl_arr[21]~q ;
wire \tdl_arr[23]~q ;
wire \tdl_arr[24]~q ;


dffeas \tdl_arr[4] (
	.clk(clk),
	.d(tdl_arr_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_4),
	.prn(vcc));
defparam \tdl_arr[4] .is_wysiwyg = "true";
defparam \tdl_arr[4] .power_up = "low";

dffeas \tdl_arr[3] (
	.clk(clk),
	.d(\tdl_arr[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_3),
	.prn(vcc));
defparam \tdl_arr[3] .is_wysiwyg = "true";
defparam \tdl_arr[3] .power_up = "low";

dffeas \tdl_arr[22] (
	.clk(clk),
	.d(\tdl_arr[21]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_22),
	.prn(vcc));
defparam \tdl_arr[22] .is_wysiwyg = "true";
defparam \tdl_arr[22] .power_up = "low";

dffeas \tdl_arr[25] (
	.clk(clk),
	.d(\tdl_arr[24]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_25),
	.prn(vcc));
defparam \tdl_arr[25] .is_wysiwyg = "true";
defparam \tdl_arr[25] .power_up = "low";

dffeas \tdl_arr[0] (
	.clk(clk),
	.d(data_in),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0]~q ),
	.prn(vcc));
defparam \tdl_arr[0] .is_wysiwyg = "true";
defparam \tdl_arr[0] .power_up = "low";

dffeas \tdl_arr[1] (
	.clk(clk),
	.d(\tdl_arr[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[1]~q ),
	.prn(vcc));
defparam \tdl_arr[1] .is_wysiwyg = "true";
defparam \tdl_arr[1] .power_up = "low";

dffeas \tdl_arr[2] (
	.clk(clk),
	.d(\tdl_arr[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[2]~q ),
	.prn(vcc));
defparam \tdl_arr[2] .is_wysiwyg = "true";
defparam \tdl_arr[2] .power_up = "low";

dffeas \tdl_arr[5] (
	.clk(clk),
	.d(tdl_arr_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[5]~q ),
	.prn(vcc));
defparam \tdl_arr[5] .is_wysiwyg = "true";
defparam \tdl_arr[5] .power_up = "low";

dffeas \tdl_arr[6] (
	.clk(clk),
	.d(\tdl_arr[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[6]~q ),
	.prn(vcc));
defparam \tdl_arr[6] .is_wysiwyg = "true";
defparam \tdl_arr[6] .power_up = "low";

dffeas \tdl_arr[7] (
	.clk(clk),
	.d(\tdl_arr[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[7]~q ),
	.prn(vcc));
defparam \tdl_arr[7] .is_wysiwyg = "true";
defparam \tdl_arr[7] .power_up = "low";

dffeas \tdl_arr[8] (
	.clk(clk),
	.d(\tdl_arr[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[8]~q ),
	.prn(vcc));
defparam \tdl_arr[8] .is_wysiwyg = "true";
defparam \tdl_arr[8] .power_up = "low";

dffeas \tdl_arr[9] (
	.clk(clk),
	.d(\tdl_arr[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[9]~q ),
	.prn(vcc));
defparam \tdl_arr[9] .is_wysiwyg = "true";
defparam \tdl_arr[9] .power_up = "low";

dffeas \tdl_arr[10] (
	.clk(clk),
	.d(\tdl_arr[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[10]~q ),
	.prn(vcc));
defparam \tdl_arr[10] .is_wysiwyg = "true";
defparam \tdl_arr[10] .power_up = "low";

dffeas \tdl_arr[11] (
	.clk(clk),
	.d(\tdl_arr[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[11]~q ),
	.prn(vcc));
defparam \tdl_arr[11] .is_wysiwyg = "true";
defparam \tdl_arr[11] .power_up = "low";

dffeas \tdl_arr[12] (
	.clk(clk),
	.d(\tdl_arr[11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[12]~q ),
	.prn(vcc));
defparam \tdl_arr[12] .is_wysiwyg = "true";
defparam \tdl_arr[12] .power_up = "low";

dffeas \tdl_arr[13] (
	.clk(clk),
	.d(\tdl_arr[12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[13]~q ),
	.prn(vcc));
defparam \tdl_arr[13] .is_wysiwyg = "true";
defparam \tdl_arr[13] .power_up = "low";

dffeas \tdl_arr[14] (
	.clk(clk),
	.d(\tdl_arr[13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[14]~q ),
	.prn(vcc));
defparam \tdl_arr[14] .is_wysiwyg = "true";
defparam \tdl_arr[14] .power_up = "low";

dffeas \tdl_arr[15] (
	.clk(clk),
	.d(\tdl_arr[14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[15]~q ),
	.prn(vcc));
defparam \tdl_arr[15] .is_wysiwyg = "true";
defparam \tdl_arr[15] .power_up = "low";

dffeas \tdl_arr[16] (
	.clk(clk),
	.d(\tdl_arr[15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[16]~q ),
	.prn(vcc));
defparam \tdl_arr[16] .is_wysiwyg = "true";
defparam \tdl_arr[16] .power_up = "low";

dffeas \tdl_arr[17] (
	.clk(clk),
	.d(\tdl_arr[16]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[17]~q ),
	.prn(vcc));
defparam \tdl_arr[17] .is_wysiwyg = "true";
defparam \tdl_arr[17] .power_up = "low";

dffeas \tdl_arr[18] (
	.clk(clk),
	.d(\tdl_arr[17]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[18]~q ),
	.prn(vcc));
defparam \tdl_arr[18] .is_wysiwyg = "true";
defparam \tdl_arr[18] .power_up = "low";

dffeas \tdl_arr[19] (
	.clk(clk),
	.d(\tdl_arr[18]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[19]~q ),
	.prn(vcc));
defparam \tdl_arr[19] .is_wysiwyg = "true";
defparam \tdl_arr[19] .power_up = "low";

dffeas \tdl_arr[20] (
	.clk(clk),
	.d(\tdl_arr[19]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[20]~q ),
	.prn(vcc));
defparam \tdl_arr[20] .is_wysiwyg = "true";
defparam \tdl_arr[20] .power_up = "low";

dffeas \tdl_arr[21] (
	.clk(clk),
	.d(\tdl_arr[20]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[21]~q ),
	.prn(vcc));
defparam \tdl_arr[21] .is_wysiwyg = "true";
defparam \tdl_arr[21] .power_up = "low";

dffeas \tdl_arr[23] (
	.clk(clk),
	.d(tdl_arr_22),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[23]~q ),
	.prn(vcc));
defparam \tdl_arr[23] .is_wysiwyg = "true";
defparam \tdl_arr[23] .power_up = "low";

dffeas \tdl_arr[24] (
	.clk(clk),
	.d(\tdl_arr[23]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[24]~q ),
	.prn(vcc));
defparam \tdl_arr[24] .is_wysiwyg = "true";
defparam \tdl_arr[24] .power_up = "low";

endmodule

module fft_asj_fft_in_write_sgl_fft_120 (
	data_rdy_int1,
	wren_0,
	wren_1,
	wren_2,
	wren_3,
	core_real_in_2,
	core_real_in_6,
	core_real_in_4,
	core_real_in_3,
	core_real_in_5,
	core_real_in_1,
	core_real_in_0,
	core_real_in_7,
	core_imag_in_7,
	core_imag_in_3,
	core_imag_in_5,
	core_imag_in_4,
	core_imag_in_6,
	core_imag_in_2,
	core_imag_in_1,
	core_imag_in_0,
	anb1,
	send_sop_s,
	global_clock_enable,
	next_block1,
	data_in_r_2,
	wr_address_i_int_0,
	wr_address_i_int_1,
	wr_address_i_int_2,
	wr_address_i_int_3,
	wr_address_i_int_4,
	wr_address_i_int_5,
	wr_address_i_int_6,
	data_in_r_6,
	data_in_r_4,
	data_in_r_3,
	data_in_r_5,
	data_in_r_1,
	data_in_r_0,
	data_in_r_7,
	data_in_i_7,
	data_in_i_3,
	data_in_i_5,
	data_in_i_4,
	data_in_i_6,
	data_in_i_2,
	data_in_i_1,
	data_in_i_0,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	data_rdy_int1;
output 	wren_0;
output 	wren_1;
output 	wren_2;
output 	wren_3;
input 	core_real_in_2;
input 	core_real_in_6;
input 	core_real_in_4;
input 	core_real_in_3;
input 	core_real_in_5;
input 	core_real_in_1;
input 	core_real_in_0;
input 	core_real_in_7;
input 	core_imag_in_7;
input 	core_imag_in_3;
input 	core_imag_in_5;
input 	core_imag_in_4;
input 	core_imag_in_6;
input 	core_imag_in_2;
input 	core_imag_in_1;
input 	core_imag_in_0;
output 	anb1;
input 	send_sop_s;
input 	global_clock_enable;
output 	next_block1;
output 	data_in_r_2;
output 	wr_address_i_int_0;
output 	wr_address_i_int_1;
output 	wr_address_i_int_2;
output 	wr_address_i_int_3;
output 	wr_address_i_int_4;
output 	wr_address_i_int_5;
output 	wr_address_i_int_6;
output 	data_in_r_6;
output 	data_in_r_4;
output 	data_in_r_3;
output 	data_in_r_5;
output 	data_in_r_1;
output 	data_in_r_0;
output 	data_in_r_7;
output 	data_in_i_7;
output 	data_in_i_3;
output 	data_in_i_5;
output 	data_in_i_4;
output 	data_in_i_6;
output 	data_in_i_2;
output 	data_in_i_1;
output 	data_in_i_0;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \str_count_en~q ;
wire \Equal0~2_combout ;
wire \str_count_en~0_combout ;
wire \count[0]~9_combout ;
wire \counter_i~0_combout ;
wire \count[0]~q ;
wire \count[0]~10 ;
wire \count[1]~12 ;
wire \count[2]~14 ;
wire \count[3]~16 ;
wire \count[4]~18 ;
wire \count[5]~20 ;
wire \count[6]~22 ;
wire \count[7]~23_combout ;
wire \count[7]~q ;
wire \count[2]~13_combout ;
wire \count[2]~q ;
wire \Equal0~0_combout ;
wire \count[7]~24 ;
wire \count[8]~25_combout ;
wire \count[8]~q ;
wire \count[4]~17_combout ;
wire \count[4]~q ;
wire \count[5]~19_combout ;
wire \count[5]~q ;
wire \count[6]~21_combout ;
wire \count[6]~q ;
wire \Equal0~1_combout ;
wire \data_rdy_int~0_combout ;
wire \count[1]~11_combout ;
wire \count[1]~q ;
wire \Add2~0_combout ;
wire \sw[0]~q ;
wire \Add2~1_combout ;
wire \Add2~2_combout ;
wire \sw[1]~q ;
wire \Mux3~0_combout ;
wire \Mux1~0_combout ;
wire \Mux1~1_combout ;
wire \Mux1~2_combout ;
wire \anb~0_combout ;
wire \next_block~0_combout ;
wire \data_in_r~0_combout ;
wire \wr_addr[0]~q ;
wire \wr_address_i_int~0_combout ;
wire \wr_addr[1]~q ;
wire \wr_address_i_int~1_combout ;
wire \count[3]~15_combout ;
wire \count[3]~q ;
wire \wr_addr[2]~q ;
wire \wr_address_i_int~2_combout ;
wire \wr_addr[3]~q ;
wire \wr_address_i_int~3_combout ;
wire \wr_addr[4]~q ;
wire \wr_address_i_int~4_combout ;
wire \wr_addr[5]~q ;
wire \wr_address_i_int~5_combout ;
wire \wr_addr[6]~q ;
wire \wr_address_i_int~6_combout ;
wire \data_in_r~1_combout ;
wire \data_in_r~2_combout ;
wire \data_in_r~3_combout ;
wire \data_in_r~4_combout ;
wire \data_in_r~5_combout ;
wire \data_in_r~6_combout ;
wire \data_in_r~7_combout ;
wire \data_in_i~0_combout ;
wire \data_in_i~1_combout ;
wire \data_in_i~2_combout ;
wire \data_in_i~3_combout ;
wire \data_in_i~4_combout ;
wire \data_in_i~5_combout ;
wire \data_in_i~6_combout ;
wire \data_in_i~7_combout ;


dffeas str_count_en(
	.clk(clk),
	.d(\str_count_en~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\str_count_en~q ),
	.prn(vcc));
defparam str_count_en.is_wysiwyg = "true";
defparam str_count_en.power_up = "low";

cycloneiii_lcell_comb \Equal0~2 (
	.dataa(\Equal0~0_combout ),
	.datab(\count[8]~q ),
	.datac(\Equal0~1_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Equal0~2_combout ),
	.cout());
defparam \Equal0~2 .lut_mask = 16'hFEFE;
defparam \Equal0~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \str_count_en~0 (
	.dataa(send_sop_s),
	.datab(\str_count_en~q ),
	.datac(gnd),
	.datad(\Equal0~2_combout ),
	.cin(gnd),
	.combout(\str_count_en~0_combout ),
	.cout());
defparam \str_count_en~0 .lut_mask = 16'hEEFF;
defparam \str_count_en~0 .sum_lutc_input = "datac";

dffeas data_rdy_int(
	.clk(clk),
	.d(\data_rdy_int~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_rdy_int1),
	.prn(vcc));
defparam data_rdy_int.is_wysiwyg = "true";
defparam data_rdy_int.power_up = "low";

dffeas \wren[0] (
	.clk(clk),
	.d(\Mux3~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wren_0),
	.prn(vcc));
defparam \wren[0] .is_wysiwyg = "true";
defparam \wren[0] .power_up = "low";

dffeas \wren[1] (
	.clk(clk),
	.d(\Mux1~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wren_1),
	.prn(vcc));
defparam \wren[1] .is_wysiwyg = "true";
defparam \wren[1] .power_up = "low";

dffeas \wren[2] (
	.clk(clk),
	.d(\Mux1~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wren_2),
	.prn(vcc));
defparam \wren[2] .is_wysiwyg = "true";
defparam \wren[2] .power_up = "low";

dffeas \wren[3] (
	.clk(clk),
	.d(\Mux1~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wren_3),
	.prn(vcc));
defparam \wren[3] .is_wysiwyg = "true";
defparam \wren[3] .power_up = "low";

dffeas anb(
	.clk(clk),
	.d(\anb~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(global_clock_enable),
	.q(anb1),
	.prn(vcc));
defparam anb.is_wysiwyg = "true";
defparam anb.power_up = "low";

dffeas next_block(
	.clk(clk),
	.d(\next_block~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(next_block1),
	.prn(vcc));
defparam next_block.is_wysiwyg = "true";
defparam next_block.power_up = "low";

dffeas \data_in_r[2] (
	.clk(clk),
	.d(\data_in_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_r_2),
	.prn(vcc));
defparam \data_in_r[2] .is_wysiwyg = "true";
defparam \data_in_r[2] .power_up = "low";

dffeas \wr_address_i_int[0] (
	.clk(clk),
	.d(\wr_address_i_int~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wr_address_i_int_0),
	.prn(vcc));
defparam \wr_address_i_int[0] .is_wysiwyg = "true";
defparam \wr_address_i_int[0] .power_up = "low";

dffeas \wr_address_i_int[1] (
	.clk(clk),
	.d(\wr_address_i_int~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wr_address_i_int_1),
	.prn(vcc));
defparam \wr_address_i_int[1] .is_wysiwyg = "true";
defparam \wr_address_i_int[1] .power_up = "low";

dffeas \wr_address_i_int[2] (
	.clk(clk),
	.d(\wr_address_i_int~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wr_address_i_int_2),
	.prn(vcc));
defparam \wr_address_i_int[2] .is_wysiwyg = "true";
defparam \wr_address_i_int[2] .power_up = "low";

dffeas \wr_address_i_int[3] (
	.clk(clk),
	.d(\wr_address_i_int~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wr_address_i_int_3),
	.prn(vcc));
defparam \wr_address_i_int[3] .is_wysiwyg = "true";
defparam \wr_address_i_int[3] .power_up = "low";

dffeas \wr_address_i_int[4] (
	.clk(clk),
	.d(\wr_address_i_int~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wr_address_i_int_4),
	.prn(vcc));
defparam \wr_address_i_int[4] .is_wysiwyg = "true";
defparam \wr_address_i_int[4] .power_up = "low";

dffeas \wr_address_i_int[5] (
	.clk(clk),
	.d(\wr_address_i_int~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wr_address_i_int_5),
	.prn(vcc));
defparam \wr_address_i_int[5] .is_wysiwyg = "true";
defparam \wr_address_i_int[5] .power_up = "low";

dffeas \wr_address_i_int[6] (
	.clk(clk),
	.d(\wr_address_i_int~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wr_address_i_int_6),
	.prn(vcc));
defparam \wr_address_i_int[6] .is_wysiwyg = "true";
defparam \wr_address_i_int[6] .power_up = "low";

dffeas \data_in_r[6] (
	.clk(clk),
	.d(\data_in_r~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_r_6),
	.prn(vcc));
defparam \data_in_r[6] .is_wysiwyg = "true";
defparam \data_in_r[6] .power_up = "low";

dffeas \data_in_r[4] (
	.clk(clk),
	.d(\data_in_r~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_r_4),
	.prn(vcc));
defparam \data_in_r[4] .is_wysiwyg = "true";
defparam \data_in_r[4] .power_up = "low";

dffeas \data_in_r[3] (
	.clk(clk),
	.d(\data_in_r~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_r_3),
	.prn(vcc));
defparam \data_in_r[3] .is_wysiwyg = "true";
defparam \data_in_r[3] .power_up = "low";

dffeas \data_in_r[5] (
	.clk(clk),
	.d(\data_in_r~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_r_5),
	.prn(vcc));
defparam \data_in_r[5] .is_wysiwyg = "true";
defparam \data_in_r[5] .power_up = "low";

dffeas \data_in_r[1] (
	.clk(clk),
	.d(\data_in_r~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_r_1),
	.prn(vcc));
defparam \data_in_r[1] .is_wysiwyg = "true";
defparam \data_in_r[1] .power_up = "low";

dffeas \data_in_r[0] (
	.clk(clk),
	.d(\data_in_r~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_r_0),
	.prn(vcc));
defparam \data_in_r[0] .is_wysiwyg = "true";
defparam \data_in_r[0] .power_up = "low";

dffeas \data_in_r[7] (
	.clk(clk),
	.d(\data_in_r~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_r_7),
	.prn(vcc));
defparam \data_in_r[7] .is_wysiwyg = "true";
defparam \data_in_r[7] .power_up = "low";

dffeas \data_in_i[7] (
	.clk(clk),
	.d(\data_in_i~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_i_7),
	.prn(vcc));
defparam \data_in_i[7] .is_wysiwyg = "true";
defparam \data_in_i[7] .power_up = "low";

dffeas \data_in_i[3] (
	.clk(clk),
	.d(\data_in_i~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_i_3),
	.prn(vcc));
defparam \data_in_i[3] .is_wysiwyg = "true";
defparam \data_in_i[3] .power_up = "low";

dffeas \data_in_i[5] (
	.clk(clk),
	.d(\data_in_i~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_i_5),
	.prn(vcc));
defparam \data_in_i[5] .is_wysiwyg = "true";
defparam \data_in_i[5] .power_up = "low";

dffeas \data_in_i[4] (
	.clk(clk),
	.d(\data_in_i~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_i_4),
	.prn(vcc));
defparam \data_in_i[4] .is_wysiwyg = "true";
defparam \data_in_i[4] .power_up = "low";

dffeas \data_in_i[6] (
	.clk(clk),
	.d(\data_in_i~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_i_6),
	.prn(vcc));
defparam \data_in_i[6] .is_wysiwyg = "true";
defparam \data_in_i[6] .power_up = "low";

dffeas \data_in_i[2] (
	.clk(clk),
	.d(\data_in_i~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_i_2),
	.prn(vcc));
defparam \data_in_i[2] .is_wysiwyg = "true";
defparam \data_in_i[2] .power_up = "low";

dffeas \data_in_i[1] (
	.clk(clk),
	.d(\data_in_i~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_i_1),
	.prn(vcc));
defparam \data_in_i[1] .is_wysiwyg = "true";
defparam \data_in_i[1] .power_up = "low";

dffeas \data_in_i[0] (
	.clk(clk),
	.d(\data_in_i~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_i_0),
	.prn(vcc));
defparam \data_in_i[0] .is_wysiwyg = "true";
defparam \data_in_i[0] .power_up = "low";

cycloneiii_lcell_comb \count[0]~9 (
	.dataa(\str_count_en~q ),
	.datab(\count[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\count[0]~9_combout ),
	.cout(\count[0]~10 ));
defparam \count[0]~9 .lut_mask = 16'h66EE;
defparam \count[0]~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \counter_i~0 (
	.dataa(send_sop_s),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\counter_i~0_combout ),
	.cout());
defparam \counter_i~0 .lut_mask = 16'hAAFF;
defparam \counter_i~0 .sum_lutc_input = "datac";

dffeas \count[0] (
	.clk(clk),
	.d(\count[0]~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\counter_i~0_combout ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\count[0]~q ),
	.prn(vcc));
defparam \count[0] .is_wysiwyg = "true";
defparam \count[0] .power_up = "low";

cycloneiii_lcell_comb \count[1]~11 (
	.dataa(\count[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[0]~10 ),
	.combout(\count[1]~11_combout ),
	.cout(\count[1]~12 ));
defparam \count[1]~11 .lut_mask = 16'h5A5F;
defparam \count[1]~11 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \count[2]~13 (
	.dataa(\count[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[1]~12 ),
	.combout(\count[2]~13_combout ),
	.cout(\count[2]~14 ));
defparam \count[2]~13 .lut_mask = 16'h5AAF;
defparam \count[2]~13 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \count[3]~15 (
	.dataa(\count[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[2]~14 ),
	.combout(\count[3]~15_combout ),
	.cout(\count[3]~16 ));
defparam \count[3]~15 .lut_mask = 16'h5A5F;
defparam \count[3]~15 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \count[4]~17 (
	.dataa(\count[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[3]~16 ),
	.combout(\count[4]~17_combout ),
	.cout(\count[4]~18 ));
defparam \count[4]~17 .lut_mask = 16'h5AAF;
defparam \count[4]~17 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \count[5]~19 (
	.dataa(\count[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[4]~18 ),
	.combout(\count[5]~19_combout ),
	.cout(\count[5]~20 ));
defparam \count[5]~19 .lut_mask = 16'h5A5F;
defparam \count[5]~19 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \count[6]~21 (
	.dataa(\count[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[5]~20 ),
	.combout(\count[6]~21_combout ),
	.cout(\count[6]~22 ));
defparam \count[6]~21 .lut_mask = 16'h5AAF;
defparam \count[6]~21 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \count[7]~23 (
	.dataa(\count[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[6]~22 ),
	.combout(\count[7]~23_combout ),
	.cout(\count[7]~24 ));
defparam \count[7]~23 .lut_mask = 16'h5A5F;
defparam \count[7]~23 .sum_lutc_input = "cin";

dffeas \count[7] (
	.clk(clk),
	.d(\count[7]~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\counter_i~0_combout ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\count[7]~q ),
	.prn(vcc));
defparam \count[7] .is_wysiwyg = "true";
defparam \count[7] .power_up = "low";

dffeas \count[2] (
	.clk(clk),
	.d(\count[2]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\counter_i~0_combout ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\count[2]~q ),
	.prn(vcc));
defparam \count[2] .is_wysiwyg = "true";
defparam \count[2] .power_up = "low";

cycloneiii_lcell_comb \Equal0~0 (
	.dataa(\count[1]~q ),
	.datab(\count[7]~q ),
	.datac(\count[0]~q ),
	.datad(\count[2]~q ),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
defparam \Equal0~0 .lut_mask = 16'hFFFE;
defparam \Equal0~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \count[8]~25 (
	.dataa(\count[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\count[7]~24 ),
	.combout(\count[8]~25_combout ),
	.cout());
defparam \count[8]~25 .lut_mask = 16'h5A5A;
defparam \count[8]~25 .sum_lutc_input = "cin";

dffeas \count[8] (
	.clk(clk),
	.d(\count[8]~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\counter_i~0_combout ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\count[8]~q ),
	.prn(vcc));
defparam \count[8] .is_wysiwyg = "true";
defparam \count[8] .power_up = "low";

dffeas \count[4] (
	.clk(clk),
	.d(\count[4]~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\counter_i~0_combout ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\count[4]~q ),
	.prn(vcc));
defparam \count[4] .is_wysiwyg = "true";
defparam \count[4] .power_up = "low";

dffeas \count[5] (
	.clk(clk),
	.d(\count[5]~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\counter_i~0_combout ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\count[5]~q ),
	.prn(vcc));
defparam \count[5] .is_wysiwyg = "true";
defparam \count[5] .power_up = "low";

dffeas \count[6] (
	.clk(clk),
	.d(\count[6]~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\counter_i~0_combout ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\count[6]~q ),
	.prn(vcc));
defparam \count[6] .is_wysiwyg = "true";
defparam \count[6] .power_up = "low";

cycloneiii_lcell_comb \Equal0~1 (
	.dataa(\count[3]~q ),
	.datab(\count[4]~q ),
	.datac(\count[5]~q ),
	.datad(\count[6]~q ),
	.cin(gnd),
	.combout(\Equal0~1_combout ),
	.cout());
defparam \Equal0~1 .lut_mask = 16'hFFFE;
defparam \Equal0~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \data_rdy_int~0 (
	.dataa(data_rdy_int1),
	.datab(\Equal0~0_combout ),
	.datac(\count[8]~q ),
	.datad(\Equal0~1_combout ),
	.cin(gnd),
	.combout(\data_rdy_int~0_combout ),
	.cout());
defparam \data_rdy_int~0 .lut_mask = 16'hFFFE;
defparam \data_rdy_int~0 .sum_lutc_input = "datac";

dffeas \count[1] (
	.clk(clk),
	.d(\count[1]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\counter_i~0_combout ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\count[1]~q ),
	.prn(vcc));
defparam \count[1] .is_wysiwyg = "true";
defparam \count[1] .power_up = "low";

cycloneiii_lcell_comb \Add2~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\count[1]~q ),
	.datad(\count[7]~q ),
	.cin(gnd),
	.combout(\Add2~0_combout ),
	.cout());
defparam \Add2~0 .lut_mask = 16'h0FF0;
defparam \Add2~0 .sum_lutc_input = "datac";

dffeas \sw[0] (
	.clk(clk),
	.d(\Add2~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sw[0]~q ),
	.prn(vcc));
defparam \sw[0] .is_wysiwyg = "true";
defparam \sw[0] .power_up = "low";

cycloneiii_lcell_comb \Add2~1 (
	.dataa(\count[1]~q ),
	.datab(\count[7]~q ),
	.datac(\count[0]~q ),
	.datad(\count[2]~q ),
	.cin(gnd),
	.combout(\Add2~1_combout ),
	.cout());
defparam \Add2~1 .lut_mask = 16'h6996;
defparam \Add2~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add2~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\count[8]~q ),
	.datad(\Add2~1_combout ),
	.cin(gnd),
	.combout(\Add2~2_combout ),
	.cout());
defparam \Add2~2 .lut_mask = 16'h0FF0;
defparam \Add2~2 .sum_lutc_input = "datac";

dffeas \sw[1] (
	.clk(clk),
	.d(\Add2~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sw[1]~q ),
	.prn(vcc));
defparam \sw[1] .is_wysiwyg = "true";
defparam \sw[1] .power_up = "low";

cycloneiii_lcell_comb \Mux3~0 (
	.dataa(\sw[0]~q ),
	.datab(\sw[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux3~0_combout ),
	.cout());
defparam \Mux3~0 .lut_mask = 16'h7777;
defparam \Mux3~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux1~0 (
	.dataa(\sw[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\sw[1]~q ),
	.cin(gnd),
	.combout(\Mux1~0_combout ),
	.cout());
defparam \Mux1~0 .lut_mask = 16'hAAFF;
defparam \Mux1~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux1~1 (
	.dataa(\sw[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\sw[0]~q ),
	.cin(gnd),
	.combout(\Mux1~1_combout ),
	.cout());
defparam \Mux1~1 .lut_mask = 16'hAAFF;
defparam \Mux1~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux1~2 (
	.dataa(\sw[0]~q ),
	.datab(\sw[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux1~2_combout ),
	.cout());
defparam \Mux1~2 .lut_mask = 16'hEEEE;
defparam \Mux1~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \anb~0 (
	.dataa(anb1),
	.datab(\Equal0~0_combout ),
	.datac(\count[8]~q ),
	.datad(\Equal0~1_combout ),
	.cin(gnd),
	.combout(\anb~0_combout ),
	.cout());
defparam \anb~0 .lut_mask = 16'h6996;
defparam \anb~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \next_block~0 (
	.dataa(reset_n),
	.datab(\Equal0~0_combout ),
	.datac(\count[8]~q ),
	.datad(\Equal0~1_combout ),
	.cin(gnd),
	.combout(\next_block~0_combout ),
	.cout());
defparam \next_block~0 .lut_mask = 16'hFFFE;
defparam \next_block~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \data_in_r~0 (
	.dataa(reset_n),
	.datab(core_real_in_2),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_r~0_combout ),
	.cout());
defparam \data_in_r~0 .lut_mask = 16'hEEEE;
defparam \data_in_r~0 .sum_lutc_input = "datac";

dffeas \wr_addr[0] (
	.clk(clk),
	.d(\count[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\wr_addr[0]~q ),
	.prn(vcc));
defparam \wr_addr[0] .is_wysiwyg = "true";
defparam \wr_addr[0] .power_up = "low";

cycloneiii_lcell_comb \wr_address_i_int~0 (
	.dataa(reset_n),
	.datab(\wr_addr[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wr_address_i_int~0_combout ),
	.cout());
defparam \wr_address_i_int~0 .lut_mask = 16'hEEEE;
defparam \wr_address_i_int~0 .sum_lutc_input = "datac";

dffeas \wr_addr[1] (
	.clk(clk),
	.d(\count[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\wr_addr[1]~q ),
	.prn(vcc));
defparam \wr_addr[1] .is_wysiwyg = "true";
defparam \wr_addr[1] .power_up = "low";

cycloneiii_lcell_comb \wr_address_i_int~1 (
	.dataa(reset_n),
	.datab(\wr_addr[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wr_address_i_int~1_combout ),
	.cout());
defparam \wr_address_i_int~1 .lut_mask = 16'hEEEE;
defparam \wr_address_i_int~1 .sum_lutc_input = "datac";

dffeas \count[3] (
	.clk(clk),
	.d(\count[3]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\counter_i~0_combout ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\count[3]~q ),
	.prn(vcc));
defparam \count[3] .is_wysiwyg = "true";
defparam \count[3] .power_up = "low";

dffeas \wr_addr[2] (
	.clk(clk),
	.d(\count[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\wr_addr[2]~q ),
	.prn(vcc));
defparam \wr_addr[2] .is_wysiwyg = "true";
defparam \wr_addr[2] .power_up = "low";

cycloneiii_lcell_comb \wr_address_i_int~2 (
	.dataa(reset_n),
	.datab(\wr_addr[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wr_address_i_int~2_combout ),
	.cout());
defparam \wr_address_i_int~2 .lut_mask = 16'hEEEE;
defparam \wr_address_i_int~2 .sum_lutc_input = "datac";

dffeas \wr_addr[3] (
	.clk(clk),
	.d(\count[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\wr_addr[3]~q ),
	.prn(vcc));
defparam \wr_addr[3] .is_wysiwyg = "true";
defparam \wr_addr[3] .power_up = "low";

cycloneiii_lcell_comb \wr_address_i_int~3 (
	.dataa(reset_n),
	.datab(\wr_addr[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wr_address_i_int~3_combout ),
	.cout());
defparam \wr_address_i_int~3 .lut_mask = 16'hEEEE;
defparam \wr_address_i_int~3 .sum_lutc_input = "datac";

dffeas \wr_addr[4] (
	.clk(clk),
	.d(\count[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\wr_addr[4]~q ),
	.prn(vcc));
defparam \wr_addr[4] .is_wysiwyg = "true";
defparam \wr_addr[4] .power_up = "low";

cycloneiii_lcell_comb \wr_address_i_int~4 (
	.dataa(reset_n),
	.datab(\wr_addr[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wr_address_i_int~4_combout ),
	.cout());
defparam \wr_address_i_int~4 .lut_mask = 16'hEEEE;
defparam \wr_address_i_int~4 .sum_lutc_input = "datac";

dffeas \wr_addr[5] (
	.clk(clk),
	.d(\count[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\wr_addr[5]~q ),
	.prn(vcc));
defparam \wr_addr[5] .is_wysiwyg = "true";
defparam \wr_addr[5] .power_up = "low";

cycloneiii_lcell_comb \wr_address_i_int~5 (
	.dataa(reset_n),
	.datab(\wr_addr[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wr_address_i_int~5_combout ),
	.cout());
defparam \wr_address_i_int~5 .lut_mask = 16'hEEEE;
defparam \wr_address_i_int~5 .sum_lutc_input = "datac";

dffeas \wr_addr[6] (
	.clk(clk),
	.d(\count[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\wr_addr[6]~q ),
	.prn(vcc));
defparam \wr_addr[6] .is_wysiwyg = "true";
defparam \wr_addr[6] .power_up = "low";

cycloneiii_lcell_comb \wr_address_i_int~6 (
	.dataa(reset_n),
	.datab(\wr_addr[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wr_address_i_int~6_combout ),
	.cout());
defparam \wr_address_i_int~6 .lut_mask = 16'hEEEE;
defparam \wr_address_i_int~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \data_in_r~1 (
	.dataa(reset_n),
	.datab(core_real_in_6),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_r~1_combout ),
	.cout());
defparam \data_in_r~1 .lut_mask = 16'hEEEE;
defparam \data_in_r~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \data_in_r~2 (
	.dataa(reset_n),
	.datab(core_real_in_4),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_r~2_combout ),
	.cout());
defparam \data_in_r~2 .lut_mask = 16'hEEEE;
defparam \data_in_r~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \data_in_r~3 (
	.dataa(reset_n),
	.datab(core_real_in_3),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_r~3_combout ),
	.cout());
defparam \data_in_r~3 .lut_mask = 16'hEEEE;
defparam \data_in_r~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \data_in_r~4 (
	.dataa(reset_n),
	.datab(core_real_in_5),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_r~4_combout ),
	.cout());
defparam \data_in_r~4 .lut_mask = 16'hEEEE;
defparam \data_in_r~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \data_in_r~5 (
	.dataa(reset_n),
	.datab(core_real_in_1),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_r~5_combout ),
	.cout());
defparam \data_in_r~5 .lut_mask = 16'hEEEE;
defparam \data_in_r~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \data_in_r~6 (
	.dataa(reset_n),
	.datab(core_real_in_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_r~6_combout ),
	.cout());
defparam \data_in_r~6 .lut_mask = 16'hEEEE;
defparam \data_in_r~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \data_in_r~7 (
	.dataa(reset_n),
	.datab(core_real_in_7),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_r~7_combout ),
	.cout());
defparam \data_in_r~7 .lut_mask = 16'hEEEE;
defparam \data_in_r~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \data_in_i~0 (
	.dataa(reset_n),
	.datab(core_imag_in_7),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_i~0_combout ),
	.cout());
defparam \data_in_i~0 .lut_mask = 16'hEEEE;
defparam \data_in_i~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \data_in_i~1 (
	.dataa(reset_n),
	.datab(core_imag_in_3),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_i~1_combout ),
	.cout());
defparam \data_in_i~1 .lut_mask = 16'hEEEE;
defparam \data_in_i~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \data_in_i~2 (
	.dataa(reset_n),
	.datab(core_imag_in_5),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_i~2_combout ),
	.cout());
defparam \data_in_i~2 .lut_mask = 16'hEEEE;
defparam \data_in_i~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \data_in_i~3 (
	.dataa(reset_n),
	.datab(core_imag_in_4),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_i~3_combout ),
	.cout());
defparam \data_in_i~3 .lut_mask = 16'hEEEE;
defparam \data_in_i~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \data_in_i~4 (
	.dataa(reset_n),
	.datab(core_imag_in_6),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_i~4_combout ),
	.cout());
defparam \data_in_i~4 .lut_mask = 16'hEEEE;
defparam \data_in_i~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \data_in_i~5 (
	.dataa(reset_n),
	.datab(core_imag_in_2),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_i~5_combout ),
	.cout());
defparam \data_in_i~5 .lut_mask = 16'hEEEE;
defparam \data_in_i~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \data_in_i~6 (
	.dataa(reset_n),
	.datab(core_imag_in_1),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_i~6_combout ),
	.cout());
defparam \data_in_i~6 .lut_mask = 16'hEEEE;
defparam \data_in_i~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \data_in_i~7 (
	.dataa(reset_n),
	.datab(core_imag_in_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_i~7_combout ),
	.cout());
defparam \data_in_i~7 .lut_mask = 16'hEEEE;
defparam \data_in_i~7 .sum_lutc_input = "datac";

endmodule

module fft_asj_fft_lpp_serial_r2_fft_120 (
	lpp_ram_data_out_sw_1_1,
	lpp_ram_data_out_sw_1_0,
	lpp_ram_data_out_sw_0_1,
	lpp_ram_data_out_sw_0_0,
	lpp_ram_data_out_sw_7_1,
	lpp_ram_data_out_sw_7_0,
	lpp_ram_data_out_sw_6_1,
	lpp_ram_data_out_sw_6_0,
	lpp_ram_data_out_sw_5_1,
	lpp_ram_data_out_sw_5_0,
	lpp_ram_data_out_sw_4_1,
	lpp_ram_data_out_sw_4_0,
	lpp_ram_data_out_sw_3_1,
	lpp_ram_data_out_sw_3_0,
	lpp_ram_data_out_sw_2_1,
	lpp_ram_data_out_sw_2_0,
	lpp_ram_data_out_sw_9_1,
	lpp_ram_data_out_sw_9_0,
	lpp_ram_data_out_sw_8_1,
	lpp_ram_data_out_sw_8_0,
	lpp_ram_data_out_sw_15_1,
	lpp_ram_data_out_sw_15_0,
	lpp_ram_data_out_sw_14_1,
	lpp_ram_data_out_sw_14_0,
	lpp_ram_data_out_sw_13_1,
	lpp_ram_data_out_sw_13_0,
	lpp_ram_data_out_sw_12_1,
	lpp_ram_data_out_sw_12_0,
	lpp_ram_data_out_sw_11_1,
	lpp_ram_data_out_sw_11_0,
	lpp_ram_data_out_sw_10_1,
	lpp_ram_data_out_sw_10_0,
	source_valid_ctrl_sop,
	stall_reg,
	source_stall_int_d,
	global_clock_enable,
	data_imag_o_0,
	data_real_o_0,
	data_imag_o_1,
	data_real_o_1,
	data_imag_o_2,
	data_real_o_2,
	data_imag_o_3,
	data_real_o_3,
	data_imag_o_4,
	data_real_o_4,
	data_imag_o_5,
	data_real_o_5,
	data_imag_o_6,
	data_real_o_6,
	data_imag_o_7,
	data_real_o_7,
	tdl_arr_4,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	lpp_ram_data_out_sw_1_1;
input 	lpp_ram_data_out_sw_1_0;
input 	lpp_ram_data_out_sw_0_1;
input 	lpp_ram_data_out_sw_0_0;
input 	lpp_ram_data_out_sw_7_1;
input 	lpp_ram_data_out_sw_7_0;
input 	lpp_ram_data_out_sw_6_1;
input 	lpp_ram_data_out_sw_6_0;
input 	lpp_ram_data_out_sw_5_1;
input 	lpp_ram_data_out_sw_5_0;
input 	lpp_ram_data_out_sw_4_1;
input 	lpp_ram_data_out_sw_4_0;
input 	lpp_ram_data_out_sw_3_1;
input 	lpp_ram_data_out_sw_3_0;
input 	lpp_ram_data_out_sw_2_1;
input 	lpp_ram_data_out_sw_2_0;
input 	lpp_ram_data_out_sw_9_1;
input 	lpp_ram_data_out_sw_9_0;
input 	lpp_ram_data_out_sw_8_1;
input 	lpp_ram_data_out_sw_8_0;
input 	lpp_ram_data_out_sw_15_1;
input 	lpp_ram_data_out_sw_15_0;
input 	lpp_ram_data_out_sw_14_1;
input 	lpp_ram_data_out_sw_14_0;
input 	lpp_ram_data_out_sw_13_1;
input 	lpp_ram_data_out_sw_13_0;
input 	lpp_ram_data_out_sw_12_1;
input 	lpp_ram_data_out_sw_12_0;
input 	lpp_ram_data_out_sw_11_1;
input 	lpp_ram_data_out_sw_11_0;
input 	lpp_ram_data_out_sw_10_1;
input 	lpp_ram_data_out_sw_10_0;
input 	source_valid_ctrl_sop;
input 	stall_reg;
input 	source_stall_int_d;
input 	global_clock_enable;
output 	data_imag_o_0;
output 	data_real_o_0;
output 	data_imag_o_1;
output 	data_real_o_1;
output 	data_imag_o_2;
output 	data_real_o_2;
output 	data_imag_o_3;
output 	data_real_o_3;
output 	data_imag_o_4;
output 	data_real_o_4;
output 	data_imag_o_5;
output 	data_real_o_5;
output 	data_imag_o_6;
output 	data_real_o_6;
output 	data_imag_o_7;
output 	data_real_o_7;
input 	tdl_arr_4;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~q ;
wire \gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~q ;
wire \gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ;
wire \gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ;
wire \gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ;
wire \gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ;
wire \gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ;
wire \gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ;
wire \gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ;
wire \gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ;
wire \gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ;
wire \gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ;
wire \gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ;
wire \gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ;
wire \gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ;
wire \gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ;
wire \output_i[1]~q ;
wire \output_i[8]~q ;
wire \output_i[0]~q ;
wire \output_r[1]~q ;
wire \output_r[8]~q ;
wire \output_r[0]~q ;
wire \output_i[2]~q ;
wire \output_r[2]~q ;
wire \output_i[3]~q ;
wire \output_r[3]~q ;
wire \output_i[4]~q ;
wire \output_r[4]~q ;
wire \output_i[5]~q ;
wire \output_r[5]~q ;
wire \output_i[6]~q ;
wire \output_r[6]~q ;
wire \output_i[7]~q ;
wire \output_r[7]~q ;
wire \output_i[0]~10_cout ;
wire \output_i[0]~12 ;
wire \output_i[0]~11_combout ;
wire \output_i[1]~14 ;
wire \output_i[1]~13_combout ;
wire \output_i[2]~16 ;
wire \output_i[2]~15_combout ;
wire \output_i[3]~18 ;
wire \output_i[3]~17_combout ;
wire \output_i[4]~20 ;
wire \output_i[4]~19_combout ;
wire \output_i[5]~22 ;
wire \output_i[5]~21_combout ;
wire \output_i[6]~24 ;
wire \output_i[6]~23_combout ;
wire \output_i[7]~26 ;
wire \output_i[7]~25_combout ;
wire \output_i[8]~27_combout ;
wire \output_r[0]~10_cout ;
wire \output_r[0]~12 ;
wire \output_r[0]~11_combout ;
wire \output_r[1]~14 ;
wire \output_r[1]~13_combout ;
wire \output_r[2]~16 ;
wire \output_r[2]~15_combout ;
wire \output_r[3]~18 ;
wire \output_r[3]~17_combout ;
wire \output_r[4]~20 ;
wire \output_r[4]~19_combout ;
wire \output_r[5]~22 ;
wire \output_r[5]~21_combout ;
wire \output_r[6]~24 ;
wire \output_r[6]~23_combout ;
wire \output_r[7]~26 ;
wire \output_r[7]~25_combout ;
wire \output_r[8]~27_combout ;
wire \offset_counter[8]~q ;
wire \offset_counter[7]~q ;
wire \offset_counter[6]~q ;
wire \offset_counter[5]~q ;
wire \offset_counter[4]~q ;
wire \offset_counter[3]~q ;
wire \offset_counter[2]~q ;
wire \offset_counter[1]~q ;
wire \offset_counter[0]~q ;
wire \offset_counter[0]~10 ;
wire \offset_counter[0]~9_combout ;
wire \offset_counter[1]~12 ;
wire \offset_counter[1]~11_combout ;
wire \offset_counter[2]~14 ;
wire \offset_counter[2]~13_combout ;
wire \offset_counter[3]~16 ;
wire \offset_counter[3]~15_combout ;
wire \offset_counter[4]~18 ;
wire \offset_counter[4]~17_combout ;
wire \offset_counter[5]~20 ;
wire \offset_counter[5]~19_combout ;
wire \offset_counter[6]~22 ;
wire \offset_counter[6]~21_combout ;
wire \offset_counter[7]~24 ;
wire \offset_counter[7]~23_combout ;
wire \offset_counter[8]~25_combout ;
wire \sign_sel~q ;
wire \Add2~1_combout ;
wire \Add2~2_combout ;
wire \Add2~3_combout ;
wire \Add2~4_combout ;
wire \Add2~5_combout ;
wire \Add2~6_combout ;
wire \Add2~7_combout ;
wire \Add2~8_combout ;
wire \Add1~1_combout ;
wire \Add1~2_combout ;
wire \Add1~3_combout ;
wire \Add1~4_combout ;
wire \Add1~5_combout ;
wire \Add1~6_combout ;
wire \Add1~7_combout ;
wire \Add1~8_combout ;
wire \sign_sel_tmp~q ;
wire \offset_counter[0]~27_combout ;
wire \sign_sel_tmp~0_combout ;
wire \data_imag_o[0]~0_combout ;
wire \data_real_o~0_combout ;
wire \data_real_o~1_combout ;
wire \data_real_o~2_combout ;
wire \data_real_o~3_combout ;
wire \data_real_o~4_combout ;
wire \data_real_o~5_combout ;
wire \data_real_o~6_combout ;
wire \data_real_o~7_combout ;


fft_asj_fft_pround_fft_120_15 \gen_full_rnd:u1 (
	.pipeline_dffe_1(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_2(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.output_i_1(\output_i[1]~q ),
	.output_i_8(\output_i[8]~q ),
	.output_i_0(\output_i[0]~q ),
	.output_i_2(\output_i[2]~q ),
	.output_i_3(\output_i[3]~q ),
	.output_i_4(\output_i[4]~q ),
	.output_i_5(\output_i[5]~q ),
	.output_i_6(\output_i[6]~q ),
	.output_i_7(\output_i[7]~q ),
	.global_clock_enable(global_clock_enable),
	.clk(clk));

fft_asj_fft_pround_fft_120_14 \gen_full_rnd:u0 (
	.pipeline_dffe_1(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_2(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.output_r_1(\output_r[1]~q ),
	.output_r_8(\output_r[8]~q ),
	.output_r_0(\output_r[0]~q ),
	.output_r_2(\output_r[2]~q ),
	.output_r_3(\output_r[3]~q ),
	.output_r_4(\output_r[4]~q ),
	.output_r_5(\output_r[5]~q ),
	.output_r_6(\output_r[6]~q ),
	.output_r_7(\output_r[7]~q ),
	.global_clock_enable(global_clock_enable),
	.clk(clk));

dffeas \output_i[1] (
	.clk(clk),
	.d(\output_i[1]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\output_i[1]~q ),
	.prn(vcc));
defparam \output_i[1] .is_wysiwyg = "true";
defparam \output_i[1] .power_up = "low";

dffeas \output_i[8] (
	.clk(clk),
	.d(\output_i[8]~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\output_i[8]~q ),
	.prn(vcc));
defparam \output_i[8] .is_wysiwyg = "true";
defparam \output_i[8] .power_up = "low";

dffeas \output_i[0] (
	.clk(clk),
	.d(\output_i[0]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\output_i[0]~q ),
	.prn(vcc));
defparam \output_i[0] .is_wysiwyg = "true";
defparam \output_i[0] .power_up = "low";

dffeas \output_r[1] (
	.clk(clk),
	.d(\output_r[1]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\output_r[1]~q ),
	.prn(vcc));
defparam \output_r[1] .is_wysiwyg = "true";
defparam \output_r[1] .power_up = "low";

dffeas \output_r[8] (
	.clk(clk),
	.d(\output_r[8]~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\output_r[8]~q ),
	.prn(vcc));
defparam \output_r[8] .is_wysiwyg = "true";
defparam \output_r[8] .power_up = "low";

dffeas \output_r[0] (
	.clk(clk),
	.d(\output_r[0]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\output_r[0]~q ),
	.prn(vcc));
defparam \output_r[0] .is_wysiwyg = "true";
defparam \output_r[0] .power_up = "low";

dffeas \output_i[2] (
	.clk(clk),
	.d(\output_i[2]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\output_i[2]~q ),
	.prn(vcc));
defparam \output_i[2] .is_wysiwyg = "true";
defparam \output_i[2] .power_up = "low";

dffeas \output_r[2] (
	.clk(clk),
	.d(\output_r[2]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\output_r[2]~q ),
	.prn(vcc));
defparam \output_r[2] .is_wysiwyg = "true";
defparam \output_r[2] .power_up = "low";

dffeas \output_i[3] (
	.clk(clk),
	.d(\output_i[3]~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\output_i[3]~q ),
	.prn(vcc));
defparam \output_i[3] .is_wysiwyg = "true";
defparam \output_i[3] .power_up = "low";

dffeas \output_r[3] (
	.clk(clk),
	.d(\output_r[3]~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\output_r[3]~q ),
	.prn(vcc));
defparam \output_r[3] .is_wysiwyg = "true";
defparam \output_r[3] .power_up = "low";

dffeas \output_i[4] (
	.clk(clk),
	.d(\output_i[4]~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\output_i[4]~q ),
	.prn(vcc));
defparam \output_i[4] .is_wysiwyg = "true";
defparam \output_i[4] .power_up = "low";

dffeas \output_r[4] (
	.clk(clk),
	.d(\output_r[4]~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\output_r[4]~q ),
	.prn(vcc));
defparam \output_r[4] .is_wysiwyg = "true";
defparam \output_r[4] .power_up = "low";

dffeas \output_i[5] (
	.clk(clk),
	.d(\output_i[5]~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\output_i[5]~q ),
	.prn(vcc));
defparam \output_i[5] .is_wysiwyg = "true";
defparam \output_i[5] .power_up = "low";

dffeas \output_r[5] (
	.clk(clk),
	.d(\output_r[5]~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\output_r[5]~q ),
	.prn(vcc));
defparam \output_r[5] .is_wysiwyg = "true";
defparam \output_r[5] .power_up = "low";

dffeas \output_i[6] (
	.clk(clk),
	.d(\output_i[6]~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\output_i[6]~q ),
	.prn(vcc));
defparam \output_i[6] .is_wysiwyg = "true";
defparam \output_i[6] .power_up = "low";

dffeas \output_r[6] (
	.clk(clk),
	.d(\output_r[6]~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\output_r[6]~q ),
	.prn(vcc));
defparam \output_r[6] .is_wysiwyg = "true";
defparam \output_r[6] .power_up = "low";

dffeas \output_i[7] (
	.clk(clk),
	.d(\output_i[7]~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\output_i[7]~q ),
	.prn(vcc));
defparam \output_i[7] .is_wysiwyg = "true";
defparam \output_i[7] .power_up = "low";

dffeas \output_r[7] (
	.clk(clk),
	.d(\output_r[7]~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\output_r[7]~q ),
	.prn(vcc));
defparam \output_r[7] .is_wysiwyg = "true";
defparam \output_r[7] .power_up = "low";

cycloneiii_lcell_comb \output_i[0]~10 (
	.dataa(\sign_sel~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\output_i[0]~10_cout ));
defparam \output_i[0]~10 .lut_mask = 16'h0055;
defparam \output_i[0]~10 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \output_i[0]~11 (
	.dataa(\Add2~2_combout ),
	.datab(lpp_ram_data_out_sw_0_0),
	.datac(gnd),
	.datad(vcc),
	.cin(\output_i[0]~10_cout ),
	.combout(\output_i[0]~11_combout ),
	.cout(\output_i[0]~12 ));
defparam \output_i[0]~11 .lut_mask = 16'h96BF;
defparam \output_i[0]~11 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \output_i[1]~13 (
	.dataa(\Add2~1_combout ),
	.datab(lpp_ram_data_out_sw_1_0),
	.datac(gnd),
	.datad(vcc),
	.cin(\output_i[0]~12 ),
	.combout(\output_i[1]~13_combout ),
	.cout(\output_i[1]~14 ));
defparam \output_i[1]~13 .lut_mask = 16'h96DF;
defparam \output_i[1]~13 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \output_i[2]~15 (
	.dataa(\Add2~8_combout ),
	.datab(lpp_ram_data_out_sw_2_0),
	.datac(gnd),
	.datad(vcc),
	.cin(\output_i[1]~14 ),
	.combout(\output_i[2]~15_combout ),
	.cout(\output_i[2]~16 ));
defparam \output_i[2]~15 .lut_mask = 16'h96BF;
defparam \output_i[2]~15 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \output_i[3]~17 (
	.dataa(\Add2~7_combout ),
	.datab(lpp_ram_data_out_sw_3_0),
	.datac(gnd),
	.datad(vcc),
	.cin(\output_i[2]~16 ),
	.combout(\output_i[3]~17_combout ),
	.cout(\output_i[3]~18 ));
defparam \output_i[3]~17 .lut_mask = 16'h96DF;
defparam \output_i[3]~17 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \output_i[4]~19 (
	.dataa(\Add2~6_combout ),
	.datab(lpp_ram_data_out_sw_4_0),
	.datac(gnd),
	.datad(vcc),
	.cin(\output_i[3]~18 ),
	.combout(\output_i[4]~19_combout ),
	.cout(\output_i[4]~20 ));
defparam \output_i[4]~19 .lut_mask = 16'h96BF;
defparam \output_i[4]~19 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \output_i[5]~21 (
	.dataa(\Add2~5_combout ),
	.datab(lpp_ram_data_out_sw_5_0),
	.datac(gnd),
	.datad(vcc),
	.cin(\output_i[4]~20 ),
	.combout(\output_i[5]~21_combout ),
	.cout(\output_i[5]~22 ));
defparam \output_i[5]~21 .lut_mask = 16'h96DF;
defparam \output_i[5]~21 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \output_i[6]~23 (
	.dataa(\Add2~4_combout ),
	.datab(lpp_ram_data_out_sw_6_0),
	.datac(gnd),
	.datad(vcc),
	.cin(\output_i[5]~22 ),
	.combout(\output_i[6]~23_combout ),
	.cout(\output_i[6]~24 ));
defparam \output_i[6]~23 .lut_mask = 16'h96BF;
defparam \output_i[6]~23 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \output_i[7]~25 (
	.dataa(\Add2~3_combout ),
	.datab(lpp_ram_data_out_sw_7_0),
	.datac(gnd),
	.datad(vcc),
	.cin(\output_i[6]~24 ),
	.combout(\output_i[7]~25_combout ),
	.cout(\output_i[7]~26 ));
defparam \output_i[7]~25 .lut_mask = 16'h96DF;
defparam \output_i[7]~25 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \output_i[8]~27 (
	.dataa(\Add2~3_combout ),
	.datab(lpp_ram_data_out_sw_7_0),
	.datac(gnd),
	.datad(gnd),
	.cin(\output_i[7]~26 ),
	.combout(\output_i[8]~27_combout ),
	.cout());
defparam \output_i[8]~27 .lut_mask = 16'h9696;
defparam \output_i[8]~27 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \output_r[0]~10 (
	.dataa(\sign_sel~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\output_r[0]~10_cout ));
defparam \output_r[0]~10 .lut_mask = 16'h0055;
defparam \output_r[0]~10 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \output_r[0]~11 (
	.dataa(\Add1~2_combout ),
	.datab(lpp_ram_data_out_sw_8_0),
	.datac(gnd),
	.datad(vcc),
	.cin(\output_r[0]~10_cout ),
	.combout(\output_r[0]~11_combout ),
	.cout(\output_r[0]~12 ));
defparam \output_r[0]~11 .lut_mask = 16'h96BF;
defparam \output_r[0]~11 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \output_r[1]~13 (
	.dataa(\Add1~1_combout ),
	.datab(lpp_ram_data_out_sw_9_0),
	.datac(gnd),
	.datad(vcc),
	.cin(\output_r[0]~12 ),
	.combout(\output_r[1]~13_combout ),
	.cout(\output_r[1]~14 ));
defparam \output_r[1]~13 .lut_mask = 16'h96DF;
defparam \output_r[1]~13 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \output_r[2]~15 (
	.dataa(\Add1~8_combout ),
	.datab(lpp_ram_data_out_sw_10_0),
	.datac(gnd),
	.datad(vcc),
	.cin(\output_r[1]~14 ),
	.combout(\output_r[2]~15_combout ),
	.cout(\output_r[2]~16 ));
defparam \output_r[2]~15 .lut_mask = 16'h96BF;
defparam \output_r[2]~15 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \output_r[3]~17 (
	.dataa(\Add1~7_combout ),
	.datab(lpp_ram_data_out_sw_11_0),
	.datac(gnd),
	.datad(vcc),
	.cin(\output_r[2]~16 ),
	.combout(\output_r[3]~17_combout ),
	.cout(\output_r[3]~18 ));
defparam \output_r[3]~17 .lut_mask = 16'h96DF;
defparam \output_r[3]~17 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \output_r[4]~19 (
	.dataa(\Add1~6_combout ),
	.datab(lpp_ram_data_out_sw_12_0),
	.datac(gnd),
	.datad(vcc),
	.cin(\output_r[3]~18 ),
	.combout(\output_r[4]~19_combout ),
	.cout(\output_r[4]~20 ));
defparam \output_r[4]~19 .lut_mask = 16'h96BF;
defparam \output_r[4]~19 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \output_r[5]~21 (
	.dataa(\Add1~5_combout ),
	.datab(lpp_ram_data_out_sw_13_0),
	.datac(gnd),
	.datad(vcc),
	.cin(\output_r[4]~20 ),
	.combout(\output_r[5]~21_combout ),
	.cout(\output_r[5]~22 ));
defparam \output_r[5]~21 .lut_mask = 16'h96DF;
defparam \output_r[5]~21 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \output_r[6]~23 (
	.dataa(\Add1~4_combout ),
	.datab(lpp_ram_data_out_sw_14_0),
	.datac(gnd),
	.datad(vcc),
	.cin(\output_r[5]~22 ),
	.combout(\output_r[6]~23_combout ),
	.cout(\output_r[6]~24 ));
defparam \output_r[6]~23 .lut_mask = 16'h96BF;
defparam \output_r[6]~23 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \output_r[7]~25 (
	.dataa(\Add1~3_combout ),
	.datab(lpp_ram_data_out_sw_15_0),
	.datac(gnd),
	.datad(vcc),
	.cin(\output_r[6]~24 ),
	.combout(\output_r[7]~25_combout ),
	.cout(\output_r[7]~26 ));
defparam \output_r[7]~25 .lut_mask = 16'h96DF;
defparam \output_r[7]~25 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \output_r[8]~27 (
	.dataa(\Add1~3_combout ),
	.datab(lpp_ram_data_out_sw_15_0),
	.datac(gnd),
	.datad(gnd),
	.cin(\output_r[7]~26 ),
	.combout(\output_r[8]~27_combout ),
	.cout());
defparam \output_r[8]~27 .lut_mask = 16'h9696;
defparam \output_r[8]~27 .sum_lutc_input = "cin";

dffeas \offset_counter[8] (
	.clk(clk),
	.d(\offset_counter[8]~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\offset_counter[0]~27_combout ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\offset_counter[8]~q ),
	.prn(vcc));
defparam \offset_counter[8] .is_wysiwyg = "true";
defparam \offset_counter[8] .power_up = "low";

dffeas \offset_counter[7] (
	.clk(clk),
	.d(\offset_counter[7]~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\offset_counter[0]~27_combout ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\offset_counter[7]~q ),
	.prn(vcc));
defparam \offset_counter[7] .is_wysiwyg = "true";
defparam \offset_counter[7] .power_up = "low";

dffeas \offset_counter[6] (
	.clk(clk),
	.d(\offset_counter[6]~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\offset_counter[0]~27_combout ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\offset_counter[6]~q ),
	.prn(vcc));
defparam \offset_counter[6] .is_wysiwyg = "true";
defparam \offset_counter[6] .power_up = "low";

dffeas \offset_counter[5] (
	.clk(clk),
	.d(\offset_counter[5]~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\offset_counter[0]~27_combout ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\offset_counter[5]~q ),
	.prn(vcc));
defparam \offset_counter[5] .is_wysiwyg = "true";
defparam \offset_counter[5] .power_up = "low";

dffeas \offset_counter[4] (
	.clk(clk),
	.d(\offset_counter[4]~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\offset_counter[0]~27_combout ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\offset_counter[4]~q ),
	.prn(vcc));
defparam \offset_counter[4] .is_wysiwyg = "true";
defparam \offset_counter[4] .power_up = "low";

dffeas \offset_counter[3] (
	.clk(clk),
	.d(\offset_counter[3]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\offset_counter[0]~27_combout ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\offset_counter[3]~q ),
	.prn(vcc));
defparam \offset_counter[3] .is_wysiwyg = "true";
defparam \offset_counter[3] .power_up = "low";

dffeas \offset_counter[2] (
	.clk(clk),
	.d(\offset_counter[2]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\offset_counter[0]~27_combout ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\offset_counter[2]~q ),
	.prn(vcc));
defparam \offset_counter[2] .is_wysiwyg = "true";
defparam \offset_counter[2] .power_up = "low";

dffeas \offset_counter[1] (
	.clk(clk),
	.d(\offset_counter[1]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\offset_counter[0]~27_combout ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\offset_counter[1]~q ),
	.prn(vcc));
defparam \offset_counter[1] .is_wysiwyg = "true";
defparam \offset_counter[1] .power_up = "low";

dffeas \offset_counter[0] (
	.clk(clk),
	.d(\offset_counter[0]~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\offset_counter[0]~27_combout ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\offset_counter[0]~q ),
	.prn(vcc));
defparam \offset_counter[0] .is_wysiwyg = "true";
defparam \offset_counter[0] .power_up = "low";

cycloneiii_lcell_comb \offset_counter[0]~9 (
	.dataa(\offset_counter[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\offset_counter[0]~9_combout ),
	.cout(\offset_counter[0]~10 ));
defparam \offset_counter[0]~9 .lut_mask = 16'h55AA;
defparam \offset_counter[0]~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \offset_counter[1]~11 (
	.dataa(\offset_counter[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\offset_counter[0]~10 ),
	.combout(\offset_counter[1]~11_combout ),
	.cout(\offset_counter[1]~12 ));
defparam \offset_counter[1]~11 .lut_mask = 16'h5A5F;
defparam \offset_counter[1]~11 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \offset_counter[2]~13 (
	.dataa(\offset_counter[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\offset_counter[1]~12 ),
	.combout(\offset_counter[2]~13_combout ),
	.cout(\offset_counter[2]~14 ));
defparam \offset_counter[2]~13 .lut_mask = 16'h5AAF;
defparam \offset_counter[2]~13 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \offset_counter[3]~15 (
	.dataa(\offset_counter[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\offset_counter[2]~14 ),
	.combout(\offset_counter[3]~15_combout ),
	.cout(\offset_counter[3]~16 ));
defparam \offset_counter[3]~15 .lut_mask = 16'h5A5F;
defparam \offset_counter[3]~15 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \offset_counter[4]~17 (
	.dataa(\offset_counter[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\offset_counter[3]~16 ),
	.combout(\offset_counter[4]~17_combout ),
	.cout(\offset_counter[4]~18 ));
defparam \offset_counter[4]~17 .lut_mask = 16'h5AAF;
defparam \offset_counter[4]~17 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \offset_counter[5]~19 (
	.dataa(\offset_counter[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\offset_counter[4]~18 ),
	.combout(\offset_counter[5]~19_combout ),
	.cout(\offset_counter[5]~20 ));
defparam \offset_counter[5]~19 .lut_mask = 16'h5A5F;
defparam \offset_counter[5]~19 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \offset_counter[6]~21 (
	.dataa(\offset_counter[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\offset_counter[5]~20 ),
	.combout(\offset_counter[6]~21_combout ),
	.cout(\offset_counter[6]~22 ));
defparam \offset_counter[6]~21 .lut_mask = 16'h5AAF;
defparam \offset_counter[6]~21 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \offset_counter[7]~23 (
	.dataa(\offset_counter[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\offset_counter[6]~22 ),
	.combout(\offset_counter[7]~23_combout ),
	.cout(\offset_counter[7]~24 ));
defparam \offset_counter[7]~23 .lut_mask = 16'h5A5F;
defparam \offset_counter[7]~23 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \offset_counter[8]~25 (
	.dataa(\offset_counter[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\offset_counter[7]~24 ),
	.combout(\offset_counter[8]~25_combout ),
	.cout());
defparam \offset_counter[8]~25 .lut_mask = 16'h5A5A;
defparam \offset_counter[8]~25 .sum_lutc_input = "cin";

dffeas sign_sel(
	.clk(clk),
	.d(\sign_sel_tmp~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sign_sel~q ),
	.prn(vcc));
defparam sign_sel.is_wysiwyg = "true";
defparam sign_sel.power_up = "low";

cycloneiii_lcell_comb \Add2~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sign_sel~q ),
	.datad(lpp_ram_data_out_sw_1_1),
	.cin(gnd),
	.combout(\Add2~1_combout ),
	.cout());
defparam \Add2~1 .lut_mask = 16'h0FF0;
defparam \Add2~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add2~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sign_sel~q ),
	.datad(lpp_ram_data_out_sw_0_1),
	.cin(gnd),
	.combout(\Add2~2_combout ),
	.cout());
defparam \Add2~2 .lut_mask = 16'h0FF0;
defparam \Add2~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add2~3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sign_sel~q ),
	.datad(lpp_ram_data_out_sw_7_1),
	.cin(gnd),
	.combout(\Add2~3_combout ),
	.cout());
defparam \Add2~3 .lut_mask = 16'h0FF0;
defparam \Add2~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add2~4 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sign_sel~q ),
	.datad(lpp_ram_data_out_sw_6_1),
	.cin(gnd),
	.combout(\Add2~4_combout ),
	.cout());
defparam \Add2~4 .lut_mask = 16'h0FF0;
defparam \Add2~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add2~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sign_sel~q ),
	.datad(lpp_ram_data_out_sw_5_1),
	.cin(gnd),
	.combout(\Add2~5_combout ),
	.cout());
defparam \Add2~5 .lut_mask = 16'h0FF0;
defparam \Add2~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add2~6 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sign_sel~q ),
	.datad(lpp_ram_data_out_sw_4_1),
	.cin(gnd),
	.combout(\Add2~6_combout ),
	.cout());
defparam \Add2~6 .lut_mask = 16'h0FF0;
defparam \Add2~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add2~7 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sign_sel~q ),
	.datad(lpp_ram_data_out_sw_3_1),
	.cin(gnd),
	.combout(\Add2~7_combout ),
	.cout());
defparam \Add2~7 .lut_mask = 16'h0FF0;
defparam \Add2~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add2~8 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sign_sel~q ),
	.datad(lpp_ram_data_out_sw_2_1),
	.cin(gnd),
	.combout(\Add2~8_combout ),
	.cout());
defparam \Add2~8 .lut_mask = 16'h0FF0;
defparam \Add2~8 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sign_sel~q ),
	.datad(lpp_ram_data_out_sw_9_1),
	.cin(gnd),
	.combout(\Add1~1_combout ),
	.cout());
defparam \Add1~1 .lut_mask = 16'h0FF0;
defparam \Add1~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add1~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sign_sel~q ),
	.datad(lpp_ram_data_out_sw_8_1),
	.cin(gnd),
	.combout(\Add1~2_combout ),
	.cout());
defparam \Add1~2 .lut_mask = 16'h0FF0;
defparam \Add1~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add1~3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sign_sel~q ),
	.datad(lpp_ram_data_out_sw_15_1),
	.cin(gnd),
	.combout(\Add1~3_combout ),
	.cout());
defparam \Add1~3 .lut_mask = 16'h0FF0;
defparam \Add1~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add1~4 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sign_sel~q ),
	.datad(lpp_ram_data_out_sw_14_1),
	.cin(gnd),
	.combout(\Add1~4_combout ),
	.cout());
defparam \Add1~4 .lut_mask = 16'h0FF0;
defparam \Add1~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sign_sel~q ),
	.datad(lpp_ram_data_out_sw_13_1),
	.cin(gnd),
	.combout(\Add1~5_combout ),
	.cout());
defparam \Add1~5 .lut_mask = 16'h0FF0;
defparam \Add1~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add1~6 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sign_sel~q ),
	.datad(lpp_ram_data_out_sw_12_1),
	.cin(gnd),
	.combout(\Add1~6_combout ),
	.cout());
defparam \Add1~6 .lut_mask = 16'h0FF0;
defparam \Add1~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add1~7 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sign_sel~q ),
	.datad(lpp_ram_data_out_sw_11_1),
	.cin(gnd),
	.combout(\Add1~7_combout ),
	.cout());
defparam \Add1~7 .lut_mask = 16'h0FF0;
defparam \Add1~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add1~8 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sign_sel~q ),
	.datad(lpp_ram_data_out_sw_10_1),
	.cin(gnd),
	.combout(\Add1~8_combout ),
	.cout());
defparam \Add1~8 .lut_mask = 16'h0FF0;
defparam \Add1~8 .sum_lutc_input = "datac";

dffeas sign_sel_tmp(
	.clk(clk),
	.d(\sign_sel_tmp~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sign_sel_tmp~q ),
	.prn(vcc));
defparam sign_sel_tmp.is_wysiwyg = "true";
defparam sign_sel_tmp.power_up = "low";

cycloneiii_lcell_comb \offset_counter[0]~27 (
	.dataa(reset_n),
	.datab(gnd),
	.datac(gnd),
	.datad(tdl_arr_4),
	.cin(gnd),
	.combout(\offset_counter[0]~27_combout ),
	.cout());
defparam \offset_counter[0]~27 .lut_mask = 16'hFF55;
defparam \offset_counter[0]~27 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sign_sel_tmp~0 (
	.dataa(\offset_counter[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sign_sel_tmp~0_combout ),
	.cout());
defparam \sign_sel_tmp~0 .lut_mask = 16'h5555;
defparam \sign_sel_tmp~0 .sum_lutc_input = "datac";

dffeas \data_imag_o[0] (
	.clk(clk),
	.d(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_imag_o[0]~0_combout ),
	.q(data_imag_o_0),
	.prn(vcc));
defparam \data_imag_o[0] .is_wysiwyg = "true";
defparam \data_imag_o[0] .power_up = "low";

dffeas \data_real_o[0] (
	.clk(clk),
	.d(\data_real_o~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_real_o_0),
	.prn(vcc));
defparam \data_real_o[0] .is_wysiwyg = "true";
defparam \data_real_o[0] .power_up = "low";

dffeas \data_imag_o[1] (
	.clk(clk),
	.d(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_imag_o[0]~0_combout ),
	.q(data_imag_o_1),
	.prn(vcc));
defparam \data_imag_o[1] .is_wysiwyg = "true";
defparam \data_imag_o[1] .power_up = "low";

dffeas \data_real_o[1] (
	.clk(clk),
	.d(\data_real_o~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_real_o_1),
	.prn(vcc));
defparam \data_real_o[1] .is_wysiwyg = "true";
defparam \data_real_o[1] .power_up = "low";

dffeas \data_imag_o[2] (
	.clk(clk),
	.d(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_imag_o[0]~0_combout ),
	.q(data_imag_o_2),
	.prn(vcc));
defparam \data_imag_o[2] .is_wysiwyg = "true";
defparam \data_imag_o[2] .power_up = "low";

dffeas \data_real_o[2] (
	.clk(clk),
	.d(\data_real_o~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_real_o_2),
	.prn(vcc));
defparam \data_real_o[2] .is_wysiwyg = "true";
defparam \data_real_o[2] .power_up = "low";

dffeas \data_imag_o[3] (
	.clk(clk),
	.d(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_imag_o[0]~0_combout ),
	.q(data_imag_o_3),
	.prn(vcc));
defparam \data_imag_o[3] .is_wysiwyg = "true";
defparam \data_imag_o[3] .power_up = "low";

dffeas \data_real_o[3] (
	.clk(clk),
	.d(\data_real_o~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_real_o_3),
	.prn(vcc));
defparam \data_real_o[3] .is_wysiwyg = "true";
defparam \data_real_o[3] .power_up = "low";

dffeas \data_imag_o[4] (
	.clk(clk),
	.d(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_imag_o[0]~0_combout ),
	.q(data_imag_o_4),
	.prn(vcc));
defparam \data_imag_o[4] .is_wysiwyg = "true";
defparam \data_imag_o[4] .power_up = "low";

dffeas \data_real_o[4] (
	.clk(clk),
	.d(\data_real_o~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_real_o_4),
	.prn(vcc));
defparam \data_real_o[4] .is_wysiwyg = "true";
defparam \data_real_o[4] .power_up = "low";

dffeas \data_imag_o[5] (
	.clk(clk),
	.d(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_imag_o[0]~0_combout ),
	.q(data_imag_o_5),
	.prn(vcc));
defparam \data_imag_o[5] .is_wysiwyg = "true";
defparam \data_imag_o[5] .power_up = "low";

dffeas \data_real_o[5] (
	.clk(clk),
	.d(\data_real_o~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_real_o_5),
	.prn(vcc));
defparam \data_real_o[5] .is_wysiwyg = "true";
defparam \data_real_o[5] .power_up = "low";

dffeas \data_imag_o[6] (
	.clk(clk),
	.d(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_imag_o[0]~0_combout ),
	.q(data_imag_o_6),
	.prn(vcc));
defparam \data_imag_o[6] .is_wysiwyg = "true";
defparam \data_imag_o[6] .power_up = "low";

dffeas \data_real_o[6] (
	.clk(clk),
	.d(\data_real_o~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_real_o_6),
	.prn(vcc));
defparam \data_real_o[6] .is_wysiwyg = "true";
defparam \data_real_o[6] .power_up = "low";

dffeas \data_imag_o[7] (
	.clk(clk),
	.d(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_imag_o[0]~0_combout ),
	.q(data_imag_o_7),
	.prn(vcc));
defparam \data_imag_o[7] .is_wysiwyg = "true";
defparam \data_imag_o[7] .power_up = "low";

dffeas \data_real_o[7] (
	.clk(clk),
	.d(\data_real_o~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_real_o_7),
	.prn(vcc));
defparam \data_real_o[7] .is_wysiwyg = "true";
defparam \data_real_o[7] .power_up = "low";

cycloneiii_lcell_comb \data_imag_o[0]~0 (
	.dataa(reset_n),
	.datab(stall_reg),
	.datac(source_valid_ctrl_sop),
	.datad(source_stall_int_d),
	.cin(gnd),
	.combout(\data_imag_o[0]~0_combout ),
	.cout());
defparam \data_imag_o[0]~0 .lut_mask = 16'hACFF;
defparam \data_imag_o[0]~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \data_real_o~0 (
	.dataa(reset_n),
	.datab(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_real_o~0_combout ),
	.cout());
defparam \data_real_o~0 .lut_mask = 16'hEEEE;
defparam \data_real_o~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \data_real_o~1 (
	.dataa(reset_n),
	.datab(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_real_o~1_combout ),
	.cout());
defparam \data_real_o~1 .lut_mask = 16'hEEEE;
defparam \data_real_o~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \data_real_o~2 (
	.dataa(reset_n),
	.datab(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_real_o~2_combout ),
	.cout());
defparam \data_real_o~2 .lut_mask = 16'hEEEE;
defparam \data_real_o~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \data_real_o~3 (
	.dataa(reset_n),
	.datab(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_real_o~3_combout ),
	.cout());
defparam \data_real_o~3 .lut_mask = 16'hEEEE;
defparam \data_real_o~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \data_real_o~4 (
	.dataa(reset_n),
	.datab(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_real_o~4_combout ),
	.cout());
defparam \data_real_o~4 .lut_mask = 16'hEEEE;
defparam \data_real_o~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \data_real_o~5 (
	.dataa(reset_n),
	.datab(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_real_o~5_combout ),
	.cout());
defparam \data_real_o~5 .lut_mask = 16'hEEEE;
defparam \data_real_o~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \data_real_o~6 (
	.dataa(reset_n),
	.datab(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_real_o~6_combout ),
	.cout());
defparam \data_real_o~6 .lut_mask = 16'hEEEE;
defparam \data_real_o~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \data_real_o~7 (
	.dataa(reset_n),
	.datab(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_real_o~7_combout ),
	.cout());
defparam \data_real_o~7 .lut_mask = 16'hEEEE;
defparam \data_real_o~7 .sum_lutc_input = "datac";

endmodule

module fft_asj_fft_pround_fft_120_14 (
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	output_r_1,
	output_r_8,
	output_r_0,
	output_r_2,
	output_r_3,
	output_r_4,
	output_r_5,
	output_r_6,
	output_r_7,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
input 	output_r_1;
input 	output_r_8;
input 	output_r_0;
input 	output_r_2;
input 	output_r_3;
input 	output_r_4;
input 	output_r_5;
input 	output_r_6;
input 	output_r_7;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_LPM_ADD_SUB_15 \gbrnd:nev:gp:lpm_add_sub_component (
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.output_r_1(output_r_1),
	.output_r_8(output_r_8),
	.output_r_0(output_r_0),
	.output_r_2(output_r_2),
	.output_r_3(output_r_3),
	.output_r_4(output_r_4),
	.output_r_5(output_r_5),
	.output_r_6(output_r_6),
	.output_r_7(output_r_7),
	.clken(global_clock_enable),
	.clock(clk));

endmodule

module fft_LPM_ADD_SUB_15 (
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	output_r_1,
	output_r_8,
	output_r_0,
	output_r_2,
	output_r_3,
	output_r_4,
	output_r_5,
	output_r_6,
	output_r_7,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
input 	output_r_1;
input 	output_r_8;
input 	output_r_0;
input 	output_r_2;
input 	output_r_3;
input 	output_r_4;
input 	output_r_5;
input 	output_r_6;
input 	output_r_7;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_add_sub_g2k auto_generated(
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.output_r_1(output_r_1),
	.output_r_8(output_r_8),
	.output_r_0(output_r_0),
	.output_r_2(output_r_2),
	.output_r_3(output_r_3),
	.output_r_4(output_r_4),
	.output_r_5(output_r_5),
	.output_r_6(output_r_6),
	.output_r_7(output_r_7),
	.clken(clken),
	.clock(clock));

endmodule

module fft_add_sub_g2k (
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	output_r_1,
	output_r_8,
	output_r_0,
	output_r_2,
	output_r_3,
	output_r_4,
	output_r_5,
	output_r_6,
	output_r_7,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
input 	output_r_1;
input 	output_r_8;
input 	output_r_0;
input 	output_r_2;
input 	output_r_3;
input 	output_r_4;
input 	output_r_5;
input 	output_r_6;
input 	output_r_7;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~9_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~10_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~11 ;
wire \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~12_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 ;
wire \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~14_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~15 ;
wire \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~16_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~17 ;
wire \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~18_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~19 ;
wire \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~20_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~21 ;
wire \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~22_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~23 ;
wire \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~24_combout ;


dffeas \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[1] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_1),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[1] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[1] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .power_up = "low";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~9 (
	.dataa(output_r_8),
	.datab(output_r_0),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~9_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~9 .lut_mask = 16'h00DD;
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~10 (
	.dataa(output_r_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~9_cout ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~10_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~11 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~10 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~10 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~12 (
	.dataa(output_r_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~11 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~12_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~12 .lut_mask = 16'h5AAF;
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~12 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~14 (
	.dataa(output_r_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~14_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~15 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~14 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~14 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~16 (
	.dataa(output_r_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~15 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~16_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~17 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~16 .lut_mask = 16'h5AAF;
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~16 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~18 (
	.dataa(output_r_5),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~17 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~18_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~19 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~18 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~18 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~20 (
	.dataa(output_r_6),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~19 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~20_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~21 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~20 .lut_mask = 16'h5AAF;
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~20 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~22 (
	.dataa(output_r_7),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~21 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~22_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~23 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~22 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~22 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~24 (
	.dataa(output_r_8),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~23 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~24_combout ),
	.cout());
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~24 .lut_mask = 16'h5A5A;
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~24 .sum_lutc_input = "cin";

endmodule

module fft_asj_fft_pround_fft_120_15 (
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	output_i_1,
	output_i_8,
	output_i_0,
	output_i_2,
	output_i_3,
	output_i_4,
	output_i_5,
	output_i_6,
	output_i_7,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
input 	output_i_1;
input 	output_i_8;
input 	output_i_0;
input 	output_i_2;
input 	output_i_3;
input 	output_i_4;
input 	output_i_5;
input 	output_i_6;
input 	output_i_7;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_LPM_ADD_SUB_16 \gbrnd:nev:gp:lpm_add_sub_component (
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.output_i_1(output_i_1),
	.output_i_8(output_i_8),
	.output_i_0(output_i_0),
	.output_i_2(output_i_2),
	.output_i_3(output_i_3),
	.output_i_4(output_i_4),
	.output_i_5(output_i_5),
	.output_i_6(output_i_6),
	.output_i_7(output_i_7),
	.clken(global_clock_enable),
	.clock(clk));

endmodule

module fft_LPM_ADD_SUB_16 (
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	output_i_1,
	output_i_8,
	output_i_0,
	output_i_2,
	output_i_3,
	output_i_4,
	output_i_5,
	output_i_6,
	output_i_7,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
input 	output_i_1;
input 	output_i_8;
input 	output_i_0;
input 	output_i_2;
input 	output_i_3;
input 	output_i_4;
input 	output_i_5;
input 	output_i_6;
input 	output_i_7;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_add_sub_g2k_1 auto_generated(
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.output_i_1(output_i_1),
	.output_i_8(output_i_8),
	.output_i_0(output_i_0),
	.output_i_2(output_i_2),
	.output_i_3(output_i_3),
	.output_i_4(output_i_4),
	.output_i_5(output_i_5),
	.output_i_6(output_i_6),
	.output_i_7(output_i_7),
	.clken(clken),
	.clock(clock));

endmodule

module fft_add_sub_g2k_1 (
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	output_i_1,
	output_i_8,
	output_i_0,
	output_i_2,
	output_i_3,
	output_i_4,
	output_i_5,
	output_i_6,
	output_i_7,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
input 	output_i_1;
input 	output_i_8;
input 	output_i_0;
input 	output_i_2;
input 	output_i_3;
input 	output_i_4;
input 	output_i_5;
input 	output_i_6;
input 	output_i_7;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~9_cout ;
wire \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~10_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~11 ;
wire \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~12_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 ;
wire \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~14_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~15 ;
wire \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~16_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~17 ;
wire \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~18_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~19 ;
wire \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~20_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~21 ;
wire \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~22_combout ;
wire \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~23 ;
wire \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~24_combout ;


dffeas \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[1] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_1),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[1] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[1] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .power_up = "low";

dffeas \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] (
	.clk(clock),
	.d(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .is_wysiwyg = "true";
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .power_up = "low";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~9 (
	.dataa(output_i_8),
	.datab(output_i_0),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~9_cout ));
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~9 .lut_mask = 16'h00DD;
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~10 (
	.dataa(output_i_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~9_cout ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~10_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~11 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~10 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~10 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~12 (
	.dataa(output_i_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~11 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~12_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~12 .lut_mask = 16'h5AAF;
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~12 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~14 (
	.dataa(output_i_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~14_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~15 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~14 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~14 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~16 (
	.dataa(output_i_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~15 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~16_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~17 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~16 .lut_mask = 16'h5AAF;
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~16 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~18 (
	.dataa(output_i_5),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~17 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~18_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~19 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~18 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~18 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~20 (
	.dataa(output_i_6),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~19 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~20_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~21 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~20 .lut_mask = 16'h5AAF;
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~20 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~22 (
	.dataa(output_i_7),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~21 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~22_combout ),
	.cout(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~23 ));
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~22 .lut_mask = 16'h5A5F;
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~22 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~24 (
	.dataa(output_i_8),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~23 ),
	.combout(\asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~24_combout ),
	.cout());
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~24 .lut_mask = 16'h5A5A;
defparam \asj_fft_sglstream_fft_120_inst|gen_radix_2_last_pass:lpp_r2|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~24 .sum_lutc_input = "cin";

endmodule

module fft_asj_fft_lpprdadr2gen_fft_120 (
	sw_0,
	global_clock_enable,
	tdl_arr_4,
	tdl_arr_0_4,
	tdl_arr_1_4,
	tdl_arr_19,
	rd_addr_b_0,
	rd_addr_b_1,
	rd_addr_b_2,
	rd_addr_b_3,
	rd_addr_b_4,
	rd_addr_b_5,
	rd_addr_b_6,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	sw_0;
input 	global_clock_enable;
output 	tdl_arr_4;
output 	tdl_arr_0_4;
output 	tdl_arr_1_4;
input 	tdl_arr_19;
output 	rd_addr_b_0;
output 	rd_addr_b_1;
output 	rd_addr_b_2;
output 	rd_addr_b_3;
output 	rd_addr_b_4;
output 	rd_addr_b_5;
output 	rd_addr_b_6;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \en_i~q ;
wire \sw[0]~5 ;
wire \sw[1]~q ;
wire \count[1]~q ;
wire \count[1]~11_combout ;
wire \sw[1]~6_combout ;
wire \en_d~q ;
wire \en_i~0_combout ;
wire \en_d~0_combout ;
wire \Add1~1_combout ;
wire \Add2~1_combout ;
wire \count[0]~10 ;
wire \count[1]~12 ;
wire \count[2]~13_combout ;
wire \counter~0_combout ;
wire \count[2]~q ;
wire \count[0]~9_combout ;
wire \count[0]~q ;
wire \Add1~0_combout ;
wire \count[2]~14 ;
wire \count[3]~16 ;
wire \count[4]~17_combout ;
wire \count[4]~q ;
wire \count[4]~18 ;
wire \count[5]~20 ;
wire \count[6]~21_combout ;
wire \count[6]~q ;
wire \Add2~0_combout ;
wire \sw[0]~3_cout ;
wire \sw[0]~4_combout ;
wire \count[3]~15_combout ;
wire \count[3]~q ;
wire \count[5]~19_combout ;
wire \count[5]~q ;
wire \count[6]~22 ;
wire \count[7]~23_combout ;
wire \count[7]~q ;
wire \count[7]~24 ;
wire \count[8]~25_combout ;
wire \count[8]~q ;
wire \rd_addr_b[6]~0_combout ;


fft_asj_fft_tdl_rst_fft_120 \gen_M4K:delay_swd (
	.sw_0(sw_0),
	.sw_1(\sw[1]~q ),
	.global_clock_enable(global_clock_enable),
	.tdl_arr_0_4(tdl_arr_0_4),
	.tdl_arr_1_4(tdl_arr_1_4),
	.clk(clk),
	.reset_n(reset_n));

fft_asj_fft_tdl_bit_rst_fft_120_2 delay_en(
	.en_i(\en_i~q ),
	.global_clock_enable(global_clock_enable),
	.tdl_arr_4(tdl_arr_4),
	.clk(clk),
	.reset_n(reset_n));

dffeas en_i(
	.clk(clk),
	.d(\en_i~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\en_i~q ),
	.prn(vcc));
defparam en_i.is_wysiwyg = "true";
defparam en_i.power_up = "low";

cycloneiii_lcell_comb \sw[0]~4 (
	.dataa(\Add1~0_combout ),
	.datab(\Add2~0_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\sw[0]~3_cout ),
	.combout(\sw[0]~4_combout ),
	.cout(\sw[0]~5 ));
defparam \sw[0]~4 .lut_mask = 16'h967F;
defparam \sw[0]~4 .sum_lutc_input = "cin";

dffeas \sw[1] (
	.clk(clk),
	.d(\sw[1]~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sw[1]~q ),
	.prn(vcc));
defparam \sw[1] .is_wysiwyg = "true";
defparam \sw[1] .power_up = "low";

dffeas \count[1] (
	.clk(clk),
	.d(\count[1]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\counter~0_combout ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\count[1]~q ),
	.prn(vcc));
defparam \count[1] .is_wysiwyg = "true";
defparam \count[1] .power_up = "low";

cycloneiii_lcell_comb \count[1]~11 (
	.dataa(\count[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[0]~10 ),
	.combout(\count[1]~11_combout ),
	.cout(\count[1]~12 ));
defparam \count[1]~11 .lut_mask = 16'h5A5F;
defparam \count[1]~11 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \sw[1]~6 (
	.dataa(\Add1~1_combout ),
	.datab(\Add2~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(\sw[0]~5 ),
	.combout(\sw[1]~6_combout ),
	.cout());
defparam \sw[1]~6 .lut_mask = 16'h9696;
defparam \sw[1]~6 .sum_lutc_input = "cin";

dffeas en_d(
	.clk(clk),
	.d(\en_d~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\en_d~q ),
	.prn(vcc));
defparam en_d.is_wysiwyg = "true";
defparam en_d.power_up = "low";

cycloneiii_lcell_comb \en_i~0 (
	.dataa(tdl_arr_19),
	.datab(gnd),
	.datac(gnd),
	.datad(\en_d~q ),
	.cin(gnd),
	.combout(\en_i~0_combout ),
	.cout());
defparam \en_i~0 .lut_mask = 16'hAAFF;
defparam \en_i~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \en_d~0 (
	.dataa(tdl_arr_19),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\en_d~0_combout ),
	.cout());
defparam \en_d~0 .lut_mask = 16'hAAFF;
defparam \en_d~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add1~1 (
	.dataa(\count[2]~q ),
	.datab(\count[0]~q ),
	.datac(\count[3]~q ),
	.datad(\count[1]~q ),
	.cin(gnd),
	.combout(\Add1~1_combout ),
	.cout());
defparam \Add1~1 .lut_mask = 16'h6996;
defparam \Add1~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add2~1 (
	.dataa(\count[4]~q ),
	.datab(\count[6]~q ),
	.datac(\count[5]~q ),
	.datad(\count[7]~q ),
	.cin(gnd),
	.combout(\Add2~1_combout ),
	.cout());
defparam \Add2~1 .lut_mask = 16'h6996;
defparam \Add2~1 .sum_lutc_input = "datac";

dffeas \sw[0] (
	.clk(clk),
	.d(\sw[0]~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(sw_0),
	.prn(vcc));
defparam \sw[0] .is_wysiwyg = "true";
defparam \sw[0] .power_up = "low";

dffeas \rd_addr_b[0] (
	.clk(clk),
	.d(\count[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_b_0),
	.prn(vcc));
defparam \rd_addr_b[0] .is_wysiwyg = "true";
defparam \rd_addr_b[0] .power_up = "low";

dffeas \rd_addr_b[1] (
	.clk(clk),
	.d(\count[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_b_1),
	.prn(vcc));
defparam \rd_addr_b[1] .is_wysiwyg = "true";
defparam \rd_addr_b[1] .power_up = "low";

dffeas \rd_addr_b[2] (
	.clk(clk),
	.d(\count[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_b_2),
	.prn(vcc));
defparam \rd_addr_b[2] .is_wysiwyg = "true";
defparam \rd_addr_b[2] .power_up = "low";

dffeas \rd_addr_b[3] (
	.clk(clk),
	.d(\count[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_b_3),
	.prn(vcc));
defparam \rd_addr_b[3] .is_wysiwyg = "true";
defparam \rd_addr_b[3] .power_up = "low";

dffeas \rd_addr_b[4] (
	.clk(clk),
	.d(\count[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_b_4),
	.prn(vcc));
defparam \rd_addr_b[4] .is_wysiwyg = "true";
defparam \rd_addr_b[4] .power_up = "low";

dffeas \rd_addr_b[5] (
	.clk(clk),
	.d(\count[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_b_5),
	.prn(vcc));
defparam \rd_addr_b[5] .is_wysiwyg = "true";
defparam \rd_addr_b[5] .power_up = "low";

dffeas \rd_addr_b[6] (
	.clk(clk),
	.d(\rd_addr_b[6]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_b_6),
	.prn(vcc));
defparam \rd_addr_b[6] .is_wysiwyg = "true";
defparam \rd_addr_b[6] .power_up = "low";

cycloneiii_lcell_comb \count[0]~9 (
	.dataa(\count[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\count[0]~9_combout ),
	.cout(\count[0]~10 ));
defparam \count[0]~9 .lut_mask = 16'h55AA;
defparam \count[0]~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \count[2]~13 (
	.dataa(\count[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[1]~12 ),
	.combout(\count[2]~13_combout ),
	.cout(\count[2]~14 ));
defparam \count[2]~13 .lut_mask = 16'h5AAF;
defparam \count[2]~13 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \counter~0 (
	.dataa(\en_i~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\counter~0_combout ),
	.cout());
defparam \counter~0 .lut_mask = 16'hAAFF;
defparam \counter~0 .sum_lutc_input = "datac";

dffeas \count[2] (
	.clk(clk),
	.d(\count[2]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\counter~0_combout ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\count[2]~q ),
	.prn(vcc));
defparam \count[2] .is_wysiwyg = "true";
defparam \count[2] .power_up = "low";

dffeas \count[0] (
	.clk(clk),
	.d(\count[0]~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\counter~0_combout ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\count[0]~q ),
	.prn(vcc));
defparam \count[0] .is_wysiwyg = "true";
defparam \count[0] .power_up = "low";

cycloneiii_lcell_comb \Add1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\count[2]~q ),
	.datad(\count[0]~q ),
	.cin(gnd),
	.combout(\Add1~0_combout ),
	.cout());
defparam \Add1~0 .lut_mask = 16'h0FF0;
defparam \Add1~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \count[3]~15 (
	.dataa(\count[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[2]~14 ),
	.combout(\count[3]~15_combout ),
	.cout(\count[3]~16 ));
defparam \count[3]~15 .lut_mask = 16'h5A5F;
defparam \count[3]~15 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \count[4]~17 (
	.dataa(\count[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[3]~16 ),
	.combout(\count[4]~17_combout ),
	.cout(\count[4]~18 ));
defparam \count[4]~17 .lut_mask = 16'h5AAF;
defparam \count[4]~17 .sum_lutc_input = "cin";

dffeas \count[4] (
	.clk(clk),
	.d(\count[4]~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\counter~0_combout ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\count[4]~q ),
	.prn(vcc));
defparam \count[4] .is_wysiwyg = "true";
defparam \count[4] .power_up = "low";

cycloneiii_lcell_comb \count[5]~19 (
	.dataa(\count[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[4]~18 ),
	.combout(\count[5]~19_combout ),
	.cout(\count[5]~20 ));
defparam \count[5]~19 .lut_mask = 16'h5A5F;
defparam \count[5]~19 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \count[6]~21 (
	.dataa(\count[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[5]~20 ),
	.combout(\count[6]~21_combout ),
	.cout(\count[6]~22 ));
defparam \count[6]~21 .lut_mask = 16'h5AAF;
defparam \count[6]~21 .sum_lutc_input = "cin";

dffeas \count[6] (
	.clk(clk),
	.d(\count[6]~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\counter~0_combout ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\count[6]~q ),
	.prn(vcc));
defparam \count[6] .is_wysiwyg = "true";
defparam \count[6] .power_up = "low";

cycloneiii_lcell_comb \Add2~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\count[4]~q ),
	.datad(\count[6]~q ),
	.cin(gnd),
	.combout(\Add2~0_combout ),
	.cout());
defparam \Add2~0 .lut_mask = 16'h0FF0;
defparam \Add2~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sw[0]~3 (
	.dataa(\count[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\sw[0]~3_cout ));
defparam \sw[0]~3 .lut_mask = 16'h00AA;
defparam \sw[0]~3 .sum_lutc_input = "datac";

dffeas \count[3] (
	.clk(clk),
	.d(\count[3]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\counter~0_combout ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\count[3]~q ),
	.prn(vcc));
defparam \count[3] .is_wysiwyg = "true";
defparam \count[3] .power_up = "low";

dffeas \count[5] (
	.clk(clk),
	.d(\count[5]~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\counter~0_combout ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\count[5]~q ),
	.prn(vcc));
defparam \count[5] .is_wysiwyg = "true";
defparam \count[5] .power_up = "low";

cycloneiii_lcell_comb \count[7]~23 (
	.dataa(\count[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[6]~22 ),
	.combout(\count[7]~23_combout ),
	.cout(\count[7]~24 ));
defparam \count[7]~23 .lut_mask = 16'h5A5F;
defparam \count[7]~23 .sum_lutc_input = "cin";

dffeas \count[7] (
	.clk(clk),
	.d(\count[7]~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\counter~0_combout ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\count[7]~q ),
	.prn(vcc));
defparam \count[7] .is_wysiwyg = "true";
defparam \count[7] .power_up = "low";

cycloneiii_lcell_comb \count[8]~25 (
	.dataa(\count[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\count[7]~24 ),
	.combout(\count[8]~25_combout ),
	.cout());
defparam \count[8]~25 .lut_mask = 16'h5A5A;
defparam \count[8]~25 .sum_lutc_input = "cin";

dffeas \count[8] (
	.clk(clk),
	.d(\count[8]~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\counter~0_combout ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\count[8]~q ),
	.prn(vcc));
defparam \count[8] .is_wysiwyg = "true";
defparam \count[8] .power_up = "low";

cycloneiii_lcell_comb \rd_addr_b[6]~0 (
	.dataa(\count[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\rd_addr_b[6]~0_combout ),
	.cout());
defparam \rd_addr_b[6]~0 .lut_mask = 16'h5555;
defparam \rd_addr_b[6]~0 .sum_lutc_input = "datac";

endmodule

module fft_asj_fft_tdl_bit_rst_fft_120_2 (
	en_i,
	global_clock_enable,
	tdl_arr_4,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	en_i;
input 	global_clock_enable;
output 	tdl_arr_4;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \tdl_arr~4_combout ;
wire \tdl_arr[0]~q ;
wire \tdl_arr~3_combout ;
wire \tdl_arr[1]~q ;
wire \tdl_arr~2_combout ;
wire \tdl_arr[2]~q ;
wire \tdl_arr~1_combout ;
wire \tdl_arr[3]~q ;
wire \tdl_arr~0_combout ;


dffeas \tdl_arr[4] (
	.clk(clk),
	.d(\tdl_arr~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_4),
	.prn(vcc));
defparam \tdl_arr[4] .is_wysiwyg = "true";
defparam \tdl_arr[4] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~4 (
	.dataa(reset_n),
	.datab(en_i),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~4_combout ),
	.cout());
defparam \tdl_arr~4 .lut_mask = 16'hEEEE;
defparam \tdl_arr~4 .sum_lutc_input = "datac";

dffeas \tdl_arr[0] (
	.clk(clk),
	.d(\tdl_arr~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0]~q ),
	.prn(vcc));
defparam \tdl_arr[0] .is_wysiwyg = "true";
defparam \tdl_arr[0] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~3 (
	.dataa(reset_n),
	.datab(\tdl_arr[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~3_combout ),
	.cout());
defparam \tdl_arr~3 .lut_mask = 16'hEEEE;
defparam \tdl_arr~3 .sum_lutc_input = "datac";

dffeas \tdl_arr[1] (
	.clk(clk),
	.d(\tdl_arr~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[1]~q ),
	.prn(vcc));
defparam \tdl_arr[1] .is_wysiwyg = "true";
defparam \tdl_arr[1] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~2 (
	.dataa(reset_n),
	.datab(\tdl_arr[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~2_combout ),
	.cout());
defparam \tdl_arr~2 .lut_mask = 16'hEEEE;
defparam \tdl_arr~2 .sum_lutc_input = "datac";

dffeas \tdl_arr[2] (
	.clk(clk),
	.d(\tdl_arr~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[2]~q ),
	.prn(vcc));
defparam \tdl_arr[2] .is_wysiwyg = "true";
defparam \tdl_arr[2] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~1 (
	.dataa(reset_n),
	.datab(\tdl_arr[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~1_combout ),
	.cout());
defparam \tdl_arr~1 .lut_mask = 16'hEEEE;
defparam \tdl_arr~1 .sum_lutc_input = "datac";

dffeas \tdl_arr[3] (
	.clk(clk),
	.d(\tdl_arr~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[3]~q ),
	.prn(vcc));
defparam \tdl_arr[3] .is_wysiwyg = "true";
defparam \tdl_arr[3] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~0 (
	.dataa(reset_n),
	.datab(\tdl_arr[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~0_combout ),
	.cout());
defparam \tdl_arr~0 .lut_mask = 16'hEEEE;
defparam \tdl_arr~0 .sum_lutc_input = "datac";

endmodule

module fft_asj_fft_tdl_rst_fft_120 (
	sw_0,
	sw_1,
	global_clock_enable,
	tdl_arr_0_4,
	tdl_arr_1_4,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	sw_0;
input 	sw_1;
input 	global_clock_enable;
output 	tdl_arr_0_4;
output 	tdl_arr_1_4;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \tdl_arr~8_combout ;
wire \tdl_arr[0][0]~q ;
wire \tdl_arr~6_combout ;
wire \tdl_arr[1][0]~q ;
wire \tdl_arr~4_combout ;
wire \tdl_arr[2][0]~q ;
wire \tdl_arr~2_combout ;
wire \tdl_arr[3][0]~q ;
wire \tdl_arr~0_combout ;
wire \tdl_arr~9_combout ;
wire \tdl_arr[0][1]~q ;
wire \tdl_arr~7_combout ;
wire \tdl_arr[1][1]~q ;
wire \tdl_arr~5_combout ;
wire \tdl_arr[2][1]~q ;
wire \tdl_arr~3_combout ;
wire \tdl_arr[3][1]~q ;
wire \tdl_arr~1_combout ;


dffeas \tdl_arr[4][0] (
	.clk(clk),
	.d(\tdl_arr~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_0_4),
	.prn(vcc));
defparam \tdl_arr[4][0] .is_wysiwyg = "true";
defparam \tdl_arr[4][0] .power_up = "low";

dffeas \tdl_arr[4][1] (
	.clk(clk),
	.d(\tdl_arr~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_1_4),
	.prn(vcc));
defparam \tdl_arr[4][1] .is_wysiwyg = "true";
defparam \tdl_arr[4][1] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~8 (
	.dataa(reset_n),
	.datab(sw_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~8_combout ),
	.cout());
defparam \tdl_arr~8 .lut_mask = 16'hEEEE;
defparam \tdl_arr~8 .sum_lutc_input = "datac";

dffeas \tdl_arr[0][0] (
	.clk(clk),
	.d(\tdl_arr~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][0]~q ),
	.prn(vcc));
defparam \tdl_arr[0][0] .is_wysiwyg = "true";
defparam \tdl_arr[0][0] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~6 (
	.dataa(reset_n),
	.datab(\tdl_arr[0][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~6_combout ),
	.cout());
defparam \tdl_arr~6 .lut_mask = 16'hEEEE;
defparam \tdl_arr~6 .sum_lutc_input = "datac";

dffeas \tdl_arr[1][0] (
	.clk(clk),
	.d(\tdl_arr~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[1][0]~q ),
	.prn(vcc));
defparam \tdl_arr[1][0] .is_wysiwyg = "true";
defparam \tdl_arr[1][0] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~4 (
	.dataa(reset_n),
	.datab(\tdl_arr[1][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~4_combout ),
	.cout());
defparam \tdl_arr~4 .lut_mask = 16'hEEEE;
defparam \tdl_arr~4 .sum_lutc_input = "datac";

dffeas \tdl_arr[2][0] (
	.clk(clk),
	.d(\tdl_arr~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[2][0]~q ),
	.prn(vcc));
defparam \tdl_arr[2][0] .is_wysiwyg = "true";
defparam \tdl_arr[2][0] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~2 (
	.dataa(reset_n),
	.datab(\tdl_arr[2][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~2_combout ),
	.cout());
defparam \tdl_arr~2 .lut_mask = 16'hEEEE;
defparam \tdl_arr~2 .sum_lutc_input = "datac";

dffeas \tdl_arr[3][0] (
	.clk(clk),
	.d(\tdl_arr~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[3][0]~q ),
	.prn(vcc));
defparam \tdl_arr[3][0] .is_wysiwyg = "true";
defparam \tdl_arr[3][0] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~0 (
	.dataa(reset_n),
	.datab(\tdl_arr[3][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~0_combout ),
	.cout());
defparam \tdl_arr~0 .lut_mask = 16'hEEEE;
defparam \tdl_arr~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \tdl_arr~9 (
	.dataa(reset_n),
	.datab(sw_1),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~9_combout ),
	.cout());
defparam \tdl_arr~9 .lut_mask = 16'hEEEE;
defparam \tdl_arr~9 .sum_lutc_input = "datac";

dffeas \tdl_arr[0][1] (
	.clk(clk),
	.d(\tdl_arr~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][1]~q ),
	.prn(vcc));
defparam \tdl_arr[0][1] .is_wysiwyg = "true";
defparam \tdl_arr[0][1] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~7 (
	.dataa(reset_n),
	.datab(\tdl_arr[0][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~7_combout ),
	.cout());
defparam \tdl_arr~7 .lut_mask = 16'hEEEE;
defparam \tdl_arr~7 .sum_lutc_input = "datac";

dffeas \tdl_arr[1][1] (
	.clk(clk),
	.d(\tdl_arr~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[1][1]~q ),
	.prn(vcc));
defparam \tdl_arr[1][1] .is_wysiwyg = "true";
defparam \tdl_arr[1][1] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~5 (
	.dataa(reset_n),
	.datab(\tdl_arr[1][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~5_combout ),
	.cout());
defparam \tdl_arr~5 .lut_mask = 16'hEEEE;
defparam \tdl_arr~5 .sum_lutc_input = "datac";

dffeas \tdl_arr[2][1] (
	.clk(clk),
	.d(\tdl_arr~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[2][1]~q ),
	.prn(vcc));
defparam \tdl_arr[2][1] .is_wysiwyg = "true";
defparam \tdl_arr[2][1] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~3 (
	.dataa(reset_n),
	.datab(\tdl_arr[2][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~3_combout ),
	.cout());
defparam \tdl_arr~3 .lut_mask = 16'hEEEE;
defparam \tdl_arr~3 .sum_lutc_input = "datac";

dffeas \tdl_arr[3][1] (
	.clk(clk),
	.d(\tdl_arr~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[3][1]~q ),
	.prn(vcc));
defparam \tdl_arr[3][1] .is_wysiwyg = "true";
defparam \tdl_arr[3][1] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~1 (
	.dataa(reset_n),
	.datab(\tdl_arr[3][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~1_combout ),
	.cout());
defparam \tdl_arr~1 .lut_mask = 16'hEEEE;
defparam \tdl_arr~1 .sum_lutc_input = "datac";

endmodule

module fft_asj_fft_m_k_counter_fft_120 (
	blk_done_int1,
	source_valid_ctrl_sop,
	stall_reg,
	source_stall_int_d,
	global_clock_enable,
	p_2,
	p_0,
	p_1,
	tdl_arr_4,
	data_rdy_vec_4,
	next_pass_i1,
	Equal0,
	tdl_arr_3,
	k_count_0,
	k_count_2,
	k_count_4,
	k_count_1,
	k_count_3,
	k_count_5,
	k_count_6,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	blk_done_int1;
input 	source_valid_ctrl_sop;
input 	stall_reg;
input 	source_stall_int_d;
input 	global_clock_enable;
output 	p_2;
output 	p_0;
output 	p_1;
input 	tdl_arr_4;
input 	data_rdy_vec_4;
output 	next_pass_i1;
output 	Equal0;
input 	tdl_arr_3;
output 	k_count_0;
output 	k_count_2;
output 	k_count_4;
output 	k_count_1;
output 	k_count_3;
output 	k_count_5;
output 	k_count_6;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Equal1~0_combout ;
wire \k_state.HOLD~q ;
wire \Selector1~0_combout ;
wire \Selector0~0_combout ;
wire \k[0]~8 ;
wire \k[1]~10 ;
wire \k[2]~14 ;
wire \k[3]~16 ;
wire \k[4]~17_combout ;
wire \cnt_k~0_combout ;
wire \fsm~0_combout ;
wire \k_state.IDLE~0_combout ;
wire \k_state.IDLE~q ;
wire \k[0]~11_combout ;
wire \k[0]~12_combout ;
wire \k[4]~q ;
wire \k[4]~18 ;
wire \k[5]~19_combout ;
wire \k[5]~q ;
wire \k[5]~20 ;
wire \k[6]~21_combout ;
wire \k[6]~q ;
wire \Equal1~1_combout ;
wire \Selector1~1_combout ;
wire \Selector1~2_combout ;
wire \k_state.RUN_CNT~q ;
wire \k_state~8_combout ;
wire \k_state.NEXT_PASS_UPD~q ;
wire \blk_done_int~0_combout ;
wire \p[0]~4_combout ;
wire \p~5_combout ;
wire \p[0]~6_combout ;
wire \p~7_combout ;
wire \p~8_combout ;
wire \next_pass_i~0_combout ;
wire \k[0]~7_combout ;
wire \k[0]~q ;
wire \k[2]~13_combout ;
wire \k[2]~q ;
wire \k[1]~9_combout ;
wire \k[1]~q ;
wire \k[3]~15_combout ;
wire \k[3]~q ;


cycloneiii_lcell_comb \Equal1~0 (
	.dataa(\k[1]~q ),
	.datab(\k[2]~q ),
	.datac(\k[3]~q ),
	.datad(\k[0]~q ),
	.cin(gnd),
	.combout(\Equal1~0_combout ),
	.cout());
defparam \Equal1~0 .lut_mask = 16'hFEFF;
defparam \Equal1~0 .sum_lutc_input = "datac";

dffeas \k_state.HOLD (
	.clk(clk),
	.d(\next_pass_i~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\k_state.HOLD~q ),
	.prn(vcc));
defparam \k_state.HOLD .is_wysiwyg = "true";
defparam \k_state.HOLD .power_up = "low";

cycloneiii_lcell_comb \Selector1~0 (
	.dataa(\k_state.HOLD~q ),
	.datab(next_pass_i1),
	.datac(Equal0),
	.datad(\fsm~0_combout ),
	.cin(gnd),
	.combout(\Selector1~0_combout ),
	.cout());
defparam \Selector1~0 .lut_mask = 16'hACFF;
defparam \Selector1~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector0~0 (
	.dataa(\k_state.HOLD~q ),
	.datab(\fsm~0_combout ),
	.datac(Equal0),
	.datad(next_pass_i1),
	.cin(gnd),
	.combout(\Selector0~0_combout ),
	.cout());
defparam \Selector0~0 .lut_mask = 16'hACFF;
defparam \Selector0~0 .sum_lutc_input = "datac";

dffeas blk_done_int(
	.clk(clk),
	.d(\blk_done_int~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(blk_done_int1),
	.prn(vcc));
defparam blk_done_int.is_wysiwyg = "true";
defparam blk_done_int.power_up = "low";

dffeas \p[2] (
	.clk(clk),
	.d(\p~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\p[0]~6_combout ),
	.q(p_2),
	.prn(vcc));
defparam \p[2] .is_wysiwyg = "true";
defparam \p[2] .power_up = "low";

dffeas \p[0] (
	.clk(clk),
	.d(\p~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\p[0]~6_combout ),
	.q(p_0),
	.prn(vcc));
defparam \p[0] .is_wysiwyg = "true";
defparam \p[0] .power_up = "low";

dffeas \p[1] (
	.clk(clk),
	.d(\p~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\p[0]~6_combout ),
	.q(p_1),
	.prn(vcc));
defparam \p[1] .is_wysiwyg = "true";
defparam \p[1] .power_up = "low";

dffeas next_pass_i(
	.clk(clk),
	.d(\next_pass_i~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(next_pass_i1),
	.prn(vcc));
defparam next_pass_i.is_wysiwyg = "true";
defparam next_pass_i.power_up = "low";

cycloneiii_lcell_comb \Equal0~0 (
	.dataa(p_2),
	.datab(gnd),
	.datac(p_0),
	.datad(p_1),
	.cin(gnd),
	.combout(Equal0),
	.cout());
defparam \Equal0~0 .lut_mask = 16'hAFFF;
defparam \Equal0~0 .sum_lutc_input = "datac";

dffeas \k_count[0] (
	.clk(clk),
	.d(\k[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(k_count_0),
	.prn(vcc));
defparam \k_count[0] .is_wysiwyg = "true";
defparam \k_count[0] .power_up = "low";

dffeas \k_count[2] (
	.clk(clk),
	.d(\k[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(k_count_2),
	.prn(vcc));
defparam \k_count[2] .is_wysiwyg = "true";
defparam \k_count[2] .power_up = "low";

dffeas \k_count[4] (
	.clk(clk),
	.d(\k[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(k_count_4),
	.prn(vcc));
defparam \k_count[4] .is_wysiwyg = "true";
defparam \k_count[4] .power_up = "low";

dffeas \k_count[1] (
	.clk(clk),
	.d(\k[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(k_count_1),
	.prn(vcc));
defparam \k_count[1] .is_wysiwyg = "true";
defparam \k_count[1] .power_up = "low";

dffeas \k_count[3] (
	.clk(clk),
	.d(\k[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(k_count_3),
	.prn(vcc));
defparam \k_count[3] .is_wysiwyg = "true";
defparam \k_count[3] .power_up = "low";

dffeas \k_count[5] (
	.clk(clk),
	.d(\k[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(k_count_5),
	.prn(vcc));
defparam \k_count[5] .is_wysiwyg = "true";
defparam \k_count[5] .power_up = "low";

dffeas \k_count[6] (
	.clk(clk),
	.d(\k[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(k_count_6),
	.prn(vcc));
defparam \k_count[6] .is_wysiwyg = "true";
defparam \k_count[6] .power_up = "low";

cycloneiii_lcell_comb \k[0]~7 (
	.dataa(\k[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\k[0]~7_combout ),
	.cout(\k[0]~8 ));
defparam \k[0]~7 .lut_mask = 16'h55AA;
defparam \k[0]~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \k[1]~9 (
	.dataa(\k[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\k[0]~8 ),
	.combout(\k[1]~9_combout ),
	.cout(\k[1]~10 ));
defparam \k[1]~9 .lut_mask = 16'h5A5F;
defparam \k[1]~9 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \k[2]~13 (
	.dataa(\k[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\k[1]~10 ),
	.combout(\k[2]~13_combout ),
	.cout(\k[2]~14 ));
defparam \k[2]~13 .lut_mask = 16'h5AAF;
defparam \k[2]~13 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \k[3]~15 (
	.dataa(\k[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\k[2]~14 ),
	.combout(\k[3]~15_combout ),
	.cout(\k[3]~16 ));
defparam \k[3]~15 .lut_mask = 16'h5A5F;
defparam \k[3]~15 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \k[4]~17 (
	.dataa(\k[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\k[3]~16 ),
	.combout(\k[4]~17_combout ),
	.cout(\k[4]~18 ));
defparam \k[4]~17 .lut_mask = 16'h5AAF;
defparam \k[4]~17 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \cnt_k~0 (
	.dataa(tdl_arr_3),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\cnt_k~0_combout ),
	.cout());
defparam \cnt_k~0 .lut_mask = 16'hAAFF;
defparam \cnt_k~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \fsm~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(tdl_arr_4),
	.datad(tdl_arr_3),
	.cin(gnd),
	.combout(\fsm~0_combout ),
	.cout());
defparam \fsm~0 .lut_mask = 16'h0FFF;
defparam \fsm~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \k_state.IDLE~0 (
	.dataa(\Selector0~0_combout ),
	.datab(\fsm~0_combout ),
	.datac(\k_state.IDLE~q ),
	.datad(reset_n),
	.cin(gnd),
	.combout(\k_state.IDLE~0_combout ),
	.cout());
defparam \k_state.IDLE~0 .lut_mask = 16'hFFF7;
defparam \k_state.IDLE~0 .sum_lutc_input = "datac";

dffeas \k_state.IDLE (
	.clk(clk),
	.d(\k_state.IDLE~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\k_state.IDLE~q ),
	.prn(vcc));
defparam \k_state.IDLE .is_wysiwyg = "true";
defparam \k_state.IDLE .power_up = "low";

cycloneiii_lcell_comb \k[0]~11 (
	.dataa(tdl_arr_3),
	.datab(\k_state.IDLE~q ),
	.datac(reset_n),
	.datad(gnd),
	.cin(gnd),
	.combout(\k[0]~11_combout ),
	.cout());
defparam \k[0]~11 .lut_mask = 16'hEFEF;
defparam \k[0]~11 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \k[0]~12 (
	.dataa(source_stall_int_d),
	.datab(source_valid_ctrl_sop),
	.datac(stall_reg),
	.datad(\k[0]~11_combout ),
	.cin(gnd),
	.combout(\k[0]~12_combout ),
	.cout());
defparam \k[0]~12 .lut_mask = 16'hF7D5;
defparam \k[0]~12 .sum_lutc_input = "datac";

dffeas \k[4] (
	.clk(clk),
	.d(\k[4]~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\cnt_k~0_combout ),
	.sload(gnd),
	.ena(\k[0]~12_combout ),
	.q(\k[4]~q ),
	.prn(vcc));
defparam \k[4] .is_wysiwyg = "true";
defparam \k[4] .power_up = "low";

cycloneiii_lcell_comb \k[5]~19 (
	.dataa(\k[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\k[4]~18 ),
	.combout(\k[5]~19_combout ),
	.cout(\k[5]~20 ));
defparam \k[5]~19 .lut_mask = 16'h5A5F;
defparam \k[5]~19 .sum_lutc_input = "cin";

dffeas \k[5] (
	.clk(clk),
	.d(\k[5]~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\cnt_k~0_combout ),
	.sload(gnd),
	.ena(\k[0]~12_combout ),
	.q(\k[5]~q ),
	.prn(vcc));
defparam \k[5] .is_wysiwyg = "true";
defparam \k[5] .power_up = "low";

cycloneiii_lcell_comb \k[6]~21 (
	.dataa(\k[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\k[5]~20 ),
	.combout(\k[6]~21_combout ),
	.cout());
defparam \k[6]~21 .lut_mask = 16'h5A5A;
defparam \k[6]~21 .sum_lutc_input = "cin";

dffeas \k[6] (
	.clk(clk),
	.d(\k[6]~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\cnt_k~0_combout ),
	.sload(gnd),
	.ena(\k[0]~12_combout ),
	.q(\k[6]~q ),
	.prn(vcc));
defparam \k[6] .is_wysiwyg = "true";
defparam \k[6] .power_up = "low";

cycloneiii_lcell_comb \Equal1~1 (
	.dataa(\Equal1~0_combout ),
	.datab(\k[4]~q ),
	.datac(\k[5]~q ),
	.datad(\k[6]~q ),
	.cin(gnd),
	.combout(\Equal1~1_combout ),
	.cout());
defparam \Equal1~1 .lut_mask = 16'hFFFE;
defparam \Equal1~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector1~1 (
	.dataa(tdl_arr_4),
	.datab(tdl_arr_3),
	.datac(gnd),
	.datad(\k_state.IDLE~q ),
	.cin(gnd),
	.combout(\Selector1~1_combout ),
	.cout());
defparam \Selector1~1 .lut_mask = 16'hEEFF;
defparam \Selector1~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector1~2 (
	.dataa(\Selector1~0_combout ),
	.datab(\Selector1~1_combout ),
	.datac(\k_state.RUN_CNT~q ),
	.datad(\Equal1~1_combout ),
	.cin(gnd),
	.combout(\Selector1~2_combout ),
	.cout());
defparam \Selector1~2 .lut_mask = 16'hFEFF;
defparam \Selector1~2 .sum_lutc_input = "datac";

dffeas \k_state.RUN_CNT (
	.clk(clk),
	.d(\Selector1~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\k_state.RUN_CNT~q ),
	.prn(vcc));
defparam \k_state.RUN_CNT .is_wysiwyg = "true";
defparam \k_state.RUN_CNT .power_up = "low";

cycloneiii_lcell_comb \k_state~8 (
	.dataa(reset_n),
	.datab(\Equal1~1_combout ),
	.datac(\k_state.RUN_CNT~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\k_state~8_combout ),
	.cout());
defparam \k_state~8 .lut_mask = 16'hFEFE;
defparam \k_state~8 .sum_lutc_input = "datac";

dffeas \k_state.NEXT_PASS_UPD (
	.clk(clk),
	.d(\k_state~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\k_state.NEXT_PASS_UPD~q ),
	.prn(vcc));
defparam \k_state.NEXT_PASS_UPD .is_wysiwyg = "true";
defparam \k_state.NEXT_PASS_UPD .power_up = "low";

cycloneiii_lcell_comb \blk_done_int~0 (
	.dataa(\k_state.NEXT_PASS_UPD~q ),
	.datab(p_2),
	.datac(p_0),
	.datad(p_1),
	.cin(gnd),
	.combout(\blk_done_int~0_combout ),
	.cout());
defparam \blk_done_int~0 .lut_mask = 16'hEFFF;
defparam \blk_done_int~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \p[0]~4 (
	.dataa(reset_n),
	.datab(gnd),
	.datac(gnd),
	.datad(tdl_arr_4),
	.cin(gnd),
	.combout(\p[0]~4_combout ),
	.cout());
defparam \p[0]~4 .lut_mask = 16'hAAFF;
defparam \p[0]~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \p~5 (
	.dataa(\p[0]~4_combout ),
	.datab(p_0),
	.datac(p_1),
	.datad(p_2),
	.cin(gnd),
	.combout(\p~5_combout ),
	.cout());
defparam \p~5 .lut_mask = 16'hEBBE;
defparam \p~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \p[0]~6 (
	.dataa(global_clock_enable),
	.datab(\p[0]~4_combout ),
	.datac(data_rdy_vec_4),
	.datad(next_pass_i1),
	.cin(gnd),
	.combout(\p[0]~6_combout ),
	.cout());
defparam \p[0]~6 .lut_mask = 16'hFFFB;
defparam \p[0]~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \p~7 (
	.dataa(reset_n),
	.datab(tdl_arr_4),
	.datac(gnd),
	.datad(p_0),
	.cin(gnd),
	.combout(\p~7_combout ),
	.cout());
defparam \p~7 .lut_mask = 16'hEEFF;
defparam \p~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \p~8 (
	.dataa(reset_n),
	.datab(tdl_arr_4),
	.datac(p_0),
	.datad(p_1),
	.cin(gnd),
	.combout(\p~8_combout ),
	.cout());
defparam \p~8 .lut_mask = 16'hBFFB;
defparam \p~8 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \next_pass_i~0 (
	.dataa(reset_n),
	.datab(\k_state.NEXT_PASS_UPD~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\next_pass_i~0_combout ),
	.cout());
defparam \next_pass_i~0 .lut_mask = 16'hEEEE;
defparam \next_pass_i~0 .sum_lutc_input = "datac";

dffeas \k[0] (
	.clk(clk),
	.d(\k[0]~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\cnt_k~0_combout ),
	.sload(gnd),
	.ena(\k[0]~12_combout ),
	.q(\k[0]~q ),
	.prn(vcc));
defparam \k[0] .is_wysiwyg = "true";
defparam \k[0] .power_up = "low";

dffeas \k[2] (
	.clk(clk),
	.d(\k[2]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\cnt_k~0_combout ),
	.sload(gnd),
	.ena(\k[0]~12_combout ),
	.q(\k[2]~q ),
	.prn(vcc));
defparam \k[2] .is_wysiwyg = "true";
defparam \k[2] .power_up = "low";

dffeas \k[1] (
	.clk(clk),
	.d(\k[1]~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\cnt_k~0_combout ),
	.sload(gnd),
	.ena(\k[0]~12_combout ),
	.q(\k[1]~q ),
	.prn(vcc));
defparam \k[1] .is_wysiwyg = "true";
defparam \k[1] .power_up = "low";

dffeas \k[3] (
	.clk(clk),
	.d(\k[3]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\cnt_k~0_combout ),
	.sload(gnd),
	.ena(\k[0]~12_combout ),
	.q(\k[3]~q ),
	.prn(vcc));
defparam \k[3] .is_wysiwyg = "true";
defparam \k[3] .power_up = "low";

endmodule

module fft_asj_fft_tdl_bit_fft_120_4 (
	global_clock_enable,
	tdl_arr_4,
	rd_addr_b_6,
	clk)/* synthesis synthesis_greybox=1 */;
input 	global_clock_enable;
output 	tdl_arr_4;
input 	rd_addr_b_6;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \tdl_arr[0]~0_combout ;
wire \tdl_arr[0]~q ;
wire \tdl_arr[1]~q ;
wire \tdl_arr[2]~q ;
wire \tdl_arr[3]~q ;


dffeas \tdl_arr[4] (
	.clk(clk),
	.d(\tdl_arr[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_4),
	.prn(vcc));
defparam \tdl_arr[4] .is_wysiwyg = "true";
defparam \tdl_arr[4] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr[0]~0 (
	.dataa(rd_addr_b_6),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr[0]~0_combout ),
	.cout());
defparam \tdl_arr[0]~0 .lut_mask = 16'h5555;
defparam \tdl_arr[0]~0 .sum_lutc_input = "datac";

dffeas \tdl_arr[0] (
	.clk(clk),
	.d(\tdl_arr[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0]~q ),
	.prn(vcc));
defparam \tdl_arr[0] .is_wysiwyg = "true";
defparam \tdl_arr[0] .power_up = "low";

dffeas \tdl_arr[1] (
	.clk(clk),
	.d(\tdl_arr[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[1]~q ),
	.prn(vcc));
defparam \tdl_arr[1] .is_wysiwyg = "true";
defparam \tdl_arr[1] .power_up = "low";

dffeas \tdl_arr[2] (
	.clk(clk),
	.d(\tdl_arr[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[2]~q ),
	.prn(vcc));
defparam \tdl_arr[2] .is_wysiwyg = "true";
defparam \tdl_arr[2] .power_up = "low";

dffeas \tdl_arr[3] (
	.clk(clk),
	.d(\tdl_arr[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[3]~q ),
	.prn(vcc));
defparam \tdl_arr[3] .is_wysiwyg = "true";
defparam \tdl_arr[3] .power_up = "low";

endmodule

module fft_asj_fft_tdl_bit_rst_fft_120_3 (
	blk_done_int,
	global_clock_enable,
	tdl_arr_11,
	blk_done_vec_2,
	tdl_arr_5,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	blk_done_int;
input 	global_clock_enable;
output 	tdl_arr_11;
input 	blk_done_vec_2;
output 	tdl_arr_5;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \tdl_arr~2_combout ;
wire \tdl_arr[9]~q ;
wire \tdl_arr~1_combout ;
wire \tdl_arr[10]~q ;
wire \tdl_arr~0_combout ;
wire \tdl_arr~8_combout ;
wire \tdl_arr[0]~q ;
wire \tdl_arr~7_combout ;
wire \tdl_arr[1]~q ;
wire \tdl_arr~6_combout ;
wire \tdl_arr[2]~q ;
wire \tdl_arr~5_combout ;
wire \tdl_arr[3]~q ;
wire \tdl_arr~4_combout ;
wire \tdl_arr[4]~q ;
wire \tdl_arr~3_combout ;


dffeas \tdl_arr[11] (
	.clk(clk),
	.d(\tdl_arr~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_11),
	.prn(vcc));
defparam \tdl_arr[11] .is_wysiwyg = "true";
defparam \tdl_arr[11] .power_up = "low";

dffeas \tdl_arr[5] (
	.clk(clk),
	.d(\tdl_arr~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_5),
	.prn(vcc));
defparam \tdl_arr[5] .is_wysiwyg = "true";
defparam \tdl_arr[5] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~2 (
	.dataa(reset_n),
	.datab(blk_done_vec_2),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~2_combout ),
	.cout());
defparam \tdl_arr~2 .lut_mask = 16'hEEEE;
defparam \tdl_arr~2 .sum_lutc_input = "datac";

dffeas \tdl_arr[9] (
	.clk(clk),
	.d(\tdl_arr~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[9]~q ),
	.prn(vcc));
defparam \tdl_arr[9] .is_wysiwyg = "true";
defparam \tdl_arr[9] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~1 (
	.dataa(reset_n),
	.datab(\tdl_arr[9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~1_combout ),
	.cout());
defparam \tdl_arr~1 .lut_mask = 16'hEEEE;
defparam \tdl_arr~1 .sum_lutc_input = "datac";

dffeas \tdl_arr[10] (
	.clk(clk),
	.d(\tdl_arr~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[10]~q ),
	.prn(vcc));
defparam \tdl_arr[10] .is_wysiwyg = "true";
defparam \tdl_arr[10] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~0 (
	.dataa(reset_n),
	.datab(\tdl_arr[10]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~0_combout ),
	.cout());
defparam \tdl_arr~0 .lut_mask = 16'hEEEE;
defparam \tdl_arr~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \tdl_arr~8 (
	.dataa(reset_n),
	.datab(blk_done_int),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~8_combout ),
	.cout());
defparam \tdl_arr~8 .lut_mask = 16'hEEEE;
defparam \tdl_arr~8 .sum_lutc_input = "datac";

dffeas \tdl_arr[0] (
	.clk(clk),
	.d(\tdl_arr~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0]~q ),
	.prn(vcc));
defparam \tdl_arr[0] .is_wysiwyg = "true";
defparam \tdl_arr[0] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~7 (
	.dataa(reset_n),
	.datab(\tdl_arr[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~7_combout ),
	.cout());
defparam \tdl_arr~7 .lut_mask = 16'hEEEE;
defparam \tdl_arr~7 .sum_lutc_input = "datac";

dffeas \tdl_arr[1] (
	.clk(clk),
	.d(\tdl_arr~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[1]~q ),
	.prn(vcc));
defparam \tdl_arr[1] .is_wysiwyg = "true";
defparam \tdl_arr[1] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~6 (
	.dataa(reset_n),
	.datab(\tdl_arr[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~6_combout ),
	.cout());
defparam \tdl_arr~6 .lut_mask = 16'hEEEE;
defparam \tdl_arr~6 .sum_lutc_input = "datac";

dffeas \tdl_arr[2] (
	.clk(clk),
	.d(\tdl_arr~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[2]~q ),
	.prn(vcc));
defparam \tdl_arr[2] .is_wysiwyg = "true";
defparam \tdl_arr[2] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~5 (
	.dataa(reset_n),
	.datab(\tdl_arr[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~5_combout ),
	.cout());
defparam \tdl_arr~5 .lut_mask = 16'hEEEE;
defparam \tdl_arr~5 .sum_lutc_input = "datac";

dffeas \tdl_arr[3] (
	.clk(clk),
	.d(\tdl_arr~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[3]~q ),
	.prn(vcc));
defparam \tdl_arr[3] .is_wysiwyg = "true";
defparam \tdl_arr[3] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~4 (
	.dataa(reset_n),
	.datab(\tdl_arr[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~4_combout ),
	.cout());
defparam \tdl_arr~4 .lut_mask = 16'hEEEE;
defparam \tdl_arr~4 .sum_lutc_input = "datac";

dffeas \tdl_arr[4] (
	.clk(clk),
	.d(\tdl_arr~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[4]~q ),
	.prn(vcc));
defparam \tdl_arr[4] .is_wysiwyg = "true";
defparam \tdl_arr[4] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~3 (
	.dataa(reset_n),
	.datab(\tdl_arr[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~3_combout ),
	.cout());
defparam \tdl_arr~3 .lut_mask = 16'hEEEE;
defparam \tdl_arr~3 .sum_lutc_input = "datac";

endmodule

module fft_asj_fft_tdl_bit_rst_fft_120_4 (
	global_clock_enable,
	tdl_arr_11,
	tdl_arr_19,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	global_clock_enable;
input 	tdl_arr_11;
output 	tdl_arr_19;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \tdl_arr~19_combout ;
wire \tdl_arr[0]~q ;
wire \tdl_arr~18_combout ;
wire \tdl_arr[1]~q ;
wire \tdl_arr~17_combout ;
wire \tdl_arr[2]~q ;
wire \tdl_arr~16_combout ;
wire \tdl_arr[3]~q ;
wire \tdl_arr~15_combout ;
wire \tdl_arr[4]~q ;
wire \tdl_arr~14_combout ;
wire \tdl_arr[5]~q ;
wire \tdl_arr~13_combout ;
wire \tdl_arr[6]~q ;
wire \tdl_arr~12_combout ;
wire \tdl_arr[7]~q ;
wire \tdl_arr~11_combout ;
wire \tdl_arr[8]~q ;
wire \tdl_arr~10_combout ;
wire \tdl_arr[9]~q ;
wire \tdl_arr~9_combout ;
wire \tdl_arr[10]~q ;
wire \tdl_arr~8_combout ;
wire \tdl_arr[11]~q ;
wire \tdl_arr~7_combout ;
wire \tdl_arr[12]~q ;
wire \tdl_arr~6_combout ;
wire \tdl_arr[13]~q ;
wire \tdl_arr~5_combout ;
wire \tdl_arr[14]~q ;
wire \tdl_arr~4_combout ;
wire \tdl_arr[15]~q ;
wire \tdl_arr~3_combout ;
wire \tdl_arr[16]~q ;
wire \tdl_arr~2_combout ;
wire \tdl_arr[17]~q ;
wire \tdl_arr~1_combout ;
wire \tdl_arr[18]~q ;
wire \tdl_arr~0_combout ;


dffeas \tdl_arr[19] (
	.clk(clk),
	.d(\tdl_arr~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_19),
	.prn(vcc));
defparam \tdl_arr[19] .is_wysiwyg = "true";
defparam \tdl_arr[19] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~19 (
	.dataa(reset_n),
	.datab(tdl_arr_11),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~19_combout ),
	.cout());
defparam \tdl_arr~19 .lut_mask = 16'hEEEE;
defparam \tdl_arr~19 .sum_lutc_input = "datac";

dffeas \tdl_arr[0] (
	.clk(clk),
	.d(\tdl_arr~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0]~q ),
	.prn(vcc));
defparam \tdl_arr[0] .is_wysiwyg = "true";
defparam \tdl_arr[0] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~18 (
	.dataa(reset_n),
	.datab(\tdl_arr[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~18_combout ),
	.cout());
defparam \tdl_arr~18 .lut_mask = 16'hEEEE;
defparam \tdl_arr~18 .sum_lutc_input = "datac";

dffeas \tdl_arr[1] (
	.clk(clk),
	.d(\tdl_arr~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[1]~q ),
	.prn(vcc));
defparam \tdl_arr[1] .is_wysiwyg = "true";
defparam \tdl_arr[1] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~17 (
	.dataa(reset_n),
	.datab(\tdl_arr[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~17_combout ),
	.cout());
defparam \tdl_arr~17 .lut_mask = 16'hEEEE;
defparam \tdl_arr~17 .sum_lutc_input = "datac";

dffeas \tdl_arr[2] (
	.clk(clk),
	.d(\tdl_arr~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[2]~q ),
	.prn(vcc));
defparam \tdl_arr[2] .is_wysiwyg = "true";
defparam \tdl_arr[2] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~16 (
	.dataa(reset_n),
	.datab(\tdl_arr[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~16_combout ),
	.cout());
defparam \tdl_arr~16 .lut_mask = 16'hEEEE;
defparam \tdl_arr~16 .sum_lutc_input = "datac";

dffeas \tdl_arr[3] (
	.clk(clk),
	.d(\tdl_arr~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[3]~q ),
	.prn(vcc));
defparam \tdl_arr[3] .is_wysiwyg = "true";
defparam \tdl_arr[3] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~15 (
	.dataa(reset_n),
	.datab(\tdl_arr[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~15_combout ),
	.cout());
defparam \tdl_arr~15 .lut_mask = 16'hEEEE;
defparam \tdl_arr~15 .sum_lutc_input = "datac";

dffeas \tdl_arr[4] (
	.clk(clk),
	.d(\tdl_arr~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[4]~q ),
	.prn(vcc));
defparam \tdl_arr[4] .is_wysiwyg = "true";
defparam \tdl_arr[4] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~14 (
	.dataa(reset_n),
	.datab(\tdl_arr[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~14_combout ),
	.cout());
defparam \tdl_arr~14 .lut_mask = 16'hEEEE;
defparam \tdl_arr~14 .sum_lutc_input = "datac";

dffeas \tdl_arr[5] (
	.clk(clk),
	.d(\tdl_arr~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[5]~q ),
	.prn(vcc));
defparam \tdl_arr[5] .is_wysiwyg = "true";
defparam \tdl_arr[5] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~13 (
	.dataa(reset_n),
	.datab(\tdl_arr[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~13_combout ),
	.cout());
defparam \tdl_arr~13 .lut_mask = 16'hEEEE;
defparam \tdl_arr~13 .sum_lutc_input = "datac";

dffeas \tdl_arr[6] (
	.clk(clk),
	.d(\tdl_arr~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[6]~q ),
	.prn(vcc));
defparam \tdl_arr[6] .is_wysiwyg = "true";
defparam \tdl_arr[6] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~12 (
	.dataa(reset_n),
	.datab(\tdl_arr[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~12_combout ),
	.cout());
defparam \tdl_arr~12 .lut_mask = 16'hEEEE;
defparam \tdl_arr~12 .sum_lutc_input = "datac";

dffeas \tdl_arr[7] (
	.clk(clk),
	.d(\tdl_arr~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[7]~q ),
	.prn(vcc));
defparam \tdl_arr[7] .is_wysiwyg = "true";
defparam \tdl_arr[7] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~11 (
	.dataa(reset_n),
	.datab(\tdl_arr[7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~11_combout ),
	.cout());
defparam \tdl_arr~11 .lut_mask = 16'hEEEE;
defparam \tdl_arr~11 .sum_lutc_input = "datac";

dffeas \tdl_arr[8] (
	.clk(clk),
	.d(\tdl_arr~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[8]~q ),
	.prn(vcc));
defparam \tdl_arr[8] .is_wysiwyg = "true";
defparam \tdl_arr[8] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~10 (
	.dataa(reset_n),
	.datab(\tdl_arr[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~10_combout ),
	.cout());
defparam \tdl_arr~10 .lut_mask = 16'hEEEE;
defparam \tdl_arr~10 .sum_lutc_input = "datac";

dffeas \tdl_arr[9] (
	.clk(clk),
	.d(\tdl_arr~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[9]~q ),
	.prn(vcc));
defparam \tdl_arr[9] .is_wysiwyg = "true";
defparam \tdl_arr[9] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~9 (
	.dataa(reset_n),
	.datab(\tdl_arr[9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~9_combout ),
	.cout());
defparam \tdl_arr~9 .lut_mask = 16'hEEEE;
defparam \tdl_arr~9 .sum_lutc_input = "datac";

dffeas \tdl_arr[10] (
	.clk(clk),
	.d(\tdl_arr~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[10]~q ),
	.prn(vcc));
defparam \tdl_arr[10] .is_wysiwyg = "true";
defparam \tdl_arr[10] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~8 (
	.dataa(reset_n),
	.datab(\tdl_arr[10]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~8_combout ),
	.cout());
defparam \tdl_arr~8 .lut_mask = 16'hEEEE;
defparam \tdl_arr~8 .sum_lutc_input = "datac";

dffeas \tdl_arr[11] (
	.clk(clk),
	.d(\tdl_arr~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[11]~q ),
	.prn(vcc));
defparam \tdl_arr[11] .is_wysiwyg = "true";
defparam \tdl_arr[11] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~7 (
	.dataa(reset_n),
	.datab(\tdl_arr[11]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~7_combout ),
	.cout());
defparam \tdl_arr~7 .lut_mask = 16'hEEEE;
defparam \tdl_arr~7 .sum_lutc_input = "datac";

dffeas \tdl_arr[12] (
	.clk(clk),
	.d(\tdl_arr~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[12]~q ),
	.prn(vcc));
defparam \tdl_arr[12] .is_wysiwyg = "true";
defparam \tdl_arr[12] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~6 (
	.dataa(reset_n),
	.datab(\tdl_arr[12]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~6_combout ),
	.cout());
defparam \tdl_arr~6 .lut_mask = 16'hEEEE;
defparam \tdl_arr~6 .sum_lutc_input = "datac";

dffeas \tdl_arr[13] (
	.clk(clk),
	.d(\tdl_arr~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[13]~q ),
	.prn(vcc));
defparam \tdl_arr[13] .is_wysiwyg = "true";
defparam \tdl_arr[13] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~5 (
	.dataa(reset_n),
	.datab(\tdl_arr[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~5_combout ),
	.cout());
defparam \tdl_arr~5 .lut_mask = 16'hEEEE;
defparam \tdl_arr~5 .sum_lutc_input = "datac";

dffeas \tdl_arr[14] (
	.clk(clk),
	.d(\tdl_arr~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[14]~q ),
	.prn(vcc));
defparam \tdl_arr[14] .is_wysiwyg = "true";
defparam \tdl_arr[14] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~4 (
	.dataa(reset_n),
	.datab(\tdl_arr[14]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~4_combout ),
	.cout());
defparam \tdl_arr~4 .lut_mask = 16'hEEEE;
defparam \tdl_arr~4 .sum_lutc_input = "datac";

dffeas \tdl_arr[15] (
	.clk(clk),
	.d(\tdl_arr~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[15]~q ),
	.prn(vcc));
defparam \tdl_arr[15] .is_wysiwyg = "true";
defparam \tdl_arr[15] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~3 (
	.dataa(reset_n),
	.datab(\tdl_arr[15]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~3_combout ),
	.cout());
defparam \tdl_arr~3 .lut_mask = 16'hEEEE;
defparam \tdl_arr~3 .sum_lutc_input = "datac";

dffeas \tdl_arr[16] (
	.clk(clk),
	.d(\tdl_arr~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[16]~q ),
	.prn(vcc));
defparam \tdl_arr[16] .is_wysiwyg = "true";
defparam \tdl_arr[16] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~2 (
	.dataa(reset_n),
	.datab(\tdl_arr[16]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~2_combout ),
	.cout());
defparam \tdl_arr~2 .lut_mask = 16'hEEEE;
defparam \tdl_arr~2 .sum_lutc_input = "datac";

dffeas \tdl_arr[17] (
	.clk(clk),
	.d(\tdl_arr~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[17]~q ),
	.prn(vcc));
defparam \tdl_arr[17] .is_wysiwyg = "true";
defparam \tdl_arr[17] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~1 (
	.dataa(reset_n),
	.datab(\tdl_arr[17]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~1_combout ),
	.cout());
defparam \tdl_arr~1 .lut_mask = 16'hEEEE;
defparam \tdl_arr~1 .sum_lutc_input = "datac";

dffeas \tdl_arr[18] (
	.clk(clk),
	.d(\tdl_arr~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[18]~q ),
	.prn(vcc));
defparam \tdl_arr[18] .is_wysiwyg = "true";
defparam \tdl_arr[18] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~0 (
	.dataa(reset_n),
	.datab(\tdl_arr[18]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~0_combout ),
	.cout());
defparam \tdl_arr~0 .lut_mask = 16'hEEEE;
defparam \tdl_arr~0 .sum_lutc_input = "datac";

endmodule

module fft_asj_fft_tdl_bit_rst_fft_120_6 (
	global_clock_enable,
	next_pass_i,
	tdl_arr_5,
	next_pass_vec_2,
	tdl_arr_9,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	global_clock_enable;
input 	next_pass_i;
output 	tdl_arr_5;
input 	next_pass_vec_2;
output 	tdl_arr_9;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \tdl_arr~5_combout ;
wire \tdl_arr[0]~q ;
wire \tdl_arr~4_combout ;
wire \tdl_arr[1]~q ;
wire \tdl_arr~3_combout ;
wire \tdl_arr[2]~q ;
wire \tdl_arr~2_combout ;
wire \tdl_arr[3]~q ;
wire \tdl_arr~1_combout ;
wire \tdl_arr[4]~q ;
wire \tdl_arr~0_combout ;
wire \tdl_arr~6_combout ;


dffeas \tdl_arr[5] (
	.clk(clk),
	.d(\tdl_arr~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_5),
	.prn(vcc));
defparam \tdl_arr[5] .is_wysiwyg = "true";
defparam \tdl_arr[5] .power_up = "low";

dffeas \tdl_arr[9] (
	.clk(clk),
	.d(\tdl_arr~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_9),
	.prn(vcc));
defparam \tdl_arr[9] .is_wysiwyg = "true";
defparam \tdl_arr[9] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~5 (
	.dataa(reset_n),
	.datab(next_pass_i),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~5_combout ),
	.cout());
defparam \tdl_arr~5 .lut_mask = 16'hEEEE;
defparam \tdl_arr~5 .sum_lutc_input = "datac";

dffeas \tdl_arr[0] (
	.clk(clk),
	.d(\tdl_arr~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0]~q ),
	.prn(vcc));
defparam \tdl_arr[0] .is_wysiwyg = "true";
defparam \tdl_arr[0] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~4 (
	.dataa(reset_n),
	.datab(\tdl_arr[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~4_combout ),
	.cout());
defparam \tdl_arr~4 .lut_mask = 16'hEEEE;
defparam \tdl_arr~4 .sum_lutc_input = "datac";

dffeas \tdl_arr[1] (
	.clk(clk),
	.d(\tdl_arr~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[1]~q ),
	.prn(vcc));
defparam \tdl_arr[1] .is_wysiwyg = "true";
defparam \tdl_arr[1] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~3 (
	.dataa(reset_n),
	.datab(\tdl_arr[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~3_combout ),
	.cout());
defparam \tdl_arr~3 .lut_mask = 16'hEEEE;
defparam \tdl_arr~3 .sum_lutc_input = "datac";

dffeas \tdl_arr[2] (
	.clk(clk),
	.d(\tdl_arr~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[2]~q ),
	.prn(vcc));
defparam \tdl_arr[2] .is_wysiwyg = "true";
defparam \tdl_arr[2] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~2 (
	.dataa(reset_n),
	.datab(\tdl_arr[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~2_combout ),
	.cout());
defparam \tdl_arr~2 .lut_mask = 16'hEEEE;
defparam \tdl_arr~2 .sum_lutc_input = "datac";

dffeas \tdl_arr[3] (
	.clk(clk),
	.d(\tdl_arr~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[3]~q ),
	.prn(vcc));
defparam \tdl_arr[3] .is_wysiwyg = "true";
defparam \tdl_arr[3] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~1 (
	.dataa(reset_n),
	.datab(\tdl_arr[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~1_combout ),
	.cout());
defparam \tdl_arr~1 .lut_mask = 16'hEEEE;
defparam \tdl_arr~1 .sum_lutc_input = "datac";

dffeas \tdl_arr[4] (
	.clk(clk),
	.d(\tdl_arr~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[4]~q ),
	.prn(vcc));
defparam \tdl_arr[4] .is_wysiwyg = "true";
defparam \tdl_arr[4] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~0 (
	.dataa(reset_n),
	.datab(\tdl_arr[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~0_combout ),
	.cout());
defparam \tdl_arr~0 .lut_mask = 16'hEEEE;
defparam \tdl_arr~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \tdl_arr~6 (
	.dataa(reset_n),
	.datab(next_pass_vec_2),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~6_combout ),
	.cout());
defparam \tdl_arr~6 .lut_mask = 16'hEEEE;
defparam \tdl_arr~6 .sum_lutc_input = "datac";

endmodule

module fft_asj_fft_tdl_bit_rst_fft_120_7 (
	global_clock_enable,
	tdl_arr_3,
	tdl_arr_4,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	global_clock_enable;
output 	tdl_arr_3;
input 	tdl_arr_4;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \tdl_arr~3_combout ;
wire \tdl_arr[0]~q ;
wire \tdl_arr~2_combout ;
wire \tdl_arr[1]~q ;
wire \tdl_arr~1_combout ;
wire \tdl_arr[2]~q ;
wire \tdl_arr~0_combout ;


dffeas \tdl_arr[3] (
	.clk(clk),
	.d(\tdl_arr~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_3),
	.prn(vcc));
defparam \tdl_arr[3] .is_wysiwyg = "true";
defparam \tdl_arr[3] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~3 (
	.dataa(reset_n),
	.datab(tdl_arr_4),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~3_combout ),
	.cout());
defparam \tdl_arr~3 .lut_mask = 16'hEEEE;
defparam \tdl_arr~3 .sum_lutc_input = "datac";

dffeas \tdl_arr[0] (
	.clk(clk),
	.d(\tdl_arr~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0]~q ),
	.prn(vcc));
defparam \tdl_arr[0] .is_wysiwyg = "true";
defparam \tdl_arr[0] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~2 (
	.dataa(reset_n),
	.datab(\tdl_arr[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~2_combout ),
	.cout());
defparam \tdl_arr~2 .lut_mask = 16'hEEEE;
defparam \tdl_arr~2 .sum_lutc_input = "datac";

dffeas \tdl_arr[1] (
	.clk(clk),
	.d(\tdl_arr~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[1]~q ),
	.prn(vcc));
defparam \tdl_arr[1] .is_wysiwyg = "true";
defparam \tdl_arr[1] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~1 (
	.dataa(reset_n),
	.datab(\tdl_arr[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~1_combout ),
	.cout());
defparam \tdl_arr~1 .lut_mask = 16'hEEEE;
defparam \tdl_arr~1 .sum_lutc_input = "datac";

dffeas \tdl_arr[2] (
	.clk(clk),
	.d(\tdl_arr~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[2]~q ),
	.prn(vcc));
defparam \tdl_arr[2] .is_wysiwyg = "true";
defparam \tdl_arr[2] .power_up = "low";

cycloneiii_lcell_comb \tdl_arr~0 (
	.dataa(reset_n),
	.datab(\tdl_arr[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~0_combout ),
	.cout());
defparam \tdl_arr~0 .lut_mask = 16'hEEEE;
defparam \tdl_arr~0 .sum_lutc_input = "datac";

endmodule

module fft_asj_fft_tdl_fft_120 (
	global_clock_enable,
	tdl_arr_4_20,
	tdl_arr_6_20,
	tdl_arr_0_20,
	tdl_arr_2_20,
	tdl_arr_1_20,
	tdl_arr_3_20,
	tdl_arr_5_20,
	tdl_arr_6_1,
	data_in,
	clk)/* synthesis synthesis_greybox=1 */;
input 	global_clock_enable;
output 	tdl_arr_4_20;
output 	tdl_arr_6_20;
output 	tdl_arr_0_20;
output 	tdl_arr_2_20;
output 	tdl_arr_1_20;
output 	tdl_arr_3_20;
output 	tdl_arr_5_20;
output 	tdl_arr_6_1;
input 	[6:0] data_in;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \tdl_arr[0][4]~q ;
wire \tdl_arr[1][4]~q ;
wire \tdl_arr[2][4]~q ;
wire \tdl_arr[3][4]~q ;
wire \tdl_arr[4][4]~q ;
wire \tdl_arr[5][4]~q ;
wire \tdl_arr[6][4]~q ;
wire \tdl_arr[7][4]~q ;
wire \tdl_arr[8][4]~q ;
wire \tdl_arr[9][4]~q ;
wire \tdl_arr[10][4]~q ;
wire \tdl_arr[11][4]~q ;
wire \tdl_arr[12][4]~q ;
wire \tdl_arr[13][4]~q ;
wire \tdl_arr[14][4]~q ;
wire \tdl_arr[15][4]~q ;
wire \tdl_arr[16][4]~q ;
wire \tdl_arr[17][4]~q ;
wire \tdl_arr[18][4]~q ;
wire \tdl_arr[19][4]~q ;
wire \tdl_arr[2][6]~q ;
wire \tdl_arr[3][6]~q ;
wire \tdl_arr[4][6]~q ;
wire \tdl_arr[5][6]~q ;
wire \tdl_arr[6][6]~q ;
wire \tdl_arr[7][6]~q ;
wire \tdl_arr[8][6]~q ;
wire \tdl_arr[9][6]~q ;
wire \tdl_arr[10][6]~q ;
wire \tdl_arr[11][6]~q ;
wire \tdl_arr[12][6]~q ;
wire \tdl_arr[13][6]~q ;
wire \tdl_arr[14][6]~q ;
wire \tdl_arr[15][6]~q ;
wire \tdl_arr[16][6]~q ;
wire \tdl_arr[17][6]~q ;
wire \tdl_arr[18][6]~q ;
wire \tdl_arr[19][6]~q ;
wire \tdl_arr[0][0]~q ;
wire \tdl_arr[1][0]~q ;
wire \tdl_arr[2][0]~q ;
wire \tdl_arr[3][0]~q ;
wire \tdl_arr[4][0]~q ;
wire \tdl_arr[5][0]~q ;
wire \tdl_arr[6][0]~q ;
wire \tdl_arr[7][0]~q ;
wire \tdl_arr[8][0]~q ;
wire \tdl_arr[9][0]~q ;
wire \tdl_arr[10][0]~q ;
wire \tdl_arr[11][0]~q ;
wire \tdl_arr[12][0]~q ;
wire \tdl_arr[13][0]~q ;
wire \tdl_arr[14][0]~q ;
wire \tdl_arr[15][0]~q ;
wire \tdl_arr[16][0]~q ;
wire \tdl_arr[17][0]~q ;
wire \tdl_arr[18][0]~q ;
wire \tdl_arr[19][0]~q ;
wire \tdl_arr[0][2]~q ;
wire \tdl_arr[1][2]~q ;
wire \tdl_arr[2][2]~q ;
wire \tdl_arr[3][2]~q ;
wire \tdl_arr[4][2]~q ;
wire \tdl_arr[5][2]~q ;
wire \tdl_arr[6][2]~q ;
wire \tdl_arr[7][2]~q ;
wire \tdl_arr[8][2]~q ;
wire \tdl_arr[9][2]~q ;
wire \tdl_arr[10][2]~q ;
wire \tdl_arr[11][2]~q ;
wire \tdl_arr[12][2]~q ;
wire \tdl_arr[13][2]~q ;
wire \tdl_arr[14][2]~q ;
wire \tdl_arr[15][2]~q ;
wire \tdl_arr[16][2]~q ;
wire \tdl_arr[17][2]~q ;
wire \tdl_arr[18][2]~q ;
wire \tdl_arr[19][2]~q ;
wire \tdl_arr[0][1]~q ;
wire \tdl_arr[1][1]~q ;
wire \tdl_arr[2][1]~q ;
wire \tdl_arr[3][1]~q ;
wire \tdl_arr[4][1]~q ;
wire \tdl_arr[5][1]~q ;
wire \tdl_arr[6][1]~q ;
wire \tdl_arr[7][1]~q ;
wire \tdl_arr[8][1]~q ;
wire \tdl_arr[9][1]~q ;
wire \tdl_arr[10][1]~q ;
wire \tdl_arr[11][1]~q ;
wire \tdl_arr[12][1]~q ;
wire \tdl_arr[13][1]~q ;
wire \tdl_arr[14][1]~q ;
wire \tdl_arr[15][1]~q ;
wire \tdl_arr[16][1]~q ;
wire \tdl_arr[17][1]~q ;
wire \tdl_arr[18][1]~q ;
wire \tdl_arr[19][1]~q ;
wire \tdl_arr[0][3]~q ;
wire \tdl_arr[1][3]~q ;
wire \tdl_arr[2][3]~q ;
wire \tdl_arr[3][3]~q ;
wire \tdl_arr[4][3]~q ;
wire \tdl_arr[5][3]~q ;
wire \tdl_arr[6][3]~q ;
wire \tdl_arr[7][3]~q ;
wire \tdl_arr[8][3]~q ;
wire \tdl_arr[9][3]~q ;
wire \tdl_arr[10][3]~q ;
wire \tdl_arr[11][3]~q ;
wire \tdl_arr[12][3]~q ;
wire \tdl_arr[13][3]~q ;
wire \tdl_arr[14][3]~q ;
wire \tdl_arr[15][3]~q ;
wire \tdl_arr[16][3]~q ;
wire \tdl_arr[17][3]~q ;
wire \tdl_arr[18][3]~q ;
wire \tdl_arr[19][3]~q ;
wire \tdl_arr[0][5]~q ;
wire \tdl_arr[1][5]~q ;
wire \tdl_arr[2][5]~q ;
wire \tdl_arr[3][5]~q ;
wire \tdl_arr[4][5]~q ;
wire \tdl_arr[5][5]~q ;
wire \tdl_arr[6][5]~q ;
wire \tdl_arr[7][5]~q ;
wire \tdl_arr[8][5]~q ;
wire \tdl_arr[9][5]~q ;
wire \tdl_arr[10][5]~q ;
wire \tdl_arr[11][5]~q ;
wire \tdl_arr[12][5]~q ;
wire \tdl_arr[13][5]~q ;
wire \tdl_arr[14][5]~q ;
wire \tdl_arr[15][5]~q ;
wire \tdl_arr[16][5]~q ;
wire \tdl_arr[17][5]~q ;
wire \tdl_arr[18][5]~q ;
wire \tdl_arr[19][5]~q ;
wire \tdl_arr[0][6]~q ;


dffeas \tdl_arr[20][4] (
	.clk(clk),
	.d(\tdl_arr[19][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_4_20),
	.prn(vcc));
defparam \tdl_arr[20][4] .is_wysiwyg = "true";
defparam \tdl_arr[20][4] .power_up = "low";

dffeas \tdl_arr[20][6] (
	.clk(clk),
	.d(\tdl_arr[19][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_6_20),
	.prn(vcc));
defparam \tdl_arr[20][6] .is_wysiwyg = "true";
defparam \tdl_arr[20][6] .power_up = "low";

dffeas \tdl_arr[20][0] (
	.clk(clk),
	.d(\tdl_arr[19][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_0_20),
	.prn(vcc));
defparam \tdl_arr[20][0] .is_wysiwyg = "true";
defparam \tdl_arr[20][0] .power_up = "low";

dffeas \tdl_arr[20][2] (
	.clk(clk),
	.d(\tdl_arr[19][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_2_20),
	.prn(vcc));
defparam \tdl_arr[20][2] .is_wysiwyg = "true";
defparam \tdl_arr[20][2] .power_up = "low";

dffeas \tdl_arr[20][1] (
	.clk(clk),
	.d(\tdl_arr[19][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_1_20),
	.prn(vcc));
defparam \tdl_arr[20][1] .is_wysiwyg = "true";
defparam \tdl_arr[20][1] .power_up = "low";

dffeas \tdl_arr[20][3] (
	.clk(clk),
	.d(\tdl_arr[19][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_3_20),
	.prn(vcc));
defparam \tdl_arr[20][3] .is_wysiwyg = "true";
defparam \tdl_arr[20][3] .power_up = "low";

dffeas \tdl_arr[20][5] (
	.clk(clk),
	.d(\tdl_arr[19][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_5_20),
	.prn(vcc));
defparam \tdl_arr[20][5] .is_wysiwyg = "true";
defparam \tdl_arr[20][5] .power_up = "low";

dffeas \tdl_arr[1][6] (
	.clk(clk),
	.d(\tdl_arr[0][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_6_1),
	.prn(vcc));
defparam \tdl_arr[1][6] .is_wysiwyg = "true";
defparam \tdl_arr[1][6] .power_up = "low";

dffeas \tdl_arr[0][4] (
	.clk(clk),
	.d(data_in[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][4]~q ),
	.prn(vcc));
defparam \tdl_arr[0][4] .is_wysiwyg = "true";
defparam \tdl_arr[0][4] .power_up = "low";

dffeas \tdl_arr[1][4] (
	.clk(clk),
	.d(\tdl_arr[0][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[1][4]~q ),
	.prn(vcc));
defparam \tdl_arr[1][4] .is_wysiwyg = "true";
defparam \tdl_arr[1][4] .power_up = "low";

dffeas \tdl_arr[2][4] (
	.clk(clk),
	.d(\tdl_arr[1][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[2][4]~q ),
	.prn(vcc));
defparam \tdl_arr[2][4] .is_wysiwyg = "true";
defparam \tdl_arr[2][4] .power_up = "low";

dffeas \tdl_arr[3][4] (
	.clk(clk),
	.d(\tdl_arr[2][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[3][4]~q ),
	.prn(vcc));
defparam \tdl_arr[3][4] .is_wysiwyg = "true";
defparam \tdl_arr[3][4] .power_up = "low";

dffeas \tdl_arr[4][4] (
	.clk(clk),
	.d(\tdl_arr[3][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[4][4]~q ),
	.prn(vcc));
defparam \tdl_arr[4][4] .is_wysiwyg = "true";
defparam \tdl_arr[4][4] .power_up = "low";

dffeas \tdl_arr[5][4] (
	.clk(clk),
	.d(\tdl_arr[4][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[5][4]~q ),
	.prn(vcc));
defparam \tdl_arr[5][4] .is_wysiwyg = "true";
defparam \tdl_arr[5][4] .power_up = "low";

dffeas \tdl_arr[6][4] (
	.clk(clk),
	.d(\tdl_arr[5][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[6][4]~q ),
	.prn(vcc));
defparam \tdl_arr[6][4] .is_wysiwyg = "true";
defparam \tdl_arr[6][4] .power_up = "low";

dffeas \tdl_arr[7][4] (
	.clk(clk),
	.d(\tdl_arr[6][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[7][4]~q ),
	.prn(vcc));
defparam \tdl_arr[7][4] .is_wysiwyg = "true";
defparam \tdl_arr[7][4] .power_up = "low";

dffeas \tdl_arr[8][4] (
	.clk(clk),
	.d(\tdl_arr[7][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[8][4]~q ),
	.prn(vcc));
defparam \tdl_arr[8][4] .is_wysiwyg = "true";
defparam \tdl_arr[8][4] .power_up = "low";

dffeas \tdl_arr[9][4] (
	.clk(clk),
	.d(\tdl_arr[8][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[9][4]~q ),
	.prn(vcc));
defparam \tdl_arr[9][4] .is_wysiwyg = "true";
defparam \tdl_arr[9][4] .power_up = "low";

dffeas \tdl_arr[10][4] (
	.clk(clk),
	.d(\tdl_arr[9][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[10][4]~q ),
	.prn(vcc));
defparam \tdl_arr[10][4] .is_wysiwyg = "true";
defparam \tdl_arr[10][4] .power_up = "low";

dffeas \tdl_arr[11][4] (
	.clk(clk),
	.d(\tdl_arr[10][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[11][4]~q ),
	.prn(vcc));
defparam \tdl_arr[11][4] .is_wysiwyg = "true";
defparam \tdl_arr[11][4] .power_up = "low";

dffeas \tdl_arr[12][4] (
	.clk(clk),
	.d(\tdl_arr[11][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[12][4]~q ),
	.prn(vcc));
defparam \tdl_arr[12][4] .is_wysiwyg = "true";
defparam \tdl_arr[12][4] .power_up = "low";

dffeas \tdl_arr[13][4] (
	.clk(clk),
	.d(\tdl_arr[12][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[13][4]~q ),
	.prn(vcc));
defparam \tdl_arr[13][4] .is_wysiwyg = "true";
defparam \tdl_arr[13][4] .power_up = "low";

dffeas \tdl_arr[14][4] (
	.clk(clk),
	.d(\tdl_arr[13][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[14][4]~q ),
	.prn(vcc));
defparam \tdl_arr[14][4] .is_wysiwyg = "true";
defparam \tdl_arr[14][4] .power_up = "low";

dffeas \tdl_arr[15][4] (
	.clk(clk),
	.d(\tdl_arr[14][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[15][4]~q ),
	.prn(vcc));
defparam \tdl_arr[15][4] .is_wysiwyg = "true";
defparam \tdl_arr[15][4] .power_up = "low";

dffeas \tdl_arr[16][4] (
	.clk(clk),
	.d(\tdl_arr[15][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[16][4]~q ),
	.prn(vcc));
defparam \tdl_arr[16][4] .is_wysiwyg = "true";
defparam \tdl_arr[16][4] .power_up = "low";

dffeas \tdl_arr[17][4] (
	.clk(clk),
	.d(\tdl_arr[16][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[17][4]~q ),
	.prn(vcc));
defparam \tdl_arr[17][4] .is_wysiwyg = "true";
defparam \tdl_arr[17][4] .power_up = "low";

dffeas \tdl_arr[18][4] (
	.clk(clk),
	.d(\tdl_arr[17][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[18][4]~q ),
	.prn(vcc));
defparam \tdl_arr[18][4] .is_wysiwyg = "true";
defparam \tdl_arr[18][4] .power_up = "low";

dffeas \tdl_arr[19][4] (
	.clk(clk),
	.d(\tdl_arr[18][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[19][4]~q ),
	.prn(vcc));
defparam \tdl_arr[19][4] .is_wysiwyg = "true";
defparam \tdl_arr[19][4] .power_up = "low";

dffeas \tdl_arr[2][6] (
	.clk(clk),
	.d(tdl_arr_6_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[2][6]~q ),
	.prn(vcc));
defparam \tdl_arr[2][6] .is_wysiwyg = "true";
defparam \tdl_arr[2][6] .power_up = "low";

dffeas \tdl_arr[3][6] (
	.clk(clk),
	.d(\tdl_arr[2][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[3][6]~q ),
	.prn(vcc));
defparam \tdl_arr[3][6] .is_wysiwyg = "true";
defparam \tdl_arr[3][6] .power_up = "low";

dffeas \tdl_arr[4][6] (
	.clk(clk),
	.d(\tdl_arr[3][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[4][6]~q ),
	.prn(vcc));
defparam \tdl_arr[4][6] .is_wysiwyg = "true";
defparam \tdl_arr[4][6] .power_up = "low";

dffeas \tdl_arr[5][6] (
	.clk(clk),
	.d(\tdl_arr[4][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[5][6]~q ),
	.prn(vcc));
defparam \tdl_arr[5][6] .is_wysiwyg = "true";
defparam \tdl_arr[5][6] .power_up = "low";

dffeas \tdl_arr[6][6] (
	.clk(clk),
	.d(\tdl_arr[5][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[6][6]~q ),
	.prn(vcc));
defparam \tdl_arr[6][6] .is_wysiwyg = "true";
defparam \tdl_arr[6][6] .power_up = "low";

dffeas \tdl_arr[7][6] (
	.clk(clk),
	.d(\tdl_arr[6][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[7][6]~q ),
	.prn(vcc));
defparam \tdl_arr[7][6] .is_wysiwyg = "true";
defparam \tdl_arr[7][6] .power_up = "low";

dffeas \tdl_arr[8][6] (
	.clk(clk),
	.d(\tdl_arr[7][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[8][6]~q ),
	.prn(vcc));
defparam \tdl_arr[8][6] .is_wysiwyg = "true";
defparam \tdl_arr[8][6] .power_up = "low";

dffeas \tdl_arr[9][6] (
	.clk(clk),
	.d(\tdl_arr[8][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[9][6]~q ),
	.prn(vcc));
defparam \tdl_arr[9][6] .is_wysiwyg = "true";
defparam \tdl_arr[9][6] .power_up = "low";

dffeas \tdl_arr[10][6] (
	.clk(clk),
	.d(\tdl_arr[9][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[10][6]~q ),
	.prn(vcc));
defparam \tdl_arr[10][6] .is_wysiwyg = "true";
defparam \tdl_arr[10][6] .power_up = "low";

dffeas \tdl_arr[11][6] (
	.clk(clk),
	.d(\tdl_arr[10][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[11][6]~q ),
	.prn(vcc));
defparam \tdl_arr[11][6] .is_wysiwyg = "true";
defparam \tdl_arr[11][6] .power_up = "low";

dffeas \tdl_arr[12][6] (
	.clk(clk),
	.d(\tdl_arr[11][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[12][6]~q ),
	.prn(vcc));
defparam \tdl_arr[12][6] .is_wysiwyg = "true";
defparam \tdl_arr[12][6] .power_up = "low";

dffeas \tdl_arr[13][6] (
	.clk(clk),
	.d(\tdl_arr[12][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[13][6]~q ),
	.prn(vcc));
defparam \tdl_arr[13][6] .is_wysiwyg = "true";
defparam \tdl_arr[13][6] .power_up = "low";

dffeas \tdl_arr[14][6] (
	.clk(clk),
	.d(\tdl_arr[13][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[14][6]~q ),
	.prn(vcc));
defparam \tdl_arr[14][6] .is_wysiwyg = "true";
defparam \tdl_arr[14][6] .power_up = "low";

dffeas \tdl_arr[15][6] (
	.clk(clk),
	.d(\tdl_arr[14][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[15][6]~q ),
	.prn(vcc));
defparam \tdl_arr[15][6] .is_wysiwyg = "true";
defparam \tdl_arr[15][6] .power_up = "low";

dffeas \tdl_arr[16][6] (
	.clk(clk),
	.d(\tdl_arr[15][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[16][6]~q ),
	.prn(vcc));
defparam \tdl_arr[16][6] .is_wysiwyg = "true";
defparam \tdl_arr[16][6] .power_up = "low";

dffeas \tdl_arr[17][6] (
	.clk(clk),
	.d(\tdl_arr[16][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[17][6]~q ),
	.prn(vcc));
defparam \tdl_arr[17][6] .is_wysiwyg = "true";
defparam \tdl_arr[17][6] .power_up = "low";

dffeas \tdl_arr[18][6] (
	.clk(clk),
	.d(\tdl_arr[17][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[18][6]~q ),
	.prn(vcc));
defparam \tdl_arr[18][6] .is_wysiwyg = "true";
defparam \tdl_arr[18][6] .power_up = "low";

dffeas \tdl_arr[19][6] (
	.clk(clk),
	.d(\tdl_arr[18][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[19][6]~q ),
	.prn(vcc));
defparam \tdl_arr[19][6] .is_wysiwyg = "true";
defparam \tdl_arr[19][6] .power_up = "low";

dffeas \tdl_arr[0][0] (
	.clk(clk),
	.d(data_in[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][0]~q ),
	.prn(vcc));
defparam \tdl_arr[0][0] .is_wysiwyg = "true";
defparam \tdl_arr[0][0] .power_up = "low";

dffeas \tdl_arr[1][0] (
	.clk(clk),
	.d(\tdl_arr[0][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[1][0]~q ),
	.prn(vcc));
defparam \tdl_arr[1][0] .is_wysiwyg = "true";
defparam \tdl_arr[1][0] .power_up = "low";

dffeas \tdl_arr[2][0] (
	.clk(clk),
	.d(\tdl_arr[1][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[2][0]~q ),
	.prn(vcc));
defparam \tdl_arr[2][0] .is_wysiwyg = "true";
defparam \tdl_arr[2][0] .power_up = "low";

dffeas \tdl_arr[3][0] (
	.clk(clk),
	.d(\tdl_arr[2][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[3][0]~q ),
	.prn(vcc));
defparam \tdl_arr[3][0] .is_wysiwyg = "true";
defparam \tdl_arr[3][0] .power_up = "low";

dffeas \tdl_arr[4][0] (
	.clk(clk),
	.d(\tdl_arr[3][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[4][0]~q ),
	.prn(vcc));
defparam \tdl_arr[4][0] .is_wysiwyg = "true";
defparam \tdl_arr[4][0] .power_up = "low";

dffeas \tdl_arr[5][0] (
	.clk(clk),
	.d(\tdl_arr[4][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[5][0]~q ),
	.prn(vcc));
defparam \tdl_arr[5][0] .is_wysiwyg = "true";
defparam \tdl_arr[5][0] .power_up = "low";

dffeas \tdl_arr[6][0] (
	.clk(clk),
	.d(\tdl_arr[5][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[6][0]~q ),
	.prn(vcc));
defparam \tdl_arr[6][0] .is_wysiwyg = "true";
defparam \tdl_arr[6][0] .power_up = "low";

dffeas \tdl_arr[7][0] (
	.clk(clk),
	.d(\tdl_arr[6][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[7][0]~q ),
	.prn(vcc));
defparam \tdl_arr[7][0] .is_wysiwyg = "true";
defparam \tdl_arr[7][0] .power_up = "low";

dffeas \tdl_arr[8][0] (
	.clk(clk),
	.d(\tdl_arr[7][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[8][0]~q ),
	.prn(vcc));
defparam \tdl_arr[8][0] .is_wysiwyg = "true";
defparam \tdl_arr[8][0] .power_up = "low";

dffeas \tdl_arr[9][0] (
	.clk(clk),
	.d(\tdl_arr[8][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[9][0]~q ),
	.prn(vcc));
defparam \tdl_arr[9][0] .is_wysiwyg = "true";
defparam \tdl_arr[9][0] .power_up = "low";

dffeas \tdl_arr[10][0] (
	.clk(clk),
	.d(\tdl_arr[9][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[10][0]~q ),
	.prn(vcc));
defparam \tdl_arr[10][0] .is_wysiwyg = "true";
defparam \tdl_arr[10][0] .power_up = "low";

dffeas \tdl_arr[11][0] (
	.clk(clk),
	.d(\tdl_arr[10][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[11][0]~q ),
	.prn(vcc));
defparam \tdl_arr[11][0] .is_wysiwyg = "true";
defparam \tdl_arr[11][0] .power_up = "low";

dffeas \tdl_arr[12][0] (
	.clk(clk),
	.d(\tdl_arr[11][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[12][0]~q ),
	.prn(vcc));
defparam \tdl_arr[12][0] .is_wysiwyg = "true";
defparam \tdl_arr[12][0] .power_up = "low";

dffeas \tdl_arr[13][0] (
	.clk(clk),
	.d(\tdl_arr[12][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[13][0]~q ),
	.prn(vcc));
defparam \tdl_arr[13][0] .is_wysiwyg = "true";
defparam \tdl_arr[13][0] .power_up = "low";

dffeas \tdl_arr[14][0] (
	.clk(clk),
	.d(\tdl_arr[13][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[14][0]~q ),
	.prn(vcc));
defparam \tdl_arr[14][0] .is_wysiwyg = "true";
defparam \tdl_arr[14][0] .power_up = "low";

dffeas \tdl_arr[15][0] (
	.clk(clk),
	.d(\tdl_arr[14][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[15][0]~q ),
	.prn(vcc));
defparam \tdl_arr[15][0] .is_wysiwyg = "true";
defparam \tdl_arr[15][0] .power_up = "low";

dffeas \tdl_arr[16][0] (
	.clk(clk),
	.d(\tdl_arr[15][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[16][0]~q ),
	.prn(vcc));
defparam \tdl_arr[16][0] .is_wysiwyg = "true";
defparam \tdl_arr[16][0] .power_up = "low";

dffeas \tdl_arr[17][0] (
	.clk(clk),
	.d(\tdl_arr[16][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[17][0]~q ),
	.prn(vcc));
defparam \tdl_arr[17][0] .is_wysiwyg = "true";
defparam \tdl_arr[17][0] .power_up = "low";

dffeas \tdl_arr[18][0] (
	.clk(clk),
	.d(\tdl_arr[17][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[18][0]~q ),
	.prn(vcc));
defparam \tdl_arr[18][0] .is_wysiwyg = "true";
defparam \tdl_arr[18][0] .power_up = "low";

dffeas \tdl_arr[19][0] (
	.clk(clk),
	.d(\tdl_arr[18][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[19][0]~q ),
	.prn(vcc));
defparam \tdl_arr[19][0] .is_wysiwyg = "true";
defparam \tdl_arr[19][0] .power_up = "low";

dffeas \tdl_arr[0][2] (
	.clk(clk),
	.d(data_in[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][2]~q ),
	.prn(vcc));
defparam \tdl_arr[0][2] .is_wysiwyg = "true";
defparam \tdl_arr[0][2] .power_up = "low";

dffeas \tdl_arr[1][2] (
	.clk(clk),
	.d(\tdl_arr[0][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[1][2]~q ),
	.prn(vcc));
defparam \tdl_arr[1][2] .is_wysiwyg = "true";
defparam \tdl_arr[1][2] .power_up = "low";

dffeas \tdl_arr[2][2] (
	.clk(clk),
	.d(\tdl_arr[1][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[2][2]~q ),
	.prn(vcc));
defparam \tdl_arr[2][2] .is_wysiwyg = "true";
defparam \tdl_arr[2][2] .power_up = "low";

dffeas \tdl_arr[3][2] (
	.clk(clk),
	.d(\tdl_arr[2][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[3][2]~q ),
	.prn(vcc));
defparam \tdl_arr[3][2] .is_wysiwyg = "true";
defparam \tdl_arr[3][2] .power_up = "low";

dffeas \tdl_arr[4][2] (
	.clk(clk),
	.d(\tdl_arr[3][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[4][2]~q ),
	.prn(vcc));
defparam \tdl_arr[4][2] .is_wysiwyg = "true";
defparam \tdl_arr[4][2] .power_up = "low";

dffeas \tdl_arr[5][2] (
	.clk(clk),
	.d(\tdl_arr[4][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[5][2]~q ),
	.prn(vcc));
defparam \tdl_arr[5][2] .is_wysiwyg = "true";
defparam \tdl_arr[5][2] .power_up = "low";

dffeas \tdl_arr[6][2] (
	.clk(clk),
	.d(\tdl_arr[5][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[6][2]~q ),
	.prn(vcc));
defparam \tdl_arr[6][2] .is_wysiwyg = "true";
defparam \tdl_arr[6][2] .power_up = "low";

dffeas \tdl_arr[7][2] (
	.clk(clk),
	.d(\tdl_arr[6][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[7][2]~q ),
	.prn(vcc));
defparam \tdl_arr[7][2] .is_wysiwyg = "true";
defparam \tdl_arr[7][2] .power_up = "low";

dffeas \tdl_arr[8][2] (
	.clk(clk),
	.d(\tdl_arr[7][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[8][2]~q ),
	.prn(vcc));
defparam \tdl_arr[8][2] .is_wysiwyg = "true";
defparam \tdl_arr[8][2] .power_up = "low";

dffeas \tdl_arr[9][2] (
	.clk(clk),
	.d(\tdl_arr[8][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[9][2]~q ),
	.prn(vcc));
defparam \tdl_arr[9][2] .is_wysiwyg = "true";
defparam \tdl_arr[9][2] .power_up = "low";

dffeas \tdl_arr[10][2] (
	.clk(clk),
	.d(\tdl_arr[9][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[10][2]~q ),
	.prn(vcc));
defparam \tdl_arr[10][2] .is_wysiwyg = "true";
defparam \tdl_arr[10][2] .power_up = "low";

dffeas \tdl_arr[11][2] (
	.clk(clk),
	.d(\tdl_arr[10][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[11][2]~q ),
	.prn(vcc));
defparam \tdl_arr[11][2] .is_wysiwyg = "true";
defparam \tdl_arr[11][2] .power_up = "low";

dffeas \tdl_arr[12][2] (
	.clk(clk),
	.d(\tdl_arr[11][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[12][2]~q ),
	.prn(vcc));
defparam \tdl_arr[12][2] .is_wysiwyg = "true";
defparam \tdl_arr[12][2] .power_up = "low";

dffeas \tdl_arr[13][2] (
	.clk(clk),
	.d(\tdl_arr[12][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[13][2]~q ),
	.prn(vcc));
defparam \tdl_arr[13][2] .is_wysiwyg = "true";
defparam \tdl_arr[13][2] .power_up = "low";

dffeas \tdl_arr[14][2] (
	.clk(clk),
	.d(\tdl_arr[13][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[14][2]~q ),
	.prn(vcc));
defparam \tdl_arr[14][2] .is_wysiwyg = "true";
defparam \tdl_arr[14][2] .power_up = "low";

dffeas \tdl_arr[15][2] (
	.clk(clk),
	.d(\tdl_arr[14][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[15][2]~q ),
	.prn(vcc));
defparam \tdl_arr[15][2] .is_wysiwyg = "true";
defparam \tdl_arr[15][2] .power_up = "low";

dffeas \tdl_arr[16][2] (
	.clk(clk),
	.d(\tdl_arr[15][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[16][2]~q ),
	.prn(vcc));
defparam \tdl_arr[16][2] .is_wysiwyg = "true";
defparam \tdl_arr[16][2] .power_up = "low";

dffeas \tdl_arr[17][2] (
	.clk(clk),
	.d(\tdl_arr[16][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[17][2]~q ),
	.prn(vcc));
defparam \tdl_arr[17][2] .is_wysiwyg = "true";
defparam \tdl_arr[17][2] .power_up = "low";

dffeas \tdl_arr[18][2] (
	.clk(clk),
	.d(\tdl_arr[17][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[18][2]~q ),
	.prn(vcc));
defparam \tdl_arr[18][2] .is_wysiwyg = "true";
defparam \tdl_arr[18][2] .power_up = "low";

dffeas \tdl_arr[19][2] (
	.clk(clk),
	.d(\tdl_arr[18][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[19][2]~q ),
	.prn(vcc));
defparam \tdl_arr[19][2] .is_wysiwyg = "true";
defparam \tdl_arr[19][2] .power_up = "low";

dffeas \tdl_arr[0][1] (
	.clk(clk),
	.d(data_in[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][1]~q ),
	.prn(vcc));
defparam \tdl_arr[0][1] .is_wysiwyg = "true";
defparam \tdl_arr[0][1] .power_up = "low";

dffeas \tdl_arr[1][1] (
	.clk(clk),
	.d(\tdl_arr[0][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[1][1]~q ),
	.prn(vcc));
defparam \tdl_arr[1][1] .is_wysiwyg = "true";
defparam \tdl_arr[1][1] .power_up = "low";

dffeas \tdl_arr[2][1] (
	.clk(clk),
	.d(\tdl_arr[1][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[2][1]~q ),
	.prn(vcc));
defparam \tdl_arr[2][1] .is_wysiwyg = "true";
defparam \tdl_arr[2][1] .power_up = "low";

dffeas \tdl_arr[3][1] (
	.clk(clk),
	.d(\tdl_arr[2][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[3][1]~q ),
	.prn(vcc));
defparam \tdl_arr[3][1] .is_wysiwyg = "true";
defparam \tdl_arr[3][1] .power_up = "low";

dffeas \tdl_arr[4][1] (
	.clk(clk),
	.d(\tdl_arr[3][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[4][1]~q ),
	.prn(vcc));
defparam \tdl_arr[4][1] .is_wysiwyg = "true";
defparam \tdl_arr[4][1] .power_up = "low";

dffeas \tdl_arr[5][1] (
	.clk(clk),
	.d(\tdl_arr[4][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[5][1]~q ),
	.prn(vcc));
defparam \tdl_arr[5][1] .is_wysiwyg = "true";
defparam \tdl_arr[5][1] .power_up = "low";

dffeas \tdl_arr[6][1] (
	.clk(clk),
	.d(\tdl_arr[5][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[6][1]~q ),
	.prn(vcc));
defparam \tdl_arr[6][1] .is_wysiwyg = "true";
defparam \tdl_arr[6][1] .power_up = "low";

dffeas \tdl_arr[7][1] (
	.clk(clk),
	.d(\tdl_arr[6][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[7][1]~q ),
	.prn(vcc));
defparam \tdl_arr[7][1] .is_wysiwyg = "true";
defparam \tdl_arr[7][1] .power_up = "low";

dffeas \tdl_arr[8][1] (
	.clk(clk),
	.d(\tdl_arr[7][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[8][1]~q ),
	.prn(vcc));
defparam \tdl_arr[8][1] .is_wysiwyg = "true";
defparam \tdl_arr[8][1] .power_up = "low";

dffeas \tdl_arr[9][1] (
	.clk(clk),
	.d(\tdl_arr[8][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[9][1]~q ),
	.prn(vcc));
defparam \tdl_arr[9][1] .is_wysiwyg = "true";
defparam \tdl_arr[9][1] .power_up = "low";

dffeas \tdl_arr[10][1] (
	.clk(clk),
	.d(\tdl_arr[9][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[10][1]~q ),
	.prn(vcc));
defparam \tdl_arr[10][1] .is_wysiwyg = "true";
defparam \tdl_arr[10][1] .power_up = "low";

dffeas \tdl_arr[11][1] (
	.clk(clk),
	.d(\tdl_arr[10][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[11][1]~q ),
	.prn(vcc));
defparam \tdl_arr[11][1] .is_wysiwyg = "true";
defparam \tdl_arr[11][1] .power_up = "low";

dffeas \tdl_arr[12][1] (
	.clk(clk),
	.d(\tdl_arr[11][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[12][1]~q ),
	.prn(vcc));
defparam \tdl_arr[12][1] .is_wysiwyg = "true";
defparam \tdl_arr[12][1] .power_up = "low";

dffeas \tdl_arr[13][1] (
	.clk(clk),
	.d(\tdl_arr[12][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[13][1]~q ),
	.prn(vcc));
defparam \tdl_arr[13][1] .is_wysiwyg = "true";
defparam \tdl_arr[13][1] .power_up = "low";

dffeas \tdl_arr[14][1] (
	.clk(clk),
	.d(\tdl_arr[13][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[14][1]~q ),
	.prn(vcc));
defparam \tdl_arr[14][1] .is_wysiwyg = "true";
defparam \tdl_arr[14][1] .power_up = "low";

dffeas \tdl_arr[15][1] (
	.clk(clk),
	.d(\tdl_arr[14][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[15][1]~q ),
	.prn(vcc));
defparam \tdl_arr[15][1] .is_wysiwyg = "true";
defparam \tdl_arr[15][1] .power_up = "low";

dffeas \tdl_arr[16][1] (
	.clk(clk),
	.d(\tdl_arr[15][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[16][1]~q ),
	.prn(vcc));
defparam \tdl_arr[16][1] .is_wysiwyg = "true";
defparam \tdl_arr[16][1] .power_up = "low";

dffeas \tdl_arr[17][1] (
	.clk(clk),
	.d(\tdl_arr[16][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[17][1]~q ),
	.prn(vcc));
defparam \tdl_arr[17][1] .is_wysiwyg = "true";
defparam \tdl_arr[17][1] .power_up = "low";

dffeas \tdl_arr[18][1] (
	.clk(clk),
	.d(\tdl_arr[17][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[18][1]~q ),
	.prn(vcc));
defparam \tdl_arr[18][1] .is_wysiwyg = "true";
defparam \tdl_arr[18][1] .power_up = "low";

dffeas \tdl_arr[19][1] (
	.clk(clk),
	.d(\tdl_arr[18][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[19][1]~q ),
	.prn(vcc));
defparam \tdl_arr[19][1] .is_wysiwyg = "true";
defparam \tdl_arr[19][1] .power_up = "low";

dffeas \tdl_arr[0][3] (
	.clk(clk),
	.d(data_in[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][3]~q ),
	.prn(vcc));
defparam \tdl_arr[0][3] .is_wysiwyg = "true";
defparam \tdl_arr[0][3] .power_up = "low";

dffeas \tdl_arr[1][3] (
	.clk(clk),
	.d(\tdl_arr[0][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[1][3]~q ),
	.prn(vcc));
defparam \tdl_arr[1][3] .is_wysiwyg = "true";
defparam \tdl_arr[1][3] .power_up = "low";

dffeas \tdl_arr[2][3] (
	.clk(clk),
	.d(\tdl_arr[1][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[2][3]~q ),
	.prn(vcc));
defparam \tdl_arr[2][3] .is_wysiwyg = "true";
defparam \tdl_arr[2][3] .power_up = "low";

dffeas \tdl_arr[3][3] (
	.clk(clk),
	.d(\tdl_arr[2][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[3][3]~q ),
	.prn(vcc));
defparam \tdl_arr[3][3] .is_wysiwyg = "true";
defparam \tdl_arr[3][3] .power_up = "low";

dffeas \tdl_arr[4][3] (
	.clk(clk),
	.d(\tdl_arr[3][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[4][3]~q ),
	.prn(vcc));
defparam \tdl_arr[4][3] .is_wysiwyg = "true";
defparam \tdl_arr[4][3] .power_up = "low";

dffeas \tdl_arr[5][3] (
	.clk(clk),
	.d(\tdl_arr[4][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[5][3]~q ),
	.prn(vcc));
defparam \tdl_arr[5][3] .is_wysiwyg = "true";
defparam \tdl_arr[5][3] .power_up = "low";

dffeas \tdl_arr[6][3] (
	.clk(clk),
	.d(\tdl_arr[5][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[6][3]~q ),
	.prn(vcc));
defparam \tdl_arr[6][3] .is_wysiwyg = "true";
defparam \tdl_arr[6][3] .power_up = "low";

dffeas \tdl_arr[7][3] (
	.clk(clk),
	.d(\tdl_arr[6][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[7][3]~q ),
	.prn(vcc));
defparam \tdl_arr[7][3] .is_wysiwyg = "true";
defparam \tdl_arr[7][3] .power_up = "low";

dffeas \tdl_arr[8][3] (
	.clk(clk),
	.d(\tdl_arr[7][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[8][3]~q ),
	.prn(vcc));
defparam \tdl_arr[8][3] .is_wysiwyg = "true";
defparam \tdl_arr[8][3] .power_up = "low";

dffeas \tdl_arr[9][3] (
	.clk(clk),
	.d(\tdl_arr[8][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[9][3]~q ),
	.prn(vcc));
defparam \tdl_arr[9][3] .is_wysiwyg = "true";
defparam \tdl_arr[9][3] .power_up = "low";

dffeas \tdl_arr[10][3] (
	.clk(clk),
	.d(\tdl_arr[9][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[10][3]~q ),
	.prn(vcc));
defparam \tdl_arr[10][3] .is_wysiwyg = "true";
defparam \tdl_arr[10][3] .power_up = "low";

dffeas \tdl_arr[11][3] (
	.clk(clk),
	.d(\tdl_arr[10][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[11][3]~q ),
	.prn(vcc));
defparam \tdl_arr[11][3] .is_wysiwyg = "true";
defparam \tdl_arr[11][3] .power_up = "low";

dffeas \tdl_arr[12][3] (
	.clk(clk),
	.d(\tdl_arr[11][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[12][3]~q ),
	.prn(vcc));
defparam \tdl_arr[12][3] .is_wysiwyg = "true";
defparam \tdl_arr[12][3] .power_up = "low";

dffeas \tdl_arr[13][3] (
	.clk(clk),
	.d(\tdl_arr[12][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[13][3]~q ),
	.prn(vcc));
defparam \tdl_arr[13][3] .is_wysiwyg = "true";
defparam \tdl_arr[13][3] .power_up = "low";

dffeas \tdl_arr[14][3] (
	.clk(clk),
	.d(\tdl_arr[13][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[14][3]~q ),
	.prn(vcc));
defparam \tdl_arr[14][3] .is_wysiwyg = "true";
defparam \tdl_arr[14][3] .power_up = "low";

dffeas \tdl_arr[15][3] (
	.clk(clk),
	.d(\tdl_arr[14][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[15][3]~q ),
	.prn(vcc));
defparam \tdl_arr[15][3] .is_wysiwyg = "true";
defparam \tdl_arr[15][3] .power_up = "low";

dffeas \tdl_arr[16][3] (
	.clk(clk),
	.d(\tdl_arr[15][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[16][3]~q ),
	.prn(vcc));
defparam \tdl_arr[16][3] .is_wysiwyg = "true";
defparam \tdl_arr[16][3] .power_up = "low";

dffeas \tdl_arr[17][3] (
	.clk(clk),
	.d(\tdl_arr[16][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[17][3]~q ),
	.prn(vcc));
defparam \tdl_arr[17][3] .is_wysiwyg = "true";
defparam \tdl_arr[17][3] .power_up = "low";

dffeas \tdl_arr[18][3] (
	.clk(clk),
	.d(\tdl_arr[17][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[18][3]~q ),
	.prn(vcc));
defparam \tdl_arr[18][3] .is_wysiwyg = "true";
defparam \tdl_arr[18][3] .power_up = "low";

dffeas \tdl_arr[19][3] (
	.clk(clk),
	.d(\tdl_arr[18][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[19][3]~q ),
	.prn(vcc));
defparam \tdl_arr[19][3] .is_wysiwyg = "true";
defparam \tdl_arr[19][3] .power_up = "low";

dffeas \tdl_arr[0][5] (
	.clk(clk),
	.d(data_in[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][5]~q ),
	.prn(vcc));
defparam \tdl_arr[0][5] .is_wysiwyg = "true";
defparam \tdl_arr[0][5] .power_up = "low";

dffeas \tdl_arr[1][5] (
	.clk(clk),
	.d(\tdl_arr[0][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[1][5]~q ),
	.prn(vcc));
defparam \tdl_arr[1][5] .is_wysiwyg = "true";
defparam \tdl_arr[1][5] .power_up = "low";

dffeas \tdl_arr[2][5] (
	.clk(clk),
	.d(\tdl_arr[1][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[2][5]~q ),
	.prn(vcc));
defparam \tdl_arr[2][5] .is_wysiwyg = "true";
defparam \tdl_arr[2][5] .power_up = "low";

dffeas \tdl_arr[3][5] (
	.clk(clk),
	.d(\tdl_arr[2][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[3][5]~q ),
	.prn(vcc));
defparam \tdl_arr[3][5] .is_wysiwyg = "true";
defparam \tdl_arr[3][5] .power_up = "low";

dffeas \tdl_arr[4][5] (
	.clk(clk),
	.d(\tdl_arr[3][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[4][5]~q ),
	.prn(vcc));
defparam \tdl_arr[4][5] .is_wysiwyg = "true";
defparam \tdl_arr[4][5] .power_up = "low";

dffeas \tdl_arr[5][5] (
	.clk(clk),
	.d(\tdl_arr[4][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[5][5]~q ),
	.prn(vcc));
defparam \tdl_arr[5][5] .is_wysiwyg = "true";
defparam \tdl_arr[5][5] .power_up = "low";

dffeas \tdl_arr[6][5] (
	.clk(clk),
	.d(\tdl_arr[5][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[6][5]~q ),
	.prn(vcc));
defparam \tdl_arr[6][5] .is_wysiwyg = "true";
defparam \tdl_arr[6][5] .power_up = "low";

dffeas \tdl_arr[7][5] (
	.clk(clk),
	.d(\tdl_arr[6][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[7][5]~q ),
	.prn(vcc));
defparam \tdl_arr[7][5] .is_wysiwyg = "true";
defparam \tdl_arr[7][5] .power_up = "low";

dffeas \tdl_arr[8][5] (
	.clk(clk),
	.d(\tdl_arr[7][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[8][5]~q ),
	.prn(vcc));
defparam \tdl_arr[8][5] .is_wysiwyg = "true";
defparam \tdl_arr[8][5] .power_up = "low";

dffeas \tdl_arr[9][5] (
	.clk(clk),
	.d(\tdl_arr[8][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[9][5]~q ),
	.prn(vcc));
defparam \tdl_arr[9][5] .is_wysiwyg = "true";
defparam \tdl_arr[9][5] .power_up = "low";

dffeas \tdl_arr[10][5] (
	.clk(clk),
	.d(\tdl_arr[9][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[10][5]~q ),
	.prn(vcc));
defparam \tdl_arr[10][5] .is_wysiwyg = "true";
defparam \tdl_arr[10][5] .power_up = "low";

dffeas \tdl_arr[11][5] (
	.clk(clk),
	.d(\tdl_arr[10][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[11][5]~q ),
	.prn(vcc));
defparam \tdl_arr[11][5] .is_wysiwyg = "true";
defparam \tdl_arr[11][5] .power_up = "low";

dffeas \tdl_arr[12][5] (
	.clk(clk),
	.d(\tdl_arr[11][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[12][5]~q ),
	.prn(vcc));
defparam \tdl_arr[12][5] .is_wysiwyg = "true";
defparam \tdl_arr[12][5] .power_up = "low";

dffeas \tdl_arr[13][5] (
	.clk(clk),
	.d(\tdl_arr[12][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[13][5]~q ),
	.prn(vcc));
defparam \tdl_arr[13][5] .is_wysiwyg = "true";
defparam \tdl_arr[13][5] .power_up = "low";

dffeas \tdl_arr[14][5] (
	.clk(clk),
	.d(\tdl_arr[13][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[14][5]~q ),
	.prn(vcc));
defparam \tdl_arr[14][5] .is_wysiwyg = "true";
defparam \tdl_arr[14][5] .power_up = "low";

dffeas \tdl_arr[15][5] (
	.clk(clk),
	.d(\tdl_arr[14][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[15][5]~q ),
	.prn(vcc));
defparam \tdl_arr[15][5] .is_wysiwyg = "true";
defparam \tdl_arr[15][5] .power_up = "low";

dffeas \tdl_arr[16][5] (
	.clk(clk),
	.d(\tdl_arr[15][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[16][5]~q ),
	.prn(vcc));
defparam \tdl_arr[16][5] .is_wysiwyg = "true";
defparam \tdl_arr[16][5] .power_up = "low";

dffeas \tdl_arr[17][5] (
	.clk(clk),
	.d(\tdl_arr[16][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[17][5]~q ),
	.prn(vcc));
defparam \tdl_arr[17][5] .is_wysiwyg = "true";
defparam \tdl_arr[17][5] .power_up = "low";

dffeas \tdl_arr[18][5] (
	.clk(clk),
	.d(\tdl_arr[17][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[18][5]~q ),
	.prn(vcc));
defparam \tdl_arr[18][5] .is_wysiwyg = "true";
defparam \tdl_arr[18][5] .power_up = "low";

dffeas \tdl_arr[19][5] (
	.clk(clk),
	.d(\tdl_arr[18][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[19][5]~q ),
	.prn(vcc));
defparam \tdl_arr[19][5] .is_wysiwyg = "true";
defparam \tdl_arr[19][5] .power_up = "low";

dffeas \tdl_arr[0][6] (
	.clk(clk),
	.d(data_in[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][6]~q ),
	.prn(vcc));
defparam \tdl_arr[0][6] .is_wysiwyg = "true";
defparam \tdl_arr[0][6] .power_up = "low";

endmodule

module fft_asj_fft_tdl_fft_120_1 (
	global_clock_enable,
	tdl_arr_0_1,
	tdl_arr_2_1,
	tdl_arr_1_1,
	data_in,
	clk)/* synthesis synthesis_greybox=1 */;
input 	global_clock_enable;
output 	tdl_arr_0_1;
output 	tdl_arr_2_1;
output 	tdl_arr_1_1;
input 	[6:0] data_in;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \tdl_arr[0][0]~q ;
wire \tdl_arr[0][2]~q ;
wire \tdl_arr[0][1]~q ;


dffeas \tdl_arr[1][0] (
	.clk(clk),
	.d(\tdl_arr[0][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_0_1),
	.prn(vcc));
defparam \tdl_arr[1][0] .is_wysiwyg = "true";
defparam \tdl_arr[1][0] .power_up = "low";

dffeas \tdl_arr[1][2] (
	.clk(clk),
	.d(\tdl_arr[0][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_2_1),
	.prn(vcc));
defparam \tdl_arr[1][2] .is_wysiwyg = "true";
defparam \tdl_arr[1][2] .power_up = "low";

dffeas \tdl_arr[1][1] (
	.clk(clk),
	.d(\tdl_arr[0][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_1_1),
	.prn(vcc));
defparam \tdl_arr[1][1] .is_wysiwyg = "true";
defparam \tdl_arr[1][1] .power_up = "low";

dffeas \tdl_arr[0][0] (
	.clk(clk),
	.d(data_in[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][0]~q ),
	.prn(vcc));
defparam \tdl_arr[0][0] .is_wysiwyg = "true";
defparam \tdl_arr[0][0] .power_up = "low";

dffeas \tdl_arr[0][2] (
	.clk(clk),
	.d(data_in[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][2]~q ),
	.prn(vcc));
defparam \tdl_arr[0][2] .is_wysiwyg = "true";
defparam \tdl_arr[0][2] .power_up = "low";

dffeas \tdl_arr[0][1] (
	.clk(clk),
	.d(data_in[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][1]~q ),
	.prn(vcc));
defparam \tdl_arr[0][1] .is_wysiwyg = "true";
defparam \tdl_arr[0][1] .power_up = "low";

endmodule

module fft_asj_fft_twadgen_fft_120 (
	global_clock_enable,
	p_2,
	p_0,
	p_1,
	twad_tdl_0_6,
	twad_tdl_1_6,
	twad_tdl_2_6,
	twad_tdl_3_6,
	twad_tdl_4_6,
	twad_tdl_5_6,
	twad_tdl_6_6,
	k_count_2,
	Mux7,
	Mux1,
	k_count_4,
	Mux11,
	k_count_1,
	k_count_3,
	k_count_5,
	k_count_6,
	clk)/* synthesis synthesis_greybox=1 */;
input 	global_clock_enable;
input 	p_2;
input 	p_0;
input 	p_1;
output 	twad_tdl_0_6;
output 	twad_tdl_1_6;
output 	twad_tdl_2_6;
output 	twad_tdl_3_6;
output 	twad_tdl_4_6;
output 	twad_tdl_5_6;
output 	twad_tdl_6_6;
input 	k_count_2;
input 	Mux7;
input 	Mux1;
input 	k_count_4;
input 	Mux11;
input 	k_count_1;
input 	k_count_3;
input 	k_count_5;
input 	k_count_6;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Mux4~0_combout ;
wire \Mux3~0_combout ;
wire \Mux1~0_combout ;
wire \Mux0~0_combout ;
wire \Mux6~0_combout ;
wire \twad_temp[0]~q ;
wire \twad_tdl[0][0]~q ;
wire \twad_tdl[1][0]~q ;
wire \twad_tdl[2][0]~q ;
wire \twad_tdl[3][0]~q ;
wire \twad_tdl[4][0]~q ;
wire \twad_tdl[5][0]~q ;
wire \Mux5~0_combout ;
wire \twad_temp[1]~q ;
wire \twad_tdl[0][1]~q ;
wire \twad_tdl[1][1]~q ;
wire \twad_tdl[2][1]~q ;
wire \twad_tdl[3][1]~q ;
wire \twad_tdl[4][1]~q ;
wire \twad_tdl[5][1]~q ;
wire \Mux4~1_combout ;
wire \twad_temp[2]~q ;
wire \twad_tdl[0][2]~q ;
wire \twad_tdl[1][2]~q ;
wire \twad_tdl[2][2]~q ;
wire \twad_tdl[3][2]~q ;
wire \twad_tdl[4][2]~q ;
wire \twad_tdl[5][2]~q ;
wire \Mux3~1_combout ;
wire \twad_temp[3]~q ;
wire \twad_tdl[0][3]~q ;
wire \twad_tdl[1][3]~q ;
wire \twad_tdl[2][3]~q ;
wire \twad_tdl[3][3]~q ;
wire \twad_tdl[4][3]~q ;
wire \twad_tdl[5][3]~q ;
wire \Mux2~2_combout ;
wire \Mux2~3_combout ;
wire \twad_temp[4]~q ;
wire \twad_tdl[0][4]~q ;
wire \twad_tdl[1][4]~q ;
wire \twad_tdl[2][4]~q ;
wire \twad_tdl[3][4]~q ;
wire \twad_tdl[4][4]~q ;
wire \twad_tdl[5][4]~q ;
wire \Mux1~1_combout ;
wire \twad_temp[5]~q ;
wire \twad_tdl[0][5]~q ;
wire \twad_tdl[1][5]~q ;
wire \twad_tdl[2][5]~q ;
wire \twad_tdl[3][5]~q ;
wire \twad_tdl[4][5]~q ;
wire \twad_tdl[5][5]~q ;
wire \Mux0~1_combout ;
wire \Mux0~2_combout ;
wire \twad_temp[6]~q ;
wire \twad_tdl[0][6]~q ;
wire \twad_tdl[1][6]~q ;
wire \twad_tdl[2][6]~q ;
wire \twad_tdl[3][6]~q ;
wire \twad_tdl[4][6]~q ;
wire \twad_tdl[5][6]~q ;


cycloneiii_lcell_comb \Mux4~0 (
	.dataa(k_count_6),
	.datab(k_count_5),
	.datac(p_0),
	.datad(p_1),
	.cin(gnd),
	.combout(\Mux4~0_combout ),
	.cout());
defparam \Mux4~0 .lut_mask = 16'hEFFE;
defparam \Mux4~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux3~0 (
	.dataa(k_count_4),
	.datab(k_count_2),
	.datac(p_0),
	.datad(p_1),
	.cin(gnd),
	.combout(\Mux3~0_combout ),
	.cout());
defparam \Mux3~0 .lut_mask = 16'hEFFE;
defparam \Mux3~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux1~0 (
	.dataa(p_0),
	.datab(Mux11),
	.datac(Mux1),
	.datad(p_1),
	.cin(gnd),
	.combout(\Mux1~0_combout ),
	.cout());
defparam \Mux1~0 .lut_mask = 16'hFAFC;
defparam \Mux1~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux0~0 (
	.dataa(k_count_6),
	.datab(k_count_3),
	.datac(p_1),
	.datad(p_2),
	.cin(gnd),
	.combout(\Mux0~0_combout ),
	.cout());
defparam \Mux0~0 .lut_mask = 16'hEFFE;
defparam \Mux0~0 .sum_lutc_input = "datac";

dffeas \twad_tdl[6][0] (
	.clk(clk),
	.d(\twad_tdl[5][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(twad_tdl_0_6),
	.prn(vcc));
defparam \twad_tdl[6][0] .is_wysiwyg = "true";
defparam \twad_tdl[6][0] .power_up = "low";

dffeas \twad_tdl[6][1] (
	.clk(clk),
	.d(\twad_tdl[5][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(twad_tdl_1_6),
	.prn(vcc));
defparam \twad_tdl[6][1] .is_wysiwyg = "true";
defparam \twad_tdl[6][1] .power_up = "low";

dffeas \twad_tdl[6][2] (
	.clk(clk),
	.d(\twad_tdl[5][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(twad_tdl_2_6),
	.prn(vcc));
defparam \twad_tdl[6][2] .is_wysiwyg = "true";
defparam \twad_tdl[6][2] .power_up = "low";

dffeas \twad_tdl[6][3] (
	.clk(clk),
	.d(\twad_tdl[5][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(twad_tdl_3_6),
	.prn(vcc));
defparam \twad_tdl[6][3] .is_wysiwyg = "true";
defparam \twad_tdl[6][3] .power_up = "low";

dffeas \twad_tdl[6][4] (
	.clk(clk),
	.d(\twad_tdl[5][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(twad_tdl_4_6),
	.prn(vcc));
defparam \twad_tdl[6][4] .is_wysiwyg = "true";
defparam \twad_tdl[6][4] .power_up = "low";

dffeas \twad_tdl[6][5] (
	.clk(clk),
	.d(\twad_tdl[5][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(twad_tdl_5_6),
	.prn(vcc));
defparam \twad_tdl[6][5] .is_wysiwyg = "true";
defparam \twad_tdl[6][5] .power_up = "low";

dffeas \twad_tdl[6][6] (
	.clk(clk),
	.d(\twad_tdl[5][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(twad_tdl_6_6),
	.prn(vcc));
defparam \twad_tdl[6][6] .is_wysiwyg = "true";
defparam \twad_tdl[6][6] .power_up = "low";

cycloneiii_lcell_comb \Mux6~0 (
	.dataa(p_0),
	.datab(k_count_6),
	.datac(p_1),
	.datad(p_2),
	.cin(gnd),
	.combout(\Mux6~0_combout ),
	.cout());
defparam \Mux6~0 .lut_mask = 16'hEFFF;
defparam \Mux6~0 .sum_lutc_input = "datac";

dffeas \twad_temp[0] (
	.clk(clk),
	.d(\Mux6~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\twad_temp[0]~q ),
	.prn(vcc));
defparam \twad_temp[0] .is_wysiwyg = "true";
defparam \twad_temp[0] .power_up = "low";

dffeas \twad_tdl[0][0] (
	.clk(clk),
	.d(\twad_temp[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\twad_tdl[0][0]~q ),
	.prn(vcc));
defparam \twad_tdl[0][0] .is_wysiwyg = "true";
defparam \twad_tdl[0][0] .power_up = "low";

dffeas \twad_tdl[1][0] (
	.clk(clk),
	.d(\twad_tdl[0][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\twad_tdl[1][0]~q ),
	.prn(vcc));
defparam \twad_tdl[1][0] .is_wysiwyg = "true";
defparam \twad_tdl[1][0] .power_up = "low";

dffeas \twad_tdl[2][0] (
	.clk(clk),
	.d(\twad_tdl[1][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\twad_tdl[2][0]~q ),
	.prn(vcc));
defparam \twad_tdl[2][0] .is_wysiwyg = "true";
defparam \twad_tdl[2][0] .power_up = "low";

dffeas \twad_tdl[3][0] (
	.clk(clk),
	.d(\twad_tdl[2][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\twad_tdl[3][0]~q ),
	.prn(vcc));
defparam \twad_tdl[3][0] .is_wysiwyg = "true";
defparam \twad_tdl[3][0] .power_up = "low";

dffeas \twad_tdl[4][0] (
	.clk(clk),
	.d(\twad_tdl[3][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\twad_tdl[4][0]~q ),
	.prn(vcc));
defparam \twad_tdl[4][0] .is_wysiwyg = "true";
defparam \twad_tdl[4][0] .power_up = "low";

dffeas \twad_tdl[5][0] (
	.clk(clk),
	.d(\twad_tdl[4][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\twad_tdl[5][0]~q ),
	.prn(vcc));
defparam \twad_tdl[5][0] .is_wysiwyg = "true";
defparam \twad_tdl[5][0] .power_up = "low";

cycloneiii_lcell_comb \Mux5~0 (
	.dataa(p_0),
	.datab(k_count_4),
	.datac(p_1),
	.datad(p_2),
	.cin(gnd),
	.combout(\Mux5~0_combout ),
	.cout());
defparam \Mux5~0 .lut_mask = 16'hEFFF;
defparam \Mux5~0 .sum_lutc_input = "datac";

dffeas \twad_temp[1] (
	.clk(clk),
	.d(\Mux5~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\twad_temp[1]~q ),
	.prn(vcc));
defparam \twad_temp[1] .is_wysiwyg = "true";
defparam \twad_temp[1] .power_up = "low";

dffeas \twad_tdl[0][1] (
	.clk(clk),
	.d(\twad_temp[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\twad_tdl[0][1]~q ),
	.prn(vcc));
defparam \twad_tdl[0][1] .is_wysiwyg = "true";
defparam \twad_tdl[0][1] .power_up = "low";

dffeas \twad_tdl[1][1] (
	.clk(clk),
	.d(\twad_tdl[0][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\twad_tdl[1][1]~q ),
	.prn(vcc));
defparam \twad_tdl[1][1] .is_wysiwyg = "true";
defparam \twad_tdl[1][1] .power_up = "low";

dffeas \twad_tdl[2][1] (
	.clk(clk),
	.d(\twad_tdl[1][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\twad_tdl[2][1]~q ),
	.prn(vcc));
defparam \twad_tdl[2][1] .is_wysiwyg = "true";
defparam \twad_tdl[2][1] .power_up = "low";

dffeas \twad_tdl[3][1] (
	.clk(clk),
	.d(\twad_tdl[2][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\twad_tdl[3][1]~q ),
	.prn(vcc));
defparam \twad_tdl[3][1] .is_wysiwyg = "true";
defparam \twad_tdl[3][1] .power_up = "low";

dffeas \twad_tdl[4][1] (
	.clk(clk),
	.d(\twad_tdl[3][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\twad_tdl[4][1]~q ),
	.prn(vcc));
defparam \twad_tdl[4][1] .is_wysiwyg = "true";
defparam \twad_tdl[4][1] .power_up = "low";

dffeas \twad_tdl[5][1] (
	.clk(clk),
	.d(\twad_tdl[4][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\twad_tdl[5][1]~q ),
	.prn(vcc));
defparam \twad_tdl[5][1] .is_wysiwyg = "true";
defparam \twad_tdl[5][1] .power_up = "low";

cycloneiii_lcell_comb \Mux4~1 (
	.dataa(\Mux4~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(p_2),
	.cin(gnd),
	.combout(\Mux4~1_combout ),
	.cout());
defparam \Mux4~1 .lut_mask = 16'hAAFF;
defparam \Mux4~1 .sum_lutc_input = "datac";

dffeas \twad_temp[2] (
	.clk(clk),
	.d(\Mux4~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\twad_temp[2]~q ),
	.prn(vcc));
defparam \twad_temp[2] .is_wysiwyg = "true";
defparam \twad_temp[2] .power_up = "low";

dffeas \twad_tdl[0][2] (
	.clk(clk),
	.d(\twad_temp[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\twad_tdl[0][2]~q ),
	.prn(vcc));
defparam \twad_tdl[0][2] .is_wysiwyg = "true";
defparam \twad_tdl[0][2] .power_up = "low";

dffeas \twad_tdl[1][2] (
	.clk(clk),
	.d(\twad_tdl[0][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\twad_tdl[1][2]~q ),
	.prn(vcc));
defparam \twad_tdl[1][2] .is_wysiwyg = "true";
defparam \twad_tdl[1][2] .power_up = "low";

dffeas \twad_tdl[2][2] (
	.clk(clk),
	.d(\twad_tdl[1][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\twad_tdl[2][2]~q ),
	.prn(vcc));
defparam \twad_tdl[2][2] .is_wysiwyg = "true";
defparam \twad_tdl[2][2] .power_up = "low";

dffeas \twad_tdl[3][2] (
	.clk(clk),
	.d(\twad_tdl[2][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\twad_tdl[3][2]~q ),
	.prn(vcc));
defparam \twad_tdl[3][2] .is_wysiwyg = "true";
defparam \twad_tdl[3][2] .power_up = "low";

dffeas \twad_tdl[4][2] (
	.clk(clk),
	.d(\twad_tdl[3][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\twad_tdl[4][2]~q ),
	.prn(vcc));
defparam \twad_tdl[4][2] .is_wysiwyg = "true";
defparam \twad_tdl[4][2] .power_up = "low";

dffeas \twad_tdl[5][2] (
	.clk(clk),
	.d(\twad_tdl[4][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\twad_tdl[5][2]~q ),
	.prn(vcc));
defparam \twad_tdl[5][2] .is_wysiwyg = "true";
defparam \twad_tdl[5][2] .power_up = "low";

cycloneiii_lcell_comb \Mux3~1 (
	.dataa(\Mux3~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(p_2),
	.cin(gnd),
	.combout(\Mux3~1_combout ),
	.cout());
defparam \Mux3~1 .lut_mask = 16'hAAFF;
defparam \Mux3~1 .sum_lutc_input = "datac";

dffeas \twad_temp[3] (
	.clk(clk),
	.d(\Mux3~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\twad_temp[3]~q ),
	.prn(vcc));
defparam \twad_temp[3] .is_wysiwyg = "true";
defparam \twad_temp[3] .power_up = "low";

dffeas \twad_tdl[0][3] (
	.clk(clk),
	.d(\twad_temp[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\twad_tdl[0][3]~q ),
	.prn(vcc));
defparam \twad_tdl[0][3] .is_wysiwyg = "true";
defparam \twad_tdl[0][3] .power_up = "low";

dffeas \twad_tdl[1][3] (
	.clk(clk),
	.d(\twad_tdl[0][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\twad_tdl[1][3]~q ),
	.prn(vcc));
defparam \twad_tdl[1][3] .is_wysiwyg = "true";
defparam \twad_tdl[1][3] .power_up = "low";

dffeas \twad_tdl[2][3] (
	.clk(clk),
	.d(\twad_tdl[1][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\twad_tdl[2][3]~q ),
	.prn(vcc));
defparam \twad_tdl[2][3] .is_wysiwyg = "true";
defparam \twad_tdl[2][3] .power_up = "low";

dffeas \twad_tdl[3][3] (
	.clk(clk),
	.d(\twad_tdl[2][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\twad_tdl[3][3]~q ),
	.prn(vcc));
defparam \twad_tdl[3][3] .is_wysiwyg = "true";
defparam \twad_tdl[3][3] .power_up = "low";

dffeas \twad_tdl[4][3] (
	.clk(clk),
	.d(\twad_tdl[3][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\twad_tdl[4][3]~q ),
	.prn(vcc));
defparam \twad_tdl[4][3] .is_wysiwyg = "true";
defparam \twad_tdl[4][3] .power_up = "low";

dffeas \twad_tdl[5][3] (
	.clk(clk),
	.d(\twad_tdl[4][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\twad_tdl[5][3]~q ),
	.prn(vcc));
defparam \twad_tdl[5][3] .is_wysiwyg = "true";
defparam \twad_tdl[5][3] .power_up = "low";

cycloneiii_lcell_comb \Mux2~2 (
	.dataa(p_0),
	.datab(k_count_6),
	.datac(k_count_3),
	.datad(p_1),
	.cin(gnd),
	.combout(\Mux2~2_combout ),
	.cout());
defparam \Mux2~2 .lut_mask = 16'hFAFC;
defparam \Mux2~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux2~3 (
	.dataa(p_1),
	.datab(p_0),
	.datac(\Mux2~2_combout ),
	.datad(k_count_5),
	.cin(gnd),
	.combout(\Mux2~3_combout ),
	.cout());
defparam \Mux2~3 .lut_mask = 16'hFFFB;
defparam \Mux2~3 .sum_lutc_input = "datac";

dffeas \twad_temp[4] (
	.clk(clk),
	.d(\Mux2~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(p_2),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\twad_temp[4]~q ),
	.prn(vcc));
defparam \twad_temp[4] .is_wysiwyg = "true";
defparam \twad_temp[4] .power_up = "low";

dffeas \twad_tdl[0][4] (
	.clk(clk),
	.d(\twad_temp[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\twad_tdl[0][4]~q ),
	.prn(vcc));
defparam \twad_tdl[0][4] .is_wysiwyg = "true";
defparam \twad_tdl[0][4] .power_up = "low";

dffeas \twad_tdl[1][4] (
	.clk(clk),
	.d(\twad_tdl[0][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\twad_tdl[1][4]~q ),
	.prn(vcc));
defparam \twad_tdl[1][4] .is_wysiwyg = "true";
defparam \twad_tdl[1][4] .power_up = "low";

dffeas \twad_tdl[2][4] (
	.clk(clk),
	.d(\twad_tdl[1][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\twad_tdl[2][4]~q ),
	.prn(vcc));
defparam \twad_tdl[2][4] .is_wysiwyg = "true";
defparam \twad_tdl[2][4] .power_up = "low";

dffeas \twad_tdl[3][4] (
	.clk(clk),
	.d(\twad_tdl[2][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\twad_tdl[3][4]~q ),
	.prn(vcc));
defparam \twad_tdl[3][4] .is_wysiwyg = "true";
defparam \twad_tdl[3][4] .power_up = "low";

dffeas \twad_tdl[4][4] (
	.clk(clk),
	.d(\twad_tdl[3][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\twad_tdl[4][4]~q ),
	.prn(vcc));
defparam \twad_tdl[4][4] .is_wysiwyg = "true";
defparam \twad_tdl[4][4] .power_up = "low";

dffeas \twad_tdl[5][4] (
	.clk(clk),
	.d(\twad_tdl[4][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\twad_tdl[5][4]~q ),
	.prn(vcc));
defparam \twad_tdl[5][4] .is_wysiwyg = "true";
defparam \twad_tdl[5][4] .power_up = "low";

cycloneiii_lcell_comb \Mux1~1 (
	.dataa(\Mux1~0_combout ),
	.datab(k_count_2),
	.datac(Mux7),
	.datad(p_2),
	.cin(gnd),
	.combout(\Mux1~1_combout ),
	.cout());
defparam \Mux1~1 .lut_mask = 16'hFEFF;
defparam \Mux1~1 .sum_lutc_input = "datac";

dffeas \twad_temp[5] (
	.clk(clk),
	.d(\Mux1~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\twad_temp[5]~q ),
	.prn(vcc));
defparam \twad_temp[5] .is_wysiwyg = "true";
defparam \twad_temp[5] .power_up = "low";

dffeas \twad_tdl[0][5] (
	.clk(clk),
	.d(\twad_temp[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\twad_tdl[0][5]~q ),
	.prn(vcc));
defparam \twad_tdl[0][5] .is_wysiwyg = "true";
defparam \twad_tdl[0][5] .power_up = "low";

dffeas \twad_tdl[1][5] (
	.clk(clk),
	.d(\twad_tdl[0][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\twad_tdl[1][5]~q ),
	.prn(vcc));
defparam \twad_tdl[1][5] .is_wysiwyg = "true";
defparam \twad_tdl[1][5] .power_up = "low";

dffeas \twad_tdl[2][5] (
	.clk(clk),
	.d(\twad_tdl[1][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\twad_tdl[2][5]~q ),
	.prn(vcc));
defparam \twad_tdl[2][5] .is_wysiwyg = "true";
defparam \twad_tdl[2][5] .power_up = "low";

dffeas \twad_tdl[3][5] (
	.clk(clk),
	.d(\twad_tdl[2][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\twad_tdl[3][5]~q ),
	.prn(vcc));
defparam \twad_tdl[3][5] .is_wysiwyg = "true";
defparam \twad_tdl[3][5] .power_up = "low";

dffeas \twad_tdl[4][5] (
	.clk(clk),
	.d(\twad_tdl[3][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\twad_tdl[4][5]~q ),
	.prn(vcc));
defparam \twad_tdl[4][5] .is_wysiwyg = "true";
defparam \twad_tdl[4][5] .power_up = "low";

dffeas \twad_tdl[5][5] (
	.clk(clk),
	.d(\twad_tdl[4][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\twad_tdl[5][5]~q ),
	.prn(vcc));
defparam \twad_tdl[5][5] .is_wysiwyg = "true";
defparam \twad_tdl[5][5] .power_up = "low";

cycloneiii_lcell_comb \Mux0~1 (
	.dataa(k_count_5),
	.datab(k_count_1),
	.datac(gnd),
	.datad(p_1),
	.cin(gnd),
	.combout(\Mux0~1_combout ),
	.cout());
defparam \Mux0~1 .lut_mask = 16'hAACC;
defparam \Mux0~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux0~2 (
	.dataa(\Mux0~0_combout ),
	.datab(\Mux0~1_combout ),
	.datac(p_0),
	.datad(p_2),
	.cin(gnd),
	.combout(\Mux0~2_combout ),
	.cout());
defparam \Mux0~2 .lut_mask = 16'hACFF;
defparam \Mux0~2 .sum_lutc_input = "datac";

dffeas \twad_temp[6] (
	.clk(clk),
	.d(\Mux0~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\twad_temp[6]~q ),
	.prn(vcc));
defparam \twad_temp[6] .is_wysiwyg = "true";
defparam \twad_temp[6] .power_up = "low";

dffeas \twad_tdl[0][6] (
	.clk(clk),
	.d(\twad_temp[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\twad_tdl[0][6]~q ),
	.prn(vcc));
defparam \twad_tdl[0][6] .is_wysiwyg = "true";
defparam \twad_tdl[0][6] .power_up = "low";

dffeas \twad_tdl[1][6] (
	.clk(clk),
	.d(\twad_tdl[0][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\twad_tdl[1][6]~q ),
	.prn(vcc));
defparam \twad_tdl[1][6] .is_wysiwyg = "true";
defparam \twad_tdl[1][6] .power_up = "low";

dffeas \twad_tdl[2][6] (
	.clk(clk),
	.d(\twad_tdl[1][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\twad_tdl[2][6]~q ),
	.prn(vcc));
defparam \twad_tdl[2][6] .is_wysiwyg = "true";
defparam \twad_tdl[2][6] .power_up = "low";

dffeas \twad_tdl[3][6] (
	.clk(clk),
	.d(\twad_tdl[2][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\twad_tdl[3][6]~q ),
	.prn(vcc));
defparam \twad_tdl[3][6] .is_wysiwyg = "true";
defparam \twad_tdl[3][6] .power_up = "low";

dffeas \twad_tdl[4][6] (
	.clk(clk),
	.d(\twad_tdl[3][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\twad_tdl[4][6]~q ),
	.prn(vcc));
defparam \twad_tdl[4][6] .is_wysiwyg = "true";
defparam \twad_tdl[4][6] .power_up = "low";

dffeas \twad_tdl[5][6] (
	.clk(clk),
	.d(\twad_tdl[4][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\twad_tdl[5][6]~q ),
	.prn(vcc));
defparam \twad_tdl[5][6] .is_wysiwyg = "true";
defparam \twad_tdl[5][6] .power_up = "low";

endmodule

module fft_asj_fft_wrengen_fft_120 (
	global_clock_enable,
	wc_i1,
	wd_i1,
	ram_a_not_b_vec_26,
	p_cd_en_2,
	p_cd_en_0,
	p_cd_en_1,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	global_clock_enable;
output 	wc_i1;
output 	wd_i1;
input 	ram_a_not_b_vec_26;
input 	p_cd_en_2;
input 	p_cd_en_0;
input 	p_cd_en_1;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wd_i~0_combout ;
wire \wc_i~0_combout ;
wire \wd_i~1_combout ;


dffeas wc_i(
	.clk(clk),
	.d(\wc_i~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wc_i1),
	.prn(vcc));
defparam wc_i.is_wysiwyg = "true";
defparam wc_i.power_up = "low";

dffeas wd_i(
	.clk(clk),
	.d(\wd_i~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wd_i1),
	.prn(vcc));
defparam wd_i.is_wysiwyg = "true";
defparam wd_i.power_up = "low";

cycloneiii_lcell_comb \wd_i~0 (
	.dataa(reset_n),
	.datab(p_cd_en_2),
	.datac(p_cd_en_0),
	.datad(p_cd_en_1),
	.cin(gnd),
	.combout(\wd_i~0_combout ),
	.cout());
defparam \wd_i~0 .lut_mask = 16'hEFFF;
defparam \wd_i~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wc_i~0 (
	.dataa(ram_a_not_b_vec_26),
	.datab(gnd),
	.datac(gnd),
	.datad(\wd_i~0_combout ),
	.cin(gnd),
	.combout(\wc_i~0_combout ),
	.cout());
defparam \wc_i~0 .lut_mask = 16'hFF55;
defparam \wc_i~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wd_i~1 (
	.dataa(ram_a_not_b_vec_26),
	.datab(\wd_i~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wd_i~1_combout ),
	.cout());
defparam \wd_i~1 .lut_mask = 16'hEEEE;
defparam \wd_i~1 .sum_lutc_input = "datac";

endmodule

module fft_asj_fft_wrswgen_fft_120 (
	global_clock_enable,
	swa_tdl_0_0,
	swa_tdl_1_0,
	tdl_arr_4_20,
	tdl_arr_6_20,
	tdl_arr_0_20,
	tdl_arr_2_20,
	tdl_arr_0_1,
	tdl_arr_2_1,
	tdl_arr_1_1,
	tdl_arr_1_20,
	tdl_arr_3_20,
	tdl_arr_5_20,
	clk)/* synthesis synthesis_greybox=1 */;
input 	global_clock_enable;
output 	swa_tdl_0_0;
output 	swa_tdl_1_0;
input 	tdl_arr_4_20;
input 	tdl_arr_6_20;
input 	tdl_arr_0_20;
input 	tdl_arr_2_20;
input 	tdl_arr_0_1;
input 	tdl_arr_2_1;
input 	tdl_arr_1_1;
input 	tdl_arr_1_20;
input 	tdl_arr_3_20;
input 	tdl_arr_5_20;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add2~0_combout ;
wire \Add1~0_combout ;
wire \Mux1~0_combout ;
wire \swd[0]~0_combout ;
wire \swd[0]~1_combout ;
wire \Mux1~1_combout ;
wire \swd[0]~2_combout ;
wire \Add0~0_combout ;
wire \Mux1~2_combout ;
wire \swd[0]~q ;
wire \Add0~1_combout ;
wire \Mux0~0_combout ;
wire \Mux0~1_combout ;
wire \Mux0~2_combout ;
wire \Mux0~3_combout ;
wire \swd[1]~q ;


cycloneiii_lcell_comb \Add2~0 (
	.dataa(tdl_arr_4_20),
	.datab(tdl_arr_6_20),
	.datac(tdl_arr_0_20),
	.datad(tdl_arr_2_20),
	.cin(gnd),
	.combout(\Add2~0_combout ),
	.cout());
defparam \Add2~0 .lut_mask = 16'h6996;
defparam \Add2~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add1~0 (
	.dataa(tdl_arr_4_20),
	.datab(\Add0~0_combout ),
	.datac(\Add0~1_combout ),
	.datad(tdl_arr_5_20),
	.cin(gnd),
	.combout(\Add1~0_combout ),
	.cout());
defparam \Add1~0 .lut_mask = 16'h6996;
defparam \Add1~0 .sum_lutc_input = "datac";

dffeas \swa_tdl[0][0] (
	.clk(clk),
	.d(\swd[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(swa_tdl_0_0),
	.prn(vcc));
defparam \swa_tdl[0][0] .is_wysiwyg = "true";
defparam \swa_tdl[0][0] .power_up = "low";

dffeas \swa_tdl[0][1] (
	.clk(clk),
	.d(\swd[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(swa_tdl_1_0),
	.prn(vcc));
defparam \swa_tdl[0][1] .is_wysiwyg = "true";
defparam \swa_tdl[0][1] .power_up = "low";

cycloneiii_lcell_comb \Mux1~0 (
	.dataa(tdl_arr_0_20),
	.datab(tdl_arr_0_1),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux1~0_combout ),
	.cout());
defparam \Mux1~0 .lut_mask = 16'hEEEE;
defparam \Mux1~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \swd[0]~0 (
	.dataa(gnd),
	.datab(tdl_arr_0_1),
	.datac(tdl_arr_2_1),
	.datad(tdl_arr_1_1),
	.cin(gnd),
	.combout(\swd[0]~0_combout ),
	.cout());
defparam \swd[0]~0 .lut_mask = 16'h3FFF;
defparam \swd[0]~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \swd[0]~1 (
	.dataa(tdl_arr_2_1),
	.datab(tdl_arr_0_1),
	.datac(tdl_arr_1_1),
	.datad(gnd),
	.cin(gnd),
	.combout(\swd[0]~1_combout ),
	.cout());
defparam \swd[0]~1 .lut_mask = 16'hFEFE;
defparam \swd[0]~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux1~1 (
	.dataa(\Add2~0_combout ),
	.datab(\Mux1~0_combout ),
	.datac(\swd[0]~0_combout ),
	.datad(\swd[0]~1_combout ),
	.cin(gnd),
	.combout(\Mux1~1_combout ),
	.cout());
defparam \Mux1~1 .lut_mask = 16'hEFFE;
defparam \Mux1~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \swd[0]~2 (
	.dataa(tdl_arr_1_1),
	.datab(gnd),
	.datac(gnd),
	.datad(tdl_arr_2_1),
	.cin(gnd),
	.combout(\swd[0]~2_combout ),
	.cout());
defparam \swd[0]~2 .lut_mask = 16'hAAFF;
defparam \swd[0]~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add0~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(tdl_arr_0_20),
	.datad(tdl_arr_2_20),
	.cin(gnd),
	.combout(\Add0~0_combout ),
	.cout());
defparam \Add0~0 .lut_mask = 16'h0FF0;
defparam \Add0~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux1~2 (
	.dataa(tdl_arr_4_20),
	.datab(\Mux1~1_combout ),
	.datac(\swd[0]~2_combout ),
	.datad(\Add0~0_combout ),
	.cin(gnd),
	.combout(\Mux1~2_combout ),
	.cout());
defparam \Mux1~2 .lut_mask = 16'h6996;
defparam \Mux1~2 .sum_lutc_input = "datac";

dffeas \swd[0] (
	.clk(clk),
	.d(\Mux1~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\swd[0]~q ),
	.prn(vcc));
defparam \swd[0] .is_wysiwyg = "true";
defparam \swd[0] .power_up = "low";

cycloneiii_lcell_comb \Add0~1 (
	.dataa(tdl_arr_0_20),
	.datab(tdl_arr_2_20),
	.datac(tdl_arr_1_20),
	.datad(tdl_arr_3_20),
	.cin(gnd),
	.combout(\Add0~1_combout ),
	.cout());
defparam \Add0~1 .lut_mask = 16'h6996;
defparam \Add0~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux0~0 (
	.dataa(tdl_arr_4_20),
	.datab(\Add0~0_combout ),
	.datac(tdl_arr_5_20),
	.datad(tdl_arr_6_20),
	.cin(gnd),
	.combout(\Mux0~0_combout ),
	.cout());
defparam \Mux0~0 .lut_mask = 16'h6996;
defparam \Mux0~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux0~1 (
	.dataa(tdl_arr_0_1),
	.datab(tdl_arr_1_20),
	.datac(\swd[0]~0_combout ),
	.datad(\swd[0]~1_combout ),
	.cin(gnd),
	.combout(\Mux0~1_combout ),
	.cout());
defparam \Mux0~1 .lut_mask = 16'hFFF7;
defparam \Mux0~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux0~2 (
	.dataa(\Add0~1_combout ),
	.datab(\Mux0~0_combout ),
	.datac(\swd[0]~1_combout ),
	.datad(\Mux0~1_combout ),
	.cin(gnd),
	.combout(\Mux0~2_combout ),
	.cout());
defparam \Mux0~2 .lut_mask = 16'h6996;
defparam \Mux0~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux0~3 (
	.dataa(\Add1~0_combout ),
	.datab(\Add0~1_combout ),
	.datac(\swd[0]~2_combout ),
	.datad(\Mux0~2_combout ),
	.cin(gnd),
	.combout(\Mux0~3_combout ),
	.cout());
defparam \Mux0~3 .lut_mask = 16'hEFFE;
defparam \Mux0~3 .sum_lutc_input = "datac";

dffeas \swd[1] (
	.clk(clk),
	.d(\Mux0~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\swd[1]~q ),
	.prn(vcc));
defparam \swd[1] .is_wysiwyg = "true";
defparam \swd[1] .power_up = "low";

endmodule

module fft_auk_dspip_avalon_streaming_controller_fft_120 (
	at_source_valid_s,
	source_packet_error_0,
	source_packet_error_1,
	valid_ctrl_int,
	master_sink_ena,
	source_stall_reg1,
	sink_stall_reg1,
	sink_ready_ctrl,
	sink_stall,
	packet_error_s_0,
	packet_error_s_1,
	Mux3,
	stall_reg1,
	Mux0,
	Mux01,
	clk,
	reset_n,
	source_ready)/* synthesis synthesis_greybox=1 */;
input 	at_source_valid_s;
output 	source_packet_error_0;
output 	source_packet_error_1;
input 	valid_ctrl_int;
input 	master_sink_ena;
output 	source_stall_reg1;
output 	sink_stall_reg1;
output 	sink_ready_ctrl;
input 	sink_stall;
input 	packet_error_s_0;
input 	packet_error_s_1;
input 	Mux3;
output 	stall_reg1;
input 	Mux0;
input 	Mux01;
input 	clk;
input 	reset_n;
input 	source_ready;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \source_stall_reg~0_combout ;
wire \sink_stall_reg~0_combout ;
wire \stall_int~2_combout ;
wire \stall_int~combout ;


dffeas \source_packet_error[0] (
	.clk(clk),
	.d(packet_error_s_0),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(source_packet_error_0),
	.prn(vcc));
defparam \source_packet_error[0] .is_wysiwyg = "true";
defparam \source_packet_error[0] .power_up = "low";

dffeas \source_packet_error[1] (
	.clk(clk),
	.d(packet_error_s_1),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(source_packet_error_1),
	.prn(vcc));
defparam \source_packet_error[1] .is_wysiwyg = "true";
defparam \source_packet_error[1] .power_up = "low";

dffeas source_stall_reg(
	.clk(clk),
	.d(\source_stall_reg~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(source_stall_reg1),
	.prn(vcc));
defparam source_stall_reg.is_wysiwyg = "true";
defparam source_stall_reg.power_up = "low";

dffeas sink_stall_reg(
	.clk(clk),
	.d(\sink_stall_reg~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sink_stall_reg1),
	.prn(vcc));
defparam sink_stall_reg.is_wysiwyg = "true";
defparam sink_stall_reg.power_up = "low";

cycloneiii_lcell_comb \sink_ready_ctrl~0 (
	.dataa(master_sink_ena),
	.datab(source_stall_reg1),
	.datac(gnd),
	.datad(sink_stall_reg1),
	.cin(gnd),
	.combout(sink_ready_ctrl),
	.cout());
defparam \sink_ready_ctrl~0 .lut_mask = 16'hEEFF;
defparam \sink_ready_ctrl~0 .sum_lutc_input = "datac";

dffeas stall_reg(
	.clk(clk),
	.d(\stall_int~combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(stall_reg1),
	.prn(vcc));
defparam stall_reg.is_wysiwyg = "true";
defparam stall_reg.power_up = "low";

cycloneiii_lcell_comb \source_stall_reg~0 (
	.dataa(Mux01),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\source_stall_reg~0_combout ),
	.cout());
defparam \source_stall_reg~0 .lut_mask = 16'h5555;
defparam \source_stall_reg~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sink_stall_reg~0 (
	.dataa(sink_stall),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sink_stall_reg~0_combout ),
	.cout());
defparam \sink_stall_reg~0 .lut_mask = 16'h5555;
defparam \sink_stall_reg~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \stall_int~2 (
	.dataa(at_source_valid_s),
	.datab(source_ready),
	.datac(valid_ctrl_int),
	.datad(Mux0),
	.cin(gnd),
	.combout(\stall_int~2_combout ),
	.cout());
defparam \stall_int~2 .lut_mask = 16'hFFBF;
defparam \stall_int~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb stall_int(
	.dataa(sink_stall),
	.datab(Mux0),
	.datac(Mux3),
	.datad(\stall_int~2_combout ),
	.cin(gnd),
	.combout(\stall_int~combout ),
	.cout());
defparam stall_int.lut_mask = 16'h7FFF;
defparam stall_int.sum_lutc_input = "datac";

endmodule

module fft_auk_dspip_avalon_streaming_sink_fft_120 (
	q_b_2,
	q_b_10,
	q_b_6,
	q_b_14,
	q_b_4,
	q_b_12,
	q_b_3,
	q_b_11,
	q_b_5,
	q_b_13,
	q_b_1,
	q_b_9,
	q_b_0,
	q_b_8,
	q_b_7,
	q_b_15,
	at_sink_ready_s1,
	sink_ready_ctrl,
	sink_stall1,
	packet_error_s_0,
	packet_error_s_1,
	send_sop_s1,
	send_eop_s1,
	clk,
	reset_n,
	sink_error_0,
	sink_error_1,
	sink_valid,
	sink_sop,
	sink_eop,
	at_sink_data)/* synthesis synthesis_greybox=1 */;
output 	q_b_2;
output 	q_b_10;
output 	q_b_6;
output 	q_b_14;
output 	q_b_4;
output 	q_b_12;
output 	q_b_3;
output 	q_b_11;
output 	q_b_5;
output 	q_b_13;
output 	q_b_1;
output 	q_b_9;
output 	q_b_0;
output 	q_b_8;
output 	q_b_7;
output 	q_b_15;
output 	at_sink_ready_s1;
input 	sink_ready_ctrl;
output 	sink_stall1;
output 	packet_error_s_0;
output 	packet_error_s_1;
output 	send_sop_s1;
output 	send_eop_s1;
input 	clk;
input 	reset_n;
input 	sink_error_0;
input 	sink_error_1;
input 	sink_valid;
input 	sink_sop;
input 	sink_eop;
input 	[15:0] at_sink_data;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \out_cnt[0]~q ;
wire \out_cnt[4]~q ;
wire \count[1]~q ;
wire \count[2]~q ;
wire \count[3]~q ;
wire \count[0]~q ;
wire \count[4]~q ;
wire \out_cnt[0]~9_combout ;
wire \out_cnt[4]~17_combout ;
wire \count[0]~11_combout ;
wire \count[1]~13_combout ;
wire \count[2]~18_combout ;
wire \count[3]~20_combout ;
wire \count[4]~22_combout ;
wire \normal_fifo:fifo_eab_on:in_fifo|auto_generated|dffe_af~q ;
wire \normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|empty_dff~q ;
wire \normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|usedw_counter|counter_reg_bit[0]~q ;
wire \Selector2~3_combout ;
wire \sink_state.start~q ;
wire \max_reached~0_combout ;
wire \Selector0~0_combout ;
wire \Selector0~1_combout ;
wire \LessThan0~0_combout ;
wire \at_sink_data_int[2]~q ;
wire \at_sink_data_int[10]~q ;
wire \at_sink_data_int[6]~q ;
wire \at_sink_data_int[14]~q ;
wire \at_sink_data_int[4]~q ;
wire \at_sink_data_int[12]~q ;
wire \at_sink_data_int[3]~q ;
wire \at_sink_data_int[11]~q ;
wire \at_sink_data_int[5]~q ;
wire \at_sink_data_int[13]~q ;
wire \at_sink_data_int[1]~q ;
wire \at_sink_data_int[9]~q ;
wire \at_sink_data_int[0]~q ;
wire \at_sink_data_int[8]~q ;
wire \at_sink_data_int[7]~q ;
wire \at_sink_data_int[15]~q ;
wire \data_take~combout ;
wire \fifo_wrreq~0_wirecell_combout ;
wire \at_sink_ready_s~0_combout ;
wire \sink_start~0_combout ;
wire \sink_start~q ;
wire \Selector2~2_combout ;
wire \sink_comb_update_2~4_combout ;
wire \sink_next_state~1_combout ;
wire \Selector1~0_combout ;
wire \sink_state.stall~q ;
wire \count[0]~12 ;
wire \count[1]~14 ;
wire \count[2]~19 ;
wire \count[3]~21 ;
wire \count[4]~23 ;
wire \count[5]~25 ;
wire \count[6]~27 ;
wire \count[7]~29 ;
wire \count[8]~30_combout ;
wire \sink_comb_update_2~1_combout ;
wire \Selector4~0_combout ;
wire \sink_state.end1~q ;
wire \Selector4~1_combout ;
wire \Selector3~7_combout ;
wire \Selector3~6_combout ;
wire \sink_state.st_err~q ;
wire \Selector5~0_combout ;
wire \Selector3~5_combout ;
wire \count[1]~32_combout ;
wire \count[1]~15_combout ;
wire \sink_comb_update_2~0_combout ;
wire \Selector2~4_combout ;
wire \Selector2~5_combout ;
wire \count[1]~16_combout ;
wire \count[1]~17_combout ;
wire \count[8]~q ;
wire \count[5]~24_combout ;
wire \count[5]~q ;
wire \count[6]~26_combout ;
wire \count[6]~q ;
wire \count[7]~28_combout ;
wire \count[7]~q ;
wire \max_reached~1_combout ;
wire \max_reached~2_combout ;
wire \data_take~4_combout ;
wire \max_reached~3_combout ;
wire \max_reached~q ;
wire \sink_comb_update_2~3_combout ;
wire \Selector6~2_combout ;
wire \Selector6~6_combout ;
wire \Selector3~2_combout ;
wire \Selector6~3_combout ;
wire \Selector6~4_combout ;
wire \Selector6~5_combout ;
wire \sink_comb_update_2~2_combout ;
wire \Selector2~6_combout ;
wire \sink_state.run1~q ;
wire \fifo_wrreq~0_combout ;
wire \Selector5~1_combout ;
wire \Selector3~3_combout ;
wire \Selector3~4_combout ;
wire \Selector5~2_combout ;
wire \Selector5~3_combout ;
wire \out_cnt[0]~10 ;
wire \out_cnt[1]~11_combout ;
wire \out_cnt[1]~12 ;
wire \out_cnt[2]~14 ;
wire \out_cnt[3]~16 ;
wire \out_cnt[4]~18 ;
wire \out_cnt[5]~19_combout ;
wire \sink_stall_s~q ;
wire \Selector8~0_combout ;
wire \sink_out_state.normal~q ;
wire \Selector7~0_combout ;
wire \out_cnt[5]~q ;
wire \out_cnt[5]~20 ;
wire \out_cnt[6]~21_combout ;
wire \out_cnt[6]~q ;
wire \out_cnt[6]~22 ;
wire \out_cnt[7]~23_combout ;
wire \out_cnt[7]~q ;
wire \LessThan0~1_combout ;
wire \out_cnt[7]~24 ;
wire \out_cnt[8]~25_combout ;
wire \out_cnt[8]~q ;
wire \LessThan0~2_combout ;
wire \out_cnt[1]~q ;
wire \out_cnt[2]~13_combout ;
wire \out_cnt[2]~q ;
wire \out_cnt[3]~15_combout ;
wire \out_cnt[3]~q ;
wire \Equal1~0_combout ;
wire \Equal1~1_combout ;
wire \Equal1~2_combout ;
wire \Selector10~2_combout ;
wire \Selector10~3_combout ;
wire \sink_out_state.empty_and_ready~q ;
wire \send_sop_eop_p~0_combout ;


fft_scfifo_1 \normal_fifo:fifo_eab_on:in_fifo (
	.q({q_unconnected_wire_17,q_unconnected_wire_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.dffe_af(\normal_fifo:fifo_eab_on:in_fifo|auto_generated|dffe_af~q ),
	.sink_out_stateempty_and_ready(\sink_out_state.empty_and_ready~q ),
	.sink_ready_ctrl(sink_ready_ctrl),
	.sink_out_statenormal(\sink_out_state.normal~q ),
	.sink_start(\sink_start~q ),
	.empty_dff(\normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|empty_dff~q ),
	.sink_stall(sink_stall1),
	.rdreq(\Selector7~0_combout ),
	.sink_staterun1(\sink_state.run1~q ),
	.sink_stateend1(\sink_state.end1~q ),
	.wrreq(\fifo_wrreq~0_combout ),
	.counter_reg_bit_0(\normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|usedw_counter|counter_reg_bit[0]~q ),
	.data({gnd,gnd,\at_sink_data_int[15]~q ,\at_sink_data_int[14]~q ,\at_sink_data_int[13]~q ,\at_sink_data_int[12]~q ,\at_sink_data_int[11]~q ,\at_sink_data_int[10]~q ,\at_sink_data_int[9]~q ,\at_sink_data_int[8]~q ,\at_sink_data_int[7]~q ,\at_sink_data_int[6]~q ,
\at_sink_data_int[5]~q ,\at_sink_data_int[4]~q ,\at_sink_data_int[3]~q ,\at_sink_data_int[2]~q ,\at_sink_data_int[1]~q ,\at_sink_data_int[0]~q }),
	.fifo_wrreq(\fifo_wrreq~0_wirecell_combout ),
	.clock(clk),
	.reset_n(reset_n));

dffeas \out_cnt[0] (
	.clk(clk),
	.d(\out_cnt[0]~9_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\LessThan0~2_combout ),
	.sload(gnd),
	.ena(\Selector7~0_combout ),
	.q(\out_cnt[0]~q ),
	.prn(vcc));
defparam \out_cnt[0] .is_wysiwyg = "true";
defparam \out_cnt[0] .power_up = "low";

dffeas \out_cnt[4] (
	.clk(clk),
	.d(\out_cnt[4]~17_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\LessThan0~2_combout ),
	.sload(gnd),
	.ena(\Selector7~0_combout ),
	.q(\out_cnt[4]~q ),
	.prn(vcc));
defparam \out_cnt[4] .is_wysiwyg = "true";
defparam \out_cnt[4] .power_up = "low";

dffeas \count[1] (
	.clk(clk),
	.d(\count[1]~13_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\count[1]~15_combout ),
	.sload(gnd),
	.ena(\count[1]~17_combout ),
	.q(\count[1]~q ),
	.prn(vcc));
defparam \count[1] .is_wysiwyg = "true";
defparam \count[1] .power_up = "low";

dffeas \count[2] (
	.clk(clk),
	.d(\count[2]~18_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\count[1]~15_combout ),
	.sload(gnd),
	.ena(\count[1]~17_combout ),
	.q(\count[2]~q ),
	.prn(vcc));
defparam \count[2] .is_wysiwyg = "true";
defparam \count[2] .power_up = "low";

dffeas \count[3] (
	.clk(clk),
	.d(\count[3]~20_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\count[1]~15_combout ),
	.sload(gnd),
	.ena(\count[1]~17_combout ),
	.q(\count[3]~q ),
	.prn(vcc));
defparam \count[3] .is_wysiwyg = "true";
defparam \count[3] .power_up = "low";

dffeas \count[0] (
	.clk(clk),
	.d(\count[0]~11_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\count[1]~15_combout ),
	.sload(gnd),
	.ena(\count[1]~17_combout ),
	.q(\count[0]~q ),
	.prn(vcc));
defparam \count[0] .is_wysiwyg = "true";
defparam \count[0] .power_up = "low";

dffeas \count[4] (
	.clk(clk),
	.d(\count[4]~22_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\count[1]~15_combout ),
	.sload(gnd),
	.ena(\count[1]~17_combout ),
	.q(\count[4]~q ),
	.prn(vcc));
defparam \count[4] .is_wysiwyg = "true";
defparam \count[4] .power_up = "low";

cycloneiii_lcell_comb \out_cnt[0]~9 (
	.dataa(\out_cnt[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\out_cnt[0]~9_combout ),
	.cout(\out_cnt[0]~10 ));
defparam \out_cnt[0]~9 .lut_mask = 16'h55AA;
defparam \out_cnt[0]~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \out_cnt[4]~17 (
	.dataa(\out_cnt[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\out_cnt[3]~16 ),
	.combout(\out_cnt[4]~17_combout ),
	.cout(\out_cnt[4]~18 ));
defparam \out_cnt[4]~17 .lut_mask = 16'h5AAF;
defparam \out_cnt[4]~17 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \count[0]~11 (
	.dataa(\count[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\count[0]~11_combout ),
	.cout(\count[0]~12 ));
defparam \count[0]~11 .lut_mask = 16'h55AA;
defparam \count[0]~11 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \count[1]~13 (
	.dataa(\count[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[0]~12 ),
	.combout(\count[1]~13_combout ),
	.cout(\count[1]~14 ));
defparam \count[1]~13 .lut_mask = 16'h5A5F;
defparam \count[1]~13 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \count[2]~18 (
	.dataa(\count[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[1]~14 ),
	.combout(\count[2]~18_combout ),
	.cout(\count[2]~19 ));
defparam \count[2]~18 .lut_mask = 16'h5AAF;
defparam \count[2]~18 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \count[3]~20 (
	.dataa(\count[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[2]~19 ),
	.combout(\count[3]~20_combout ),
	.cout(\count[3]~21 ));
defparam \count[3]~20 .lut_mask = 16'h5A5F;
defparam \count[3]~20 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \count[4]~22 (
	.dataa(\count[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[3]~21 ),
	.combout(\count[4]~22_combout ),
	.cout(\count[4]~23 ));
defparam \count[4]~22 .lut_mask = 16'h5AAF;
defparam \count[4]~22 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Selector2~3 (
	.dataa(\sink_state.run1~q ),
	.datab(\sink_state.stall~q ),
	.datac(sink_valid),
	.datad(sink_sop),
	.cin(gnd),
	.combout(\Selector2~3_combout ),
	.cout());
defparam \Selector2~3 .lut_mask = 16'hEFFF;
defparam \Selector2~3 .sum_lutc_input = "datac";

dffeas \sink_state.start (
	.clk(clk),
	.d(\Selector0~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sink_state.start~q ),
	.prn(vcc));
defparam \sink_state.start .is_wysiwyg = "true";
defparam \sink_state.start .power_up = "low";

cycloneiii_lcell_comb \max_reached~0 (
	.dataa(\count[1]~q ),
	.datab(\count[2]~q ),
	.datac(\count[3]~q ),
	.datad(\count[0]~q ),
	.cin(gnd),
	.combout(\max_reached~0_combout ),
	.cout());
defparam \max_reached~0 .lut_mask = 16'hFEFF;
defparam \max_reached~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector0~0 (
	.dataa(\sink_state.end1~q ),
	.datab(sink_sop),
	.datac(at_sink_ready_s1),
	.datad(sink_valid),
	.cin(gnd),
	.combout(\Selector0~0_combout ),
	.cout());
defparam \Selector0~0 .lut_mask = 16'hEFFF;
defparam \Selector0~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector0~1 (
	.dataa(\Selector2~2_combout ),
	.datab(\Selector0~0_combout ),
	.datac(\sink_comb_update_2~0_combout ),
	.datad(\Selector5~0_combout ),
	.cin(gnd),
	.combout(\Selector0~1_combout ),
	.cout());
defparam \Selector0~1 .lut_mask = 16'hFFF7;
defparam \Selector0~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \LessThan0~0 (
	.dataa(\out_cnt[0]~q ),
	.datab(\out_cnt[1]~q ),
	.datac(\out_cnt[2]~q ),
	.datad(\out_cnt[3]~q ),
	.cin(gnd),
	.combout(\LessThan0~0_combout ),
	.cout());
defparam \LessThan0~0 .lut_mask = 16'h7FFF;
defparam \LessThan0~0 .sum_lutc_input = "datac";

dffeas \at_sink_data_int[2] (
	.clk(clk),
	.d(at_sink_data[2]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[2]~q ),
	.prn(vcc));
defparam \at_sink_data_int[2] .is_wysiwyg = "true";
defparam \at_sink_data_int[2] .power_up = "low";

dffeas \at_sink_data_int[10] (
	.clk(clk),
	.d(at_sink_data[10]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[10]~q ),
	.prn(vcc));
defparam \at_sink_data_int[10] .is_wysiwyg = "true";
defparam \at_sink_data_int[10] .power_up = "low";

dffeas \at_sink_data_int[6] (
	.clk(clk),
	.d(at_sink_data[6]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[6]~q ),
	.prn(vcc));
defparam \at_sink_data_int[6] .is_wysiwyg = "true";
defparam \at_sink_data_int[6] .power_up = "low";

dffeas \at_sink_data_int[14] (
	.clk(clk),
	.d(at_sink_data[14]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[14]~q ),
	.prn(vcc));
defparam \at_sink_data_int[14] .is_wysiwyg = "true";
defparam \at_sink_data_int[14] .power_up = "low";

dffeas \at_sink_data_int[4] (
	.clk(clk),
	.d(at_sink_data[4]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[4]~q ),
	.prn(vcc));
defparam \at_sink_data_int[4] .is_wysiwyg = "true";
defparam \at_sink_data_int[4] .power_up = "low";

dffeas \at_sink_data_int[12] (
	.clk(clk),
	.d(at_sink_data[12]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[12]~q ),
	.prn(vcc));
defparam \at_sink_data_int[12] .is_wysiwyg = "true";
defparam \at_sink_data_int[12] .power_up = "low";

dffeas \at_sink_data_int[3] (
	.clk(clk),
	.d(at_sink_data[3]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[3]~q ),
	.prn(vcc));
defparam \at_sink_data_int[3] .is_wysiwyg = "true";
defparam \at_sink_data_int[3] .power_up = "low";

dffeas \at_sink_data_int[11] (
	.clk(clk),
	.d(at_sink_data[11]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[11]~q ),
	.prn(vcc));
defparam \at_sink_data_int[11] .is_wysiwyg = "true";
defparam \at_sink_data_int[11] .power_up = "low";

dffeas \at_sink_data_int[5] (
	.clk(clk),
	.d(at_sink_data[5]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[5]~q ),
	.prn(vcc));
defparam \at_sink_data_int[5] .is_wysiwyg = "true";
defparam \at_sink_data_int[5] .power_up = "low";

dffeas \at_sink_data_int[13] (
	.clk(clk),
	.d(at_sink_data[13]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[13]~q ),
	.prn(vcc));
defparam \at_sink_data_int[13] .is_wysiwyg = "true";
defparam \at_sink_data_int[13] .power_up = "low";

dffeas \at_sink_data_int[1] (
	.clk(clk),
	.d(at_sink_data[1]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[1]~q ),
	.prn(vcc));
defparam \at_sink_data_int[1] .is_wysiwyg = "true";
defparam \at_sink_data_int[1] .power_up = "low";

dffeas \at_sink_data_int[9] (
	.clk(clk),
	.d(at_sink_data[9]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[9]~q ),
	.prn(vcc));
defparam \at_sink_data_int[9] .is_wysiwyg = "true";
defparam \at_sink_data_int[9] .power_up = "low";

dffeas \at_sink_data_int[0] (
	.clk(clk),
	.d(at_sink_data[0]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[0]~q ),
	.prn(vcc));
defparam \at_sink_data_int[0] .is_wysiwyg = "true";
defparam \at_sink_data_int[0] .power_up = "low";

dffeas \at_sink_data_int[8] (
	.clk(clk),
	.d(at_sink_data[8]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[8]~q ),
	.prn(vcc));
defparam \at_sink_data_int[8] .is_wysiwyg = "true";
defparam \at_sink_data_int[8] .power_up = "low";

dffeas \at_sink_data_int[7] (
	.clk(clk),
	.d(at_sink_data[7]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[7]~q ),
	.prn(vcc));
defparam \at_sink_data_int[7] .is_wysiwyg = "true";
defparam \at_sink_data_int[7] .power_up = "low";

dffeas \at_sink_data_int[15] (
	.clk(clk),
	.d(at_sink_data[15]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[15]~q ),
	.prn(vcc));
defparam \at_sink_data_int[15] .is_wysiwyg = "true";
defparam \at_sink_data_int[15] .power_up = "low";

cycloneiii_lcell_comb data_take(
	.dataa(\sink_state.run1~q ),
	.datab(\sink_state.end1~q ),
	.datac(\Selector2~6_combout ),
	.datad(\Selector4~0_combout ),
	.cin(gnd),
	.combout(\data_take~combout ),
	.cout());
defparam data_take.lut_mask = 16'hFFFE;
defparam data_take.sum_lutc_input = "datac";

cycloneiii_lcell_comb \fifo_wrreq~0_wirecell (
	.dataa(\fifo_wrreq~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_wrreq~0_wirecell_combout ),
	.cout());
defparam \fifo_wrreq~0_wirecell .lut_mask = 16'h5555;
defparam \fifo_wrreq~0_wirecell .sum_lutc_input = "datac";

dffeas at_sink_ready_s(
	.clk(clk),
	.d(\at_sink_ready_s~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(at_sink_ready_s1),
	.prn(vcc));
defparam at_sink_ready_s.is_wysiwyg = "true";
defparam at_sink_ready_s.power_up = "low";

cycloneiii_lcell_comb sink_stall(
	.dataa(gnd),
	.datab(gnd),
	.datac(\sink_start~q ),
	.datad(\normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|empty_dff~q ),
	.cin(gnd),
	.combout(sink_stall1),
	.cout());
defparam sink_stall.lut_mask = 16'h0FFF;
defparam sink_stall.sum_lutc_input = "datac";

dffeas \packet_error_s[0] (
	.clk(clk),
	.d(\Selector6~5_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(packet_error_s_0),
	.prn(vcc));
defparam \packet_error_s[0] .is_wysiwyg = "true";
defparam \packet_error_s[0] .power_up = "low";

dffeas \packet_error_s[1] (
	.clk(clk),
	.d(\Selector5~3_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(packet_error_s_1),
	.prn(vcc));
defparam \packet_error_s[1] .is_wysiwyg = "true";
defparam \packet_error_s[1] .power_up = "low";

dffeas send_sop_s(
	.clk(clk),
	.d(\Equal1~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\send_sop_eop_p~0_combout ),
	.q(send_sop_s1),
	.prn(vcc));
defparam send_sop_s.is_wysiwyg = "true";
defparam send_sop_s.power_up = "low";

dffeas send_eop_s(
	.clk(clk),
	.d(\LessThan0~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\send_sop_eop_p~0_combout ),
	.q(send_eop_s1),
	.prn(vcc));
defparam send_eop_s.is_wysiwyg = "true";
defparam send_eop_s.power_up = "low";

cycloneiii_lcell_comb \at_sink_ready_s~0 (
	.dataa(\normal_fifo:fifo_eab_on:in_fifo|auto_generated|dffe_af~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\at_sink_ready_s~0_combout ),
	.cout());
defparam \at_sink_ready_s~0 .lut_mask = 16'h5555;
defparam \at_sink_ready_s~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sink_start~0 (
	.dataa(\sink_start~q ),
	.datab(\normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|usedw_counter|counter_reg_bit[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sink_start~0_combout ),
	.cout());
defparam \sink_start~0 .lut_mask = 16'hEEEE;
defparam \sink_start~0 .sum_lutc_input = "datac";

dffeas sink_start(
	.clk(clk),
	.d(\sink_start~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sink_start~q ),
	.prn(vcc));
defparam sink_start.is_wysiwyg = "true";
defparam sink_start.power_up = "low";

cycloneiii_lcell_comb \Selector2~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(sink_error_0),
	.datad(sink_error_1),
	.cin(gnd),
	.combout(\Selector2~2_combout ),
	.cout());
defparam \Selector2~2 .lut_mask = 16'h0FFF;
defparam \Selector2~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sink_comb_update_2~4 (
	.dataa(\max_reached~q ),
	.datab(gnd),
	.datac(sink_eop),
	.datad(at_sink_ready_s1),
	.cin(gnd),
	.combout(\sink_comb_update_2~4_combout ),
	.cout());
defparam \sink_comb_update_2~4 .lut_mask = 16'hAFFF;
defparam \sink_comb_update_2~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sink_next_state~1 (
	.dataa(sink_valid),
	.datab(gnd),
	.datac(gnd),
	.datad(at_sink_ready_s1),
	.cin(gnd),
	.combout(\sink_next_state~1_combout ),
	.cout());
defparam \sink_next_state~1 .lut_mask = 16'hAAFF;
defparam \sink_next_state~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector1~0 (
	.dataa(\Selector2~3_combout ),
	.datab(\Selector2~2_combout ),
	.datac(\sink_comb_update_2~4_combout ),
	.datad(\sink_next_state~1_combout ),
	.cin(gnd),
	.combout(\Selector1~0_combout ),
	.cout());
defparam \Selector1~0 .lut_mask = 16'hFEFF;
defparam \Selector1~0 .sum_lutc_input = "datac";

dffeas \sink_state.stall (
	.clk(clk),
	.d(\Selector1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sink_state.stall~q ),
	.prn(vcc));
defparam \sink_state.stall .is_wysiwyg = "true";
defparam \sink_state.stall .power_up = "low";

cycloneiii_lcell_comb \count[5]~24 (
	.dataa(\count[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[4]~23 ),
	.combout(\count[5]~24_combout ),
	.cout(\count[5]~25 ));
defparam \count[5]~24 .lut_mask = 16'h5A5F;
defparam \count[5]~24 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \count[6]~26 (
	.dataa(\count[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[5]~25 ),
	.combout(\count[6]~26_combout ),
	.cout(\count[6]~27 ));
defparam \count[6]~26 .lut_mask = 16'h5AAF;
defparam \count[6]~26 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \count[7]~28 (
	.dataa(\count[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[6]~27 ),
	.combout(\count[7]~28_combout ),
	.cout(\count[7]~29 ));
defparam \count[7]~28 .lut_mask = 16'h5A5F;
defparam \count[7]~28 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \count[8]~30 (
	.dataa(\count[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\count[7]~29 ),
	.combout(\count[8]~30_combout ),
	.cout());
defparam \count[8]~30 .lut_mask = 16'h5A5A;
defparam \count[8]~30 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \sink_comb_update_2~1 (
	.dataa(at_sink_ready_s1),
	.datab(sink_valid),
	.datac(sink_eop),
	.datad(\max_reached~q ),
	.cin(gnd),
	.combout(\sink_comb_update_2~1_combout ),
	.cout());
defparam \sink_comb_update_2~1 .lut_mask = 16'hFFFE;
defparam \sink_comb_update_2~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector4~0 (
	.dataa(\Selector2~3_combout ),
	.datab(\sink_comb_update_2~1_combout ),
	.datac(sink_error_0),
	.datad(sink_error_1),
	.cin(gnd),
	.combout(\Selector4~0_combout ),
	.cout());
defparam \Selector4~0 .lut_mask = 16'hEFFF;
defparam \Selector4~0 .sum_lutc_input = "datac";

dffeas \sink_state.end1 (
	.clk(clk),
	.d(\Selector4~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sink_state.end1~q ),
	.prn(vcc));
defparam \sink_state.end1 .is_wysiwyg = "true";
defparam \sink_state.end1 .power_up = "low";

cycloneiii_lcell_comb \Selector4~1 (
	.dataa(\sink_state.run1~q ),
	.datab(\sink_state.stall~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector4~1_combout ),
	.cout());
defparam \Selector4~1 .lut_mask = 16'hEEEE;
defparam \Selector4~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector3~7 (
	.dataa(sink_valid),
	.datab(sink_sop),
	.datac(\Selector4~1_combout ),
	.datad(\sink_comb_update_2~3_combout ),
	.cin(gnd),
	.combout(\Selector3~7_combout ),
	.cout());
defparam \Selector3~7 .lut_mask = 16'hFFFE;
defparam \Selector3~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector3~6 (
	.dataa(\Selector3~4_combout ),
	.datab(\Selector3~5_combout ),
	.datac(\Selector3~7_combout ),
	.datad(\Selector2~2_combout ),
	.cin(gnd),
	.combout(\Selector3~6_combout ),
	.cout());
defparam \Selector3~6 .lut_mask = 16'hFEFF;
defparam \Selector3~6 .sum_lutc_input = "datac";

dffeas \sink_state.st_err (
	.clk(clk),
	.d(\Selector3~6_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sink_state.st_err~q ),
	.prn(vcc));
defparam \sink_state.st_err .is_wysiwyg = "true";
defparam \sink_state.st_err .power_up = "low";

cycloneiii_lcell_comb \Selector5~0 (
	.dataa(\sink_state.start~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\sink_state.st_err~q ),
	.cin(gnd),
	.combout(\Selector5~0_combout ),
	.cout());
defparam \Selector5~0 .lut_mask = 16'hAAFF;
defparam \Selector5~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector3~5 (
	.dataa(\Selector3~2_combout ),
	.datab(\sink_state.end1~q ),
	.datac(at_sink_ready_s1),
	.datad(\Selector5~0_combout ),
	.cin(gnd),
	.combout(\Selector3~5_combout ),
	.cout());
defparam \Selector3~5 .lut_mask = 16'hFEFF;
defparam \Selector3~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \count[1]~32 (
	.dataa(sink_error_0),
	.datab(sink_error_1),
	.datac(\max_reached~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\count[1]~32_combout ),
	.cout());
defparam \count[1]~32 .lut_mask = 16'hFEFE;
defparam \count[1]~32 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \count[1]~15 (
	.dataa(\Selector3~4_combout ),
	.datab(\Selector3~5_combout ),
	.datac(\Selector3~7_combout ),
	.datad(\count[1]~32_combout ),
	.cin(gnd),
	.combout(\count[1]~15_combout ),
	.cout());
defparam \count[1]~15 .lut_mask = 16'hFFFE;
defparam \count[1]~15 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sink_comb_update_2~0 (
	.dataa(at_sink_ready_s1),
	.datab(sink_valid),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sink_comb_update_2~0_combout ),
	.cout());
defparam \sink_comb_update_2~0 .lut_mask = 16'hEEEE;
defparam \sink_comb_update_2~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector2~4 (
	.dataa(\Selector2~3_combout ),
	.datab(\sink_comb_update_2~0_combout ),
	.datac(sink_eop),
	.datad(\max_reached~q ),
	.cin(gnd),
	.combout(\Selector2~4_combout ),
	.cout());
defparam \Selector2~4 .lut_mask = 16'hEFFF;
defparam \Selector2~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector2~5 (
	.dataa(sink_sop),
	.datab(\sink_comb_update_2~0_combout ),
	.datac(\sink_state.end1~q ),
	.datad(\Selector5~0_combout ),
	.cin(gnd),
	.combout(\Selector2~5_combout ),
	.cout());
defparam \Selector2~5 .lut_mask = 16'hFEFF;
defparam \Selector2~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \count[1]~16 (
	.dataa(\Selector3~5_combout ),
	.datab(\Selector2~2_combout ),
	.datac(\Selector2~5_combout ),
	.datad(\Selector4~0_combout ),
	.cin(gnd),
	.combout(\count[1]~16_combout ),
	.cout());
defparam \count[1]~16 .lut_mask = 16'hFFFB;
defparam \count[1]~16 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \count[1]~17 (
	.dataa(\Selector3~4_combout ),
	.datab(\Selector3~7_combout ),
	.datac(\Selector2~4_combout ),
	.datad(\count[1]~16_combout ),
	.cin(gnd),
	.combout(\count[1]~17_combout ),
	.cout());
defparam \count[1]~17 .lut_mask = 16'hFFFE;
defparam \count[1]~17 .sum_lutc_input = "datac";

dffeas \count[8] (
	.clk(clk),
	.d(\count[8]~30_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\count[1]~15_combout ),
	.sload(gnd),
	.ena(\count[1]~17_combout ),
	.q(\count[8]~q ),
	.prn(vcc));
defparam \count[8] .is_wysiwyg = "true";
defparam \count[8] .power_up = "low";

dffeas \count[5] (
	.clk(clk),
	.d(\count[5]~24_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\count[1]~15_combout ),
	.sload(gnd),
	.ena(\count[1]~17_combout ),
	.q(\count[5]~q ),
	.prn(vcc));
defparam \count[5] .is_wysiwyg = "true";
defparam \count[5] .power_up = "low";

dffeas \count[6] (
	.clk(clk),
	.d(\count[6]~26_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\count[1]~15_combout ),
	.sload(gnd),
	.ena(\count[1]~17_combout ),
	.q(\count[6]~q ),
	.prn(vcc));
defparam \count[6] .is_wysiwyg = "true";
defparam \count[6] .power_up = "low";

dffeas \count[7] (
	.clk(clk),
	.d(\count[7]~28_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\count[1]~15_combout ),
	.sload(gnd),
	.ena(\count[1]~17_combout ),
	.q(\count[7]~q ),
	.prn(vcc));
defparam \count[7] .is_wysiwyg = "true";
defparam \count[7] .power_up = "low";

cycloneiii_lcell_comb \max_reached~1 (
	.dataa(\count[4]~q ),
	.datab(\count[5]~q ),
	.datac(\count[6]~q ),
	.datad(\count[7]~q ),
	.cin(gnd),
	.combout(\max_reached~1_combout ),
	.cout());
defparam \max_reached~1 .lut_mask = 16'hFFFE;
defparam \max_reached~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \max_reached~2 (
	.dataa(\max_reached~0_combout ),
	.datab(\count[8]~q ),
	.datac(\max_reached~1_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\max_reached~2_combout ),
	.cout());
defparam \max_reached~2 .lut_mask = 16'hFEFE;
defparam \max_reached~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \data_take~4 (
	.dataa(\Selector2~4_combout ),
	.datab(\Selector2~5_combout ),
	.datac(\Selector2~2_combout ),
	.datad(\Selector4~0_combout ),
	.cin(gnd),
	.combout(\data_take~4_combout ),
	.cout());
defparam \data_take~4 .lut_mask = 16'h7FFF;
defparam \data_take~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \max_reached~3 (
	.dataa(\max_reached~q ),
	.datab(\max_reached~2_combout ),
	.datac(\data_take~4_combout ),
	.datad(\Selector3~6_combout ),
	.cin(gnd),
	.combout(\max_reached~3_combout ),
	.cout());
defparam \max_reached~3 .lut_mask = 16'hEFFE;
defparam \max_reached~3 .sum_lutc_input = "datac";

dffeas max_reached(
	.clk(clk),
	.d(\max_reached~3_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\max_reached~q ),
	.prn(vcc));
defparam max_reached.is_wysiwyg = "true";
defparam max_reached.power_up = "low";

cycloneiii_lcell_comb \sink_comb_update_2~3 (
	.dataa(sink_eop),
	.datab(gnd),
	.datac(gnd),
	.datad(\max_reached~q ),
	.cin(gnd),
	.combout(\sink_comb_update_2~3_combout ),
	.cout());
defparam \sink_comb_update_2~3 .lut_mask = 16'hAAFF;
defparam \sink_comb_update_2~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector6~2 (
	.dataa(\sink_comb_update_2~2_combout ),
	.datab(\sink_next_state~1_combout ),
	.datac(\sink_comb_update_2~3_combout ),
	.datad(sink_error_1),
	.cin(gnd),
	.combout(\Selector6~2_combout ),
	.cout());
defparam \Selector6~2 .lut_mask = 16'hFEFF;
defparam \Selector6~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector6~6 (
	.dataa(\sink_state.run1~q ),
	.datab(\sink_state.stall~q ),
	.datac(sink_error_0),
	.datad(\Selector6~2_combout ),
	.cin(gnd),
	.combout(\Selector6~6_combout ),
	.cout());
defparam \Selector6~6 .lut_mask = 16'hFFFE;
defparam \Selector6~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector3~2 (
	.dataa(sink_valid),
	.datab(gnd),
	.datac(gnd),
	.datad(sink_sop),
	.cin(gnd),
	.combout(\Selector3~2_combout ),
	.cout());
defparam \Selector3~2 .lut_mask = 16'hAAFF;
defparam \Selector3~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector6~3 (
	.dataa(\sink_state.end1~q ),
	.datab(sink_error_0),
	.datac(\Selector3~2_combout ),
	.datad(sink_error_1),
	.cin(gnd),
	.combout(\Selector6~3_combout ),
	.cout());
defparam \Selector6~3 .lut_mask = 16'hFEFF;
defparam \Selector6~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector6~4 (
	.dataa(sink_error_0),
	.datab(\sink_comb_update_2~0_combout ),
	.datac(sink_sop),
	.datad(sink_error_1),
	.cin(gnd),
	.combout(\Selector6~4_combout ),
	.cout());
defparam \Selector6~4 .lut_mask = 16'hEFFF;
defparam \Selector6~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector6~5 (
	.dataa(\Selector6~6_combout ),
	.datab(\Selector6~3_combout ),
	.datac(\Selector6~4_combout ),
	.datad(\Selector5~0_combout ),
	.cin(gnd),
	.combout(\Selector6~5_combout ),
	.cout());
defparam \Selector6~5 .lut_mask = 16'hFEFF;
defparam \Selector6~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sink_comb_update_2~2 (
	.dataa(sink_valid),
	.datab(sink_sop),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sink_comb_update_2~2_combout ),
	.cout());
defparam \sink_comb_update_2~2 .lut_mask = 16'hEEEE;
defparam \sink_comb_update_2~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector2~6 (
	.dataa(sink_error_0),
	.datab(sink_error_1),
	.datac(\Selector2~4_combout ),
	.datad(\Selector2~5_combout ),
	.cin(gnd),
	.combout(\Selector2~6_combout ),
	.cout());
defparam \Selector2~6 .lut_mask = 16'hFFF7;
defparam \Selector2~6 .sum_lutc_input = "datac";

dffeas \sink_state.run1 (
	.clk(clk),
	.d(\Selector2~6_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sink_state.run1~q ),
	.prn(vcc));
defparam \sink_state.run1 .is_wysiwyg = "true";
defparam \sink_state.run1 .power_up = "low";

cycloneiii_lcell_comb \fifo_wrreq~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sink_state.run1~q ),
	.datad(\sink_state.end1~q ),
	.cin(gnd),
	.combout(\fifo_wrreq~0_combout ),
	.cout());
defparam \fifo_wrreq~0 .lut_mask = 16'hFFF0;
defparam \fifo_wrreq~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector5~1 (
	.dataa(sink_error_1),
	.datab(\sink_state.stall~q ),
	.datac(\fifo_wrreq~0_combout ),
	.datad(\Selector5~0_combout ),
	.cin(gnd),
	.combout(\Selector5~1_combout ),
	.cout());
defparam \Selector5~1 .lut_mask = 16'hFEFF;
defparam \Selector5~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector3~3 (
	.dataa(sink_valid),
	.datab(at_sink_ready_s1),
	.datac(\max_reached~q ),
	.datad(sink_eop),
	.cin(gnd),
	.combout(\Selector3~3_combout ),
	.cout());
defparam \Selector3~3 .lut_mask = 16'h6996;
defparam \Selector3~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector3~4 (
	.dataa(\sink_state.stall~q ),
	.datab(\sink_state.run1~q ),
	.datac(\Selector3~3_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector3~4_combout ),
	.cout());
defparam \Selector3~4 .lut_mask = 16'hFEFE;
defparam \Selector3~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector5~2 (
	.dataa(sink_valid),
	.datab(\Selector4~1_combout ),
	.datac(\sink_comb_update_2~3_combout ),
	.datad(\Selector3~4_combout ),
	.cin(gnd),
	.combout(\Selector5~2_combout ),
	.cout());
defparam \Selector5~2 .lut_mask = 16'hFFFE;
defparam \Selector5~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector5~3 (
	.dataa(\sink_comb_update_2~2_combout ),
	.datab(sink_error_0),
	.datac(\Selector5~1_combout ),
	.datad(\Selector5~2_combout ),
	.cin(gnd),
	.combout(\Selector5~3_combout ),
	.cout());
defparam \Selector5~3 .lut_mask = 16'hFFF7;
defparam \Selector5~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \out_cnt[1]~11 (
	.dataa(\out_cnt[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\out_cnt[0]~10 ),
	.combout(\out_cnt[1]~11_combout ),
	.cout(\out_cnt[1]~12 ));
defparam \out_cnt[1]~11 .lut_mask = 16'h5A5F;
defparam \out_cnt[1]~11 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \out_cnt[2]~13 (
	.dataa(\out_cnt[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\out_cnt[1]~12 ),
	.combout(\out_cnt[2]~13_combout ),
	.cout(\out_cnt[2]~14 ));
defparam \out_cnt[2]~13 .lut_mask = 16'h5AAF;
defparam \out_cnt[2]~13 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \out_cnt[3]~15 (
	.dataa(\out_cnt[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\out_cnt[2]~14 ),
	.combout(\out_cnt[3]~15_combout ),
	.cout(\out_cnt[3]~16 ));
defparam \out_cnt[3]~15 .lut_mask = 16'h5A5F;
defparam \out_cnt[3]~15 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \out_cnt[5]~19 (
	.dataa(\out_cnt[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\out_cnt[4]~18 ),
	.combout(\out_cnt[5]~19_combout ),
	.cout(\out_cnt[5]~20 ));
defparam \out_cnt[5]~19 .lut_mask = 16'h5A5F;
defparam \out_cnt[5]~19 .sum_lutc_input = "cin";

dffeas sink_stall_s(
	.clk(clk),
	.d(sink_stall1),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sink_stall_s~q ),
	.prn(vcc));
defparam sink_stall_s.is_wysiwyg = "true";
defparam sink_stall_s.power_up = "low";

cycloneiii_lcell_comb \Selector8~0 (
	.dataa(sink_ready_ctrl),
	.datab(\sink_stall_s~q ),
	.datac(\sink_out_state.normal~q ),
	.datad(sink_stall1),
	.cin(gnd),
	.combout(\Selector8~0_combout ),
	.cout());
defparam \Selector8~0 .lut_mask = 16'hFFF7;
defparam \Selector8~0 .sum_lutc_input = "datac";

dffeas \sink_out_state.normal (
	.clk(clk),
	.d(\Selector8~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sink_out_state.normal~q ),
	.prn(vcc));
defparam \sink_out_state.normal .is_wysiwyg = "true";
defparam \sink_out_state.normal .power_up = "low";

cycloneiii_lcell_comb \Selector7~0 (
	.dataa(\sink_out_state.empty_and_ready~q ),
	.datab(sink_ready_ctrl),
	.datac(\sink_out_state.normal~q ),
	.datad(sink_stall1),
	.cin(gnd),
	.combout(\Selector7~0_combout ),
	.cout());
defparam \Selector7~0 .lut_mask = 16'hEFFF;
defparam \Selector7~0 .sum_lutc_input = "datac";

dffeas \out_cnt[5] (
	.clk(clk),
	.d(\out_cnt[5]~19_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\LessThan0~2_combout ),
	.sload(gnd),
	.ena(\Selector7~0_combout ),
	.q(\out_cnt[5]~q ),
	.prn(vcc));
defparam \out_cnt[5] .is_wysiwyg = "true";
defparam \out_cnt[5] .power_up = "low";

cycloneiii_lcell_comb \out_cnt[6]~21 (
	.dataa(\out_cnt[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\out_cnt[5]~20 ),
	.combout(\out_cnt[6]~21_combout ),
	.cout(\out_cnt[6]~22 ));
defparam \out_cnt[6]~21 .lut_mask = 16'h5AAF;
defparam \out_cnt[6]~21 .sum_lutc_input = "cin";

dffeas \out_cnt[6] (
	.clk(clk),
	.d(\out_cnt[6]~21_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\LessThan0~2_combout ),
	.sload(gnd),
	.ena(\Selector7~0_combout ),
	.q(\out_cnt[6]~q ),
	.prn(vcc));
defparam \out_cnt[6] .is_wysiwyg = "true";
defparam \out_cnt[6] .power_up = "low";

cycloneiii_lcell_comb \out_cnt[7]~23 (
	.dataa(\out_cnt[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\out_cnt[6]~22 ),
	.combout(\out_cnt[7]~23_combout ),
	.cout(\out_cnt[7]~24 ));
defparam \out_cnt[7]~23 .lut_mask = 16'h5A5F;
defparam \out_cnt[7]~23 .sum_lutc_input = "cin";

dffeas \out_cnt[7] (
	.clk(clk),
	.d(\out_cnt[7]~23_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\LessThan0~2_combout ),
	.sload(gnd),
	.ena(\Selector7~0_combout ),
	.q(\out_cnt[7]~q ),
	.prn(vcc));
defparam \out_cnt[7] .is_wysiwyg = "true";
defparam \out_cnt[7] .power_up = "low";

cycloneiii_lcell_comb \LessThan0~1 (
	.dataa(\out_cnt[4]~q ),
	.datab(\out_cnt[5]~q ),
	.datac(\out_cnt[6]~q ),
	.datad(\out_cnt[7]~q ),
	.cin(gnd),
	.combout(\LessThan0~1_combout ),
	.cout());
defparam \LessThan0~1 .lut_mask = 16'h7FFF;
defparam \LessThan0~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \out_cnt[8]~25 (
	.dataa(\out_cnt[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\out_cnt[7]~24 ),
	.combout(\out_cnt[8]~25_combout ),
	.cout());
defparam \out_cnt[8]~25 .lut_mask = 16'h5A5A;
defparam \out_cnt[8]~25 .sum_lutc_input = "cin";

dffeas \out_cnt[8] (
	.clk(clk),
	.d(\out_cnt[8]~25_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\LessThan0~2_combout ),
	.sload(gnd),
	.ena(\Selector7~0_combout ),
	.q(\out_cnt[8]~q ),
	.prn(vcc));
defparam \out_cnt[8] .is_wysiwyg = "true";
defparam \out_cnt[8] .power_up = "low";

cycloneiii_lcell_comb \LessThan0~2 (
	.dataa(\LessThan0~0_combout ),
	.datab(\LessThan0~1_combout ),
	.datac(gnd),
	.datad(\out_cnt[8]~q ),
	.cin(gnd),
	.combout(\LessThan0~2_combout ),
	.cout());
defparam \LessThan0~2 .lut_mask = 16'hFF77;
defparam \LessThan0~2 .sum_lutc_input = "datac";

dffeas \out_cnt[1] (
	.clk(clk),
	.d(\out_cnt[1]~11_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\LessThan0~2_combout ),
	.sload(gnd),
	.ena(\Selector7~0_combout ),
	.q(\out_cnt[1]~q ),
	.prn(vcc));
defparam \out_cnt[1] .is_wysiwyg = "true";
defparam \out_cnt[1] .power_up = "low";

dffeas \out_cnt[2] (
	.clk(clk),
	.d(\out_cnt[2]~13_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\LessThan0~2_combout ),
	.sload(gnd),
	.ena(\Selector7~0_combout ),
	.q(\out_cnt[2]~q ),
	.prn(vcc));
defparam \out_cnt[2] .is_wysiwyg = "true";
defparam \out_cnt[2] .power_up = "low";

dffeas \out_cnt[3] (
	.clk(clk),
	.d(\out_cnt[3]~15_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\LessThan0~2_combout ),
	.sload(gnd),
	.ena(\Selector7~0_combout ),
	.q(\out_cnt[3]~q ),
	.prn(vcc));
defparam \out_cnt[3] .is_wysiwyg = "true";
defparam \out_cnt[3] .power_up = "low";

cycloneiii_lcell_comb \Equal1~0 (
	.dataa(\out_cnt[0]~q ),
	.datab(\out_cnt[1]~q ),
	.datac(\out_cnt[2]~q ),
	.datad(\out_cnt[3]~q ),
	.cin(gnd),
	.combout(\Equal1~0_combout ),
	.cout());
defparam \Equal1~0 .lut_mask = 16'h7FFF;
defparam \Equal1~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Equal1~1 (
	.dataa(\out_cnt[4]~q ),
	.datab(\out_cnt[5]~q ),
	.datac(\out_cnt[6]~q ),
	.datad(\out_cnt[7]~q ),
	.cin(gnd),
	.combout(\Equal1~1_combout ),
	.cout());
defparam \Equal1~1 .lut_mask = 16'h7FFF;
defparam \Equal1~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Equal1~2 (
	.dataa(\Equal1~0_combout ),
	.datab(\Equal1~1_combout ),
	.datac(gnd),
	.datad(\out_cnt[8]~q ),
	.cin(gnd),
	.combout(\Equal1~2_combout ),
	.cout());
defparam \Equal1~2 .lut_mask = 16'hEEFF;
defparam \Equal1~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector10~2 (
	.dataa(\sink_out_state.empty_and_ready~q ),
	.datab(sink_ready_ctrl),
	.datac(\sink_stall_s~q ),
	.datad(\sink_out_state.normal~q ),
	.cin(gnd),
	.combout(\Selector10~2_combout ),
	.cout());
defparam \Selector10~2 .lut_mask = 16'hBEFF;
defparam \Selector10~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector10~3 (
	.dataa(\sink_start~q ),
	.datab(\normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|empty_dff~q ),
	.datac(\Selector10~2_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector10~3_combout ),
	.cout());
defparam \Selector10~3 .lut_mask = 16'hF7F7;
defparam \Selector10~3 .sum_lutc_input = "datac";

dffeas \sink_out_state.empty_and_ready (
	.clk(clk),
	.d(\Selector10~3_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sink_out_state.empty_and_ready~q ),
	.prn(vcc));
defparam \sink_out_state.empty_and_ready .is_wysiwyg = "true";
defparam \sink_out_state.empty_and_ready .power_up = "low";

cycloneiii_lcell_comb \send_sop_eop_p~0 (
	.dataa(sink_ready_ctrl),
	.datab(\sink_out_state.empty_and_ready~q ),
	.datac(\sink_out_state.normal~q ),
	.datad(sink_stall1),
	.cin(gnd),
	.combout(\send_sop_eop_p~0_combout ),
	.cout());
defparam \send_sop_eop_p~0 .lut_mask = 16'hEFFF;
defparam \send_sop_eop_p~0 .sum_lutc_input = "datac";

endmodule

module fft_scfifo_1 (
	q,
	dffe_af,
	sink_out_stateempty_and_ready,
	sink_ready_ctrl,
	sink_out_statenormal,
	sink_start,
	empty_dff,
	sink_stall,
	rdreq,
	sink_staterun1,
	sink_stateend1,
	wrreq,
	counter_reg_bit_0,
	data,
	fifo_wrreq,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[17:0] q;
output 	dffe_af;
input 	sink_out_stateempty_and_ready;
input 	sink_ready_ctrl;
input 	sink_out_statenormal;
input 	sink_start;
output 	empty_dff;
input 	sink_stall;
input 	rdreq;
input 	sink_staterun1;
input 	sink_stateend1;
input 	wrreq;
output 	counter_reg_bit_0;
input 	[17:0] data;
input 	fifo_wrreq;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft_scfifo_nch1 auto_generated(
	.q({q_unconnected_wire_17,q_unconnected_wire_16,q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.dffe_af1(dffe_af),
	.sink_out_stateempty_and_ready(sink_out_stateempty_and_ready),
	.sink_ready_ctrl(sink_ready_ctrl),
	.sink_out_statenormal(sink_out_statenormal),
	.sink_start(sink_start),
	.empty_dff(empty_dff),
	.sink_stall(sink_stall),
	.rdreq(rdreq),
	.sink_staterun1(sink_staterun1),
	.sink_stateend1(sink_stateend1),
	.wrreq(wrreq),
	.counter_reg_bit_0(counter_reg_bit_0),
	.data({gnd,gnd,data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.fifo_wrreq(fifo_wrreq),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module fft_scfifo_nch1 (
	q,
	dffe_af1,
	sink_out_stateempty_and_ready,
	sink_ready_ctrl,
	sink_out_statenormal,
	sink_start,
	empty_dff,
	sink_stall,
	rdreq,
	sink_staterun1,
	sink_stateend1,
	wrreq,
	counter_reg_bit_0,
	data,
	fifo_wrreq,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[17:0] q;
output 	dffe_af1;
input 	sink_out_stateempty_and_ready;
input 	sink_ready_ctrl;
input 	sink_out_statenormal;
input 	sink_start;
output 	empty_dff;
input 	sink_stall;
input 	rdreq;
input 	sink_staterun1;
input 	sink_stateend1;
input 	wrreq;
output 	counter_reg_bit_0;
input 	[17:0] data;
input 	fifo_wrreq;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \dpfifo|usedw_counter|counter_reg_bit[2]~q ;
wire \dpfifo|usedw_counter|counter_reg_bit[1]~q ;
wire \dffe_af~0_combout ;
wire \dffe_af~1_combout ;


fft_a_dpfifo_gn81 dpfifo(
	.q({q_unconnected_wire_17,q_unconnected_wire_16,q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.counter_reg_bit_2(\dpfifo|usedw_counter|counter_reg_bit[2]~q ),
	.counter_reg_bit_1(\dpfifo|usedw_counter|counter_reg_bit[1]~q ),
	.sink_out_stateempty_and_ready(sink_out_stateempty_and_ready),
	.sink_ready_ctrl(sink_ready_ctrl),
	.sink_out_statenormal(sink_out_statenormal),
	.sink_start(sink_start),
	.empty_dff1(empty_dff),
	.sink_stall(sink_stall),
	.rreq(rdreq),
	.sink_staterun1(sink_staterun1),
	.sink_stateend1(sink_stateend1),
	.wreq(wrreq),
	.counter_reg_bit_0(counter_reg_bit_0),
	.data({gnd,gnd,data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.wreq1(fifo_wrreq),
	.clock(clock),
	.reset_n(reset_n));

dffeas dffe_af(
	.clk(clock),
	.d(\dffe_af~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe_af1),
	.prn(vcc));
defparam dffe_af.is_wysiwyg = "true";
defparam dffe_af.power_up = "low";

cycloneiii_lcell_comb \dffe_af~0 (
	.dataa(rdreq),
	.datab(wrreq),
	.datac(dffe_af1),
	.datad(counter_reg_bit_0),
	.cin(gnd),
	.combout(\dffe_af~0_combout ),
	.cout());
defparam \dffe_af~0 .lut_mask = 16'hFDFF;
defparam \dffe_af~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \dffe_af~1 (
	.dataa(dffe_af1),
	.datab(\dpfifo|usedw_counter|counter_reg_bit[2]~q ),
	.datac(\dpfifo|usedw_counter|counter_reg_bit[1]~q ),
	.datad(\dffe_af~0_combout ),
	.cin(gnd),
	.combout(\dffe_af~1_combout ),
	.cout());
defparam \dffe_af~1 .lut_mask = 16'hFFBE;
defparam \dffe_af~1 .sum_lutc_input = "datac";

endmodule

module fft_a_dpfifo_gn81 (
	q,
	counter_reg_bit_2,
	counter_reg_bit_1,
	sink_out_stateempty_and_ready,
	sink_ready_ctrl,
	sink_out_statenormal,
	sink_start,
	empty_dff1,
	sink_stall,
	rreq,
	sink_staterun1,
	sink_stateend1,
	wreq,
	counter_reg_bit_0,
	data,
	wreq1,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[17:0] q;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
input 	sink_out_stateempty_and_ready;
input 	sink_ready_ctrl;
input 	sink_out_statenormal;
input 	sink_start;
output 	empty_dff1;
input 	sink_stall;
input 	rreq;
input 	sink_staterun1;
input 	sink_stateend1;
input 	wreq;
output 	counter_reg_bit_0;
input 	[17:0] data;
input 	wreq1;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \_~2_combout ;
wire \usedw_is_1_dff~q ;
wire \usedw_will_be_1~3_combout ;
wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \low_addressa[0]~q ;
wire \rd_ptr_lsb~q ;
wire \ram_read_address[0]~0_combout ;
wire \rd_ptr_msb|counter_reg_bit[0]~q ;
wire \low_addressa[1]~q ;
wire \ram_read_address[1]~1_combout ;
wire \rd_ptr_msb|counter_reg_bit[1]~q ;
wire \low_addressa[2]~q ;
wire \ram_read_address[2]~2_combout ;
wire \_~7_combout ;
wire \_~8_combout ;
wire \_~9_combout ;
wire \usedw_will_be_1~4_combout ;
wire \rd_ptr_lsb~0_combout ;
wire \usedw_is_0_dff~q ;
wire \_~3_combout ;
wire \_~4_combout ;
wire \_~5_combout ;
wire \usedw_will_be_1~2_combout ;
wire \_~6_combout ;


fft_cntr_lmb wr_ptr(
	.fifo_wrreq(wreq),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.clock(clock),
	.reset_n(reset_n));

fft_cntr_1n7 usedw_counter(
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	._(\_~2_combout ),
	.updown(wreq1),
	.clock(clock),
	.reset_n(reset_n));

fft_cntr_kmb rd_ptr_msb(
	.counter_reg_bit_0(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_msb|counter_reg_bit[1]~q ),
	._(\_~8_combout ),
	.clock(clock),
	.reset_n(reset_n));

fft_altsyncram_nrf1 FIFOram(
	.q_b({q_b_unconnected_wire_17,q_b_unconnected_wire_16,q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.clocken1(rreq),
	.wren_a(wreq),
	.data_a({gnd,gnd,data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.address_a({\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.address_b({\ram_read_address[2]~2_combout ,\ram_read_address[1]~1_combout ,\ram_read_address[0]~0_combout }),
	.clock0(clock),
	.clock1(clock));

cycloneiii_lcell_comb \_~2 (
	.dataa(wreq),
	.datab(sink_out_stateempty_and_ready),
	.datac(sink_ready_ctrl),
	.datad(\_~9_combout ),
	.cin(gnd),
	.combout(\_~2_combout ),
	.cout());
defparam \_~2 .lut_mask = 16'h6996;
defparam \_~2 .sum_lutc_input = "datac";

dffeas usedw_is_1_dff(
	.clk(clock),
	.d(\usedw_will_be_1~3_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_1_dff~q ),
	.prn(vcc));
defparam usedw_is_1_dff.is_wysiwyg = "true";
defparam usedw_is_1_dff.power_up = "low";

cycloneiii_lcell_comb \usedw_will_be_1~3 (
	.dataa(\usedw_is_1_dff~q ),
	.datab(rreq),
	.datac(wreq),
	.datad(\usedw_will_be_1~4_combout ),
	.cin(gnd),
	.combout(\usedw_will_be_1~3_combout ),
	.cout());
defparam \usedw_will_be_1~3 .lut_mask = 16'hEBBE;
defparam \usedw_will_be_1~3 .sum_lutc_input = "datac";

dffeas \low_addressa[0] (
	.clk(clock),
	.d(\ram_read_address[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[0]~q ),
	.prn(vcc));
defparam \low_addressa[0] .is_wysiwyg = "true";
defparam \low_addressa[0] .power_up = "low";

dffeas rd_ptr_lsb(
	.clk(clock),
	.d(\rd_ptr_lsb~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rreq),
	.q(\rd_ptr_lsb~q ),
	.prn(vcc));
defparam rd_ptr_lsb.is_wysiwyg = "true";
defparam rd_ptr_lsb.power_up = "low";

cycloneiii_lcell_comb \ram_read_address[0]~0 (
	.dataa(\low_addressa[0]~q ),
	.datab(gnd),
	.datac(rreq),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\ram_read_address[0]~0_combout ),
	.cout());
defparam \ram_read_address[0]~0 .lut_mask = 16'hA0AF;
defparam \ram_read_address[0]~0 .sum_lutc_input = "datac";

dffeas \low_addressa[1] (
	.clk(clock),
	.d(\ram_read_address[1]~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[1]~q ),
	.prn(vcc));
defparam \low_addressa[1] .is_wysiwyg = "true";
defparam \low_addressa[1] .power_up = "low";

cycloneiii_lcell_comb \ram_read_address[1]~1 (
	.dataa(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datab(\low_addressa[1]~q ),
	.datac(gnd),
	.datad(rreq),
	.cin(gnd),
	.combout(\ram_read_address[1]~1_combout ),
	.cout());
defparam \ram_read_address[1]~1 .lut_mask = 16'hAACC;
defparam \ram_read_address[1]~1 .sum_lutc_input = "datac";

dffeas \low_addressa[2] (
	.clk(clock),
	.d(\ram_read_address[2]~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[2]~q ),
	.prn(vcc));
defparam \low_addressa[2] .is_wysiwyg = "true";
defparam \low_addressa[2] .power_up = "low";

cycloneiii_lcell_comb \ram_read_address[2]~2 (
	.dataa(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datab(\low_addressa[2]~q ),
	.datac(gnd),
	.datad(rreq),
	.cin(gnd),
	.combout(\ram_read_address[2]~2_combout ),
	.cout());
defparam \ram_read_address[2]~2 .lut_mask = 16'hAACC;
defparam \ram_read_address[2]~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \_~7 (
	.dataa(\rd_ptr_lsb~q ),
	.datab(sink_out_stateempty_and_ready),
	.datac(sink_out_statenormal),
	.datad(gnd),
	.cin(gnd),
	.combout(\_~7_combout ),
	.cout());
defparam \_~7 .lut_mask = 16'hDFDF;
defparam \_~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \_~8 (
	.dataa(sink_out_stateempty_and_ready),
	.datab(sink_ready_ctrl),
	.datac(sink_stall),
	.datad(\_~7_combout ),
	.cin(gnd),
	.combout(\_~8_combout ),
	.cout());
defparam \_~8 .lut_mask = 16'hFFEF;
defparam \_~8 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \_~9 (
	.dataa(sink_start),
	.datab(empty_dff1),
	.datac(sink_out_stateempty_and_ready),
	.datad(sink_out_statenormal),
	.cin(gnd),
	.combout(\_~9_combout ),
	.cout());
defparam \_~9 .lut_mask = 16'hFEFF;
defparam \_~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \usedw_will_be_1~4 (
	.dataa(sink_staterun1),
	.datab(sink_stateend1),
	.datac(\_~4_combout ),
	.datad(\usedw_is_0_dff~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~4_combout ),
	.cout());
defparam \usedw_will_be_1~4 .lut_mask = 16'hFFF6;
defparam \usedw_will_be_1~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rd_ptr_lsb~0 (
	.dataa(\rd_ptr_lsb~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\rd_ptr_lsb~0_combout ),
	.cout());
defparam \rd_ptr_lsb~0 .lut_mask = 16'h5555;
defparam \rd_ptr_lsb~0 .sum_lutc_input = "datac";

dffeas empty_dff(
	.clk(clock),
	.d(\_~6_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(empty_dff1),
	.prn(vcc));
defparam empty_dff.is_wysiwyg = "true";
defparam empty_dff.power_up = "low";

dffeas usedw_is_0_dff(
	.clk(clock),
	.d(\_~3_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_0_dff~q ),
	.prn(vcc));
defparam usedw_is_0_dff.is_wysiwyg = "true";
defparam usedw_is_0_dff.power_up = "low";

cycloneiii_lcell_comb \_~3 (
	.dataa(\usedw_is_1_dff~q ),
	.datab(rreq),
	.datac(wreq),
	.datad(\usedw_is_0_dff~q ),
	.cin(gnd),
	.combout(\_~3_combout ),
	.cout());
defparam \_~3 .lut_mask = 16'hFF7D;
defparam \_~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \_~4 (
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(counter_reg_bit_0),
	.datad(counter_reg_bit_2),
	.cin(gnd),
	.combout(\_~4_combout ),
	.cout());
defparam \_~4 .lut_mask = 16'hAFFF;
defparam \_~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \_~5 (
	.dataa(rreq),
	.datab(\_~4_combout ),
	.datac(sink_staterun1),
	.datad(sink_stateend1),
	.cin(gnd),
	.combout(\_~5_combout ),
	.cout());
defparam \_~5 .lut_mask = 16'hEFFF;
defparam \_~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \usedw_will_be_1~2 (
	.dataa(\usedw_is_1_dff~q ),
	.datab(\usedw_is_0_dff~q ),
	.datac(rreq),
	.datad(wreq),
	.cin(gnd),
	.combout(\usedw_will_be_1~2_combout ),
	.cout());
defparam \usedw_will_be_1~2 .lut_mask = 16'hBFFB;
defparam \usedw_will_be_1~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \_~6 (
	.dataa(\_~3_combout ),
	.datab(\_~5_combout ),
	.datac(\usedw_will_be_1~2_combout ),
	.datad(wreq),
	.cin(gnd),
	.combout(\_~6_combout ),
	.cout());
defparam \_~6 .lut_mask = 16'hBFFF;
defparam \_~6 .sum_lutc_input = "datac";

endmodule

module fft_altsyncram_nrf1 (
	q_b,
	clocken1,
	wren_a,
	data_a,
	address_a,
	address_b,
	clock0,
	clock1)/* synthesis synthesis_greybox=1 */;
output 	[17:0] q_b;
input 	clocken1;
input 	wren_a;
input 	[17:0] data_a;
input 	[2:0] address_a;
input 	[2:0] address_b;
input 	clock0;
input 	clock1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

cycloneiii_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.clk1_output_clock_enable = "ena1";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|auk_dspip_avalon_streaming_sink_fft_120:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_nch1:auto_generated|a_dpfifo_gn81:dpfifo|altsyncram_nrf1:FIFOram|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 3;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 7;
defparam ram_block1a2.port_a_logical_ram_depth = 8;
defparam ram_block1a2.port_a_logical_ram_width = 18;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 3;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "clock1";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 7;
defparam ram_block1a2.port_b_logical_ram_depth = 8;
defparam ram_block1a2.port_b_logical_ram_width = 18;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk1_output_clock_enable = "ena1";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|auk_dspip_avalon_streaming_sink_fft_120:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_nch1:auto_generated|a_dpfifo_gn81:dpfifo|altsyncram_nrf1:FIFOram|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 3;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 7;
defparam ram_block1a10.port_a_logical_ram_depth = 8;
defparam ram_block1a10.port_a_logical_ram_width = 18;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 3;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "clock1";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 7;
defparam ram_block1a10.port_b_logical_ram_depth = 8;
defparam ram_block1a10.port_b_logical_ram_width = 18;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk1_output_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|auk_dspip_avalon_streaming_sink_fft_120:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_nch1:auto_generated|a_dpfifo_gn81:dpfifo|altsyncram_nrf1:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 3;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 7;
defparam ram_block1a6.port_a_logical_ram_depth = 8;
defparam ram_block1a6.port_a_logical_ram_width = 18;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 3;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "clock1";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 7;
defparam ram_block1a6.port_b_logical_ram_depth = 8;
defparam ram_block1a6.port_b_logical_ram_width = 18;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk1_output_clock_enable = "ena1";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|auk_dspip_avalon_streaming_sink_fft_120:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_nch1:auto_generated|a_dpfifo_gn81:dpfifo|altsyncram_nrf1:FIFOram|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 3;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 7;
defparam ram_block1a14.port_a_logical_ram_depth = 8;
defparam ram_block1a14.port_a_logical_ram_width = 18;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 3;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "clock1";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 7;
defparam ram_block1a14.port_b_logical_ram_depth = 8;
defparam ram_block1a14.port_b_logical_ram_width = 18;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.clk1_output_clock_enable = "ena1";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|auk_dspip_avalon_streaming_sink_fft_120:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_nch1:auto_generated|a_dpfifo_gn81:dpfifo|altsyncram_nrf1:FIFOram|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 3;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 7;
defparam ram_block1a4.port_a_logical_ram_depth = 8;
defparam ram_block1a4.port_a_logical_ram_width = 18;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 3;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "clock1";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 7;
defparam ram_block1a4.port_b_logical_ram_depth = 8;
defparam ram_block1a4.port_b_logical_ram_width = 18;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk1_output_clock_enable = "ena1";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|auk_dspip_avalon_streaming_sink_fft_120:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_nch1:auto_generated|a_dpfifo_gn81:dpfifo|altsyncram_nrf1:FIFOram|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 3;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 7;
defparam ram_block1a12.port_a_logical_ram_depth = 8;
defparam ram_block1a12.port_a_logical_ram_width = 18;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 3;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "clock1";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 7;
defparam ram_block1a12.port_b_logical_ram_depth = 8;
defparam ram_block1a12.port_b_logical_ram_width = 18;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.clk1_output_clock_enable = "ena1";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|auk_dspip_avalon_streaming_sink_fft_120:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_nch1:auto_generated|a_dpfifo_gn81:dpfifo|altsyncram_nrf1:FIFOram|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 3;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 7;
defparam ram_block1a3.port_a_logical_ram_depth = 8;
defparam ram_block1a3.port_a_logical_ram_width = 18;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 3;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "clock1";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 7;
defparam ram_block1a3.port_b_logical_ram_depth = 8;
defparam ram_block1a3.port_b_logical_ram_width = 18;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk1_output_clock_enable = "ena1";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|auk_dspip_avalon_streaming_sink_fft_120:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_nch1:auto_generated|a_dpfifo_gn81:dpfifo|altsyncram_nrf1:FIFOram|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 3;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 7;
defparam ram_block1a11.port_a_logical_ram_depth = 8;
defparam ram_block1a11.port_a_logical_ram_width = 18;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 3;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "clock1";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 7;
defparam ram_block1a11.port_b_logical_ram_depth = 8;
defparam ram_block1a11.port_b_logical_ram_width = 18;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk1_output_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|auk_dspip_avalon_streaming_sink_fft_120:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_nch1:auto_generated|a_dpfifo_gn81:dpfifo|altsyncram_nrf1:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 3;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 7;
defparam ram_block1a5.port_a_logical_ram_depth = 8;
defparam ram_block1a5.port_a_logical_ram_width = 18;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 3;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "clock1";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 7;
defparam ram_block1a5.port_b_logical_ram_depth = 8;
defparam ram_block1a5.port_b_logical_ram_width = 18;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk1_output_clock_enable = "ena1";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|auk_dspip_avalon_streaming_sink_fft_120:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_nch1:auto_generated|a_dpfifo_gn81:dpfifo|altsyncram_nrf1:FIFOram|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 3;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 7;
defparam ram_block1a13.port_a_logical_ram_depth = 8;
defparam ram_block1a13.port_a_logical_ram_width = 18;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 3;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "clock1";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 7;
defparam ram_block1a13.port_b_logical_ram_depth = 8;
defparam ram_block1a13.port_b_logical_ram_width = 18;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.clk1_output_clock_enable = "ena1";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|auk_dspip_avalon_streaming_sink_fft_120:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_nch1:auto_generated|a_dpfifo_gn81:dpfifo|altsyncram_nrf1:FIFOram|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 3;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 7;
defparam ram_block1a1.port_a_logical_ram_depth = 8;
defparam ram_block1a1.port_a_logical_ram_width = 18;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 3;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "clock1";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 7;
defparam ram_block1a1.port_b_logical_ram_depth = 8;
defparam ram_block1a1.port_b_logical_ram_width = 18;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk1_output_clock_enable = "ena1";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|auk_dspip_avalon_streaming_sink_fft_120:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_nch1:auto_generated|a_dpfifo_gn81:dpfifo|altsyncram_nrf1:FIFOram|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 3;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 7;
defparam ram_block1a9.port_a_logical_ram_depth = 8;
defparam ram_block1a9.port_a_logical_ram_width = 18;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 3;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "clock1";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 7;
defparam ram_block1a9.port_b_logical_ram_depth = 8;
defparam ram_block1a9.port_b_logical_ram_width = 18;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.clk1_output_clock_enable = "ena1";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|auk_dspip_avalon_streaming_sink_fft_120:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_nch1:auto_generated|a_dpfifo_gn81:dpfifo|altsyncram_nrf1:FIFOram|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 3;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 7;
defparam ram_block1a0.port_a_logical_ram_depth = 8;
defparam ram_block1a0.port_a_logical_ram_width = 18;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 3;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "clock1";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 7;
defparam ram_block1a0.port_b_logical_ram_depth = 8;
defparam ram_block1a0.port_b_logical_ram_width = 18;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk1_output_clock_enable = "ena1";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|auk_dspip_avalon_streaming_sink_fft_120:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_nch1:auto_generated|a_dpfifo_gn81:dpfifo|altsyncram_nrf1:FIFOram|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 3;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 7;
defparam ram_block1a8.port_a_logical_ram_depth = 8;
defparam ram_block1a8.port_a_logical_ram_width = 18;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 3;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "clock1";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 7;
defparam ram_block1a8.port_b_logical_ram_depth = 8;
defparam ram_block1a8.port_b_logical_ram_width = 18;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk1_output_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|auk_dspip_avalon_streaming_sink_fft_120:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_nch1:auto_generated|a_dpfifo_gn81:dpfifo|altsyncram_nrf1:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 3;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 7;
defparam ram_block1a7.port_a_logical_ram_depth = 8;
defparam ram_block1a7.port_a_logical_ram_width = 18;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 3;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "clock1";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 7;
defparam ram_block1a7.port_b_logical_ram_depth = 8;
defparam ram_block1a7.port_b_logical_ram_width = 18;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk1_output_clock_enable = "ena1";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "asj_fft_sglstream_fft_120:asj_fft_sglstream_fft_120_inst|auk_dspip_avalon_streaming_sink_fft_120:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_nch1:auto_generated|a_dpfifo_gn81:dpfifo|altsyncram_nrf1:FIFOram|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 3;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 7;
defparam ram_block1a15.port_a_logical_ram_depth = 8;
defparam ram_block1a15.port_a_logical_ram_width = 18;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 3;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "clock1";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 7;
defparam ram_block1a15.port_b_logical_ram_depth = 8;
defparam ram_block1a15.port_b_logical_ram_width = 18;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";

endmodule

module fft_cntr_1n7 (
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	_,
	updown,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
input 	_;
input 	updown;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita0~combout ;


dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

cycloneiii_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h5566;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneiii_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A6F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneiii_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout());
defparam counter_comb_bita2.lut_mask = 16'h5A5A;
defparam counter_comb_bita2.sum_lutc_input = "cin";

endmodule

module fft_cntr_kmb (
	counter_reg_bit_0,
	counter_reg_bit_1,
	_,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
input 	_;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

cycloneiii_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneiii_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout());
defparam counter_comb_bita1.lut_mask = 16'h5A5A;
defparam counter_comb_bita1.sum_lutc_input = "cin";

endmodule

module fft_cntr_lmb (
	fifo_wrreq,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	fifo_wrreq;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wrreq),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wrreq),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wrreq),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

cycloneiii_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneiii_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneiii_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout());
defparam counter_comb_bita2.lut_mask = 16'h5A5A;
defparam counter_comb_bita2.sum_lutc_input = "cin";

endmodule

module fft_auk_dspip_avalon_streaming_source_fft_120 (
	data_count,
	at_source_error_0,
	at_source_error_1,
	at_source_sop_s1,
	at_source_eop_s1,
	at_source_valid_s1,
	at_source_data_0,
	at_source_data_1,
	at_source_data_2,
	at_source_data_3,
	at_source_data_4,
	at_source_data_5,
	at_source_data_14,
	at_source_data_15,
	at_source_data_16,
	at_source_data_17,
	at_source_data_18,
	at_source_data_19,
	at_source_data_20,
	at_source_data_21,
	at_source_data_6,
	at_source_data_7,
	at_source_data_8,
	at_source_data_9,
	at_source_data_10,
	at_source_data_11,
	at_source_data_12,
	at_source_data_13,
	source_packet_error_0,
	source_packet_error_1,
	valid_ctrl_int2,
	source_stall_reg,
	master_source_ena,
	source_valid_ctrl_sop,
	Mux3,
	source_valid_ctrl_sop1,
	stall_reg,
	source_stall_int_d1,
	data,
	Mux0,
	Mux01,
	clk,
	reset_n,
	source_ready)/* synthesis synthesis_greybox=1 */;
input 	[8:0] data_count;
output 	at_source_error_0;
output 	at_source_error_1;
output 	at_source_sop_s1;
output 	at_source_eop_s1;
output 	at_source_valid_s1;
output 	at_source_data_0;
output 	at_source_data_1;
output 	at_source_data_2;
output 	at_source_data_3;
output 	at_source_data_4;
output 	at_source_data_5;
output 	at_source_data_14;
output 	at_source_data_15;
output 	at_source_data_16;
output 	at_source_data_17;
output 	at_source_data_18;
output 	at_source_data_19;
output 	at_source_data_20;
output 	at_source_data_21;
output 	at_source_data_6;
output 	at_source_data_7;
output 	at_source_data_8;
output 	at_source_data_9;
output 	at_source_data_10;
output 	at_source_data_11;
output 	at_source_data_12;
output 	at_source_data_13;
input 	source_packet_error_0;
input 	source_packet_error_1;
output 	valid_ctrl_int2;
input 	source_stall_reg;
input 	master_source_ena;
input 	source_valid_ctrl_sop;
output 	Mux3;
input 	source_valid_ctrl_sop1;
input 	stall_reg;
output 	source_stall_int_d1;
input 	[21:0] data;
output 	Mux0;
output 	Mux01;
input 	clk;
input 	reset_n;
input 	source_ready;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \data_count_int[1]~q ;
wire \count_finished~0_combout ;
wire \data_count_int1[1]~q ;
wire \count_finished~1_combout ;
wire \count_finished~2_combout ;
wire \data_count_int1[8]~q ;
wire \Selector3~0_combout ;
wire \Mux2~2_combout ;
wire \source_state.st_err~q ;
wire \Selector2~8_combout ;
wire \packet_error0~combout ;
wire \Selector1~0_combout ;
wire \Selector1~1_combout ;
wire \source_state.sop~q ;
wire \Mux3~1_combout ;
wire \data_count_int1[6]~q ;
wire \first_data~0_combout ;
wire \first_data~q ;
wire \data_select~0_combout ;
wire \Mux1~0_combout ;
wire \valid_ctrl_inter1~0_combout ;
wire \valid_ctrl_int1~q ;
wire \Mux2~3_combout ;
wire \Mux2~0_combout ;
wire \Mux2~4_combout ;
wire \data_count_int[6]~q ;
wire \data_count_int[4]~q ;
wire \data_count_int[5]~q ;
wire \count_finished~3_combout ;
wire \data_count_int1[4]~q ;
wire \data_count_int1[5]~q ;
wire \count_finished~4_combout ;
wire \count_finished~5_combout ;
wire \valid_ctrl_int_selected~0_combout ;
wire \data_count_int[8]~q ;
wire \data_count_int_selected[8]~0_combout ;
wire \count_finished~combout ;
wire \Selector1~2_combout ;
wire \Selector2~7_combout ;
wire \Selector1~5_combout ;
wire \Selector2~6_combout ;
wire \source_state.run1~q ;
wire \Selector3~1_combout ;
wire \Selector3~2_combout ;
wire \source_state.end1~q ;
wire \data_count_int1[3]~q ;
wire \data_count_int[3]~q ;
wire \data_count_int[2]~q ;
wire \data_count_int[0]~q ;
wire \source_comb_update_2~0_combout ;
wire \data_count_int1[2]~q ;
wire \data_count_int1[0]~q ;
wire \source_comb_update_2~1_combout ;
wire \source_comb_update_2~2_combout ;
wire \data_count_int[7]~q ;
wire \source_comb_update_2~3_combout ;
wire \data_count_int1[7]~q ;
wire \source_comb_update_2~4_combout ;
wire \source_comb_update_2~5_combout ;
wire \source_comb_update_2~6_combout ;
wire \Selector0~1_combout ;
wire \source_state.start~q ;
wire \Selector0~0_combout ;
wire \Selector1~3_combout ;
wire \Selector1~4_combout ;
wire \Selector5~0_combout ;
wire \Selector5~1_combout ;
wire \at_source_valid_int~0_combout ;
wire \at_source_valid_int~1_combout ;
wire \at_source_valid_int~2_combout ;
wire \at_source_valid_int~3_combout ;
wire \data_int1[0]~q ;
wire \data_int[0]~q ;
wire \data_int_selected[0]~0_combout ;
wire \data_int1[1]~q ;
wire \data_int[1]~q ;
wire \data_int_selected[1]~1_combout ;
wire \data_int1[2]~q ;
wire \data_int[2]~q ;
wire \data_int_selected[2]~2_combout ;
wire \data_int1[3]~q ;
wire \data_int[3]~q ;
wire \data_int_selected[3]~3_combout ;
wire \data_int1[4]~q ;
wire \data_int[4]~q ;
wire \data_int_selected[4]~4_combout ;
wire \data_int1[5]~q ;
wire \data_int[5]~q ;
wire \data_int_selected[5]~5_combout ;
wire \data_int1[14]~q ;
wire \data_int[14]~q ;
wire \data_int_selected[14]~6_combout ;
wire \data_int1[15]~q ;
wire \data_int[15]~q ;
wire \data_int_selected[15]~7_combout ;
wire \data_int1[16]~q ;
wire \data_int[16]~q ;
wire \data_int_selected[16]~8_combout ;
wire \data_int1[17]~q ;
wire \data_int[17]~q ;
wire \data_int_selected[17]~9_combout ;
wire \data_int1[18]~q ;
wire \data_int[18]~q ;
wire \data_int_selected[18]~10_combout ;
wire \data_int1[19]~q ;
wire \data_int[19]~q ;
wire \data_int_selected[19]~11_combout ;
wire \data_int1[20]~q ;
wire \data_int[20]~q ;
wire \data_int_selected[20]~12_combout ;
wire \data_int1[21]~q ;
wire \data_int[21]~q ;
wire \data_int_selected[21]~13_combout ;
wire \data_int1[6]~q ;
wire \data_int[6]~q ;
wire \data_int_selected[6]~14_combout ;
wire \data_int1[7]~q ;
wire \data_int[7]~q ;
wire \data_int_selected[7]~15_combout ;
wire \data_int1[8]~q ;
wire \data_int[8]~q ;
wire \data_int_selected[8]~16_combout ;
wire \data_int1[9]~q ;
wire \data_int[9]~q ;
wire \data_int_selected[9]~17_combout ;
wire \data_int1[10]~q ;
wire \data_int[10]~q ;
wire \data_int_selected[10]~18_combout ;
wire \data_int1[11]~q ;
wire \data_int[11]~q ;
wire \data_int_selected[11]~19_combout ;
wire \data_int1[12]~q ;
wire \data_int[12]~q ;
wire \data_int_selected[12]~20_combout ;
wire \data_int1[13]~q ;
wire \data_int[13]~q ;
wire \data_int_selected[13]~21_combout ;
wire \valid_ctrl_inter~0_combout ;
wire \was_stalled~0_combout ;
wire \was_stalled~1_combout ;
wire \was_stalled~q ;
wire \valid_ctrl_inter~1_combout ;
wire \Mux2~1_combout ;
wire \Mux0~1_combout ;


dffeas \data_count_int[1] (
	.clk(clk),
	.d(data_count[1]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_count_int[1]~q ),
	.prn(vcc));
defparam \data_count_int[1] .is_wysiwyg = "true";
defparam \data_count_int[1] .power_up = "low";

cycloneiii_lcell_comb \count_finished~0 (
	.dataa(\data_count_int[2]~q ),
	.datab(\data_count_int[1]~q ),
	.datac(\data_count_int[3]~q ),
	.datad(\data_count_int[0]~q ),
	.cin(gnd),
	.combout(\count_finished~0_combout ),
	.cout());
defparam \count_finished~0 .lut_mask = 16'h7FFF;
defparam \count_finished~0 .sum_lutc_input = "datac";

dffeas \data_count_int1[1] (
	.clk(clk),
	.d(data_count[1]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_count_int1[1]~q ),
	.prn(vcc));
defparam \data_count_int1[1] .is_wysiwyg = "true";
defparam \data_count_int1[1] .power_up = "low";

cycloneiii_lcell_comb \count_finished~1 (
	.dataa(\data_count_int1[2]~q ),
	.datab(\data_count_int1[1]~q ),
	.datac(\data_count_int1[0]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\count_finished~1_combout ),
	.cout());
defparam \count_finished~1 .lut_mask = 16'h7F7F;
defparam \count_finished~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \count_finished~2 (
	.dataa(\data_select~0_combout ),
	.datab(\data_count_int1[3]~q ),
	.datac(\count_finished~0_combout ),
	.datad(\count_finished~1_combout ),
	.cin(gnd),
	.combout(\count_finished~2_combout ),
	.cout());
defparam \count_finished~2 .lut_mask = 16'hF7B3;
defparam \count_finished~2 .sum_lutc_input = "datac";

dffeas \data_count_int1[8] (
	.clk(clk),
	.d(data_count[8]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_count_int1[8]~q ),
	.prn(vcc));
defparam \data_count_int1[8] .is_wysiwyg = "true";
defparam \data_count_int1[8] .power_up = "low";

cycloneiii_lcell_comb \Selector3~0 (
	.dataa(\source_state.end1~q ),
	.datab(at_source_valid_s1),
	.datac(source_ready),
	.datad(\packet_error0~combout ),
	.cin(gnd),
	.combout(\Selector3~0_combout ),
	.cout());
defparam \Selector3~0 .lut_mask = 16'hBFFF;
defparam \Selector3~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux2~2 (
	.dataa(master_source_ena),
	.datab(source_valid_ctrl_sop),
	.datac(source_stall_reg),
	.datad(\was_stalled~q ),
	.cin(gnd),
	.combout(\Mux2~2_combout ),
	.cout());
defparam \Mux2~2 .lut_mask = 16'hEFFF;
defparam \Mux2~2 .sum_lutc_input = "datac";

dffeas \source_state.st_err (
	.clk(clk),
	.d(\packet_error0~combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\source_state.st_err~q ),
	.prn(vcc));
defparam \source_state.st_err .is_wysiwyg = "true";
defparam \source_state.st_err .power_up = "low";

cycloneiii_lcell_comb \Selector2~8 (
	.dataa(source_packet_error_0),
	.datab(source_packet_error_1),
	.datac(\source_state.sop~q ),
	.datad(\count_finished~combout ),
	.cin(gnd),
	.combout(\Selector2~8_combout ),
	.cout());
defparam \Selector2~8 .lut_mask = 16'hFFF7;
defparam \Selector2~8 .sum_lutc_input = "datac";

dffeas \at_source_error[0] (
	.clk(clk),
	.d(source_packet_error_0),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(at_source_error_0),
	.prn(vcc));
defparam \at_source_error[0] .is_wysiwyg = "true";
defparam \at_source_error[0] .power_up = "low";

dffeas \at_source_error[1] (
	.clk(clk),
	.d(source_packet_error_1),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(at_source_error_1),
	.prn(vcc));
defparam \at_source_error[1] .is_wysiwyg = "true";
defparam \at_source_error[1] .power_up = "low";

dffeas at_source_sop_s(
	.clk(clk),
	.d(\Selector1~4_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(at_source_sop_s1),
	.prn(vcc));
defparam at_source_sop_s.is_wysiwyg = "true";
defparam at_source_sop_s.power_up = "low";

dffeas at_source_eop_s(
	.clk(clk),
	.d(\Selector5~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(at_source_eop_s1),
	.prn(vcc));
defparam at_source_eop_s.is_wysiwyg = "true";
defparam at_source_eop_s.power_up = "low";

dffeas at_source_valid_s(
	.clk(clk),
	.d(\at_source_valid_int~3_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(at_source_valid_s1),
	.prn(vcc));
defparam at_source_valid_s.is_wysiwyg = "true";
defparam at_source_valid_s.power_up = "low";

dffeas \at_source_data[0] (
	.clk(clk),
	.d(\data_int_selected[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_0),
	.prn(vcc));
defparam \at_source_data[0] .is_wysiwyg = "true";
defparam \at_source_data[0] .power_up = "low";

dffeas \at_source_data[1] (
	.clk(clk),
	.d(\data_int_selected[1]~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_1),
	.prn(vcc));
defparam \at_source_data[1] .is_wysiwyg = "true";
defparam \at_source_data[1] .power_up = "low";

dffeas \at_source_data[2] (
	.clk(clk),
	.d(\data_int_selected[2]~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_2),
	.prn(vcc));
defparam \at_source_data[2] .is_wysiwyg = "true";
defparam \at_source_data[2] .power_up = "low";

dffeas \at_source_data[3] (
	.clk(clk),
	.d(\data_int_selected[3]~3_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_3),
	.prn(vcc));
defparam \at_source_data[3] .is_wysiwyg = "true";
defparam \at_source_data[3] .power_up = "low";

dffeas \at_source_data[4] (
	.clk(clk),
	.d(\data_int_selected[4]~4_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_4),
	.prn(vcc));
defparam \at_source_data[4] .is_wysiwyg = "true";
defparam \at_source_data[4] .power_up = "low";

dffeas \at_source_data[5] (
	.clk(clk),
	.d(\data_int_selected[5]~5_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_5),
	.prn(vcc));
defparam \at_source_data[5] .is_wysiwyg = "true";
defparam \at_source_data[5] .power_up = "low";

dffeas \at_source_data[14] (
	.clk(clk),
	.d(\data_int_selected[14]~6_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_14),
	.prn(vcc));
defparam \at_source_data[14] .is_wysiwyg = "true";
defparam \at_source_data[14] .power_up = "low";

dffeas \at_source_data[15] (
	.clk(clk),
	.d(\data_int_selected[15]~7_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_15),
	.prn(vcc));
defparam \at_source_data[15] .is_wysiwyg = "true";
defparam \at_source_data[15] .power_up = "low";

dffeas \at_source_data[16] (
	.clk(clk),
	.d(\data_int_selected[16]~8_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_16),
	.prn(vcc));
defparam \at_source_data[16] .is_wysiwyg = "true";
defparam \at_source_data[16] .power_up = "low";

dffeas \at_source_data[17] (
	.clk(clk),
	.d(\data_int_selected[17]~9_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_17),
	.prn(vcc));
defparam \at_source_data[17] .is_wysiwyg = "true";
defparam \at_source_data[17] .power_up = "low";

dffeas \at_source_data[18] (
	.clk(clk),
	.d(\data_int_selected[18]~10_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_18),
	.prn(vcc));
defparam \at_source_data[18] .is_wysiwyg = "true";
defparam \at_source_data[18] .power_up = "low";

dffeas \at_source_data[19] (
	.clk(clk),
	.d(\data_int_selected[19]~11_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_19),
	.prn(vcc));
defparam \at_source_data[19] .is_wysiwyg = "true";
defparam \at_source_data[19] .power_up = "low";

dffeas \at_source_data[20] (
	.clk(clk),
	.d(\data_int_selected[20]~12_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_20),
	.prn(vcc));
defparam \at_source_data[20] .is_wysiwyg = "true";
defparam \at_source_data[20] .power_up = "low";

dffeas \at_source_data[21] (
	.clk(clk),
	.d(\data_int_selected[21]~13_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_21),
	.prn(vcc));
defparam \at_source_data[21] .is_wysiwyg = "true";
defparam \at_source_data[21] .power_up = "low";

dffeas \at_source_data[6] (
	.clk(clk),
	.d(\data_int_selected[6]~14_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_6),
	.prn(vcc));
defparam \at_source_data[6] .is_wysiwyg = "true";
defparam \at_source_data[6] .power_up = "low";

dffeas \at_source_data[7] (
	.clk(clk),
	.d(\data_int_selected[7]~15_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_7),
	.prn(vcc));
defparam \at_source_data[7] .is_wysiwyg = "true";
defparam \at_source_data[7] .power_up = "low";

dffeas \at_source_data[8] (
	.clk(clk),
	.d(\data_int_selected[8]~16_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_8),
	.prn(vcc));
defparam \at_source_data[8] .is_wysiwyg = "true";
defparam \at_source_data[8] .power_up = "low";

dffeas \at_source_data[9] (
	.clk(clk),
	.d(\data_int_selected[9]~17_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_9),
	.prn(vcc));
defparam \at_source_data[9] .is_wysiwyg = "true";
defparam \at_source_data[9] .power_up = "low";

dffeas \at_source_data[10] (
	.clk(clk),
	.d(\data_int_selected[10]~18_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_10),
	.prn(vcc));
defparam \at_source_data[10] .is_wysiwyg = "true";
defparam \at_source_data[10] .power_up = "low";

dffeas \at_source_data[11] (
	.clk(clk),
	.d(\data_int_selected[11]~19_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_11),
	.prn(vcc));
defparam \at_source_data[11] .is_wysiwyg = "true";
defparam \at_source_data[11] .power_up = "low";

dffeas \at_source_data[12] (
	.clk(clk),
	.d(\data_int_selected[12]~20_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_12),
	.prn(vcc));
defparam \at_source_data[12] .is_wysiwyg = "true";
defparam \at_source_data[12] .power_up = "low";

dffeas \at_source_data[13] (
	.clk(clk),
	.d(\data_int_selected[13]~21_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_13),
	.prn(vcc));
defparam \at_source_data[13] .is_wysiwyg = "true";
defparam \at_source_data[13] .power_up = "low";

dffeas valid_ctrl_int(
	.clk(clk),
	.d(\valid_ctrl_inter~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(valid_ctrl_int2),
	.prn(vcc));
defparam valid_ctrl_int.is_wysiwyg = "true";
defparam valid_ctrl_int.power_up = "low";

cycloneiii_lcell_comb \Mux3~0 (
	.dataa(\Mux2~1_combout ),
	.datab(source_valid_ctrl_sop),
	.datac(source_stall_reg),
	.datad(\valid_ctrl_int1~q ),
	.cin(gnd),
	.combout(Mux3),
	.cout());
defparam \Mux3~0 .lut_mask = 16'hEFFF;
defparam \Mux3~0 .sum_lutc_input = "datac";

dffeas source_stall_int_d(
	.clk(clk),
	.d(Mux01),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(source_stall_int_d1),
	.prn(vcc));
defparam source_stall_int_d.is_wysiwyg = "true";
defparam source_stall_int_d.power_up = "low";

cycloneiii_lcell_comb \Mux0~0 (
	.dataa(\valid_ctrl_int1~q ),
	.datab(valid_ctrl_int2),
	.datac(\first_data~q ),
	.datad(source_ready),
	.cin(gnd),
	.combout(Mux0),
	.cout());
defparam \Mux0~0 .lut_mask = 16'hEFFF;
defparam \Mux0~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux0~2 (
	.dataa(at_source_valid_s1),
	.datab(Mux0),
	.datac(Mux3),
	.datad(\Mux0~1_combout ),
	.cin(gnd),
	.combout(Mux01),
	.cout());
defparam \Mux0~2 .lut_mask = 16'hFFFE;
defparam \Mux0~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb packet_error0(
	.dataa(source_packet_error_0),
	.datab(source_packet_error_1),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\packet_error0~combout ),
	.cout());
defparam packet_error0.lut_mask = 16'hEEEE;
defparam packet_error0.sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector1~0 (
	.dataa(at_source_valid_s1),
	.datab(gnd),
	.datac(gnd),
	.datad(source_ready),
	.cin(gnd),
	.combout(\Selector1~0_combout ),
	.cout());
defparam \Selector1~0 .lut_mask = 16'hAAFF;
defparam \Selector1~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector1~1 (
	.dataa(\source_state.sop~q ),
	.datab(\Selector1~0_combout ),
	.datac(source_packet_error_0),
	.datad(source_packet_error_1),
	.cin(gnd),
	.combout(\Selector1~1_combout ),
	.cout());
defparam \Selector1~1 .lut_mask = 16'hEFFF;
defparam \Selector1~1 .sum_lutc_input = "datac";

dffeas \source_state.sop (
	.clk(clk),
	.d(\Selector1~4_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\source_state.sop~q ),
	.prn(vcc));
defparam \source_state.sop .is_wysiwyg = "true";
defparam \source_state.sop .power_up = "low";

cycloneiii_lcell_comb \Mux3~1 (
	.dataa(\Mux2~0_combout ),
	.datab(Mux3),
	.datac(gnd),
	.datad(source_ready),
	.cin(gnd),
	.combout(\Mux3~1_combout ),
	.cout());
defparam \Mux3~1 .lut_mask = 16'hEEFF;
defparam \Mux3~1 .sum_lutc_input = "datac";

dffeas \data_count_int1[6] (
	.clk(clk),
	.d(data_count[6]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_count_int1[6]~q ),
	.prn(vcc));
defparam \data_count_int1[6] .is_wysiwyg = "true";
defparam \data_count_int1[6] .power_up = "low";

cycloneiii_lcell_comb \first_data~0 (
	.dataa(\valid_ctrl_int1~q ),
	.datab(\first_data~q ),
	.datac(at_source_valid_s1),
	.datad(source_ready),
	.cin(gnd),
	.combout(\first_data~0_combout ),
	.cout());
defparam \first_data~0 .lut_mask = 16'hEBBE;
defparam \first_data~0 .sum_lutc_input = "datac";

dffeas first_data(
	.clk(clk),
	.d(\first_data~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\first_data~q ),
	.prn(vcc));
defparam first_data.is_wysiwyg = "true";
defparam first_data.power_up = "low";

cycloneiii_lcell_comb \data_select~0 (
	.dataa(at_source_valid_s1),
	.datab(\first_data~q ),
	.datac(\valid_ctrl_int1~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_select~0_combout ),
	.cout());
defparam \data_select~0 .lut_mask = 16'hFEFE;
defparam \data_select~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux1~0 (
	.dataa(source_ready),
	.datab(valid_ctrl_int2),
	.datac(\valid_ctrl_int1~q ),
	.datad(at_source_valid_s1),
	.cin(gnd),
	.combout(\Mux1~0_combout ),
	.cout());
defparam \Mux1~0 .lut_mask = 16'hFAFC;
defparam \Mux1~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \valid_ctrl_inter1~0 (
	.dataa(\Mux3~1_combout ),
	.datab(\valid_ctrl_int1~q ),
	.datac(\data_select~0_combout ),
	.datad(\Mux1~0_combout ),
	.cin(gnd),
	.combout(\valid_ctrl_inter1~0_combout ),
	.cout());
defparam \valid_ctrl_inter1~0 .lut_mask = 16'hEFFF;
defparam \valid_ctrl_inter1~0 .sum_lutc_input = "datac";

dffeas valid_ctrl_int1(
	.clk(clk),
	.d(\valid_ctrl_inter1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\valid_ctrl_int1~q ),
	.prn(vcc));
defparam valid_ctrl_int1.is_wysiwyg = "true";
defparam valid_ctrl_int1.power_up = "low";

cycloneiii_lcell_comb \Mux2~3 (
	.dataa(source_ready),
	.datab(at_source_valid_s1),
	.datac(\first_data~q ),
	.datad(\valid_ctrl_int1~q ),
	.cin(gnd),
	.combout(\Mux2~3_combout ),
	.cout());
defparam \Mux2~3 .lut_mask = 16'hFEFF;
defparam \Mux2~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux2~0 (
	.dataa(at_source_valid_s1),
	.datab(valid_ctrl_int2),
	.datac(\valid_ctrl_int1~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux2~0_combout ),
	.cout());
defparam \Mux2~0 .lut_mask = 16'hFEFE;
defparam \Mux2~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux2~4 (
	.dataa(\Mux2~2_combout ),
	.datab(\Mux2~3_combout ),
	.datac(gnd),
	.datad(\Mux2~0_combout ),
	.cin(gnd),
	.combout(\Mux2~4_combout ),
	.cout());
defparam \Mux2~4 .lut_mask = 16'hEEFF;
defparam \Mux2~4 .sum_lutc_input = "datac";

dffeas \data_count_int[6] (
	.clk(clk),
	.d(data_count[6]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_count_int[6]~q ),
	.prn(vcc));
defparam \data_count_int[6] .is_wysiwyg = "true";
defparam \data_count_int[6] .power_up = "low";

dffeas \data_count_int[4] (
	.clk(clk),
	.d(data_count[4]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_count_int[4]~q ),
	.prn(vcc));
defparam \data_count_int[4] .is_wysiwyg = "true";
defparam \data_count_int[4] .power_up = "low";

dffeas \data_count_int[5] (
	.clk(clk),
	.d(data_count[5]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_count_int[5]~q ),
	.prn(vcc));
defparam \data_count_int[5] .is_wysiwyg = "true";
defparam \data_count_int[5] .power_up = "low";

cycloneiii_lcell_comb \count_finished~3 (
	.dataa(\data_count_int[7]~q ),
	.datab(\data_count_int[6]~q ),
	.datac(\data_count_int[4]~q ),
	.datad(\data_count_int[5]~q ),
	.cin(gnd),
	.combout(\count_finished~3_combout ),
	.cout());
defparam \count_finished~3 .lut_mask = 16'h7FFF;
defparam \count_finished~3 .sum_lutc_input = "datac";

dffeas \data_count_int1[4] (
	.clk(clk),
	.d(data_count[4]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_count_int1[4]~q ),
	.prn(vcc));
defparam \data_count_int1[4] .is_wysiwyg = "true";
defparam \data_count_int1[4] .power_up = "low";

dffeas \data_count_int1[5] (
	.clk(clk),
	.d(data_count[5]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_count_int1[5]~q ),
	.prn(vcc));
defparam \data_count_int1[5] .is_wysiwyg = "true";
defparam \data_count_int1[5] .power_up = "low";

cycloneiii_lcell_comb \count_finished~4 (
	.dataa(\data_count_int1[7]~q ),
	.datab(\data_count_int1[4]~q ),
	.datac(\data_count_int1[5]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\count_finished~4_combout ),
	.cout());
defparam \count_finished~4 .lut_mask = 16'h7F7F;
defparam \count_finished~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \count_finished~5 (
	.dataa(\data_select~0_combout ),
	.datab(\data_count_int1[6]~q ),
	.datac(\count_finished~3_combout ),
	.datad(\count_finished~4_combout ),
	.cin(gnd),
	.combout(\count_finished~5_combout ),
	.cout());
defparam \count_finished~5 .lut_mask = 16'hF7B3;
defparam \count_finished~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \valid_ctrl_int_selected~0 (
	.dataa(valid_ctrl_int2),
	.datab(at_source_valid_s1),
	.datac(\first_data~q ),
	.datad(\valid_ctrl_int1~q ),
	.cin(gnd),
	.combout(\valid_ctrl_int_selected~0_combout ),
	.cout());
defparam \valid_ctrl_int_selected~0 .lut_mask = 16'hFFFE;
defparam \valid_ctrl_int_selected~0 .sum_lutc_input = "datac";

dffeas \data_count_int[8] (
	.clk(clk),
	.d(data_count[8]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_count_int[8]~q ),
	.prn(vcc));
defparam \data_count_int[8] .is_wysiwyg = "true";
defparam \data_count_int[8] .power_up = "low";

cycloneiii_lcell_comb \data_count_int_selected[8]~0 (
	.dataa(\data_count_int1[8]~q ),
	.datab(\data_count_int[8]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_count_int_selected[8]~0_combout ),
	.cout());
defparam \data_count_int_selected[8]~0 .lut_mask = 16'hAACC;
defparam \data_count_int_selected[8]~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb count_finished(
	.dataa(\count_finished~2_combout ),
	.datab(\count_finished~5_combout ),
	.datac(\valid_ctrl_int_selected~0_combout ),
	.datad(\data_count_int_selected[8]~0_combout ),
	.cin(gnd),
	.combout(\count_finished~combout ),
	.cout());
defparam count_finished.lut_mask = 16'hEFFF;
defparam count_finished.sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector1~2 (
	.dataa(at_source_valid_s1),
	.datab(\source_state.sop~q ),
	.datac(\count_finished~combout ),
	.datad(\Selector1~1_combout ),
	.cin(gnd),
	.combout(\Selector1~2_combout ),
	.cout());
defparam \Selector1~2 .lut_mask = 16'hFFD8;
defparam \Selector1~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector2~7 (
	.dataa(at_source_valid_s1),
	.datab(source_ready),
	.datac(\count_finished~combout ),
	.datad(\packet_error0~combout ),
	.cin(gnd),
	.combout(\Selector2~7_combout ),
	.cout());
defparam \Selector2~7 .lut_mask = 16'hFBFF;
defparam \Selector2~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector1~5 (
	.dataa(at_source_valid_s1),
	.datab(source_ready),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector1~5_combout ),
	.cout());
defparam \Selector1~5 .lut_mask = 16'hEEEE;
defparam \Selector1~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector2~6 (
	.dataa(\Selector2~8_combout ),
	.datab(\source_state.run1~q ),
	.datac(\Selector2~7_combout ),
	.datad(\Selector1~5_combout ),
	.cin(gnd),
	.combout(\Selector2~6_combout ),
	.cout());
defparam \Selector2~6 .lut_mask = 16'hFFFE;
defparam \Selector2~6 .sum_lutc_input = "datac";

dffeas \source_state.run1 (
	.clk(clk),
	.d(\Selector2~6_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\source_state.run1~q ),
	.prn(vcc));
defparam \source_state.run1 .is_wysiwyg = "true";
defparam \source_state.run1 .power_up = "low";

cycloneiii_lcell_comb \Selector3~1 (
	.dataa(\source_state.sop~q ),
	.datab(\source_state.run1~q ),
	.datac(source_packet_error_0),
	.datad(source_packet_error_1),
	.cin(gnd),
	.combout(\Selector3~1_combout ),
	.cout());
defparam \Selector3~1 .lut_mask = 16'hEFFF;
defparam \Selector3~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector3~2 (
	.dataa(\Selector3~0_combout ),
	.datab(\Selector3~1_combout ),
	.datac(\count_finished~combout ),
	.datad(\Selector1~0_combout ),
	.cin(gnd),
	.combout(\Selector3~2_combout ),
	.cout());
defparam \Selector3~2 .lut_mask = 16'hEFFF;
defparam \Selector3~2 .sum_lutc_input = "datac";

dffeas \source_state.end1 (
	.clk(clk),
	.d(\Selector3~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\source_state.end1~q ),
	.prn(vcc));
defparam \source_state.end1 .is_wysiwyg = "true";
defparam \source_state.end1 .power_up = "low";

dffeas \data_count_int1[3] (
	.clk(clk),
	.d(data_count[3]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_count_int1[3]~q ),
	.prn(vcc));
defparam \data_count_int1[3] .is_wysiwyg = "true";
defparam \data_count_int1[3] .power_up = "low";

dffeas \data_count_int[3] (
	.clk(clk),
	.d(data_count[3]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_count_int[3]~q ),
	.prn(vcc));
defparam \data_count_int[3] .is_wysiwyg = "true";
defparam \data_count_int[3] .power_up = "low";

dffeas \data_count_int[2] (
	.clk(clk),
	.d(data_count[2]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_count_int[2]~q ),
	.prn(vcc));
defparam \data_count_int[2] .is_wysiwyg = "true";
defparam \data_count_int[2] .power_up = "low";

dffeas \data_count_int[0] (
	.clk(clk),
	.d(data_count[0]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_count_int[0]~q ),
	.prn(vcc));
defparam \data_count_int[0] .is_wysiwyg = "true";
defparam \data_count_int[0] .power_up = "low";

cycloneiii_lcell_comb \source_comb_update_2~0 (
	.dataa(\data_count_int[1]~q ),
	.datab(\data_count_int[3]~q ),
	.datac(\data_count_int[2]~q ),
	.datad(\data_count_int[0]~q ),
	.cin(gnd),
	.combout(\source_comb_update_2~0_combout ),
	.cout());
defparam \source_comb_update_2~0 .lut_mask = 16'h7FFF;
defparam \source_comb_update_2~0 .sum_lutc_input = "datac";

dffeas \data_count_int1[2] (
	.clk(clk),
	.d(data_count[2]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_count_int1[2]~q ),
	.prn(vcc));
defparam \data_count_int1[2] .is_wysiwyg = "true";
defparam \data_count_int1[2] .power_up = "low";

dffeas \data_count_int1[0] (
	.clk(clk),
	.d(data_count[0]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_count_int1[0]~q ),
	.prn(vcc));
defparam \data_count_int1[0] .is_wysiwyg = "true";
defparam \data_count_int1[0] .power_up = "low";

cycloneiii_lcell_comb \source_comb_update_2~1 (
	.dataa(\data_count_int1[1]~q ),
	.datab(\data_count_int1[2]~q ),
	.datac(\data_count_int1[0]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\source_comb_update_2~1_combout ),
	.cout());
defparam \source_comb_update_2~1 .lut_mask = 16'h7F7F;
defparam \source_comb_update_2~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \source_comb_update_2~2 (
	.dataa(\data_select~0_combout ),
	.datab(\data_count_int1[3]~q ),
	.datac(\source_comb_update_2~0_combout ),
	.datad(\source_comb_update_2~1_combout ),
	.cin(gnd),
	.combout(\source_comb_update_2~2_combout ),
	.cout());
defparam \source_comb_update_2~2 .lut_mask = 16'hF7B3;
defparam \source_comb_update_2~2 .sum_lutc_input = "datac";

dffeas \data_count_int[7] (
	.clk(clk),
	.d(data_count[7]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_count_int[7]~q ),
	.prn(vcc));
defparam \data_count_int[7] .is_wysiwyg = "true";
defparam \data_count_int[7] .power_up = "low";

cycloneiii_lcell_comb \source_comb_update_2~3 (
	.dataa(\data_count_int[6]~q ),
	.datab(\data_count_int[4]~q ),
	.datac(\data_count_int[5]~q ),
	.datad(\data_count_int[7]~q ),
	.cin(gnd),
	.combout(\source_comb_update_2~3_combout ),
	.cout());
defparam \source_comb_update_2~3 .lut_mask = 16'h7FFF;
defparam \source_comb_update_2~3 .sum_lutc_input = "datac";

dffeas \data_count_int1[7] (
	.clk(clk),
	.d(data_count[7]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_count_int1[7]~q ),
	.prn(vcc));
defparam \data_count_int1[7] .is_wysiwyg = "true";
defparam \data_count_int1[7] .power_up = "low";

cycloneiii_lcell_comb \source_comb_update_2~4 (
	.dataa(\data_count_int1[4]~q ),
	.datab(\data_count_int1[5]~q ),
	.datac(\data_count_int1[7]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\source_comb_update_2~4_combout ),
	.cout());
defparam \source_comb_update_2~4 .lut_mask = 16'h7F7F;
defparam \source_comb_update_2~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \source_comb_update_2~5 (
	.dataa(\data_count_int1[6]~q ),
	.datab(\data_select~0_combout ),
	.datac(\source_comb_update_2~3_combout ),
	.datad(\source_comb_update_2~4_combout ),
	.cin(gnd),
	.combout(\source_comb_update_2~5_combout ),
	.cout());
defparam \source_comb_update_2~5 .lut_mask = 16'hF7D5;
defparam \source_comb_update_2~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \source_comb_update_2~6 (
	.dataa(\valid_ctrl_int_selected~0_combout ),
	.datab(\source_comb_update_2~2_combout ),
	.datac(\source_comb_update_2~5_combout ),
	.datad(\data_count_int_selected[8]~0_combout ),
	.cin(gnd),
	.combout(\source_comb_update_2~6_combout ),
	.cout());
defparam \source_comb_update_2~6 .lut_mask = 16'hFEFF;
defparam \source_comb_update_2~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector0~1 (
	.dataa(\source_state.st_err~q ),
	.datab(\Selector0~0_combout ),
	.datac(\source_comb_update_2~6_combout ),
	.datad(\packet_error0~combout ),
	.cin(gnd),
	.combout(\Selector0~1_combout ),
	.cout());
defparam \Selector0~1 .lut_mask = 16'hFFF7;
defparam \Selector0~1 .sum_lutc_input = "datac";

dffeas \source_state.start (
	.clk(clk),
	.d(\Selector0~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\source_state.start~q ),
	.prn(vcc));
defparam \source_state.start .is_wysiwyg = "true";
defparam \source_state.start .power_up = "low";

cycloneiii_lcell_comb \Selector0~0 (
	.dataa(at_source_valid_s1),
	.datab(source_ready),
	.datac(\source_state.end1~q ),
	.datad(\source_state.start~q ),
	.cin(gnd),
	.combout(\Selector0~0_combout ),
	.cout());
defparam \Selector0~0 .lut_mask = 16'hFEFF;
defparam \Selector0~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector1~3 (
	.dataa(\source_comb_update_2~6_combout ),
	.datab(\Selector0~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector1~3_combout ),
	.cout());
defparam \Selector1~3 .lut_mask = 16'hEEEE;
defparam \Selector1~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector1~4 (
	.dataa(\packet_error0~combout ),
	.datab(\Selector1~1_combout ),
	.datac(\Selector1~2_combout ),
	.datad(\Selector1~3_combout ),
	.cin(gnd),
	.combout(\Selector1~4_combout ),
	.cout());
defparam \Selector1~4 .lut_mask = 16'hFFD8;
defparam \Selector1~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector5~0 (
	.dataa(\packet_error0~combout ),
	.datab(\source_state.end1~q ),
	.datac(\source_state.start~q ),
	.datad(\Selector1~5_combout ),
	.cin(gnd),
	.combout(\Selector5~0_combout ),
	.cout());
defparam \Selector5~0 .lut_mask = 16'hEFFF;
defparam \Selector5~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector5~1 (
	.dataa(\Selector5~0_combout ),
	.datab(\source_state.sop~q ),
	.datac(\source_state.run1~q ),
	.datad(\Selector2~7_combout ),
	.cin(gnd),
	.combout(\Selector5~1_combout ),
	.cout());
defparam \Selector5~1 .lut_mask = 16'hFEFF;
defparam \Selector5~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \at_source_valid_int~0 (
	.dataa(source_packet_error_0),
	.datab(source_packet_error_1),
	.datac(source_ready),
	.datad(gnd),
	.cin(gnd),
	.combout(\at_source_valid_int~0_combout ),
	.cout());
defparam \at_source_valid_int~0 .lut_mask = 16'h7F7F;
defparam \at_source_valid_int~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \at_source_valid_int~1 (
	.dataa(\valid_ctrl_int_selected~0_combout ),
	.datab(\packet_error0~combout ),
	.datac(at_source_valid_s1),
	.datad(\at_source_valid_int~0_combout ),
	.cin(gnd),
	.combout(\at_source_valid_int~1_combout ),
	.cout());
defparam \at_source_valid_int~1 .lut_mask = 16'hFFFB;
defparam \at_source_valid_int~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \at_source_valid_int~2 (
	.dataa(at_source_valid_s1),
	.datab(\Selector3~2_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\at_source_valid_int~2_combout ),
	.cout());
defparam \at_source_valid_int~2 .lut_mask = 16'hEEEE;
defparam \at_source_valid_int~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \at_source_valid_int~3 (
	.dataa(\Selector1~4_combout ),
	.datab(\Selector2~6_combout ),
	.datac(\at_source_valid_int~1_combout ),
	.datad(\at_source_valid_int~2_combout ),
	.cin(gnd),
	.combout(\at_source_valid_int~3_combout ),
	.cout());
defparam \at_source_valid_int~3 .lut_mask = 16'hFFFE;
defparam \at_source_valid_int~3 .sum_lutc_input = "datac";

dffeas \data_int1[0] (
	.clk(clk),
	.d(data[0]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[0]~q ),
	.prn(vcc));
defparam \data_int1[0] .is_wysiwyg = "true";
defparam \data_int1[0] .power_up = "low";

dffeas \data_int[0] (
	.clk(clk),
	.d(data[0]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[0]~q ),
	.prn(vcc));
defparam \data_int[0] .is_wysiwyg = "true";
defparam \data_int[0] .power_up = "low";

cycloneiii_lcell_comb \data_int_selected[0]~0 (
	.dataa(\data_int1[0]~q ),
	.datab(\data_int[0]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[0]~0_combout ),
	.cout());
defparam \data_int_selected[0]~0 .lut_mask = 16'hAACC;
defparam \data_int_selected[0]~0 .sum_lutc_input = "datac";

dffeas \data_int1[1] (
	.clk(clk),
	.d(data[1]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[1]~q ),
	.prn(vcc));
defparam \data_int1[1] .is_wysiwyg = "true";
defparam \data_int1[1] .power_up = "low";

dffeas \data_int[1] (
	.clk(clk),
	.d(data[1]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[1]~q ),
	.prn(vcc));
defparam \data_int[1] .is_wysiwyg = "true";
defparam \data_int[1] .power_up = "low";

cycloneiii_lcell_comb \data_int_selected[1]~1 (
	.dataa(\data_int1[1]~q ),
	.datab(\data_int[1]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[1]~1_combout ),
	.cout());
defparam \data_int_selected[1]~1 .lut_mask = 16'hAACC;
defparam \data_int_selected[1]~1 .sum_lutc_input = "datac";

dffeas \data_int1[2] (
	.clk(clk),
	.d(data[2]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[2]~q ),
	.prn(vcc));
defparam \data_int1[2] .is_wysiwyg = "true";
defparam \data_int1[2] .power_up = "low";

dffeas \data_int[2] (
	.clk(clk),
	.d(data[2]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[2]~q ),
	.prn(vcc));
defparam \data_int[2] .is_wysiwyg = "true";
defparam \data_int[2] .power_up = "low";

cycloneiii_lcell_comb \data_int_selected[2]~2 (
	.dataa(\data_int1[2]~q ),
	.datab(\data_int[2]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[2]~2_combout ),
	.cout());
defparam \data_int_selected[2]~2 .lut_mask = 16'hAACC;
defparam \data_int_selected[2]~2 .sum_lutc_input = "datac";

dffeas \data_int1[3] (
	.clk(clk),
	.d(data[3]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[3]~q ),
	.prn(vcc));
defparam \data_int1[3] .is_wysiwyg = "true";
defparam \data_int1[3] .power_up = "low";

dffeas \data_int[3] (
	.clk(clk),
	.d(data[3]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[3]~q ),
	.prn(vcc));
defparam \data_int[3] .is_wysiwyg = "true";
defparam \data_int[3] .power_up = "low";

cycloneiii_lcell_comb \data_int_selected[3]~3 (
	.dataa(\data_int1[3]~q ),
	.datab(\data_int[3]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[3]~3_combout ),
	.cout());
defparam \data_int_selected[3]~3 .lut_mask = 16'hAACC;
defparam \data_int_selected[3]~3 .sum_lutc_input = "datac";

dffeas \data_int1[4] (
	.clk(clk),
	.d(data[4]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[4]~q ),
	.prn(vcc));
defparam \data_int1[4] .is_wysiwyg = "true";
defparam \data_int1[4] .power_up = "low";

dffeas \data_int[4] (
	.clk(clk),
	.d(data[4]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[4]~q ),
	.prn(vcc));
defparam \data_int[4] .is_wysiwyg = "true";
defparam \data_int[4] .power_up = "low";

cycloneiii_lcell_comb \data_int_selected[4]~4 (
	.dataa(\data_int1[4]~q ),
	.datab(\data_int[4]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[4]~4_combout ),
	.cout());
defparam \data_int_selected[4]~4 .lut_mask = 16'hAACC;
defparam \data_int_selected[4]~4 .sum_lutc_input = "datac";

dffeas \data_int1[5] (
	.clk(clk),
	.d(data[5]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[5]~q ),
	.prn(vcc));
defparam \data_int1[5] .is_wysiwyg = "true";
defparam \data_int1[5] .power_up = "low";

dffeas \data_int[5] (
	.clk(clk),
	.d(data[5]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[5]~q ),
	.prn(vcc));
defparam \data_int[5] .is_wysiwyg = "true";
defparam \data_int[5] .power_up = "low";

cycloneiii_lcell_comb \data_int_selected[5]~5 (
	.dataa(\data_int1[5]~q ),
	.datab(\data_int[5]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[5]~5_combout ),
	.cout());
defparam \data_int_selected[5]~5 .lut_mask = 16'hAACC;
defparam \data_int_selected[5]~5 .sum_lutc_input = "datac";

dffeas \data_int1[14] (
	.clk(clk),
	.d(data[14]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[14]~q ),
	.prn(vcc));
defparam \data_int1[14] .is_wysiwyg = "true";
defparam \data_int1[14] .power_up = "low";

dffeas \data_int[14] (
	.clk(clk),
	.d(data[14]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[14]~q ),
	.prn(vcc));
defparam \data_int[14] .is_wysiwyg = "true";
defparam \data_int[14] .power_up = "low";

cycloneiii_lcell_comb \data_int_selected[14]~6 (
	.dataa(\data_int1[14]~q ),
	.datab(\data_int[14]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[14]~6_combout ),
	.cout());
defparam \data_int_selected[14]~6 .lut_mask = 16'hAACC;
defparam \data_int_selected[14]~6 .sum_lutc_input = "datac";

dffeas \data_int1[15] (
	.clk(clk),
	.d(data[15]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[15]~q ),
	.prn(vcc));
defparam \data_int1[15] .is_wysiwyg = "true";
defparam \data_int1[15] .power_up = "low";

dffeas \data_int[15] (
	.clk(clk),
	.d(data[15]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[15]~q ),
	.prn(vcc));
defparam \data_int[15] .is_wysiwyg = "true";
defparam \data_int[15] .power_up = "low";

cycloneiii_lcell_comb \data_int_selected[15]~7 (
	.dataa(\data_int1[15]~q ),
	.datab(\data_int[15]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[15]~7_combout ),
	.cout());
defparam \data_int_selected[15]~7 .lut_mask = 16'hAACC;
defparam \data_int_selected[15]~7 .sum_lutc_input = "datac";

dffeas \data_int1[16] (
	.clk(clk),
	.d(data[16]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[16]~q ),
	.prn(vcc));
defparam \data_int1[16] .is_wysiwyg = "true";
defparam \data_int1[16] .power_up = "low";

dffeas \data_int[16] (
	.clk(clk),
	.d(data[16]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[16]~q ),
	.prn(vcc));
defparam \data_int[16] .is_wysiwyg = "true";
defparam \data_int[16] .power_up = "low";

cycloneiii_lcell_comb \data_int_selected[16]~8 (
	.dataa(\data_int1[16]~q ),
	.datab(\data_int[16]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[16]~8_combout ),
	.cout());
defparam \data_int_selected[16]~8 .lut_mask = 16'hAACC;
defparam \data_int_selected[16]~8 .sum_lutc_input = "datac";

dffeas \data_int1[17] (
	.clk(clk),
	.d(data[17]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[17]~q ),
	.prn(vcc));
defparam \data_int1[17] .is_wysiwyg = "true";
defparam \data_int1[17] .power_up = "low";

dffeas \data_int[17] (
	.clk(clk),
	.d(data[17]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[17]~q ),
	.prn(vcc));
defparam \data_int[17] .is_wysiwyg = "true";
defparam \data_int[17] .power_up = "low";

cycloneiii_lcell_comb \data_int_selected[17]~9 (
	.dataa(\data_int1[17]~q ),
	.datab(\data_int[17]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[17]~9_combout ),
	.cout());
defparam \data_int_selected[17]~9 .lut_mask = 16'hAACC;
defparam \data_int_selected[17]~9 .sum_lutc_input = "datac";

dffeas \data_int1[18] (
	.clk(clk),
	.d(data[18]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[18]~q ),
	.prn(vcc));
defparam \data_int1[18] .is_wysiwyg = "true";
defparam \data_int1[18] .power_up = "low";

dffeas \data_int[18] (
	.clk(clk),
	.d(data[18]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[18]~q ),
	.prn(vcc));
defparam \data_int[18] .is_wysiwyg = "true";
defparam \data_int[18] .power_up = "low";

cycloneiii_lcell_comb \data_int_selected[18]~10 (
	.dataa(\data_int1[18]~q ),
	.datab(\data_int[18]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[18]~10_combout ),
	.cout());
defparam \data_int_selected[18]~10 .lut_mask = 16'hAACC;
defparam \data_int_selected[18]~10 .sum_lutc_input = "datac";

dffeas \data_int1[19] (
	.clk(clk),
	.d(data[19]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[19]~q ),
	.prn(vcc));
defparam \data_int1[19] .is_wysiwyg = "true";
defparam \data_int1[19] .power_up = "low";

dffeas \data_int[19] (
	.clk(clk),
	.d(data[19]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[19]~q ),
	.prn(vcc));
defparam \data_int[19] .is_wysiwyg = "true";
defparam \data_int[19] .power_up = "low";

cycloneiii_lcell_comb \data_int_selected[19]~11 (
	.dataa(\data_int1[19]~q ),
	.datab(\data_int[19]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[19]~11_combout ),
	.cout());
defparam \data_int_selected[19]~11 .lut_mask = 16'hAACC;
defparam \data_int_selected[19]~11 .sum_lutc_input = "datac";

dffeas \data_int1[20] (
	.clk(clk),
	.d(data[20]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[20]~q ),
	.prn(vcc));
defparam \data_int1[20] .is_wysiwyg = "true";
defparam \data_int1[20] .power_up = "low";

dffeas \data_int[20] (
	.clk(clk),
	.d(data[20]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[20]~q ),
	.prn(vcc));
defparam \data_int[20] .is_wysiwyg = "true";
defparam \data_int[20] .power_up = "low";

cycloneiii_lcell_comb \data_int_selected[20]~12 (
	.dataa(\data_int1[20]~q ),
	.datab(\data_int[20]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[20]~12_combout ),
	.cout());
defparam \data_int_selected[20]~12 .lut_mask = 16'hAACC;
defparam \data_int_selected[20]~12 .sum_lutc_input = "datac";

dffeas \data_int1[21] (
	.clk(clk),
	.d(data[21]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[21]~q ),
	.prn(vcc));
defparam \data_int1[21] .is_wysiwyg = "true";
defparam \data_int1[21] .power_up = "low";

dffeas \data_int[21] (
	.clk(clk),
	.d(data[21]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[21]~q ),
	.prn(vcc));
defparam \data_int[21] .is_wysiwyg = "true";
defparam \data_int[21] .power_up = "low";

cycloneiii_lcell_comb \data_int_selected[21]~13 (
	.dataa(\data_int1[21]~q ),
	.datab(\data_int[21]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[21]~13_combout ),
	.cout());
defparam \data_int_selected[21]~13 .lut_mask = 16'hAACC;
defparam \data_int_selected[21]~13 .sum_lutc_input = "datac";

dffeas \data_int1[6] (
	.clk(clk),
	.d(data[6]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[6]~q ),
	.prn(vcc));
defparam \data_int1[6] .is_wysiwyg = "true";
defparam \data_int1[6] .power_up = "low";

dffeas \data_int[6] (
	.clk(clk),
	.d(data[6]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[6]~q ),
	.prn(vcc));
defparam \data_int[6] .is_wysiwyg = "true";
defparam \data_int[6] .power_up = "low";

cycloneiii_lcell_comb \data_int_selected[6]~14 (
	.dataa(\data_int1[6]~q ),
	.datab(\data_int[6]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[6]~14_combout ),
	.cout());
defparam \data_int_selected[6]~14 .lut_mask = 16'hAACC;
defparam \data_int_selected[6]~14 .sum_lutc_input = "datac";

dffeas \data_int1[7] (
	.clk(clk),
	.d(data[7]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[7]~q ),
	.prn(vcc));
defparam \data_int1[7] .is_wysiwyg = "true";
defparam \data_int1[7] .power_up = "low";

dffeas \data_int[7] (
	.clk(clk),
	.d(data[7]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[7]~q ),
	.prn(vcc));
defparam \data_int[7] .is_wysiwyg = "true";
defparam \data_int[7] .power_up = "low";

cycloneiii_lcell_comb \data_int_selected[7]~15 (
	.dataa(\data_int1[7]~q ),
	.datab(\data_int[7]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[7]~15_combout ),
	.cout());
defparam \data_int_selected[7]~15 .lut_mask = 16'hAACC;
defparam \data_int_selected[7]~15 .sum_lutc_input = "datac";

dffeas \data_int1[8] (
	.clk(clk),
	.d(data[8]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[8]~q ),
	.prn(vcc));
defparam \data_int1[8] .is_wysiwyg = "true";
defparam \data_int1[8] .power_up = "low";

dffeas \data_int[8] (
	.clk(clk),
	.d(data[8]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[8]~q ),
	.prn(vcc));
defparam \data_int[8] .is_wysiwyg = "true";
defparam \data_int[8] .power_up = "low";

cycloneiii_lcell_comb \data_int_selected[8]~16 (
	.dataa(\data_int1[8]~q ),
	.datab(\data_int[8]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[8]~16_combout ),
	.cout());
defparam \data_int_selected[8]~16 .lut_mask = 16'hAACC;
defparam \data_int_selected[8]~16 .sum_lutc_input = "datac";

dffeas \data_int1[9] (
	.clk(clk),
	.d(data[9]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[9]~q ),
	.prn(vcc));
defparam \data_int1[9] .is_wysiwyg = "true";
defparam \data_int1[9] .power_up = "low";

dffeas \data_int[9] (
	.clk(clk),
	.d(data[9]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[9]~q ),
	.prn(vcc));
defparam \data_int[9] .is_wysiwyg = "true";
defparam \data_int[9] .power_up = "low";

cycloneiii_lcell_comb \data_int_selected[9]~17 (
	.dataa(\data_int1[9]~q ),
	.datab(\data_int[9]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[9]~17_combout ),
	.cout());
defparam \data_int_selected[9]~17 .lut_mask = 16'hAACC;
defparam \data_int_selected[9]~17 .sum_lutc_input = "datac";

dffeas \data_int1[10] (
	.clk(clk),
	.d(data[10]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[10]~q ),
	.prn(vcc));
defparam \data_int1[10] .is_wysiwyg = "true";
defparam \data_int1[10] .power_up = "low";

dffeas \data_int[10] (
	.clk(clk),
	.d(data[10]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[10]~q ),
	.prn(vcc));
defparam \data_int[10] .is_wysiwyg = "true";
defparam \data_int[10] .power_up = "low";

cycloneiii_lcell_comb \data_int_selected[10]~18 (
	.dataa(\data_int1[10]~q ),
	.datab(\data_int[10]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[10]~18_combout ),
	.cout());
defparam \data_int_selected[10]~18 .lut_mask = 16'hAACC;
defparam \data_int_selected[10]~18 .sum_lutc_input = "datac";

dffeas \data_int1[11] (
	.clk(clk),
	.d(data[11]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[11]~q ),
	.prn(vcc));
defparam \data_int1[11] .is_wysiwyg = "true";
defparam \data_int1[11] .power_up = "low";

dffeas \data_int[11] (
	.clk(clk),
	.d(data[11]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[11]~q ),
	.prn(vcc));
defparam \data_int[11] .is_wysiwyg = "true";
defparam \data_int[11] .power_up = "low";

cycloneiii_lcell_comb \data_int_selected[11]~19 (
	.dataa(\data_int1[11]~q ),
	.datab(\data_int[11]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[11]~19_combout ),
	.cout());
defparam \data_int_selected[11]~19 .lut_mask = 16'hAACC;
defparam \data_int_selected[11]~19 .sum_lutc_input = "datac";

dffeas \data_int1[12] (
	.clk(clk),
	.d(data[12]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[12]~q ),
	.prn(vcc));
defparam \data_int1[12] .is_wysiwyg = "true";
defparam \data_int1[12] .power_up = "low";

dffeas \data_int[12] (
	.clk(clk),
	.d(data[12]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[12]~q ),
	.prn(vcc));
defparam \data_int[12] .is_wysiwyg = "true";
defparam \data_int[12] .power_up = "low";

cycloneiii_lcell_comb \data_int_selected[12]~20 (
	.dataa(\data_int1[12]~q ),
	.datab(\data_int[12]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[12]~20_combout ),
	.cout());
defparam \data_int_selected[12]~20 .lut_mask = 16'hAACC;
defparam \data_int_selected[12]~20 .sum_lutc_input = "datac";

dffeas \data_int1[13] (
	.clk(clk),
	.d(data[13]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[13]~q ),
	.prn(vcc));
defparam \data_int1[13] .is_wysiwyg = "true";
defparam \data_int1[13] .power_up = "low";

dffeas \data_int[13] (
	.clk(clk),
	.d(data[13]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[13]~q ),
	.prn(vcc));
defparam \data_int[13] .is_wysiwyg = "true";
defparam \data_int[13] .power_up = "low";

cycloneiii_lcell_comb \data_int_selected[13]~21 (
	.dataa(\data_int1[13]~q ),
	.datab(\data_int[13]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[13]~21_combout ),
	.cout());
defparam \data_int_selected[13]~21 .lut_mask = 16'hAACC;
defparam \data_int_selected[13]~21 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \valid_ctrl_inter~0 (
	.dataa(valid_ctrl_int2),
	.datab(\data_select~0_combout ),
	.datac(\Mux1~0_combout ),
	.datad(\packet_error0~combout ),
	.cin(gnd),
	.combout(\valid_ctrl_inter~0_combout ),
	.cout());
defparam \valid_ctrl_inter~0 .lut_mask = 16'hEFFF;
defparam \valid_ctrl_inter~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \was_stalled~0 (
	.dataa(source_valid_ctrl_sop1),
	.datab(stall_reg),
	.datac(gnd),
	.datad(source_stall_int_d1),
	.cin(gnd),
	.combout(\was_stalled~0_combout ),
	.cout());
defparam \was_stalled~0 .lut_mask = 16'hEEFF;
defparam \was_stalled~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \was_stalled~1 (
	.dataa(\was_stalled~q ),
	.datab(\Mux2~4_combout ),
	.datac(\Mux3~1_combout ),
	.datad(\was_stalled~0_combout ),
	.cin(gnd),
	.combout(\was_stalled~1_combout ),
	.cout());
defparam \was_stalled~1 .lut_mask = 16'hFEFF;
defparam \was_stalled~1 .sum_lutc_input = "datac";

dffeas was_stalled(
	.clk(clk),
	.d(\was_stalled~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\was_stalled~q ),
	.prn(vcc));
defparam was_stalled.is_wysiwyg = "true";
defparam was_stalled.power_up = "low";

cycloneiii_lcell_comb \valid_ctrl_inter~1 (
	.dataa(\valid_ctrl_inter~0_combout ),
	.datab(\Mux2~4_combout ),
	.datac(\was_stalled~q ),
	.datad(\was_stalled~0_combout ),
	.cin(gnd),
	.combout(\valid_ctrl_inter~1_combout ),
	.cout());
defparam \valid_ctrl_inter~1 .lut_mask = 16'h8BFF;
defparam \valid_ctrl_inter~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux2~1 (
	.dataa(master_source_ena),
	.datab(gnd),
	.datac(gnd),
	.datad(\was_stalled~q ),
	.cin(gnd),
	.combout(\Mux2~1_combout ),
	.cout());
defparam \Mux2~1 .lut_mask = 16'hAAFF;
defparam \Mux2~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux0~1 (
	.dataa(gnd),
	.datab(at_source_valid_s1),
	.datac(source_ready),
	.datad(valid_ctrl_int2),
	.cin(gnd),
	.combout(\Mux0~1_combout ),
	.cout());
defparam \Mux0~1 .lut_mask = 16'h3FFF;
defparam \Mux0~1 .sum_lutc_input = "datac";

endmodule
