��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\����q�?��e�I8�b�Ǽ$��"����ׯ1�V0���m�a�I/�$Q3ztl:�6�����`Ii��E���I�v�m&b�1��7�zw"�����	"��S�G� �Bvo��S�����ް���8>쁢�=R��+t����p�fT4G�m��?��-�)u:���ʘ��Ր1��ap�'Ŧ�Q�m9U�K�#�*����]4������jNcz�NNei�*��^I/ʩ����T�I�ǫ�k`�o4�|k	����C ��`�&'e���-� g-!4�wD�H��6"c[S-6�Т H���PA���Q�ب_WaXBz?l��x�.=[%�T�+� `{F�X��!�R��ވ��e�P*�[�����߄�X=��S��+�S��X����1e�;����B���<�$������,&�u����)C[� �9A�?�h�T@�؛�Y���,9���"�Ov�4��-��|ִ�!�$A��x#2��ō��#�}�.�I�0�r�8M{���X0�TE�M��H�u�۴-4�����e-��}c���&���Μ`"m���������`�'MI
1|�tg�#M��lؾT΂S�Ӿ�*��s�����Q S�0����cm �g*[�Ҷ���G�i�^UTD�*$K��nc�DvF�b�.�;Vs@���9�U��q^��O$:�%�f����!V�YW����j����#��ȹ���X�ڃ���s7�h�\�Oi@!|9_���^q�һ5D/it��u��EJҠ�
Gm
�[7O���|�/�Ze�Â��a��NO�g�9k�gY���P9�zt���(��,FZ]ߓ�i�<� ����:\�eG{�.j���W3d�t��Rz���5@��@�l���A�^k:
Il�����MTv�D
�h���Ǿ2^g�yX
P\e�(��$�9�2(��Yw:����u'X�3�jw��. �"�c�&�s��(l8S8�)BN�9�}��i.{�3R��n~�,�i��BV�kc�h�X����Ȧ	/���$���'���)U�:X/i��pso*�?�`�l����E���Q�%�ۀ����:�>
�e���3\����idK'��vӁ���,���wE� ��5��Ү��̇��<ˑڅ��p�n�8�Ņ�������,��~�ji
u��9�!|řB=�W�~s�QO�Y�HA�k��
�S>L����c]v0c�J�8���D�C^�r�&���e��s�4M�-�3 F�n�K��gF�a��<'�^��o1�J�t���,���d�8k��'�"�zD'	8����C�-0x��"H���:��&��3oa��s�l9�bk��jr�t��;!:���>����ǎ�����Έuק�Z�]�Q=�����&���	�ՠ���*�4t�[id)���9+B=�<�V��}$E��N�����p���].���rL�����*x�qV��j���D���H�¼N)��55����	�&ܤ�^�e".�j<�~�+҇��8OS�~>;$09����Bp�w�TFz�F���Fwb Q���(��_�2�}l7��o�T(a5�e��̖�g�x��s�Zq�5��qcږ
�6�3����ݔ8�����������i���0�G��������W;H5⅁�����1}�Lp�p{�*Yz#n;]?��2�V"�m��:��Pu��Զ��%��*��wg�?Z�� �ș�O���m�����du��~��� ���w��f��J�Q���K�^O�H���W��0�g�fO���uWi�v��O��Vja<m.�2��?9��W�ɟ�0#ގ�d%rA��@g� ��`�� �A�쒼�t��i��ܸA�7=3��>M��%1��w�܋%�S`���۩���7���(s6i\������j����ST��}�j��{�Ep <a��^���s� ��Jz�T�&���_���U����~������G�j��}�p:ѳl���^�(Z�ZIOh�:s�f;o������m�����DKb-p�Yv���զ�I��ي����w����xG`Err�n\b⺑���Q��h���Et��I�o���{m���H���w��̪�%KX}�A����I+��;w#ʯ��o�����O�a�Ք��6�A[��8{�Oz��zx��j�H�}��1kAn��V��I�&5�#�}�nW5.����p#!��D� ��̌��qv���jO�v�n�eL��� oL+\�VUfݑ	�;��"��D_'p-m�tg}�EDoP��%�5�燳��	�ש�8���L�C܋��n��I�?(}��]xp*����=3��*�7�Ո���K�Z�俌�rPЈ�����(TD�M���,��>ޅE &X��.9w&�2��җ6�p]_����r�0�z��=2�u�PK��SE��1�Ĵ�hrJҙ��^z��7�)��e�9� N	�K_!(E�t��>�AA;>3��DT���U�'Yr^�L�S�$��@b�����#��&���t�#������·�����FȞa�>3�s8K���^�%�S��#��'j��0���`��b�3�8E�"��=#���$܏�B��zۦB�1�?�2�6D~77�d?9@n�JME�q�Om}�(�j��M�E������N5D++�z�$u��x��\�T;�cf��u�����o�$� ��=���rA��Y_�O-�&RY-�ni������M��M�L9� !�>)ͭ���]c˻�EY�j�����6�$��}49��A�pN�L��q�����؄�9����L���=s��w�]�`�3�&�hI��Q�6)K2(���ٕ�W�^���)mv���1�t�t��%`&!>�S	O��QllH�u9��j<0�|�IF>��:5��Vů7u�͎W�P��/�i�ҳ"m�r��2���B�ZǢ��J��i@�8)~�UUz��R�V4ҝbt@X܁.*}��5��|Q �������s���^Z�=�����d�~��F� #&+���S��g��4�9�\��=��i�(�~�%@����᪬<�Gd��C ��Tju� ��{�X,�P%���94'ޛ�䁵x��k�]0�<UX�w�[���X�IN��/���<����{��o���<fE��۸�k�$�$��BKJ��с��[����[@�e[��{�4�"��;��¦��v�4�1aQ��Imx�;���h��r8�W�4�ӂ֫��y�s3M����Id{��ZM�q'[g_��M���Ŗ���-T���{hZ��rC�s�h������Z�g���'�@�~����1�.,ϔ�j_�L���I��-�����xf�^��.hRD�#iŊ02aĭ��o��-XUa� }�&�9m�-��#YK7%w2$��K:�0�Tr�j��� �s��՛��]*>��/ULNֵ�jj��7��{U�Cֽ��;�T�5�O���\��-��TΩҪK|AYP7�*$�/��]�������n߲{�i̽G \XP�[JI�j�7E[�>w��&F�}���UWC��[���FX��f�j ���`b�ُa����R�"�]c��e��t'�.@�f'ZV�h)ñ5����xM���+~M�Sm�b�1��.��e���ɖ�K.�2���Ew9�Q5��a����2�֬��J��m+��P&T@gKΓψG�Wi:>T���$�W����|4�.���H�;��>2eS@T��n�C	ʹ�P�����0��lu��Jo�b��0	t�iC^pZ��k���k3�@�� �z	N[!Ω��ݱ���=�Ӆm�~�|o�?z^�Q#c���
fYC��ui�"6M�7�w@��-`����TCn̌����%�i��as��
������~�,��L(4=(;t����l�<�^H�]bDiB 
���Sp� �c��]9��t�S�.��2	��⯣`��t}����V������<���:]�
��F��>��Il���#;F�D5�J�X�k�bӝ���E��R�g�;Uǂ�$�@�н�o�I���xj�o� ���#.�it�ǲ;��*�2_B%�M̫�&��(��N���]r��f��8�6�t֏�;F¼R�ѥsQ�	@�|Ҋ��ޠg�H��+��"7���!�|H�{-�"���iQ71�T���|d�J���<�1��
��n&�H���G�oqr�]�4�c{B��%K�3�	3�}��Q�0M:��	�Iѕ@�5����x�t&���jV��,�)5v$DcV8M���U�j��%� C\�Zj�q5�(�M�9- K4ẕ���TY���Ʌཕ�� �n$,�P�@&�A����]1�ݯ�����-���0j�Q��'�M�t�]��<�ؘ����nPX��}e���G��X�^;N��0�e�y8�Uw_���Ƕ�c�%ym^���杊�ڐh��\Է���2�y@[�c��;|��މ��?.���g���d��}������b8rG��'�_�r�BD���}�b�T�p�q$�N*�;���5h��Sa�[81�¿����3�$|3�X���mFA��4.�����ƻ�ʯ�3�l"���@���T����^|��s�����Ja��BK+t���S�uf�p��8��U	��ݧ����B��p`��9�H�3�Th��}���3rV!2��r��3�]'1��X�/�Z'f���ơ`A���bÉe��+��L�cT�� 聵_����l�a�����|}ͪ&Օm�[��{(?ׯ(jJ�Y)�JPx�����'����r`��tP��Cf$�E2��ϫ�����u!������4�}�#!������f�y��pU�=�Up2s�ڥ������@Dd��� N$ŝ���P�d����bo`��7����������7�ѧ}���*_!`��L�G�Z��l#o�+=,p��`�V��АL�O���,/R�'�~�T���>�N=q���/��b���(q��������!Z�S�6��I���al7!8��P�p�E�l�� �Aț,���g�����	K��bB�w�`��<&��S��;�"]�\����䈲�
nI���p�Ҍ?
TI'ٮ�/�p�)j�G29g>��1�b>b��q�8c p)�e��W✀��78mW-(C�֡��5�4�`�>� ��H�/^�%bNl�\05�M�M�Q���Hg׬�:c}U\oF5�qE��,7�nQ��ͺ�]ꅂD��7��9gR�ymB��SW��[�����)��`���n��=��˂6~���A��n!)7��Nn9����>f�I�\��t�]���=�G�(�����Խ&���o1{d�e����G�5`P�6��F��#��`������f �%���c{@_a�S�������� ���̖���+�b�Q�0v4���aM* �~%��ӯ~b`��)���'L��_Ǆ7��3�7�Wz����H�{��FP��aZ�{�-��e(�OϙP[��
wtD�a-GZ8�!��:[H����g�D_�߉q�9�A�x�%�6_��F�1���每��7;*G�n��s�r0� �3K�����k-kءi؅ bV���9��y�d�0O��d���4�`�_��Ľ�/
���"�.
飯)K�\@�[=�Seʇ��YK��X��Ұ(�
�<
�����i7�e;���u>�K��Z���	t�ns�¤���[�ꈥ�道6-�Kո�=6�.�>{�������C
�+���[��)&����ĝ�x�#�wM��z��I�9I��.��,�M"-4x��]��4��qW/-��A\,j�K��K���M�i|pO�œ�] ��$�|7\+�%�=����o��+h���]S>� r�os�=��]^wu�$�Ռjr���Q�oU>hzO(WÎ\#|ޔ�
iM�@�N �bW�EUv��g�����'���ѡ������Vk��T]%F�ɨ�(���j,���*^*�߀�����b�K��$h0z=����VF��\:��F�|�Y댡n$n��A�3������ {��ۦTp)� ��R6;=ւ����̡��t*K�}�r縄���'zdG}#��7՘ϊt�Ko�Ы1D�	M����p��Ob��Ϊ���d��k��9G��,5s��}K+���b.6czk��g5VYr��*��[�W�*�
DcSK�j��>�x_�:�ш�]�����LJܾx��z�)w0��N�~\֏ ��<�껪�,oCz�5�1����wߊ�$��E_��Kk1i8)��Kϔ�����W6ف{`�k�.�O�9;ds�!�`7��7(8���^3=�J��R���	��SͿ@���%K|����ѳ�٭ҽ�!�9��]�X8�	��:����ޙ�r�q(�YՕq��w��*���-������l���� ����]��/��y��#����4�����^�@𼃂�����M��f{��[�@Ek��hH�Wq�5Mr���~��*���ў���s��H	�;�Fʧ���G`��M&M�`B;��ͮ�t��
u��y?M}�JR�U��%lW��Id�qs��,��Plˏ�	���J�aˢIL_׃6&��nF���Y�Z�e��.�c%P!��)	�����l�,���$����"
W�*6����ij6���Ԕ�gJ�5��!}�Ҋe ����&��zPxJh�m�r�	���!��{p��-A�2T��)q�V���:�>B܁Y�yt�*I�p}%Ϧ~��˭t��S��+
�d�H���՛��p�����C�5
�
�	+��H�Y�'�찷�`�O%�+��W4T���a�<�� #V�!?k���0��	Kw��c��7�U�+.R`I����[=_�ɘlM���-��xM�}��hЪ�͉�`p8������:�,	X���(�Q�Nt��_�I���!4�����J�dnP��Lh[ϣz�q�QO[�[Z�p��@�쒗�E�m�=k������b6�aU/�;z���"�y�3]������Θ���8i�:�2�=�f���p%�j(`�R��h�H�E�>�y���iW)K>��Wd��E�5?���-L H]NB�^��Y@,� }�Ǭ|��.!��� �zI���y�<�#�
`���y����#���,Xď.�1���]��>yzd�l[��
��'��Qu
PHv��h��'���)[VTN�(�[3[���:)�X�n���o,���!?�i�Y��+�H��8�g�����D����B�7`^�w�� ���O)�Xp����Pw� �bj���͠>J��a��0`�C�%-���
�j~ו<bY�����B�Kueє>d+Y�H5�y^�؝� }��e�M�I��B��b&���Y�|G�1�b$½gc��=�ä�m:�'��H�x@H�*���N:�ܝB��c��4�n�/rޤ��"�5�3���@���cY�����O���#ϡ�3�� ƙ��c"�@��O�����-�E(�������وo����M]M�L>7��Ye���a���E�(��t ĜJ>�M#F�5]��w� }p����0w��a�	��J3����Ɉ��{PH@,�܁�1
�G��e�*9<��6�ƿ�u�2�u=tsqI��� G9��]��0�z�sR�w��+ax����h, ]]��b9+����?4t�X��1_��}%] ��(���P�����@��NY��6��F�5�]����	���7I�"��b�|��u�#��� !���{lE�b�.A�x�*�kǘ��5@'�a̜��ΈA���2�1�6��	�ÊFpvH�UP��Ͳ=�o�Z��z��N�֮����rW�d��Lx C
�f �:?�?�?.(v��˸�����(��T�)�������͊��L��iuG")Q%i�o�91k�c]�TP:��O9^<�*��sԺ���j6��sՍ򋾁����~h�Y�_%P�װh���`Xd�k����⊲.�Xǅ8o/"�f�����*�=}O��z�"K�z!Xn�ܮ��2cO��Ͼ4=�*�}'�F"9��	�!��8� ��owRH��8�:� �u��Y�
X2��+��D/
�8�fq{���Xz*({�m�{���1��8��=t�^(����sg�0a�B��S�F�f-|����ׁw��=2��:|O�Up��w�5@�F"�c�F��� ɾ�_=�K����y��)�1�NpV�M;���r�[ˋ����G���n����@��~�'���63�gW�l�eq���9*�T�!�� A���h��$z�m	?�`^�]�<iS�V��>C�ݙ, 59@!5���d,��ÅW����ɧ�w��W脮��H���,<��!���u^z[�Xj�㺢ߣ[�!D���E�Ϟ	@\=�.�J��������v+�@�o�ϩ�B��u�M,I��q�Jx��_A�x����:lP��-0ݯ�\�w��$�O`���~�=���"`�ӌAQ8���q�u|�� @9������֏���Rn�}6=H�l�8��yXaլu�=�Mn�:�mJ�l]�$\g�H(�+����cݾKLRp�}�H[��F�O>;��m����Y��_l����P2ڗ��ҥ��樌p]��ڿGR5��|�O_`~���Ϗ	Ī�<��"��$��Y�����t�"�����)[��ND��o;�)h`�z���v�I�k���c���a�:�W�	�l�[��I�y��0����r��j�7��q�h<�b3��љN�٭ZE��u�+���J��r�c����fg��l���"���ƍ���K_��tU����[�����@ĵ��zγ����p���*+&	���Wtp���g��o�:�q���N|�d�����(��/7u�YW}$��@��V�p��k��Y���(CM�<:�w�̄k��ayx����IP��Şj�F����7�؏���~z!q��U�����3����
����8�gL��Xb�r��,�t�k��G��D�w�>BW��r�酄��<\߄*\��-��=A{�����^5y�����Ç�f�4_��xى���ƫϰkFV��?� &�Y�Y����<�
�Zک��*�ͫ���Cz�}��;¤����5t�x8�4q��Y�U	��O�X�C���;��)C6u-�IB�j|oN���]��Bl4e��Q��:N`�OT:k7�xnX��-��6��pK�k��&O����+#'�K��9�s���΃��?a֑ܝ�����w5�B�u)#x+�Z����C�DDj���-''�#�l��.hS�@v`��O�'�M���ٶ�	�s�x�6��C�rC	��&/v�A�����_�ɏ�eB�0n���k�4�H��Վ�h��	p�$�zM#�GO��S����~)A���mt���m��aD6�<R� �r�Şb�0{Zx����9�\S��@�WN�6_)_m�\_�pv�͞�݅(a�U��\?���/�,�9ڿ�8A�@<�rM�V�ݨ�n�#v�a���tFP#��O�0W�K��J��`�xPV��l������m��� ���ė�^�D��5޽o-F�?��уv�`�)�S�Bq�r���!�-A��G�#�f���Z�Dr� �@��^H��F2��A�"��P�1/>tʧLY_6����eVȽ��ߢ�v����k�C`YY� E�H���ޅw�g��R�g�@iT�l�urPq��!��_x�YF(qc��]�sUE�Iߨ��s�G�x�o_\xK;JʝZ�!toO���.e}�^Oa������|�T�A*aT҈����H0��A�
�hj'z����C*�J���rʝ��︦���(�ĻZC�J5kT�t�V���JMϋ�x�y��n�����u�!�sPu����ꯢ"ߴ�H��H`�J~��MC#vX�0~t^��^C��/�����>�x ������!����X�g�	1�P`�&�1�]}�4Z��:���mJ�ݰk=Թ��T]�� J� /�y��?������+�=����0�n��_���v(���<�����{Dȹ����/�$G�>��Y8���
I�`7�{ixҳ��q���������t�D�&p?��?�|�:��Fe&��`�0ոzA>-]�@�_�m);�L�<�#Gh��\!ɣD��E�����G��I�F^��7Ouy��?h_/�����WFCՌ_���y�� �n,�Gt;�}(�R�Ȩ���kn��s
m2�Z��\~!�����f���qG%�sw�e��6�C%�ǿ%D%r�L���d�v�+��Ez�����ҥ�ӔF����k1
4V�J��]�V�)�C����@�a ��z�lX�}�a��G븏����PMę��+����0��Lj;W|+Oo�v�Qp���Q ܿѝJ#Ӷ�t��-A�*W\�����O7�߻���%	;��p�) {�*m1�+{�����UZm`�p>��8mX�?Ȕ/x�\h�>�(��V�ĶdXu��Sz����.mIV��p��Vs&�E{'T�u�0����^1�&���y찂j��A3��*�FNU��Œ�!)����*H����)�J1��ʁ�;��sb�\�)<��[ +d�$E����խ�����l1/;�h����)���<U�`��a惝9e�q험G(�fu��@B*���J�$����A^�A�,�	6�S��C�%aëR�j:��b�G�, @�"UWׯ�bhYI�l�ACvƑ�>㼷�!�T^�)����ťt)��h��8�����wOU�z�G����J�u���Z3�gi<E�o}�!�M���O�7k:�?>U�؉Y}�[+��(��K,���]D�CZ�{]����&]<MY-��?�Ά�`�0�\��;*&�<Q�x��&�-D�zt'У�s%���i-F6���AaY(�K�Q��
$>'\Y2��!s!������؅0����?��N�v0L�u瀣��5���a_��d��W������ ���&��ڞ�B�;,���>�w���p���h 0Tu�<\S��e=d�b���O���a�
#��7O��o9�o�HPyg����p\�O�z���a|��0p������I��]jC���~nH	�s��
�bK'�|��vAh<b�vӲ��T���ˍ��1`�+_��ʒ���7/��޵���؈��<8�r��ٸ[������������Q
�$0d�E���&jXhrtv���
ẫ���w�H����6���%�5z2PWA"h����}�~f%AQɑ]�eI�~���y�*A!2��.|��SA� ݬ��!7��n�S�R{�-���gą ��R��d����	���W(9�+�v���)�3�7�N���@z�
u��ۂާv�$�>�<��8�U�$�����,6��<8'�e5�R�=�x�^����ꝕ��4j-Ԡv8��_�8F���[��k�~;��k�\O�]�R\�%V�X�T�釞�-RHÂ9��f�j���5���$=�_R7м^���Vzޑ$U�̺h�C����>���e�t�-sHZ1}���g�7�b���4P\�%O;�3��/�|n�:+�P�i�i��à)A�2�q�wEG�:֐;0����=�3G��`P)����ie�C�~�i*~�P0�J���DLɁa�MF�?�_;�\�>����z�L�GP��_=�eu�M!���LQ��H� �����W��0�JKy4�p+�X�(��x�nD��5��[""��L�ٿm��0���9����P��Qꢡ��O��9�F�W�w3�����qwG5Z�saȺ�����i]����˳\I\��awMOz���Xg	7?��N���>�白���$s������h;�O�ݖg�� �����z?�a�8)GǑ��.!�
(�N>�U'ߌ���S���B��X�]飋m+��h~ɤ5L�+�P&��OZh7e~�Kq�Oy!�p�������\����g���ъB��n��8��z�����7N�㾔4 �I�W���}{S��������]9&O*��J��
�$�tq�i�-�V��crS�*�;�����%��+���Q�\G�0zP8h��)N[�����0{�@j��wZu���킡,EX���>��_��B��ft�AT��mҕ�N�5�.�$�)T�)���]�ɒx�/�"��\C��i{�/9Qvm���h�j�_��I8�Н���J��nr��x�K7~��Ɔ���=�`t_A�lCE��>ރ��2V5�����}�p�:���+��R��X��`Ӗw�:�)\%�a����pz�6.���Ļ�'�y�O�����I�O��Rq�`�/���[\�1��+}.��OZ�Z��F�=��y����|a�.X%�,����ԍ��ō]�ʅxH;s��~�Ux���-�i�~����u�(�
���Y�FZf����`���p�D F������j)�0��ci�6ڤ*'��}���)7MH(�W����YF�T�{�R�џ��T�䧕��r�W�r�}�o9��%�G++��_<a�٥�.

y�����`��Ԧ�*k���9�|���WIS.d�S�I^��_�����u퐿��E����:E����f	�A�2u��lPg�M��t�v�dy�?N�A	�޳�<��@!�����B>��
���U���	�IcA�M�]=���i�Ҥ^@-��_\���"K��6-4�Ɔ���C��.�G��WB�8o�8�4�]��+�>�d-�Z�N�)����·�4�-���{ˁ��<|Rp^�}���0<��i�`R�5as��I��>&���?�����De%��&QLWw�7�a/���{Y�ئ1E��lm��*���˻3W�f�.s������Ү�/�U����������.�a" q�9zI�+��?
�®X5�w�jj�^�je%�݉u�E�G}���cǺ)���	 h�G���B��7��3�b�U�GwԸ�
%�x��{or��s��a�F�&Ǿa*g���yq��j���	����%W��N	������VV���9�`f�,\PR`�/��^ 䯃t9�F�D�M��������YP���D�cHx�$.��1��ѩzu��Y��y�K���#)c�[!��Hf�z���%;���a���ȫ�x��k���e�]/��:� L���x��?��?��	>s�F[��]j3�D���'c�I��6��l��i�2��8���$�ь�?|iL��4�'���#��-�ګ��$�XU������^��Y��[v>	���@���wKE,� G�{+�h���`�=�C*�pe3��0�@~�J�� �A������NA(b)4 ky��ֳ�6A� ��G���꒝��������`X���18o�N����,��2� �=1��ױ������=�H��ĸ�|�}�{�|:!y�	�^�6�1�
 u���Y�T���E08��s�^�D�,�mx�e��6�y&�$�����q,��[(����sw�n�8��ϔ�'D�_��ur��� � �8�XuM��c��5{����!Q;��50�u��xV�,X�ED˼�ۍa�4���b4�q�%�]��B�%ѳd������#�{���������IٓL�`��pwf��4��'�Zg�ғ+�r|(��&�Q�yv a��h�m1N��)l6t�95%���L%�y�nꗌ���'#�t���R�����i�9b�k��a3%�6�[��\�HN�ݏ�5�S3����-.Xv�Ů�?��GCy�e�[�a��_��y$���
����u8���GL9��?:���#}X�J�}����񯙢�?��
UK!�[Pp�w><9}g����5/@W���]���3��;�5Z��'����ά��]�w¾?��:Qs�.h��1#���jf���G�Y�	���Ӳ3��1�9O_B�B�5z�i��F�#Ƽ�C��a=���*� H���yΪ�zb�Y�iD���=���:+�@���c�i�)2ń�]W�p� �gKlG�L���)=�j�`�4l�D/��6��c��G��U���
Jb܎���Dz���_H����8�����'3]�y�s����3o����idY����������]��Z8��h������t{�,ė�5>��oD�}mG�SFi�]r�wWHͩ�HR��zX0f#��B5� r�a��x?1Eݓ`�N��l;��$���d���8fL����;v���b��f�6�KϠC'�|��f�Qmd��� �nxJ�<ƫ���{<�W7�RH+Z1�����1�!��}F������.�t�-��w&�	d	#���WN�������?CBc��qD���᪚/ş�� ��1K�x� ��>���y��VJD�:����T�;D*}l��Z���g�ˠ��I�8��%@Լ	�����Ie����C�D��=��B�vt!�X`�a�oc5�NPj�tP�)V�fR���} Md�N�rȔm:���H��]�A&W� :7]�9mab�i(���wV�pf_�h�ԟ���(PIX�ĉR2�B�v_�͖(/ �Ng�×��+�{i*���Jb����͗�HUӪ�k�W��!n�ϔV嚱�ı�h�����V�B\�ؕa�[Y��@���b"q��/0+~sbSL��z֝%����T��#��s{[t'����$���fNԕ��G��0вP��.�ҐA2�ء�h {<L��f\��C`���t5A�ʤ�r�����ِ�B�:���{���n˂^1G�_����)W瀎����R�����d��E�slK�u8����5�H�s8�u��Ƃ8�K���ޑ���I�'���^�/�Z[

Q ��z�������� ���n�v�Y,��^.�*���3^(-rtk��9�s�8u�����Z+f��~Cޭ �(�������j*(�����j��bb���O�$��a�Kh|�h���d�_؟˪hV�kx� ��.Q�$B�u�s�[�Ԙ��`���ƋB����!ჺ����Y��C �]<w?�=����C߹��k�HOb��ib*;�o�G
�aC�V!�2���ul�b�ʾ.���^G�lJS��"���P��i��	 �����TSH&v��,��3��fs��+�E�؛w���	T�˟&c���(xG�k��#'s�[C4|Ty����0ͷ��3y$��� �9�@Х�kcss���H�*��J#g��B��Ƙ����T����SW~	�le9�s�7�0��l���˩�!߃� ���:VC��Ĵ���r/��id���M@�j��s7we�(00�_�+�t�I�A��Zc��#�!H�Ay������>"��u2��>�>�+8�mq�8WN�����*��v ��&F�6ݸx5��a���Մ�t.NN���Y�A΃�6�g���9�q�����p�h�2��$���2�ZlE�r�Q}a�][䣍�/s�Tl�ߎs�07~>�2:N8Ȉ�LRk<v�ZמiE�[�=�gvgSy��EC|�����ky,Ѻ\(�(��A�ُ��}|>����=Z��{���n=�Z(d/h�g��J>т�-�J�V�e�m�w3�d�B�v��nB���邁n �*���!XjQ�v����էt���x~����� s�a���wjt�,��̜�֬��a������>��0���u�?#uʮ9"�Q: -yĝxy��2���9�՞6iW,�c�5H6���5�v�J��K��(f�z�C�N[ݰ�P��ń��j����Y�k�0��v���O��n����_��l�I)�O�ISNj~E~�B�!��<t8�ӭW8;L\�B7�?v� ��	��	b�(��m�V/+�$���zE8p��,͂!�"�,�>�Q�Ȳ��F�i�4����?�|]���֒��+�Gji`�]�`��l~�Q�����(<r��Ѳ�2���ߦ���R<�W6?p �jT�]���X:@L�ȶ���j
o���&�j���!���/}����)Ӵ4�d�k��MGw�!(��}�k�E�*�΂��@6��aG���WV>	�������1���#�:�ܩ��$��kx���n��y�0�=Q��M�v�q,��Kn\ոShkŪFamg��L)-;�0594e�g�C���!�%�hy�O�&�Q4g�yR����T���k�i��
E���a�ۡI�����a�o�������ِ�оD���=p-�܏c�U�!�[�e��'Ȁ�|���,�Q7�N;��i=�g8��B��:��k96a��ܥ��}�����4�����^����tG	:�����L�kN����&
�$�*�K��8��}���CYd�B=��U}/������@�s6����E|.;��U��g��֋�1����^�h��JA�U�O-q��d��.�;�6I�A�[�j#Z�)~{�N����T�;#�:Iݭ��Ew������\�q>�)��6�K�a��#���*�f�:���&S+��9����:���m��Z�D��(a@�޴��Ҿ8�VS�9�M�V����@�${�3k��]<��k�2=�W�$��d���V �TH;��}Ӊ�������tP�,���;���i����q��~F���&8����o�3 ��v@�k>�f�O6�;]G�ZhP�Ec!�4���"YÑ�ZG���Ca/s�ۯ
p�ۺ��8���`�[�L!A��D�� ��M�3@aX���rÁj�Č��И�hWjp9Y_���΂�ƥ�
F:θ2��2�U����H8����t!y[G�� QIxf\[צj�s�b!�1ue@-�c�P���Q���W�i�w�D��;�U�3�,�	?{U�./��L���.� ����6}V&�����R�S`i]��X�.^rĔ�����"[׵��T�Ja�[����Zr#�9-��%����3���$���?�J��:�ö�T�p��x/Q ���H�w�z���V�����]�e�-m�OWX&����T���
1�����-�ědqՑK�<��$c.5n\�3��N������t�aOK��4�x�I��m�c�5��3$x���}�"y�������i�l��c�4��G�K�]F�.�!�c�/��F@|��&��
5g	vMo�l��T�(g��q
2ҩ"/Y�Ǖ2��1�q�@;��^�l?���yzBig"��!�C����aH�1�n0E�.	�Y
��t��a�x�W_��ʱ6i�L����2�k����BN$�sq-��E�/dv���I[��[kR{0��ò?
2z�}�/[�x�Tx<�q�-��N�9st�*��f��ɗ�Yv����,+�qŭ�\�F�'.^L�s��]���։h�Lg~��T��Se��/bQ~����WjL&���T.�{���#_�/�6^�J���RnM������Z.pVa�^Y�	0��2���Ǡ���m%~N9߁X�������	l���-.y��;[�Z�P`����Hn#�Rx��@��/9��%�;�u��h6\��GI�r[�f��I	zkl����8�2@��OW�RN�I�CX�Ib[�D��k����7�+�U�8������}f!�Xb���RWJ�0�M�� �M�IA�H��dP���L���w�Kֿ���\&g%�{wrv�-4����`��B0bx̽@�2�F�Ad9n���(�_+B�k��a��M,�l̘=�5��N���J^ �\ 3�myEh)d��['Ө8��C����<w��6��'W���cx@CW���]i��� ϻ�v/�.@��$������xΥ$5��H��ٶ2�����!7#��ګ��B�OX�mz��~O����k�������0� �II�N��iؚ���8P����-��ϙX;�OUZ�R?����1]	?�]&6�VE��L�l(w�a�l;+�J�w�� p��1~H��-��5��[B���^^C&'��j�����/@['�\���ĮB�5�7��*��{���%�`�Y�}�Z���k���n�%A��Q>[�z�k�	I���]%���w=��� $�_ݸG�8�-Yĥ:jɚ�D���F����W�"�T�����!�"���^��~�K�Վ�·�+c�-�mgwy�$���d��6�H:���f�!,�]	��u�.�����,�,����N`;b2��5uEO>�o�V�8�.7Y݈��$�<7>��6����M�������8��߈�t5�4��!o3L!c�K�K3
�
���0(h+�|�2s�'^���H��	JlyL��A�|��[m/�7t��X�Ǩ�ᅐW���ͧɝ�]���~��6'������e E���c���=��'a�rt��X�R�,`�i�#r�O�<�M4�yR�)�㵛����tm���y�.�|�>!���p����sqZ�O;=%aS;������N��kd<������u���V#�׿��;�e�yQ^��&�*O6���w�1l�hw����`4S�
���R�5�.̈:!�;p�h���|6RZs{�IP�k|��΂Ѡ��=ُ`�2)?f)��x��� 2�L�B���M}Mt3�VD������靾���9C�x<3����4�\��zEKl"���-�Cv�).��1(����0����U�6yv�h�3�?e� [�I9]��R,���,�a#�>�b� -���{o�V�����&����	��S��:y��%���_����C�!�q��스�|%���,P���!����5��`�K�����!�a�C���9��=|�i�g)��|X^�زL{t�<���5e�(߇5��D�V�sN�V���j�L$�%�*73��X�*�l�v;c0Ȭ����.y� M��|R~�>�t|zi6�z���i�����,�g�*�� ���R�JK��FeE��<\1�+f��6���#]�\X�)������ƾn<��v��*�7~�j�7{�"
o�e]@�K��j�G0]�� ?��!����Ni�c���� �������Q����:by=�ß��2+Y
:���ܟ':&�qﮅ��R[���4���מ����^7`����@}2�BM����Ct�p��W�	�<Q�tx%�H
�4c����z���5�Q�O�:�1v�@d?�{c�>�VABq�f��w�0�Z^�ݙ��C��0j���0���^�9]�2���{qC��a�����Uѥֈ:\}߾~��'P���3��c`����G!����������Ǜi�UF��X�(&��]a��P����8���E�Y*U%�ך(�~���AM�YD����V䱽�n��k��=�C��__j��)�� �V<��4PEy����Ё��O}��E��s�t~ёP2��t�"u�C�_��^� ��M�-�Z��6Z� �ƑuC)h6�+�H�5q���6h&/�5))B�J�QV-�8�Rk���9�-_�#l/+7���18������.3��e�}�U��ޙ_��b�9�ҥ�����b�As�r�O��L��p:������@�Y4��n�$��`H��#x��A��4R�[��r�Dͦz�R Oj�^���X�͊�ެ鏛��{��醭\u����(�|AN�^��jZb��N���y>U�!^T��V�ק�ugdʃ�m��!	X�n��	S���W�\��K"uv���Z�LFW�>�j�jyeG[n%m�lƘ�~qj��&ii�����9���'�2sk���5	����UD|�VS�7:��x��Л�Y�[�sV��qVuh����7�E�dUA0T�NIZ�k�=����+D���z�����C��F�:���	�|�L�>%��$lG���x�� ��-�l&�ޢ?	}��M�##'6�r���)�(�2�6����D��zA��NȢ"�*�4Xo�X�u����:�r�8*9�o������TӃ��x��pɾ��f�A��ag*�L��@c&#Lg�4��L��`��X�5ug|`�����Zdv�u:A�,��^N���p�qW�=�����+�����E�}>�c�w��x7�a�M{��
1��|�Č�KĀ�A� Μ���0�Z>*ڱ	O/]>�KjKI�k^�R̮���[j"�r�B.�C� C���:�]�!�Ì�c��_D��q�b׿�}e�4�؃{�̕�>)�xjh��t붦2?��p��kٛ役��2�U��t�{�7��ˏ�y�oY��阩M��U��%�����8�x��3Z�i�z�Wra�I���:�m��E��X�8b2��yq��-��{�e�%mԟ��hM3M��<<pb
���7�ȡ�kN�Suxɺ=�~2��(��*ѻb�6,�>����-����s�l�2_/>V��8F�h��E��;��@ȝ���iJ�I}8UJi��U�_�ĲG�%�p�43!Z�CM��d�	�`&wz}����f���L�=B���8����`��x��7s����E�u@ꂤ�Ԓłny�i���ƅ�㍅��=��b��n��.~���~��v�<R`�O�E�틓":��A=��Z^�']PNv�<A���7�������� �cг�Z���|\^����<PQ������?���ц�4L�X+0K3Hʘ�k5�N�6r5"���|�o^<��DO���kS�2Í7��R� ���b����9�F<��sw���6a��Ǜb��`�i��FŉO�}�b�X��<ױp�7��I�s���50��]�5,���p�i���c%|����j���7�u37��M������t�-Nڙ�r\��?e
��-�}�@	����� YZ#7��c��>�]gzaM>}:���6o�r�.�ǎ7"�~��gR�J	5��d� ����t����J���]�嫱���R\1�%t���Tֲ/4����SD�NB�.�i����R���z�PƮ;u}�`���fL��vLw�4�jB�椆ܞLw� ���
3�\��F�>5����1 9��^�)�C��`
yq��d'����C����J�)�,I��gדT����j�s�"�v��yYqy� ��������~��H�r���R��3"b��/!�Vq�/^*t~�@��م��o��H4SlMZ�cг��ew�cv�)�H!t�_��-��9SHV�x�YB��^�����&~�'\�6���%����%b|�[F{|��̪�`a�(�Ry�l��d%�k�͹�%�u�]:νdѮ�ǝݩ��
XB�-QGx��C�żءT�p��؈/���bR�U����m?�'ʯ���~�_�Pm�޲��j0�qN�\����ݜ��X�#Ox��N�o�t������p��'��o7����g�i�ڧV�Π֤��mi����X�v����Iq�NH�3a�;���'2��ص#���!�����Ԕp��pM�I��S#�/\e�	����1��\��I�͜��*�A�ρy�+f�8�iw;�{��0oSp��i�,�P]�=/=��E[��t��|�0#<2�x���AF���Q��b���������Π�iI��E�'g�6��IY�x�d��Nj������{��"V;o����U%�peա�X�q,��ya�£�ݞ�:���ĤB^���	N�Z����0 a���Q�qv��O{ѩqS�6��3��`�"����2r�jN��&B�H���)��CL����kk�n#����(�YX��JR�>Z�2ڏ�"���
�;h�2}�I�;���T(N����w��d^��tv��:*�>�@���6g���$G�9_���$��{9~��u�츐
��:��k7�������7��Ǔ��at��W����t�B�7�O��.綾�	{��έ�#�x);�7oo����g��ה�(�����L:ͦ0�x'�t�C�rPӨ���� QHGq�S��)9�9Tr��P쐍i�k�P���`�S����s�#42X`��S>�tg�pz�/_�;�hK����c�?P��Ada���\v�b��!�1r2���e���$r3����tG$NE�GQ�_d�*G��E$��X��W��$��P7�J@�)|�����D����ǝ.��V��j�<�,�1`��Yۉ!�b�4A��B���K��vK���7��n���>L>�nD�7 Fj��	�o��+?���L�#n�� 1�4�۟ y)�Q��4rg�&�D���:�>(dg�c�Z-��f��\��T�l�G��m��T���`�h3��k8g�%݃��a����#�����y�K�7.A:(E?(?F�ĕn-\�Q�mt9	����~�v������x�V`��|N�p��Xƞ�/�Q�D��r�y�qVdЪ델�W����.� 'g�a����zj4&9�ٳ�1DtM��#tܩ����O��E���GS�'%�����y�&�E:!q=�}�{X�!ѩ��y^�,�] �rˋ�(�1i?&�=���=`�u�{9V{��ŝG�$�ڄ�Df� m%ˎ���^Bsʌ�RəQ*K������F���	0hF¬ܟ)���ve`��+�$l��,KE-�,mͨQ�@���j]�'>5�+��@��MeB&�/*<>���lcE�}K�|@���^�-Z�'CRJ9��qQ�l��*s�� VX6շ6�zR�!<%A�Y�gdru�OІ�����lZ�FЯ�������[O0w��Ys�����>�-��2J1�
3#��'�8��1�_� }k�}�?QIŞ~��qσ���z�tf1E]p�h_���$\4[���
�!A�����T-���Z�~}����vP���q�4~V����rϩʟl7�J��yhFj̤Cx6�^�
d��v��&�>Ev�d�5"� �� ١�=�v�f3M�I��n����S
�os��:H��Y7��ި�W�(����;#�9���d��ͥUJ�%th9��}���&RҎ\�U6����~3Z�AC�����X�70=��iչ��i��w��i�`;�D��7Ǒ� 5�z�u�[��jT9��bط"?�bTf=��c])m�b4:1L�W��^m��@o&\p�gG	�R��2��3��W���I-2 �K-M9�׌�L�������u��l�rk�H�>Ɗ���s��CwZu����Ij�G�)'�1f�[�bS/�ѝ�%���ɝ�h�m�	�{��k�x��	o������j�T��LCx9�~_��7IF����ڐ�7F�0��@s؆�9���i��p��{Wqn4�w�^�d�?�Ënf�����6�M��]����`Tk���NUI� ������2�DEGg,�cX�Nw��N��L��y%�	�L�A҃��&��>vQw\�
�<Z���K�V�,˺M�����oB�M�Pdal��0�o��� Q=@u�󖋍"/C��n���(FeS�@��q�ڒF��h�t�f�Ʌ���}|P�u���b�8O?�ఁ��%�@n�O^�Q˯D���Ƚ�A�s���n%뷗�d�<ab3f'2����#�NL7����x
�^�����t�B2z�*��p�A�ks<t���p#���"���ɪ~b��� ��O��	�\ۭ)t�!�bH������ʛ|2$��ྙ� G
����}3x�-^CFZs���ZmU�NJկ��<�1H��aC�U��\��M��&6�ˍ��eI�Bg������6`hs���b#Q[�A#�� h3>L�W����'�D2�c��~�hj$Аp=h���ISA� �n��K��4�K�k�Z���C`=L;#g4���.��2��Ά3SD2.�e^�0^dp^W�v����XRk����um�!샅`l�=��(�4���-U���DcND�nːD��$E� ۽�8���]��y����t�"0�&E�=�.���׻�	n�m1`ے�B͈�� 6A�~NX��v��AGީz~�{��ARW�C�����6`u@P?�q�f�h!�����){�����;I|�t���� Mwv�"�r�0x��Z��Y&�ag���p`o·�a�j�"]N���h�J�`n��Ox"?�z`�C�|7�*�e=���Z.��;+�B��B}>��ҫ4Bߩqf�~f!p�z�]lZ o�װ=�U5`��;�.����~��]l[�B�*z"bv�0{�֌W�Hi"تL��)J7W��qn=|�Z��lJ�@�t���)�I]=b0W��=��S}���>4J�*���7K��bl�T ��x��%kf�_��2��fN:m�n4�i S�x�
�P$���3T�m���B�^�ڟ$�+�|�t��Ӭ��0ҙ����@��Ŕ��v˸mV!.qc4��$7���������9��M�RV�m�X~���n����Iӵ.�V3hG��Ɗ��j�I���/de�Ō�y��Agb>#=����:���+���G�#�r@��d���z'W���e| )������ܐ�Qh2�:�ˡ�'6&Vد����
���"u�U_�.�]ã0�E6C��Ug�o���vo�myƆu���9V)�zz�t�u ����1c�
��^y{!Ԛ᫵�|��A����n3��2��L��.Ӗi��2�h.�ڳ����3"�G��׫��(A��AJ�ݫN�RaI'b�����7���K�n�L)GB����o���Ma �t�1�+w�W7�8|�Y��F�c�T�e��z-����7zR��S@{K��g�l?��]�ÿ)#����L�)s��ص~�b;:�҉ׁ�f�<�ʋ.��67V�c*��p��lGO ����s�*l�ᛍx�k��h�uD���NvM�3=]�C��J#���r��X�%=-�	��u�oiī(*E���k\�z-�s�;N�����x������.Z�)��V`�))�� ��i�č�*�2R����@,���_`��3uZ��,	pS���8�1O,��
�
æˁa�e}24��=.�إ�kk�OU�&�0A�\�NۡBx�P*:������M��=#|*F����CD�n�t��ɢM�A&`�AwH��qrxf}���z��e-���Gɫ�*�NF������2.%�Q��n���Z*���;;�r�L��:���A��ړ=�� �"�gE��|�n7o~7���\�;�p��������6�iɪȟ�j}әBM�.0��go����ßʋ� �s�����K����LHJ(j|2>������'��U�w��>AR@L��-=�yB����lҨ���.6�و#�B�5��@uA	�M��~��fc��	MW�I�C�E.�/z@'S��}����M8��|�*�jtd�~U�O��X[�R�쮇ȣ�c��ό���]s_��M��3%' �:*r�5��F�f7�����w&,C�AH��r��Q���WP*q�"U5ڗ�j�Љ[5�H �������Y���ۄ3؇%�i`���Y��L�t���u�n(�9|��<�a�M�H�L܎�7 �Ie^��۠XxX,�)~�dt�-�O�Q��'?M2�?iu�+\��l}�w���g[Q��1��xU�P��q��6�,����M?!�?�MT���M؏�D�J�Z�!��*�s��$Տ����2����z���3(4SԋòapR,]���8�� Cƣ^0b�$P��#|!�_��w'�r�%��xU6�W���~�ܗ�}��TmZeq� ��&&H+�F:(vT[�ǖ
�m>]ݼ	NJ�� ����І����@����OQau��җ�5��Oq�QZ��F~5��28�q��s�h�Ћ�yiS��K��^�	�{����&)��)�Ү�wT �g\7�'�쨋�C��&���X��!T����v�b�p�~��F�&�.S����huƍM���ö�q?4+����:oN?��9b�L�Q�}�x�ҨdU�{�8�{�<�e��X�,2�A��餾������<���:��4�ص��e(-5�g����Sߘ�!�xcK.�q�2��M�>��u�E�2�W�e��L�;7�ӱ�f+�q��`r�����IjV%�#��/�v����	�
�Plpv�nȸ����d�e{��+�K���I�E�_����޺c���bQ$�TX	N%)"&V��;�c|�����s��������Y7��U hK�X�Pak2q�33������8� ���qa�ë�H^,�_^��&��f�%�NS�x�i7�����OU��CFd�3�ܖ	U��9��V�*�{&�n �1b1���B7�_b�1{$�^�������¸�<t�b)/m�t�6��~��SSm.c+cP�'�!!7�-QP��K���������x��#\��"U!8����E_���M�~��b�[ڼn��G�3H��E����#">֖W7m	��ڋ(��
��t��Yc-�۳U[�u��-����y���:v�%��P~�`�������u$��s��#_������=U Y�"�Jɟ�9�8�e��nY�(��J�QJ������+���R,�n��9NX��E�����9�{!m��pS��/�$��?�W���10X�#U�OP����O��K��2x��M;��z��[>>�D� ��^%���Fm�R�������sa.t����v�*.�x�N�
PW�rE
��[)E��NM=p�,��ݙ^���c��M������)BI^�Eb�+QP�N�s�#�M��Q��t��a�c]f�h]+f�����j75lo��g��.v�f
_t]Sn���q�}�# ���ͨ����5ފZ��W?`Z��L��V��$��o���Dr�^M-$�_�m�u�1���hj�J%�H�rlǪ�%s���Cee�v�bL�_����_���8��Y�����X^J�7Z_��lF1Ep�r�t�My�p����.�HA��m���(SAj�iH]���!'���d�@\��6�zZ�xo��R#r_�
u�q�3(���훇m8"-3����;��P�/���5t?�+�I�◖�]� ��{	e�n�vw��
r����\<ٸ��);��M3��e�d��-^�w�� .�C�E���T=�]$�^]�_0|���Hɶz�D�X�h����+%�Q�!z�	��֓�Y+��d��b�f�����++�}����T�0c-Jc�5�>ҹ]<:*����S��$�w{�K��m���L�	N�X�/�]�ze\�(X%x�5W�<#�* c��!�&�gҪ�����2�)Hĵ���7�PTC�Qz��ϩ��L�JZ?V,w�bAƏ�A���2��L�cs6�� ��d�[�tͨ�~G=ye�%�����ժ��VB��y�'�37z<Q0�M~��)��r�/�TH^	#!@w��ɀ�����*Z�.��A��-��C�k�Jː�!��l�լ�rn-��VS�dx�}vj�;6 �@1�A�˯pC�W�ԉ�]AV��s��OcN@��)D���`do�A�Íܐ�I�雙$�L�����{ǲ�`O[��}�MwQ�/l�^��,�� 3A|���S�Yo���$�\�#<��	��YCV�z�����Z��D�=Dנ�zԄH۰z3&!�4ss�ᐻB�9W�pp���9����Z���q�%:�9V\{QW\e�
"�E��$�E���I������M��Z�-�`�Џ!���$ec�f���2�v�Y�I�iĳ�D���W�'m$q�N惂T����.�/�� �a�m7u�x\tb1�'�58c�H*�K�p��5"l|*Z��Q���}��hj�D�i���(�'ȭ?���*��v<lJ�0�ֈ�s�2����[-�)�9v��ʖ�&,��1�����u��PO�l���8�!�Ude��5l+�Ybˢ%h��]�Z��0���6��V�Wke�,�р�p���[�4��8�����z.{��[{.�?r9�*ct�?ϭ�0��g*U8Y7v������iWF����)ġ�r��|� �Tl'�#����H9�qN��c@!������j�:Q��~�/�д���V2��C7�KG��|P`����]J�Zn�!��r�4��G�O�*�[py�6�.�E5�P����T�w/�X�� ��?�B���ݺ�`��i��ԊKNY(A�)�G�?4��r���'M�f�������<7�=���1��z�[y�|}l�A��j�D�����T�K��2
��b�8�����|)��EM1$�křg���~l�q��O࿗����e0Jk5�����Ȍ�	��Xp)m�rn7i��2��2��,�g4�n;^̾��u���g�RJz;�m�-�~���i�P�F��W)�vȉ��h���׊Xa����t5\tf`U6��%ص21��rNFw<}O8�bM%�`x�梋&�Ɲ����hԛ�"/,Ӫ���|g�k��ǂϳ]v�K��O,��6�kI�e��uxUx�����M\"т��x��tRHa��NA| N�D�����a���KR����@��׍�4��rA��k�k�c�poTnT��"�Z�iP��K�}[���R��%��Q�A��Ǆᣏ�l5v�>�j�k�BIT�g��Q���Ӿ���p�>��g5��HF26�����,��O��s������u��=�2�.]��5b�vvw�a��f����-7u�f��c	��[ő�3�&�]�87JE�Ѥ�
J=�-O�*ŐS��e�:)8Y��S`7�Tri|��-�m����L?�WY]�,5L�SK��v�ž"N;=�
S�Q�Tֱ���������J�-]5�]���aK��M�U��U��6����+�%>��ɍ�Qj.t�%� ���@e��������d��f��U��K����~�{���W/Y[ڳ`�,��ग��ڊ4A÷
�h~	(E�U}����5�r�%���i[+��?g���0���	�j��%��Wn2@��7��"R��ד�uh�3G���>dG9���n��}��N6�R@b	��l'��$C��v#�)�®��Zq��z��+��I(�2m6��/�ώ���.\�����_$1�9^'A[��t�>�{CZ���BȆ���cx�RnG"5�׀a,��ܭ��t)ӑ��D��j/�̫
�^���aeK(�tRK����M���1|1&'�6�tDl��lx�h��9,Ǻ%ò��=�n�X-���N��\��'V�iܣ!�1H�>��2�r���ik<��U����ܬT����ڨ*q��9n�[��L��V�ɚtRF����i֣Y������Q
�,�k����!�|%i�b�O��4r����
É{�"t����;�b`�5g0�8�5i]��8���:���z_��h�#� n?��t[5��� �~-�c�O����a�7!�]�2I\:�%�q����8b������� ���W��cT3Uu~)�B4��/3��G_%�&�ʩ2M[��MصG6I+���#���{F3jκ�]!p�cLv��B3; |�����X����+����,�7���0� ճu����'�cs�.�C8>oT�y���[RQ_�E�E[ �]�E?�,����%t�"��qC#K�RD�������+? �;h`]���"cö�w�%a�X:D����o8��U�[Ţ|x!��jC�񤪧
��ۯ�od��'7�����@�6J���.D���c�����'/�g�5���*l�����GE�7���;A6�5,SXq}��6�rgbO�t9G�5�`��xD|��:��3�:#���ҍw�ݹ1���G |z�#�*���v1i�9}V�׼#_/A����$���Q�mrxa�y#O�U�>��4xzVƨaZ�P�^0�c �?�
1 ���&��]'nJ�!�A��d��eﾶw��T�p{��)*V(���e\���,V��"�����e�#f�:+lBH�<i��FA�-�I4{QQ��6����枏m�Z��N�9����7�"��y�?��VS����6N���4k�AM#KCS���o�b�|{��Rhrr�R�z&=b� `N�+�ʲK��tPfg����ҫ�q[�W�l[<�ͣ�L`���8���$����H-���W��4Dh�+Oq�aI/j�U"�w;��_`�>����4��=�
\����*�KKom�sQ��\yQ�~�s4��`,D�m�sL�w�������jVZ�rOB�űY]��LaO�B*o�FL�L���S��,f@�#D��ݲfr�<�c�ʕ#�t���ñ:�J��z�,�?�tOj���65u6�S����)Z�<}�C�3l��lնK�*Ӆ1�eMEef1eQ�oZIW^{w��we���i��f3E��J���;���g����0�Ȇ�x�~�=ݘ)�Al���~#��Ql����0�6N�'_.��#m�t���������� M���J&��+d%¤�L�v�N����8�y��I�7<�@/��y��l�{hB��a8��.Cɪ�,꼙������?d��먃C�ސv�(4��i�V�ͺ���9��.�V�x�ukrQi����ɫH�Vx�)��h�޲Ӫ�D�3.Z����7���J�Y�0cG�8V�|WyC�3Y�Yr�ɬəY�qnH7l��'�4 ���������u��s^Ȼ��A�p�ß�w�~�vImU�2��'u�$|���Eَ��0V,��/ň�@]�"��2����&4�j�7�ݺ_쬡gf��~'� �n�V���H�v�C/�(����شe�@v��I��I�y+���1AoDj}�$'�p�Z�Ы'��������bReY+���I�K��o�Q�jz��9�x��bEMUG/1�+j��iג[���� �1jw��L���],�{��La9&��m�<�`h�g����=̬� �t�z|.��\V��-i��m�q�8>�����x�:�}�����>Zt\�q1�u���;�� �3����/�{=����D������N��R�$�n�N��\���w}U ��~/�B��Z<ޒ��^v����5�`�kj�=a%�1����n%�N�9'nP���������~5�u+��u��B<l�D'�^iP�^���̣n�������X5��a�1����"���&x08|�D�+- a��8{>K�Ȁk{���'��p4ˬ�ѩ����(5�[�@1�o'�!�����݉��9��Zj�в�(��ӟ~�vXEi��M^�Ϭ�C�`��z����v��x"�k�J��0�_	W��Za�UȄV)q;����&~ѐ�GE���z��E���	�G�_�Ȟ+�]3{?�[̎v�ۖ�XJP�RҊ��w.�P r��[c֙r~~.����r%5�+�Vۅ�|Z�h��,L��?�55�"�^)�/�*)��_q�쮿^��g��ˎk�5%�g�=���^J<.L�Ԛ����`��7RK�����V(��@����E�O��/=\z��~K�M��ב�Gj*����@g���t��׻�A�I��� �~���b'&a��h,�1���1DE���둬�ݺ�T �(&;��X
�R�FƜ��](2��
Lt$����4�l��~�V4,�I���&S��<�u��f���h�{VC��,�SB���0�yl�I�c�%�jmYz��Dh���g퀩��X7U�L6��$Tn�@r�:����ꪒ�O�!)��<���h��T�PG��3��g�~��5{jMH$}���=�q�ƹ4��t�f���=},/�	�1�� �h�������k�h���ߴ� �CN��0�������r;�x����s�g��c�֍�z\&/�ȏ�+��=��z���|�f��J�(>��$�d"L��U��_d��-�6"�#RÃo,d�k���آ�)��'[lI�Mg�l̀�L�䐾Y|3gϺ�Gi ���c�O��S&�t}?��c���qi����u�#Z� �M4�8�h6�ޖ���W��a�������qW�-f4T�|r�P	�3��.�3n�`}hl������Ori��d"�Q�(��pr�D�A�:Y�:3]�9Aj|�
-L�ƒ%�z[2�?;G���>Nh���LͩN��>����<R���Q���΅�eu�_KG�Ko�T,۬!0<���O$2���wORE��z�˳�yA`��z�E�TG	�X��A��?S��h��r��7�>V��=�a�P�4��ڋ]�l&S���|hcV�_�9J�'�h�:S������0��-v[���Tr���G�X�5YyJ�W�=g���o�k�q�zL���<�}�G��CN�{�]­G,��߽������!6��<��橰�\���f)CwX\ˢ^B4�R