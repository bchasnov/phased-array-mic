��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�k�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������H�W޵α���N-�`��6����ݾ�FF��eF4��_}<�ےA�[,�|{�?r+-��5K�z��!��[��S}Σ{$Gx^����c��ƀPfƆ����Ƙ�P�Kt�U.Qd�ަ(*�:Ԇ�F�jdoL:�)K�o<h�Dxeq�0�!�z7������Fr�Jİ���;���|v8mG�?��s^�D�1��}��!�H8�$��dD�x�V�3F��l��x`.� o�Jj�P�cc��|ʮ�
_1��ÂU9'^>"�p��XQ'w,y���퉆�J� bL�![^)", z�ͷ.$�"�7���4�h`S�a��n��H�=[�u�6@8.
k��=�m8�Iΰ����w@U��Z,u|��v�>�2Ua�h�p˪ߪ��g��o�w��*�I��B����?�	D�f�{��%�G5�4���ܓavx+M%d�:*�}CꃩFu�yl���:�j9�?��(Y���ҵ7���ٸ[���+R�E��z��}ie��0z7���h�3�!���
��.j�&L	����{�xh���G��!��(�^�#	�)r`sa����(��u��^�H�өQ~a�b�_O��#�7G~�#��X� �fF�&�'2r�>|*�|S&5Zʒ�G�$c+[b�Z���u!S4��+r��;R�h��+�sw)��%���b�$����o1��P��/�IɞA��Ij nV؎��mn��&}��r5}?�n�Z|Q����G�zIHHQ<�1 ��\��P��S3��uKԲꔣ�_Ŗ���} ��|NH7��r������z�_��Wz[.��̽�܁6��'p1�s�I޼�@|�#�4��9D�-UB8+W���47�����w�>-|(0���F���o:�R�dDM��5פ;��)l�hi����-��x?uw�+�9Qs�8�X�C{�����A~+�)�|� nI*h�:�YцP��i�>Ţ�K-��Y�m9h���/X�5�>�O����������C�<AR�_���u����H9[NL47��[˞��`^^r������L�_�{�I�h�)�3�����Ӻ������V�7�`�Ӕ����}�K���(v�C[[�'��j�� ��$kح�DZ8+ϧ�ǣk��A�����rӵ�۩ ̖2&�Y�u�.��D
���<Gt���"q�ì��O �V�)>�K�#qv)Tk����B��z���C��T*c��U�J�8�xŔ�C�7�x����6Lp��J��CE~l�����׎���{�s������T`8��?/�ߣ8�,b[#T/��U�}~qO�ݵ`���,��NTD
���t�"�؎kE~�<�Ě��Y?2A(��Q�_�z�hU�N��1a�	E&T�.�0���ڝa,��$tIJL6>�Ǖ7:w���_d[�B��Z���}��G����5�q0@כ�DO�9Afu���@�TJT�ҷ\�΍�x��7�(ty:��"��J�c��_��(�r�kU�cr�&־��<���@�	��
�u�d����&�ڎH\O���x����.Y��1T,8��잌ѻ���r���M���7���]߆��r��5317��u<��^�Y-Y%��4c�B��9�V�R��̧�H�T*h��?}-G a�a�H�K��h���܍�;�u􊞄�Y�usj���D�O��S��qlڣV�:R���ֵ]ג�P��rb�a�E������6��%m�^X�]@&������� <~�����i���M�F9��t
>B���Z����Mz����9�<��>����{:wrC�����v�O�Ĥ�Ƹ'A^�&(�������_��R;Ϥ�D��7_3&���"��΀Ar�Iϴ!��0Ͼ��o�M�����P�*y2�iٞM�3�Gd:�4�a	���ve�4��������d �ڦq��3�MS�;�9�b�|i�[���;Vb�(B�!��4��g�	Kr�ݘ ��djɰ�h�v����ܩB�LU`Z�.fH�X*�g1�0��bHJ��I�����J'䧬�#	� �0�B]�70�i`%�_Ŗ�j�}�H��|
&���u闿m�����Tj��ʚ[vP��]_/,ܻU�E�t�ƞ�ΛNz�c&E����U�uҮ�hy�ŝ��#PR�u#�N�0d��h"���lDf�ާ�/�������#���X���*�� MyC�A�:q6c�������-Y�blq+�ī_��0��X��ez�Ljp�����ؕ�V�{?�~v������l)���.\�����i��f�`�: ��9м:����l�y�t�D;~d�~���!W7iмT����~�TGH�E���n2bZs��,s�!=���K*����(Ф	3G�вʱA�ͭ�n/뼪�Ba'U�:����Q8�U���H}��S�������X*� �,��q��StYF�$�$Ky]����AH�C�=d�L�`)%��V+��R����"	жi>}��o�Z��F��&GWU߮]_�����^
�5�~2�\J�i�o����{처���Ru��:N���ս�م�@�����}>'�Iˀ}�w�@���_���&-y3�)u����~�>w�rO
��I���>����ǎ-n�d/�k��Y�9�3KH���n_�a��*ђ�h�\^�L\��o�L)� S��F�<��)�ܕ)�Uf�e4�Sr�I�`�X6[^�k��x���_ ����f�d��\�P�*O��N�c}�������][��,���8�6� @�D=�NJ���k�Z��"0sk��W����eכ~ZjI�2�),8m�N-tmq!�ʁg�0�3���ׅ�J#B=�0S�~�b��U�@[
P�<��+/�����%�bg�}H���HB�ٸ��q,$����%�:��>��̗�N��q