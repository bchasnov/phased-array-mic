��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|/K�^!�� �Ϊ�I.F3�h�]D���� �1x�ϓ�k�K]b�ec���9�̑�2�۰�}EW��E�aǧ�b��S��+�/Aė �d��׫�~^^��y�4�4pjTK��~<OS[�EI|�ݾ�wi���tW3|��.�OZ�1޻��w���BB�+�{S`j����0���� �Vh��5N:ը�*�R��~ǣ!�Ţ2(<�����&��M��V7o��/T*�����%��}A���*q	Q�Ӗ{��n�s��S��~��vIv^��;K%�c��0�t�H��4���9��S��=t�Or(�J�!���`��m��@��ݬ��@�ԧ�"]l��~��WH�4,} ��cc�|�,��J�X���P��h��z[���ɰ[")y��!��z���:�i'��{��\k� �gßZ�/j��߷��C8�M����|�L�-q�
џNϑG��7�]}�Q8�	&�ēQ��W�iB$��y���b=�k:I�fA/�;��� �sp����)�����Z[/ݎ7�����\���w�)�F�^s�l�3JO:c.�t���LmnJ�F�P>Ƃđ�;���,&g:@���o�1}�E�Sa9��W���_�ՐγsQ�D���>���E����t�M�QOK�59+�%"<�����᐀������f���UĮ�wH���
���ЩLH���@�H�pY�<c�RӢ�ٔ�x�*�6�s/��y��M��xK3�e8+3�^�l��o̎xM:\Gm�F#���"�N�ȶ��&���<+#��e�ݙ�'Y��N��B�M�!�3�G�l2�� @�ķ��M4(q7~�o�{|> ��<�(�fv��\Ԥ���!�?�eqG��U(-�%q�W�o����Cb,��H�AI�b�4����ά����	h�>��8��e@�5r׊��w^���ea�%�����S�\�(�챢�R��C��w�i^���8|�P�޿�e�KX��~�VQ%6(0����'�n\�O�<e¢Oq�����,��pd��n�K�T�����xsZ-���7k�DJ�Xs�^W��t^�v[�X3t#���ä�P�P��E��@������je<��1��l��V:m�|/2wHB0*��}�9�)��jV���x�N��p�\:ߌrU2��8�a�Jq��̈́�lW��b{�V%d-�9^W���a='a6����&3��P�re��=Z���ьؤ�����Ϩ��%��DvO��~.ϓ�-�t9�r�Z1U(��e36"���>�!0�S.�7'h��E���#���ri*]�T�V(�����/�c�7����� )ˋ�7\>�؟�����'D�!���N[B�?	������"h����Gu*�S���'����aW�Rrh�ĉ�5��lJ�+翠��K�-�Y��)�;E-5ұ}�PX᰷)T�3	<z�-d��f���:/���9����!%��$��<����`�F�:j���f��W/w̘ �R�w��z�;�6�z<Lơcb�ie����#j�����P)k����g���#��]*������xF4�,X��?��"�T_%�K�c�k9��Z���Y�&�ܰp�3]�Ê�+�g�y�b�d�5Z־d��k��}ZW�2������_�_���!�� ���?ǕY�f��OB�xD���F?�q�'A�\���	zKM��>VFD�'A����-�חD��� Pa��o:!�����e$g��s�5Ѷ�*'��Up-��;���ܖW�D6��'����f�mq�U�Ї���AI�i�t�-̉��ug~pipXc�Z2�E�ͫ��}i��l����U�D1�5^S���N~o\r.���w�J���Oڕ�g�� �yd�pN�j��g��D��Sp��2;k�s�[q
r��褩F#9`��WC��zLE�*O4^ӧ��������<��_��|i��1��.�����T
�zUm	��4�<�G
��w%A֧���H�΍���w�P:���-�a�Yu�ְ�+���x^mq�����ZV�`QZ�9���?�N���9�aK�B�#L���|\l|>P�5���nfz�p־=�����X4��ΰ��߭�j�����S���y����1%��h�>%���~�u�����=���u�#�;b�<T�9��=*��	��{�+��[zrQ��Li�D�������Q�Ɨ�LR/��V0Cx�ק�hE���7�4݁�����M����:AW�3Iת��ߜO���t��	�F�A��6KsO���H&m��	�ʟ�-d��iQ�7u`^_�r��K��t��q��f�c������a`�K���X�G�	��6�����o���0�RW��Y�:d�;X�ׇ��bj&�ߨ6�@�P��R���1�T��&�R���S�O!ռm��-�wK?��ku�'�t�P�>Y<|�Z���g�X��.k+16����L�uоU5�o���jqN&�(3�i��u�,E�F��S�:\�-��o��LB�d���μ?[�@'�*-]�Ɣ}&����=�d1�v���w�{���"��HA�{�j<7��i�6�	6�}�#��U�{��-3J�[�$@����������;u�:��X�xC�t����N�z���筞~��S�o�K���\o��o2k��J��^g�;�>�)k���JI�z��UOB�~�$�	���
�0
LSǍ�O���Cuӿ���Yס��(�Q76��Db=L|�c��#������z(=�6�z�v%�#֪��0_2��8����g���������1D'9�l�d����v����}t��m�Ӧݝ4G̱Sً����Y仅�T�<�neVU�dJguR����G[C��<�@�#4���fK�{˳ �yՐ\N�KⰅ�G��V�P�U�;�i�~�{�N�,3�%yS\e�@�$�)&LL'|�@�v�f�~$��l�Q�jS��okX�M&W奐!�c
J�[2 ���9����ziF����򖔶�:8`���,�v7I} �8g��5��[�i�r ��(��L7�@�	Lw�� �V	Nn��ZB7���ۏ�b ��
�W��2��BM��g=͙�ϸ)��4�����U�V�Д7�t��RS�G�7J��9�`]��7��5�����q��'��df"۵!��he��,"H�W�꺦ڵ��ϖ��x�z(���JjF����
��/rc3�^J+9\�@���\���
��]7���읍�bV��"���E�Q��������#Jh5hص�A�O_��Mqտ[�X�2��>6�9��:���!yD8LQ\D�*i��He��H��1�Gغ�X�0���ל�K ���P0�3�?�_��b�u%$�(n�k���v=R˞s8>|~��uƽP��0��/�~\>�R�$�X�����T��Z����٧F�i�t�]e��a=W�V�I��ؗ;�	�2@XV�_'�-�@=��/����A]�kR�'�+���k:�A!sG�y��	��5�1���?r�Z.,�g�\h �fj��m(bTbT��Q<�iF���K{TjW40"�7���N;gl�{�i־3e�Wю^ޔe��p�r����� t�Y	��C軈��M�E�߮}�v���b�Cptu��#�'~"W)�c���#f�l��~o����\�����`�J'�]��k�h���u�A���>�86�A����]��%X�ku4�\P����B� �=@�����U^�.��GV�+�%���[A}B) ]�W׉$L�SQ����AW5���Q~y6m�����/ښ}¨�6_0��ь�ˢ�������!�h��Y�NC���4�[����5xi�Ϥ2�@#�N�jL2z��g�Z%֝$Du�A��i�P��� ��}@.^��)��3�O}G��w�Q�sV��c��\Q?N�qN	Ed ʀ���\�?(��-��.+[ ��?��ۆ$_�R�6�z�N3��|8ZNnH���ԓY��L? ���9 Q���rO���c�K�Q7�ۆ#)md�ߤ/f�;���;�qgi�`T��ɍ�q3�-�!p(���y�c��I�I�x��)�����8���B�F3KY�ē��O�	�W��p@����(_�H�w��$vJ��Gz��DN�p��>�(���o���槟�56����s�g�&&���D(m��1*��(c,Gc��y!�y���'{rK�B��2�W����y�n�W�Xh�>T��O�$~s����p}0��{os��v�V��8��ԧ���1�"R�ߚ>�@��t�yQ�'���nI�D!ɯ�|;���4�dc�ql�?�,����|�|��U.�J�a�T��d�[ އ�B�{�^��ɡ��������2����uCcs>	��H��pg�t��x]�r�#wz�)�Z���K��5f/i��,��,PGG��	ѨU�}{Y�|O���Ɨ9�6M��ּ��P�����y�٦��	g��9�,���+��w��嗧�<�P(_8j�v�)�����?�d$�< �ޖw�5)��ܳz\N���p���I����P�L=:�s0<��/�R���8��{6�qV$��9^�;iL�@���'�c0��㸸�$�@�8\��J5��K���ĵ5W�n�XCk�5Z�(��b&�(Fǔ�e�a�C"e��A�
|"�A�K3?����x�=~R`�=�{�C�ף��ps����S�QxƏ����)fl���܀m|�3���D[��6����>%�=佶��w�l�h�.1n�1���8�Ο�x+���GĠ(vnszY���.&����|���<��7�8:��-��܄��Z����d-�O�<��;���x7��^�w�I�U"��1,c����0B��'���S�!������=.��=�U�9}���%�Ɛ���f��BC9�0R^�/*4>6l��M8�C5����7�QTKwN�t`4g��x�%S�g��HB~C��{}�7��X�M53��솲��W	�	"!ʘ��3�>���j��.]N_l����ǯ��-K����o��jX�I��w��㫅.���r����ڗ6f n�͇���ސ7�+5��8ԡ��*e=���ٹ#+3��`�@��ξȞ=<��Y�S�z���8�<?��-��W�r��"v� ��%�%�M�اX�/j�)��~/��Q0)�ҳ�A�D2�f#h�,;�w��;?�B�)��x����N�}'�8RĴ����m�J����녎Hk�)�FC�q�`;FV��9�ԏ������D"�"9E��j|Hy~��2D�f��m��_i���Qd���v��䝥r���#�~����ۙP�=�����Q��~0���~�4�܇����DK�*�7o�����˺c��te�Q��D�4���a�l��iQ�Rg�ɬ��P����xx���]���]�N���)���r��`z��mVz�Q�Lr�f���a�p�N�Аg2��d�>-ϖ�e�����a�d�}@��-_�6P7�(���D�����M�c*�h�n�����k0z�z�&v���b����<S��|���Ay��ӆ=�\�[~�f
LTp>�v�?�q]L�\�_�8G�Kz��|������W9��r m+��\�X��r�� `�؉��D+e@ ǒѥ�<ý	q<]�D����m�G��_���5ܑ�!��S�,H�`D$tfi�G�v���y4^��p��6��9\Z���_�����o����.�	�U�(	B�0�*r� ������yg=�=H7QZ��)�MJ-�r�;��⣰��4�i�ǡ���P�?���������8~kӟ�ˊ!$3�j-�N�!.|�0�/����Z�n�J��%��a���^�х���i\X�4��)h�=lѓU8֘lX��>W<� G��IҜ�}�W����.���C�w�?���:�=����1���v������J�4��B�{Z�+�D�"n!�J'i�������� ��(_f�K�@MQf��,k�#pK�0B!�[ J md�2>E�q�C���]������B� V~AS 7��n#]�@*̆Tm�\��9�^���g9��#v�;ޕ����Ln�//�k�y(�6�b�wl1��>؉o����1�յsј-����I��B�wlª�L؂`<�F��[
����( �N�Z|ʪ���𭸔�C�����_�>�S�ӿ�p��� �w�eѼ����}�������:w�n�������O5|#��*t��N��k�S���ɖ����-!���<�ڥ�=W;�m��͘��2���p(��6�{�V�>XmN��D�b�]{������%�iE� $Gi|M#*3�B�媤������(c��6_ʀ�-"RK�FT��pҊ�Ѻ��O���
���n��x{xu{2��4�!�^�S�̯����x� M�B	��El,�ۨY�~��p'��oEt���iB����5H�J�nh���ǆ�&�/*/�%��-�l��w&�+�;q9�z@�Z����O�-�Ki�!�^,��K��9�К����m�b����l�pLCe�&y��,�=�;�blK�wIp��
	���b��iB��n���M��Ց�Y�Ɋ)��6��L�sݯ-�7�]�09�i7m�)�gf4!�� ����jxS�ܐzH���3�L��N�l
��TO˖�'�E{">n^7�eF�CK��j�ˢ=����w<����{�j�����}~�w^i��)P0��U����=z�M{���[���Uj#�_�o�>R�i��!4�����ylf?<��n8`����P	'3�$�̯I��f�4ػ(��#�y-��]�-O�`Ge��������_zF}��Q���#�jh��o$����:9��R�D�̅�f��%Id)Y �Ŧp�0���a��B�TLPln=�-��+:�7IYd���[5Zl�Z�4M�~�ηH�O'k|�x�G	����������	�n8pQ��ఝm�&��� �E�l�14~�`�za_f��0Uze�b��j�o�܃ʶ��c��j�_ �O���I)����(�8�j��V�'9+_����z:�Q�<O('����M�����@�����4��tB��8Ć���/I��6��ŗ�+��ߟgͤq պ.9ѷ����z��9W�I�)�^���E��J�Qe�[��mQ���/qk��Br��%-0g�{�we��q�\4g��Y���\-.��~�]�ɕ,߄�}ߍ�ԯ�DMC`	فP��p=�+���E���uno�V��nB���8Ŷڥ0�Q�qRX�{v�6��Ita�������c���