��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\����q�?��e�I8�b�Ǽ$��"����ׯ1�V0�����/]�^H�V9�r�8��	��;���j6�Կ��(9V(:��V��s�̮{17���G5�{{-izq���ˎ�P?V��K��L.�j�"���0��E��2��l��-���	�����a|���70+~)%���՗HH�y�@5�u�
Z��uZ� m��Z mK����?�4�g\8W���p)���>&*f�q3
F+�έ����2�q���Q�w�{���F��W��db`Y嚥Q��']J����Y� ��^���?<:�EV�[�{vw48���7d�R���%	��b��0�L�1J��:��D҉��F��EB!�N)3C�e��+��a�M>1�Y�Bj8����h��e����5��)��"%�e�B�,d�{׮z.g p~S�c�<�t?Qdل����V�t���˵�+[��z�+�w᯻%�3St��22%���Υ{�L���4�����1<��M����Ę^��|��3o���D`�B���](�D}6Fu��}�on����p�O�̣`���T�^�j�O+e�a|7�}�h�����WH��hJӾuC�.}W6��SX����a�ӪI�{��gt׶�AY ���[:�:gN2qM@b�I����Iã���62{��v��[���^���i�WV8ܺ[�#��&������F�P���Z�Wߧ���0h��j5��e���[���ߓΩ�K��1|�,gx#8�eF������dWw��)_Q�wηk��i����`�V��a3���������F��|�6�����VM�;�!rL���i �r4u�YiE�'�2 b\�`����e)�w�k.�b%�3d�'yHnUfɅ����

@+��Dl�/�*��oc��ǮP��wf�5�rX�?`���uy�;I`w�A�)�T-�-9��;�剩x�����voH��e��P��G�e�5Đ��B[�2���̯�뉽�;0i$+i0܇����LFs��s D��%��>�ɼ�ЀF��-X�Q�y���i�B����o���Kd3$��yB��a�'�T��h���2��{s7e����t�Ҍ����R�����&�ͱ�L��	o����o�b`2�K�蒃��C{�*��V�	�K���Kb4��Ն���y��5�z���Z4�ڸ9$�m���C�1W����nw��ȋ��
����ZN�Ĕ��������	�Ya�X-`�0����n46&��G]�C�o#�����\P[h1mt;��mM�t�+\���L��M�A���VF=cn����$͢!��d�'�$T�M(]�6��Ͼ{�j����i5�����#?���rW��W)ِ '��V���w>Jf�~��`2����}J ��F��c9����/�ő�E����C�(]
$�qE���R���������x��l��h�9�S�`}Ϋ)�Uj�F2�Qu�7�p)%>j�e:w�4�N54�����ѵ�e��fRde�:��o�Z�3Z�E���=6�'*]{	�ɮ���I��s5@�x����. ��V�8#�Y)3��^�M�u/u*�4���%�6��aws�+�\��K�ٞ)Éw�'=a�V�0�!X�1��8�u�n�ކLi�0���%a��� �Cs7Tk�s�ۚ����晉�N_�D�3�Tꯧ8BF���O�l�# ��6P�$�?�?�GN�q�C��vnI���C���[����.��dV���fMD
2 Ч[�]���^��g�̈���g����SB�1�&P�MP�V��a[L{�oo�W \�?����Z}�(�*F.|�=xtOA0l�#mq -��:��x�P�B�GS,%�b�sF�����vZv�KlJb�Ө����o��gKډz7�����x^��7�&����8��ܯ{6Jܑ��)�v��%*r�
̀خ��k�89��7l��d����LҀJ�{��P�B��Pi"{�<�\ʢ�:��Ⱦ+�[[���֨1ra�t�.�j�w`�����0':Sr���M��@i�`Zz��&�
tٙ�e�@�V��My@�F�
��m3������`D�u����/֩��7��h�i���RfڸS\�d5̏�M�������]���H���nm2 ��������o�U���X ����1'q�N,cD���n�v� ����>V���]
������u��n�y�z���&{a<u������
���,�5��Fӆ��ҰF}ۥ�-�Ur�c������픧� yw�RE�B;-�f�D
�@�_��]�$HIB�|�KfĄ-i�rҢ��B�5�@I����N��pp9!ФH51��x%`�{�����n1�Er�B�I�'���w����(�_�8$.���k`���Rb��BA �6��da��B4f/l̼smn�"�`�v8�Js��B�[�'sg>WH�O/?x�ez��N��8J��w���w ����#:�j(*
&�@[,��zd��������9L�gLVzCr��+*�p��NR)�<��} /����Ja�#�G��iK G�)L�s�JPo�Q�	
+k��'�m��w8������l�ה).���4�)("��>h�!�a�#<d޺F�^��G�d܀{���uC�vޔGdg��*�\�9�J���;�I��.��	��ОIV'��wUf�y8����m�3���+��۔���y5j>,^u��)v�k��&&pYfwy���O������5�6�<_�y k뭟W�XXq�1�!���H����E3�Й����c wY���*�ި;����T���azt��F*j;��B�!���{��h��ˤ�Q6�9�Wl������@o�ĭ�d���WB�f�խ�wQQ�4�Ա�+a*�$t��J�~Rg�i�6S"&��U�C�1����@�=R���bţ����r��������VL0uC���9�Lf�D"�햯�i�^�����mȒ��N����!�@~�Cq�ǆV�?�:x5kA�	�3X��8����-���q�^a�+�tO������zY�1:QXj��}����y���F*�	 a4�����d
 "���3����!�U=�6`���_��b1 @vj1ٵK#�j���a�����R�t̍�W���H3�&{�,
�A��'�<0���~!��4ۏԀí�+����{� m��IB<��ҍ�w�9Yfs4����y�����7�,�0Ru�E�jȰ{!�a�c����Bf[+���LG63�Yój:�;ֈ
�3#���+��l �����H2;c��� /qs�ƾ\0���])P��.�D	\�4��H��Z�m�n��WR~Y�	S��s�����So}F��m�w�0���.�/r���`�j�e¿��ȣ@��mb��_��������~��	tܘ@���`� 4��9� 1��`���z��MBX;2L��	 "�[g�ĉS�B���[���3!�ó�Ј�TN �R��Usܺs�hDDn���ph��/�E����o�#/�6,w�����2�:n!���$`�S.�C���j�\,
�2e�"]��J-��*(�Y>xC*��'�թGYg.�~�&Jl�'V �5L�Գ�D�@�X��lg}qG����3n��7�Ɲ��䀔+�8C
�<B�n�j]fI ���c��Ȁu@+��:7�$�2�Q�i=Y�n"�6am�k�ԂU唵?��g׋E�K���k�,���֘dZ�:xvr_#����`�rX닒��:n�P�Ck��P�S</]�v}���P�vh�� �*�7'�lN�e��b���_�����.9^�xEJ����.r�o�5W�~��w�T�h3ĳ7^���A�ǝq'�j(�܃e_{.�4�n�������0Z��*6r����M~�6i{o���x�?@��O�Gm����Nq���U�2�\1@<P�!�c��)Ы��}����%�gР�K��,�N.eu�;ר�7�H]�\�G�t�Q4�D�g��n+W��ƃQ��ߛR��3�kP��ES�� ����n���ʗd7��oXlk�@2R��z�ˀ�س�S��UI:��� ά?��xSr���Q;�#��ǒ��(B�����V5n�𹓮��g���U�P�+������N��vIT�\<tH3章n3��NY�Jn���,�& &�����H��޵��FϹF,-8H��u�`i!��QB�Z���˻VsB�>cο;�{P��]hfB�[��7�O�O7����Q��x1=�/R���(L��aKEC��lE�z�b1��PS��\h���^�'��t��@V���oJ��/��Y�vs�̵�8��}�7Gϵ+5�����1�Ҏ���|!����:�^�T鸵5�I_�j�mގ��\�gk+�a�Q�$�3����Y|t�t T�y�awyY_IX Ux��	�<�Jg>�EP��
n��^����c��P.����i�,�6�a�ª���{AJ�Y��r0@�#W6�3E�Ziě:{LnW@~+�y�2֤jj�F2_����M8��j�l���T���vΑ��)Gömٜ�%��!\8��bZ����Ƿ
<&uxav[@�
\͟�����bz��P\���G�T��\G�R���V��%��O���)�Z!(٠%vm�W�����^w������~,=���ܡ5}x�G�:"�a�
��4��k���l ������+v$���j0aO�Kl��x�h�T�{iH:w7���$%�jŮ�e�CY�� S�ŷ5C9_Y��߶MN���j棍��L���j�l�I�h�
��)8%��Hn !��x��Z���1��녝P�: �L$�^�B�dj�����$��H��!	�� B��#�k{����~��,D*�H��~�>�/��,�@cZ.WNK!�e�͏�x�H�>V�f���q�i���
�w�W�]�v}ǈ�W��]���T�T���'��5�O��hww�y��1�lu��'����\+�x#w��� A�T.�<��X���/��Otg��ī�%P��7vӗ��w�\�V��M�J�l�fm���I���G�8~
��^�Go�A�fip#��Ѡ١���T��i�5�,��$K�xZw� k�2)�fK�%��u-�עYG�������X��M��8X��+It�$�U8�p'�C�B~l
S9y�� �j���>Q���~������M�"����;���?� ����G�������^�M+y�W���%ɇ�(���b��!�� �!��4Ԓ��N��ӰQ)�����Э�;dR�#�����EEH���� ½�P��L�x�1	2m��Nk�i�3� �ė����F�E{ޏuD�6�j��k}�	�K��2�-4�>o��92�ȳ��#Y�e�Q��ɬ�ÌL�dZ���T��1��V��zf��u7���@A�?���=���Tǀ#�	�ʩ�,�4� -d��������6�SYY��o[�ʶ����6�����䔅4y�5���Ӣ�}\!S�w�����[Oz��c�xr�~u��|#�������Na��F����:0g���d	G����Kb�x���!���q�Qe���*+���Y]���묇X���=l�.<{��\��~0��g[y88eL�,���㪊�b�Cھ�S�9��QE�@����aÇ��Ż����}�o���1�v놔�u�($�L�b^�a�%�)�f-�3��Ol��?Y�?�2ܲ7���9^�j3�'Q>J�,�K��O:)���4D�s�3�P��zq�M�y��}M@��u�Pf���ү�[�Oۢ�\����q,�$���M��ܖi�ZL���5)ġ�@�>�5	(֥����k^'��߲$�����w��UYP����`)^L�t��\�oFH:b�t����eZ��iS�@���vǺ�Tr�h�f�ü�r���mq�a�Ҷ�V8�����3l��ߜ� �-[�2����H�
[(U?D�`2�qes�Σz�k
!�~���}��ERd��Ɲ�����at`�i���q�E݋*�gOF-I�%x�GA�*ۈUa�<ȍ+��=�>��	=�B0�GU���z�Y�%�'p�7it^p�3����M�ǜ�	Y*�Y;V�Oj��u+���aP��/U�u�R���'�,iEyL�@�2�_*�t���qG�h[{�>��M��>����W��V����)r���Y�M������4s&�?�o��W����[1�s��"�;�~�V�`n�i�
��c�����?��;��SL��@_� 5~e^�s�ͼ��d��9e��}����z��'٨��Ұ(FRD�2��Mb���#�����ɢbBCy�޸_�ݹN�Gp�޿�g�IhF�?P���<�c溢_l�d���q��J�P�c
��
�]0]����W<���|�.Z��Om�D��@ڔX48��曘�g������v1�`E�j*�Ձ= ��=A5�
:��QW�yR��|�^�8.����k=&��X�ǍW^���W~���U���r%C��ǙZk[Y<a9\N�9������,2��_ļQ�	.z�>3@ܬw�N��H����n��n�:}���S&t��0{D�t�P���ds����赡쟈�4��m�����ɮ[���^�@	52�i��z9�����7E���N����[a�*��8�����*�����BYR��Z� (:|rɮ1�=�v���C?Ho�z���zb��4��c?��:8�G����#[�@#����
�cfyM�}�#�h
��6�5슾�?B���r�lZ ���,��Z�)_>��c��)���U�=瑮uN�	�w�Ŗ�}*�[B���VǏ&�V�������z����Ͷt�Cp��;���(�_)s�A&9%���0������RC����V���i�����9�-'���Ͽ��q��:d�+4�꽠䕅Nʃ�e֊X�	EL��]Ѫ=�i�]��A�B��)v�:������
���p�����;_T_ﾰ�=3���米Z��YaB�!��2��^�� [%5)�m07��=1���P��p��F�����ڻ=�B~��8��`���6��s�bi)��qk�$�0���
`�����3���[f���Dio��N��ֺ�,�"�v.�6��d����+2Um�9�K��Ԅ_��u�-�,Q�4_�}���*R6f�w�Qy����T��w�8,�>�0�j���w\���>Q�ȳ=֭�.a�]cJvɰ�;����e�<�r��G�.��,$�'A�k�+9��G\!�����O!�pɑ�6��6'nW�q��C��m�i�?J!yv�;��ǳPد2��O	��s��@��㩏�m�6B�z�ϘI��(4镔�p����$����5�3�E1ל�Eu�L&z���<i�I ��5�~�֮Xo���]�im�{X\�C�[ê�#�� s��L��&x�.��U��-��$�
�͚�3h�҅�!��UM�!?��v}�C��9pf�rɓ���pQG��s!��|X:�r9�-L���>sL��o��7���)��_����k��6�L�*�5B@�jVMq�����M1�gf�l�[[���C���x�7�H�W=H������l�4T�R����a�
��0���H/~x
}�^ ~*��p���/�G�l�e�
�G����34���W�X �����)&�Kc��� .�D5
�m����B�^���m�<�8>�6����?�mw��G{������ص(\%�&-�����!����^���%{'�o��Nճ̃C�U�m���N9k�)�:K �Rx��#bHtfwXn��X��u��6���[_Vod8�z`��.%x��X;¦��x�&q'+�ߥ�|#���+�R�	�sW�onp�NX��Ϲ�e'�Tq��|�~��IDr9 ���29����.p��/��:%Y8�̉�3�7Z� �Q1��O\�	5�RY�i@�k�����&0U�\��A�~�lL��n0pW`d�c��$7�U$ �S� #�ڨ�P`eД�(d�"c_��^sz���?7#��Tw��¦�6��I����gɸg���ԉ��򈽪��Om:�)�v�����	��caG�TE� 7k��2�jr���+2@K�FO2u�&��y�̉x����F����<���Ӑi,\�~kS�ƾP�n[�=�SDӲ`�Pt	5�G��p�lt�J��?n�[���ʆ��Z>�m ��Ȅ&�e0f7��g�C,^�������|M?�*R��C��F&[%��H�A��=��p�#ы���p�[�f�����u;��zd.�EV҃�i�1D����!pb����V��ʙv`��ͭ<|���f0��E�(�;_�C/]TZ���%�q�SCt�4��t3�׹����v8��8�F�c4V�[��}c�꫓]-���Yo�9}|~*W�nT����N@n ���+�^8���2�d����t,1�i�%|�¦�=��1�J� ҴC�Г�U��U�z�U���LP&��^�\bG��T�A�X���4~� D�0�?��@�8���{u�3�E�Lx�S�&��)�j�h[hT��ۯ�ـ2h�G�\�rGtphv��\��͛�s���~�'�Pİ��VS���N�����A�-��@�i,@�$"r��m�K���� �-Z�ԩ+8��O����9�q�u���l��§���؋�@[ɝ���x�Gf�% �f$��!�{+@�,�YR�բ�S`s����)�C;�Y�e�������}���9rWȭ�.���5n�$�ES���L��i��|�%�˧F��}F�)���F_kD
6��wSo*�x~S�g�U� �M�dR��Ɔ���%ή�9>�:i)�?�����d�V�c�mLhq�#*ȋ�e'���1�Og�v2���@xyʮd���W�Ef6�xq+b~d��5�¿�/�(�
O%ٽ�6���`H�)e�`@:�����J���aN��N�G�+9YB�G����h!Q�k!�����h�Jr�����Mw"2iH
{L_�*O�t�h,�l��U�ybJ;�fA�5+�Y$�B��~��*�
�]�KD���*̓r��W����*�g�2\����q��lj���OD�+��;���.��n�3��~/�
���H�t����o�硔��:�~)�}i���u#"@D���ءX��h9̙�j��X=R�OQ��R�~�?����U`����1�͖=���3�݁z�v�0�yn/�ffW"�Z_p�F���&�MJ���D����z�&m�3(<E��c��>���k�R�5V�r+��0s��N��x�?s.o?�3}.0�D@Y�(��d\}�����D�D*���<aɣ3ھ�[D0f��?��-\(�X�{��ޔݣ31��u�	��mku��ō�HM�]�:3�3��J62��JrC5�V�b:���e\"q�j��cT9���Q���jװ�nk�u@���I�/�9��s�\�yz������i�5oӪ3Q���b��rVzK1��?u��}ح��+��;�lgU�DIF�g��vu.R&�yH��y�
R�z�$:p>v�rA)1�Ö��OnW;���@��Ϙ���o�����fS*�|��s�=os+DL��渫z��5g�%��^u��5�#��}�T/�@D7�����/+Vv��M�0��y��JrNP"6!'�W�?�L�IHs_��UM���P�C�
U=
T�d�ow>Z����VTn��,C�3	��^�[`F�_�E^ӾE�A�$�&o`�)��}~�!�F�bV*ިq��AIe�GT�]������H��5�(����wQ�u��SՏ[4"��fs��(�a��z'o�������2-MIH�xA3:���)K���kW�V�#{FО�Y�!�q׎�:�|\�H�y�8%Ol�����~��[�]�����	 ��$)k}�3�8��J~m!���3���Zq�'"v�Wkҕ�TEn[O>���m��y�û�@c�.�N|�8gS0�-�g�"r��J]��NC��p
{���B�k� ȅ}"�p�|�s1'�Ww�VN]nEm�{����`��_.�?k�{/��!�|F��;�����BZp��bVm,�D�/��Vֈ^F3�2*�l1�*���c�n/ ,
�oS��:�a�˙��
3S&r���z%�:���C~�FM��`b��8�ǔHKI�9D������ޒcڲ�&��=���Y���~�������Qߒ!���6��U<���~�L�Wkʏs�'���"���7��8�;l_r#^2{�V}�)� _�՛����t'{���y�	#/gq_vj0��+P��F��Z^��b�ɲY�+�t3/��y'k�����]{�QQ���}����d�sed�F���8]7�֪�s�e|'X�U,�z¿�\A'�����d��J���ͨ�I����Չ��2� �F���? ��CM\���������0T��*��78EZ��V�F:��2�.�p
\��Ԓ���5j�z.Q�4I��@�q2�0���B_� -���J���~T�^����"K�06a��"'��=��5�!4���<����A/���/)�G������>͐s�LW�|*B���S��.1�9ڏ��5��[�%|��q��?�B�����ԧ<�"�x=�]b���g���Z���:���QP8��S�h����\m~蕳�P�!Ǎ�1���r�h���8̙����7��W�`i�?(�9�袓�ܒ#ϗ�O�} I�<3��ŧӇ��?�7h"�hRbO�wH�v�Ɗ��	xmU*~8ҥy��Q�b�j50r5Hc��E�v6� ��8�>:�|Dm�g2�B�jP�Fh��������E2|������ �1t��M�'��x�>[�v4( fV�Ϩi��:`��i����F����|�?� N�+Ot�,�џt�^����Ϳs�5����IX ���L����GN���`S��|"�0`PG��ZI�P��b8-L)�8v8׼Y:�Єw�_���k_#/��2���A�%�V_h#�;ɧ|H��ߔ14��3�$�[�+��8.i��a#KϮE������`���tf�m���	94ϯѣ�������o)���G%�T��Z�/1)�rW����MP���W�(��]��p,�V�y��L����_�S�J��Rv�`�%�p�������Lj�WfO���T��&��<#������JƉ�X6K�f�94J4þ�����-:�,�N��_��M�9��^-�N~J�g}r���
�� ��WHd����82�#j��[Zͤ"��F������7�����l<�}�c�o��~2W�q��d>�q��_���g1'��H����=Ƶg�cD�mv������y�k:aRx�<Tb��f�#%V��O�����3��ĵ�|Vf0�^w^������$2U�=��9'I���܈�
g��lyj|2�,�|I�ܤ��!���䐛��+�:D��,{�<��9G�23.���+UE�u�]@#u�n�1}� �8y�U��Գ�H��̌6Q�B��R)e.�v?�~Y������^+SHFi�=��K�L�4�=�C���v�1Q��?:�i�����uT z�oAR0���E8� ��Xbe�Ր�n��g�ǔ����:��\ ��
�n����/�����B��4CP�ZĹ*<�/{5�83[�Uqi8 ��1q-�'f^��o�91ə�g�r=�?�pܰHÕ�E0��*���l'�Qp�l*\��&������1������1Sv�ɛ����k�=���;�����=��ĽV+s�a�J����%���q����ks�"������8�#�$S��Р�&�5���*uy���Ct�P�<.�T������{�.�Ta��n����.���O��N ���j�->88�߿�w�y7�G�e)Y�����5^s,�;�8������5�����@S�<S�%K9u��.�߬�e�)���{���g⤀ɼ1�șfP��Y=*�B�����E9�v��"6]>::!�t�?��S�>.�R^���CK��o� ��b�ld<��k��C/ok�1OQ��yx���գx_ ѝʘ�*�$ݐQ���:wMcI���ag�e�v���/�D�� �ݽjDQ[�ѽ������U��������ّ9f_�:!inu�� �X�$GY��!�3ߣ�q��o��՟%�}�r*�7[ ��c�윭������:�V ��c�V����^�@�Ys)`��kĊ=x�!�;Ϛ������@p�{^�>����b������,�i#k����7�܁oj Xm���ʹ�B䅤�Gf�G_���d����h��l���6��9a��/�樼�d��O���a�`���׎�
r����IR�U��A�&�����/��X]��/.7��Q��ie�yJ�˅C'm�Ę�N �%�{�f�%��V�B�>98y��<��v�{8��G �9��M��e��ţ�`L޴怹�a�2�_@@M�6N��X|�E-9���ˌT�h��>�A	I7+�&�0ed�����?���F��R<ølfe/���u�d4�j��l�2�6Է��L�H��hѐ�.�{�͕�č$<�� ��=��S0g9�0
����odT�JR�h҄�l��t1�2w���g��6{4��6
����'b/��Jh�m�=X6J�ܷk��҆iz.��Z��czq�������$Y�����TM0�P��;����kl�u2��1m�Cſ�}�] ��	{��EP�}M-�~�a�~?���'X��uE?��c	skf\��x���}�/�����QY�#}��ߌ>�%�藶�iؽ��!^W)����H5\��<����	z��za�{���Q���J6��I \��4D3U�nɪ4�&M% ���U����J-;�AD�59��J��=+��-XɯH�?|�&۔۹5�C��큚N#n5e�p��kg��"�V�������Zm�{����_b�^�o�a�s�����?�uq3:��a��B���8�H��.$��!A_x�
�5Z=�ѓ�֜v�+jm
�+��K������b��P�^�J<�7����5p0	7۝�m��C�������۔V=|3���~ϙ�j���Ǒ�uX�R(j��������5+�+#�S�{��Kz����+�	��9I��
ӴM�&v�P1�~���k/��7��〚%"�Ҷ�Q������q��V���q��e�ƕ��%�؛�w��:��d��:����Vl�J+���JE�|�p��ߋ������sP��7�*�!�"G%�����Mb��6��ߋJ˚EK����K{�;�D��rU��i.;��}n%|1��A���`�9�JW|X�H}+q'i�|�갭8T���p��ܳ���\����韝�W2b*�*���.�����!�4�<	߲U��*�om�ߓav�&��V���$O��z��OK�aia��I�5SB
c|�t���	M�e��ҷ���.[DJ�\�*��0�ٹ0>g���)D �����!�Y<� �S�~=���}�{z5p����VdgH4Ɋ����Ii&e�˩��D�w���=���8�6R��j��hskl�C?���()w��}��AŶi�c=�6������ؠ�Ȼ�e\ެnV�eѹэ7v�J��O+�klxN>f���%!b;D<��Y窩4:���.���ax4l���ǎ8$k��������S/�����/WR�k`��%&���29�e�Զ�lD��ۻw��a�@���h�y]Gi*�|��ф�L��,8�*X�`g��b,	�g�x{H��?B�z�bT�V\�w�D�]A:^	WHӧP'���qE��mD���?� OR��"��PB��kZ�p����Rn�^�e�=�>��D�VH��g��;��p�@Í��(t��"_x
"��hD�&���k�֫����K��ol2%��Ez?@Jl�zʽ�1���r����4aN��-e	e��M�mVn�-u�؈ېw��#g1,�V䳖���͡G䅬�F&#��bn����}]!�G�h��؟���~Jo%��K����GS����VK6�L�'u�('0'���5�<�n���R�>^���\pX�d�5GZ	��H�� ;>�����"��H������C�tW%�@�Q��e�t�l�KZHK).�����e�
��ˡ�,K���C�&6U�$ŵ0��E��Go���$���~$����5-�� {��Xgi�E���l��00R�X������^j�/��ק�6pv(�I�����'+�|O�.t>���s�;Z��4M�"��8�h��"��Ղ��j�2l��a�.C�����
"�{��jL�1+d�����Ԙ��\�g;�,�%>�쪿'E+�\�4���NI؋[�\����T��b W~�8�_�n���(���S�T����'.�
�ӗ��3F!�A�#b]e���M�w����|}ה��:�M���hMЕ>�O��L)1\���B5	�ї�K�d��4r��q��^��yB�����2D��P��=��!<��26K�el����j�#N����,N��2|*IQ�1��a�V܀X0[h�<leQ�� \��c�%��B��>P�0_����ou�=����|�k��C!������.Lsr� ���ÚqQ;��r���c�f�X���2�����Q�r�O