��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�tڐ�!��Q�����xZ�H��V�� �]d��� ��h�hQ�/���o�~�կ>?�5�z�+|��"D�[�!#��.J �SJ�Ҕ�5�Y7�0�f[秡3ڕ4�O�~�	����u�Q�Q�H��)*��V�o���}m�'_z�8�y�@� K$E�R�5^R�Ԇk2�vv�#�80����I��JI,3)e�_�&䜭������=��Ӏ]g-����Q[5g�#AҤ	F���d7��(�Bh��ѣqL�#Eǯbw�Ӓ�4Cw��t�h@r�!`�=&�#(�wUB�"�)M�5*/E���(ߕ�J^�/5�P�+O>�4��ʽ|���遱->�0 �G�I�W�a��s��#�IB�^S�
�t�rǔ�-4�9��s�g�5�+�55"f�!���f��DѶ��X!���j�_�6�H:���_uwR�=:9k0�h
�`��̆�hAv<��3)���<����y�xz/>�Ht�G���D�Q�Je�UEo�"S��u���	� ��1e;A_�PKV���E���E�9^�a��%�z�B���.���
�4z�>��ƿT�]{]��X���r��$Sv&�G�Z��%�s�~�\|R�����I&M�Y~�Lc��\Y�\R�6)'I�d�cK��9	2;���HY$<i@���!r����|$ӥA����3��r�z5��3OHq^�U��sx�D�?>���<����!7��(�$�ĥ��n_$m�C�55>�5���;�~���F�
�H.
֞CAf��ﺊ80�G,�5�UԬ�;����$7�/���<4��r�H 5���
�^^H����(�Dܨ��Å5�V��dU�.'4#.ҹ�����=<}˄��_��L��<�TM#z97-�$:c:�T��7��{�X��]2z(Lq�����mO3��Om�rZ*F`{6��-��{NBE7b�{s���r�*��J8�Z�2� ��[�aJ;#(��AK���}(a
�v:��@��5Y�!�S������w�=zb���Y.�S��Zj��X$�������_��W,��X1r���w�M����W�V����¾ψN�{�I{4߂]�S}h]o)�x�m�%��A��U45"s�бѮ3d���9Lrb�٣O��?{�T��"jVD�7;�ZA����ٗ�+i٢�i�:��{rD�Lӭ!4�w�55o˄GrE���>5���'�*yk���u��:uKVnl0q@��&Э�<d�r*���EI4#�t�д�1�W��R,K�������ʋn�$+�x�dx>����DQ���1bH�@����ޏE�^����#�}p��x�"H«��"��dRԎ�GA�r�Ka�ج�5�)8�V��g�`ݸ���\Q_=��8��0�dS���Rx��5����Vr��Iy�^a��?��冎�e�	)W��F��c5�5_;��V]1nګ{�L%�),�)=p��O'�%��I+����$�?Q�F<~/�$��=Dg����t_�`O���.�|��.K1�h_P2�
,I�_�H�0�Ez;�L�]��۝+���SI�z�d���v�4�KP&c��@��3�	J[
c�9-�+��"4��|�B`|6�3��JMX� ��w��%\u�(�>��&��R�+�/1YAK}\�<��̹+�z���0�~]���C�|j����dTf#�B�o2�}1����X�=�"�A��T��]�!Cf��bmS'��=5�v�>��K��܂���}Vkl����	==���_lš:s��ʵ~ %�̓@�����p3r��pj���.h�F��c��^�r{§��Y=��rM��f�����U#ܤ7��<��>]���+�m?c���H�.t��6�����B�C���!_:"[n��q�u6�C�	c��֞��3l��������k�A41�f���1.q�S�3gF��;�½�6�RM(LS�񬓷E��1�EU;X/z��@_tDL箭v��O낭��<!�XH�\}�N�G�FVό��9��c��R���(Z�w�ʦA�b�}���g�!)�����"��;�J�0S�L��U��1b��0(��2��0$_����G���o�\;�L�hõ�4]_\?!V��g͐���w�C�ì����(�B��%䄫Ss����ú��S��=���QЂh]�0:q̓挶d��}�R�����\Ww���)�ϖ�e������В*!mz*�����=q�7f�H*�";�{��G9�+��I��D|�x�z�S�ἧ���V6	'�v�}s@w�'�=u:��B4*�_YLoP�Կ���V/��W�*�e}-t�$����ú+��U�[\��oy���RF_����(�iʎ��/V�u�{�y☺��oM�p����Yv�+M��:�˖d����^I9��k���>�^#_ޝ��\��"����E �g,h��\(��]p��|	'[WJ��"����'���au��E���n�+�>Ta��/�~ǰ�}�2���ҵ�C���§�Ժ�����9�@��Ф�%�|�\���LPCT*��A��l�+�uY�]@�����<�A��U4{�E�S����2���V��{�{1���d�-qf5�i��}���0BK�r>y�E���y&���/�����ձ6:$�32PI�+Xq2�Yt�x��>g^p��g�㗔h���a���"Q�G*�
Lxi