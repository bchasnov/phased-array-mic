��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�=�V�i����K�ވ(Uό��ի���`6�dY$;v�#c-@��z�Z�0w4�(�ࡉE��^ٽ,c�v^KeA�U-�*p[��Yj�(/������+�?��5���!�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ;l�Fv1�ϯq׆������s@���'����j����դ�P:�Cb�{�'�t�ɟ�>��(Hw-�u�� !i�^lZ��C�{��И���i�-|�|�I�Dd#����i��	�4�@$,d�������v=�3�A�pO�w�tE���M�ȼ{;��?4P:ٮ�7���F�ڦ� w0=L+=~�&P0q[��^�-\ߛw�T��e�z�"�[S��B=q��È��A7�D��]�!Tl�f�+K������<d��\�毙�����gpȷX[���;ފ@n�%%�WNr5��X�hqҶ�=PY�0��WΈ>��uX�+4 ʿ =�������5�i	��,�Hɴ���d��h�(P�pFtk_���'E.ݷ�T�q����l!�&˃S*��, �FȽ�'(�k���=J�?�>:̃�7�\���9����Px%[�C��a�d�%�}�qyh�!�ۍG��x�58��Θ�|l�zFSg�\j=)霃��f��L�U��!�@C(����U>�RRrT� ���X(�A�G���I?�/�I��"�?�Z��E�T�w>�3p�>����G�FJ`Eޑ^��&z9P4��,�N���*�
;�˰d~4�� ��'�L�͛�e��ث
|%��QLZ��s����9[S��ʝ��:W�7��������gG�^:�6���3=x;-��;
�
��_a���-�V�,+Z���N�69"|����a��tZ>�G�.�/�2�7]�Mg�S@~_m����7�ZҫӁ(�,�	2?���G\�^�����c,Sʴ� ���F�g�\OA6��-+���L�����**l�K��:H�\��B��r�A8��ѵ��1M jp��x���?S��p�k��ʷ8ώsr>!w�2�O���q'y,�g{"�b���ipD�L���#2d��!��K��VFha��_�
]{P���(���*8����N}��^�g�&��L�%j�s�è��s|�IyHP�Ao�m�mi��Nȝ�j����*�
�D�+���v�.RJe���N����1Q
�.�%x�a���t�(:��C�Q�X���C~�EY��!f�����
�A�L/�	Ha��KS�7�t��Q��L,����|�����{� ��J�����q�?��"=l���z-�-8�����l� ��W}���3�p���5�������4���B��^�n�^�5��w��C)�k$?�(��J��	�剃ل�p�]Y�������/�2�3njR��A ��3wQ"U���ش�N+oR���ɉ�ˉZ^�Rr*�
a3S��ra�<��+�t8��`=��}����F�8�p*pPC��Jp�ۊ̶n���=`�ϰ hݙ���	"+��r�0s�������=dzx�<A|�vu�l�Z�7��x��`&����ы�hP�����$��Ă2LX,]Y����!'�TGY��������Y1#�ߺ���s�=�9J�@���?�/���|+�ڧ�d݆�~��; � =PqM �[�U�S������NN�䦎���J�H�I#s���_����b�X�f�*��7�N��7���\F+n�S��žX�$�'BR4?I��V�7a�S��%��Ĥ�ÙH9�y���[��t�����kE�S�t�H���.Ǹ�2��T��'�o�ؐ	\*�3j��v���a��h�;S�R�[���_t`���h�-��$��bV�?y9�R�����Pd��C�)~�=[�h:`�Els����I5E�|ݤe���s\�c��aπD.#/G���#���.��X���o"[�%	�<O�#p���G.�(����U�;�� X��
���3G�_�nݗflU�1P�|��wv�.1f.���?��,��ұ�&&5��I2�1�`��lyTwؗz����G�2���0c$Y̑���l'\���{�-�~%T��<�O������mX�(;i�j�%��t��2p��9!��d^�qD:l����$\i�SBh>�{ړ�����[q�9�����⊢��NǓ��~�;����!�g�(6GVÀz*���!��)�_�Q���Yĥ69!i���07n]�y��<O��P��s�_˾	��Omv�����$,PR^A���4�&w .�"���� �eY�&j�)ފ�߽^���r�� �x~�LtǴuq�K4���#Ou�+�?�J!�^qr雌'X��Ն8M!l�OfQ�_݅�E68�[�������3�ms���Zך���*)� ���A�krw����Y�q�S��Q��ϊ����O�1��
���	�I�ӟ��ǋ��t03	�
�@�=�)Ze��/nzXK�Pg-���G*=����л�r_��P�|�)U�F����1��F{)�� ��tA,+��x�(@'�V��B����Y��kz�i��ݬ��Ҁ&ñ���_o{�8Q�T0g(E���e�������"�!�D��<%�g@��럳c�c�N�U+���_Uʚ۾}�~���	.r�sG���^V�)�!�dw5��P|Q���΀�t�m6'&�=�LWM#(����w�-5o��f��sJ��g����8�rJ9�f	.43gĵ[K|�w�rͷs:~:�d�?�]3��k�����ӛ�u�u������C+���='@w3������w�;";iA�p.�5C��w�m��V�L���$���\&��f)��A�?�yFb�kp����J?3R���5���h���}��� ����so}��72E��C&\��>�O�͙̊�n��^�C(r`#��t��3�����>f�5/�WN>g�D���n��.��r��:�
��O�QrWֺ��u!��
!��e����:�"����섳�*��d>t�ZU�V���w��e9��w�;?\��h�X�KAT�-��$i��9�o�[�*n�����?{	�<��NFe��P먵m���p�}���=�����Ce�Bɇ�7iQ,';?5��g�{̉�%�.)��vr?��(�����ޛ��/
��F�T�$�̟R�8�L���uB)�J��"[��mB�`�)���$9<��&�v�H�u��#U��<f<�?i�`�W�("y�����S&�c�!~8�	H>�[���f9����eW�2�Aa_�_7�ǵL���OwF>Q���}��ħ[�����	�4��,���kWr?�����&YM�n��rdt��������X���"��cy].�h�/�����g��\�򲼆�vF����ׯ�w����;�^�k���*��z�T���1rz����{;���2���ʙ c��֥�T�e����p�q�nvS�F��S,��<Oy���o�3�����d��^�xxth��'>�K(�ڊ�.Oޯ���#���s��N��lD�Y[��,8�(���إ�Ħ>��-����:���EI���N��/�7t���	P����e6$`1���6-��b�ݼ7�L/��r&Kv��5�q�e�|s����=�ʱpf�+:�Y���pD����7����%�t�VԯPa�����f�5��9��8sy5�C����=�ˇj�h1ՠ��$�K���Ä��"���v#/鄯�4�T)�O8Nbs�}Хb�cb��!��k%ء��X�i�>1�⩖�x�7���.#6��H[�������=�\Ք���Y�{�,��~,���T\:�	���/��AA�_M�	�6آ�'xNOp�����5�2A����Q�׌�}6��'�]�����=Q���$Ă��=I.�&��B��NO��rM��cbl��UKw����l8\�;��+��\�3��i���D�����&�5�YO���OI��J�lp����A����͉�4��S���
��d�����H�4c�BMa����&�F��F��X���2a^�MX�� 2��|�p�
^c9�\/)��[��x�b��5��vk]J$� �C�T.�[��A��jW"c�*e�q�M�E�?�O�ބ��!d���4��tJMg���Щ4����:~�T���p�M�|N$���}��ͿNb��GK��逡[�������a9��Ι�i�XY�-�D�ku}2�}�����Ȝa���x���ΎPʩҜ�X�r�p�n��X�k�WDeM�}���#R�����t��+����X^ab�ib�\uP�3Ѭ7Kp���ǿ�&IRXlS:��4����R����ο5��gf�3�k �ʑ7f�9����웓��/eOe6��/mԷ�e��A<&��0�,���%m;�v���H���#l 	kHB�#��!��,������&벹K�Y:�*x�sMr4�a��_{����G������|_��kU-,�ʰ�Nev$�G��	x,�7A)ͬ:��@���/�0�~7��>T1ҡ/o���?)V�/ ��7ޠ����M뿠~[��)w���-T�?��`�&kDǇG;��RVs�A����s	@y�ڻ�KRLMg v�e�a>�$9�$��>�Qhv�k�f�� ��*'V���(h�:�O�]�;�J[kOR��s�y�6$@!9�d���	�57�=�m d��N���}� q�ũA�W�&���csZƧ��T��<k�1����;���	�Ox�BW;5��\G�9�1��6��Od�.�Lv�}ы���w/-X��F�H��k.����������7��7@D����ӗ܆�m g�
�/��YԙJF�`����[�
KY�Y����۞�htK�L��R����v���Y�s��Fyo��%�CR��W�6'h�0{TW/i�4��4h�o1��Ȍ���[}����T�3rE	��z��?ٓ癔�7��T2�|�y"�^�]� Ȱu�G��G�l���d��:�0��"�c�N��J��C�~@[�{�)�"�(���}W����w�Ks�u�k�h���,siRſ���k�ƐT�B�8s��V=i�v�~����Ɋ�ϳYz�����������$F�o��t,x'82���]�8��J���}H=��-�%��%�!̬�0(�o6���@<I�m ��AP��}&zQ�Yj��d�n ��*�,W�,3Aj����>,�<U���z�T��&Ή�QLWr{g8T1V��֯X���F��㒤���������T�)����b�뀩�����lG��	����k?����pM۔��-Lw�]��4�a�Q��%K=U�{�M�Z��k!gO�1̷}b[�Ɲ�0G� �D�����/�'2�w����Y�|?*LAs�H�3)���%VP�m�����I48X��B����׎-y�8�����������&cG����)�.��1IIʆJBLQ��*�`�<֘
!2���l�*:�`��B�:oK�XO��g��Xs�IUL������m���?k�B�@���q����Q��^�I� B���k"��+S�B��H��e�r��E��-�`�C��7J E�6hB����s�pKW�gk�f����Y6.<��P���f�����U6;�]Ť��E�`��%Z���Ix�t?W6$D"Z|��<�bb>Y]�j�{�И�8�Ψ|�>�UO�s���-�=j��]�N��l�݋�_b����a�քrw�|�)���<�m\�5����[+h��x�y��Ve�4������)���_�l�em2�,K��V���!����{]�ש��Bp���s���d���@�爴�ꑳ��b;��x/��֒�Y-��'h����2����q���
A�R)���`�w��?���f�K��3��0!^tX�s�*��H����{`3�[0	����R��ډ+��?����Є���ҼO����^�Z�~ڼ]��x�z��[(�oՉ����y�'w�
�(ެL�2��!ULE�P�p5���7�jq%$1�[�*q�H?z+����C�A�k�;�ϥn��"��O%�;N�^��U�yu~���
����r�p䓟}�� �i�-��\��%����Y�)5AQ�����#@ M�I���2��Q���gp�e?�0 ڂ	��4GL�)���꼸��mc@��E�uI�@��};���yF�����v��	E�U_0�K�E9�q
��%��ʇ��<�ԧ�h){��@�����K�L�a���;~���.�s��;	"PS�e.S�RԝlѮ�;�T��|&�΍�|^��+Z��רj_�	`�:��"%N��Z�n���<���a�<�ṫ5n��x�ʅ�ìb�#�Z ֵ�c�yl��/�E�+�<n)�Uɺ���&HEd%hc�� ����M?[�#���?���������Meլo
A����l�H���ԒZCVV=2���C�����S�8>w�g�#4?�$��FXrI�ĉ�2A�Lc��mʀO,�Ze�_��~ndJqd����s���۸��9�:�U|�q�3ϘfL��
e?���+.S�e�v����;;���紶��a����&^��r�LWS�\��Y��0���~~�u��qA�U;/�b-�{up�Δ\jG̓s�QQ8r�֦�6�!��I�O���Q�~�^"E
���}��yN�T���~�%��A��tp�r^�+���A-M!�酦���S.h7:BU���mJ(��;eR	�B!��+��Xɽ����$ ���ΰ4yI!���6�
��c��I�%'x#m�K�Y1_�P=U�N�
o���7� U�r����{��2=���)e��r�С:�͟+!;��WCq�!E�t�U���'�����s������ӹb� 01�>�����'t�aq�R�d�o=i��;��g��E�`?�c��;ڼj�o2�4���]%�5�L�O�YNR����7Ρ\FN�uA��@/om���н��a7�Ʉo4X���g�`��bj��=4�)�<y��f���հK�"k����<�ʢ�#r)�0����DG�}?`�P-�mq=���~��H`���q?�a����#}=�cO�M(�O%lٻ��Q�%�0��'��|{
��bLEs`"��O�P)����б��!�=�߉r��*(Y�2&d9�����2�Z�����pOq���1�-C$�Ε���9L�{|�mnU�]S�� ���Mx� �#<�P��v�fK<󅦔�s4����	�]{�`���̷�Ac���P}_zݼ^��ŵN�q�<�r9����	�^����R��@g�V�v�R�}糙�-�S@O��~��mYʹ��[�Y��M¦1<^��&^6�POX}齨��Fb�`��
k�[3Bs�t��vd�gK:z)�oȥ���䳁����W���"�Yȣԧ� |Z�HH���9uy�n�?��,O�\��QbY�<��M+� Cx�:G��F&ş�w�yYk�YNNy��-Ρ"G�������BpCo�Mw]<[�Z�q����ܠ� ���"�R��Oq�=2�xz!!Oq�m�lВ��3�^��S�9��Ϫ�f�jHJv1�w&����p#_�����<��$�]<���t���r� S]�I"kq^9�w[ I� OC\B�ܹ�2�2��Л��~VWv�b���=eO�5x�,�����J:� +4eD������y��
Qc�$�B����(�J�=y�����=����eL�����i�����1:s�,[�Lz`]��%~}���V�.'#}b�p=�ȓ-K�.k�^���
Sk���j��� C̃��$����-�3E��d6{8fԨ���+��\��;d[�)AI�N&�Ia
�z
F�h��L<�U�n!��Q�$x�X䇄�z��E�*��v�VD t����/A^��y���'��DxJ3P���BD<�KQ�fXO:�\�ߡ\�'0�jC!���.VF!�O� x�;.�]%��*�c��M@���\l ����㨮Gz@N�h;p��'�Ҽ%�Š��T��@�|��p׀*l�/��-l=��mb�a�#e8�/��a[�3(Mx�B�T,A=�^h���Eo���?����24�sT6�U��
��}��o9�� ��3=�Aď��z�w�=�����N�����Xk�cB@��='�L�\(�|>�)a3� ��N�P��o%o"���L������6\vm��Ϫtkn���?wW�*�(�f�g��M��:Z����-��p5�~��%+�&�N�в�-'������B�E$�~a���1fB��u�d+��K�S�=j��y-U���n	m*;���*��gA���n�9x��H�?{z�j���\�e�V~�x�/vW/�	�Q�1Ws�c,��	b��k�6q�̨�5�؊�ކ���I^�k@F��)���dF}b���J�H�u��i�)��.20�6�]��D�p�n哬�w��ٵ���0H	=�u��/R_�7oD}�;����#A_cSs��{�$��hEt���:4��
{r^��$xO��E)�dNg�9�_ra�UQaG�~���n�4-��k�v�W'@�֧��̴J�T�1��$5]|W6��aک_3��*{��J�G�[�*Ɠ�T�]ld�����b�!����w��y�?(m�Hb�U�3�w{ z��9�49',��'��?�-���l�x�=��>򑃹��xU~3G���α�����֩�\�S���J����9/���O2%�W�V�m�,�����E�OE�Lᑄ��^�������� �a�A�#����)�G����T5�h�އkd3O!}��˖�ѯK,[�K?�L�������fd�ۦ��a����p����A�1��G����:훙�0OF����o{�J��J���6� \3��ퟚ��7j�1^��^F���@�A��0�� c��h�P#S�; u�H'ؓs/�bt��G+b�il�i�����!9g-",,�4�"{�߾�'�?�����%P̨9�vX�7s\�]�x��)��:e������4?u3{��|*9c�Hg�M�8,�mbm�b�]��R��t�ν�����t���+�I7�^F�S=��P�� C�=��'�b�¿Q�{�a�=����l���lh3A��	%������6���%ov�1���vHp�L�t#T֎����;K�:��5�+�O.)y�
��k�|���^��3T��3�\�����n]v��Q�ҁ-̆ʛ^0�3->�>�L����M��V�FP��{+�gW�O�z��N����Vԋ�7�C�n�K��q���V�xӄ%A��"���N��i�ɏp^?���z��eO���U���/�����,L���gI�%^?�Md�كb�� ���S��W<�

��jcD%���o�l����[5�+�u�4x��Kqb��(Zr���.6���v�)n�'IT�+p:*X��y����%\1B�}IVX��a��:�~��Ә�̣��m�������^�	,��M}�(B\h/�����vy�5oǐ��q?�ԃ�ۙ�8�OU!ag�g�����6J��[��W���t��C�laZ���έ:���9�&�!l�l/���DsʖP���2sƢ�yt���\�	�?pNhZ�M�>trlT�Eݿ6�j*�ǀep�e9��Ȏr�F�V�9�ɞ ��T�~WǡKykZ)�n�x�,�a���]oq��QI�}��I�n�*�a�*�?;�\�7Gi����3Y�y��T��ºb�FA�7�����!��3o�+)<�lo�ќ��z��<�ߨ��3�I>o�u��|�K�"�+�ܟ�swj��}���{�,3�2���`?�:��<ȗ�ߡVD��]w�!��R]�M5�)Qr�6�F�xXo�O7������pl����<�q &����t�(m%'IŰ�&��)��&#!k�ԉ��ۏ����������'ypW� +�zp%EU&�n|���ܩC��1���ΰ���yOUz��{\,���[�)��7I��! *�X�O�%H�s�ed���Y��}œ�⨕_v:���1'�h���p�������id�`�k	�+���+�9Ӷ����FS�/n��T�S��V$Uv���3��-�7M;�{jv�߬�JQ&D�4�}�WRQ�eP�������r��l+��!?c�U@�]@���w0<�h����D}w6X�<�&�
K���$��D�����,TQ�!�JЛj"6�x���H�X�*�b��L�ʁ���